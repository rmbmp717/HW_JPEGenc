module dct_2d_u8(
  input wire clk,
  input wire [511:0] x,
  output wire [511:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [15:0] smul16b_8b_x_8b (input reg [7:0] lhs, input reg [7:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [15:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul16b_8b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_6b (input reg [7:0] lhs, input reg [5:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [16:0] smul17b_8b_x_9b (input reg [7:0] lhs, input reg [8:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [16:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul17b_8b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_7b (input reg [31:0] lhs, input reg [6:0] rhs);
    begin
      umul32b_32b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [7:0] x_unflattened[0:7][0:7];
  assign x_unflattened[0][0] = x[7:0];
  assign x_unflattened[0][1] = x[15:8];
  assign x_unflattened[0][2] = x[23:16];
  assign x_unflattened[0][3] = x[31:24];
  assign x_unflattened[0][4] = x[39:32];
  assign x_unflattened[0][5] = x[47:40];
  assign x_unflattened[0][6] = x[55:48];
  assign x_unflattened[0][7] = x[63:56];
  assign x_unflattened[1][0] = x[71:64];
  assign x_unflattened[1][1] = x[79:72];
  assign x_unflattened[1][2] = x[87:80];
  assign x_unflattened[1][3] = x[95:88];
  assign x_unflattened[1][4] = x[103:96];
  assign x_unflattened[1][5] = x[111:104];
  assign x_unflattened[1][6] = x[119:112];
  assign x_unflattened[1][7] = x[127:120];
  assign x_unflattened[2][0] = x[135:128];
  assign x_unflattened[2][1] = x[143:136];
  assign x_unflattened[2][2] = x[151:144];
  assign x_unflattened[2][3] = x[159:152];
  assign x_unflattened[2][4] = x[167:160];
  assign x_unflattened[2][5] = x[175:168];
  assign x_unflattened[2][6] = x[183:176];
  assign x_unflattened[2][7] = x[191:184];
  assign x_unflattened[3][0] = x[199:192];
  assign x_unflattened[3][1] = x[207:200];
  assign x_unflattened[3][2] = x[215:208];
  assign x_unflattened[3][3] = x[223:216];
  assign x_unflattened[3][4] = x[231:224];
  assign x_unflattened[3][5] = x[239:232];
  assign x_unflattened[3][6] = x[247:240];
  assign x_unflattened[3][7] = x[255:248];
  assign x_unflattened[4][0] = x[263:256];
  assign x_unflattened[4][1] = x[271:264];
  assign x_unflattened[4][2] = x[279:272];
  assign x_unflattened[4][3] = x[287:280];
  assign x_unflattened[4][4] = x[295:288];
  assign x_unflattened[4][5] = x[303:296];
  assign x_unflattened[4][6] = x[311:304];
  assign x_unflattened[4][7] = x[319:312];
  assign x_unflattened[5][0] = x[327:320];
  assign x_unflattened[5][1] = x[335:328];
  assign x_unflattened[5][2] = x[343:336];
  assign x_unflattened[5][3] = x[351:344];
  assign x_unflattened[5][4] = x[359:352];
  assign x_unflattened[5][5] = x[367:360];
  assign x_unflattened[5][6] = x[375:368];
  assign x_unflattened[5][7] = x[383:376];
  assign x_unflattened[6][0] = x[391:384];
  assign x_unflattened[6][1] = x[399:392];
  assign x_unflattened[6][2] = x[407:400];
  assign x_unflattened[6][3] = x[415:408];
  assign x_unflattened[6][4] = x[423:416];
  assign x_unflattened[6][5] = x[431:424];
  assign x_unflattened[6][6] = x[439:432];
  assign x_unflattened[6][7] = x[447:440];
  assign x_unflattened[7][0] = x[455:448];
  assign x_unflattened[7][1] = x[463:456];
  assign x_unflattened[7][2] = x[471:464];
  assign x_unflattened[7][3] = x[479:472];
  assign x_unflattened[7][4] = x[487:480];
  assign x_unflattened[7][5] = x[495:488];
  assign x_unflattened[7][6] = x[503:496];
  assign x_unflattened[7][7] = x[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_x[0:7][0:7];
  always @ (posedge clk) begin
    p0_x[0][0] <= x_unflattened[0][0];
    p0_x[0][1] <= x_unflattened[0][1];
    p0_x[0][2] <= x_unflattened[0][2];
    p0_x[0][3] <= x_unflattened[0][3];
    p0_x[0][4] <= x_unflattened[0][4];
    p0_x[0][5] <= x_unflattened[0][5];
    p0_x[0][6] <= x_unflattened[0][6];
    p0_x[0][7] <= x_unflattened[0][7];
    p0_x[1][0] <= x_unflattened[1][0];
    p0_x[1][1] <= x_unflattened[1][1];
    p0_x[1][2] <= x_unflattened[1][2];
    p0_x[1][3] <= x_unflattened[1][3];
    p0_x[1][4] <= x_unflattened[1][4];
    p0_x[1][5] <= x_unflattened[1][5];
    p0_x[1][6] <= x_unflattened[1][6];
    p0_x[1][7] <= x_unflattened[1][7];
    p0_x[2][0] <= x_unflattened[2][0];
    p0_x[2][1] <= x_unflattened[2][1];
    p0_x[2][2] <= x_unflattened[2][2];
    p0_x[2][3] <= x_unflattened[2][3];
    p0_x[2][4] <= x_unflattened[2][4];
    p0_x[2][5] <= x_unflattened[2][5];
    p0_x[2][6] <= x_unflattened[2][6];
    p0_x[2][7] <= x_unflattened[2][7];
    p0_x[3][0] <= x_unflattened[3][0];
    p0_x[3][1] <= x_unflattened[3][1];
    p0_x[3][2] <= x_unflattened[3][2];
    p0_x[3][3] <= x_unflattened[3][3];
    p0_x[3][4] <= x_unflattened[3][4];
    p0_x[3][5] <= x_unflattened[3][5];
    p0_x[3][6] <= x_unflattened[3][6];
    p0_x[3][7] <= x_unflattened[3][7];
    p0_x[4][0] <= x_unflattened[4][0];
    p0_x[4][1] <= x_unflattened[4][1];
    p0_x[4][2] <= x_unflattened[4][2];
    p0_x[4][3] <= x_unflattened[4][3];
    p0_x[4][4] <= x_unflattened[4][4];
    p0_x[4][5] <= x_unflattened[4][5];
    p0_x[4][6] <= x_unflattened[4][6];
    p0_x[4][7] <= x_unflattened[4][7];
    p0_x[5][0] <= x_unflattened[5][0];
    p0_x[5][1] <= x_unflattened[5][1];
    p0_x[5][2] <= x_unflattened[5][2];
    p0_x[5][3] <= x_unflattened[5][3];
    p0_x[5][4] <= x_unflattened[5][4];
    p0_x[5][5] <= x_unflattened[5][5];
    p0_x[5][6] <= x_unflattened[5][6];
    p0_x[5][7] <= x_unflattened[5][7];
    p0_x[6][0] <= x_unflattened[6][0];
    p0_x[6][1] <= x_unflattened[6][1];
    p0_x[6][2] <= x_unflattened[6][2];
    p0_x[6][3] <= x_unflattened[6][3];
    p0_x[6][4] <= x_unflattened[6][4];
    p0_x[6][5] <= x_unflattened[6][5];
    p0_x[6][6] <= x_unflattened[6][6];
    p0_x[6][7] <= x_unflattened[6][7];
    p0_x[7][0] <= x_unflattened[7][0];
    p0_x[7][1] <= x_unflattened[7][1];
    p0_x[7][2] <= x_unflattened[7][2];
    p0_x[7][3] <= x_unflattened[7][3];
    p0_x[7][4] <= x_unflattened[7][4];
    p0_x[7][5] <= x_unflattened[7][5];
    p0_x[7][6] <= x_unflattened[7][6];
    p0_x[7][7] <= x_unflattened[7][7];
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_array_index_133943_comb;
  wire [7:0] p1_array_index_133944_comb;
  wire [7:0] p1_array_index_133945_comb;
  wire [7:0] p1_array_index_133946_comb;
  wire [7:0] p1_array_index_133965_comb;
  wire [7:0] p1_array_index_133966_comb;
  wire [7:0] p1_array_index_133971_comb;
  wire [7:0] p1_array_index_133972_comb;
  wire [7:0] p1_array_index_133963_comb;
  wire [7:0] p1_array_index_133968_comb;
  wire [7:0] p1_array_index_133969_comb;
  wire [7:0] p1_array_index_133974_comb;
  wire [7:0] p1_array_index_133964_comb;
  wire [7:0] p1_array_index_133967_comb;
  wire [7:0] p1_array_index_133970_comb;
  wire [7:0] p1_array_index_133973_comb;
  wire [7:0] p1_array_index_133923_comb;
  wire [7:0] p1_array_index_133924_comb;
  wire [7:0] p1_array_index_133925_comb;
  wire [7:0] p1_array_index_133926_comb;
  wire [7:0] p1_array_index_133927_comb;
  wire [7:0] p1_array_index_133928_comb;
  wire [7:0] p1_array_index_133929_comb;
  wire [7:0] p1_array_index_133930_comb;
  wire [7:0] p1_array_index_133931_comb;
  wire [7:0] p1_array_index_133932_comb;
  wire [7:0] p1_array_index_133933_comb;
  wire [7:0] p1_array_index_133934_comb;
  wire [7:0] p1_array_index_133935_comb;
  wire [7:0] p1_array_index_133936_comb;
  wire [7:0] p1_array_index_133937_comb;
  wire [7:0] p1_array_index_133938_comb;
  wire [7:0] p1_array_index_133939_comb;
  wire [7:0] p1_array_index_133940_comb;
  wire [7:0] p1_array_index_133941_comb;
  wire [7:0] p1_array_index_133942_comb;
  wire [7:0] p1_array_index_133947_comb;
  wire [7:0] p1_array_index_133948_comb;
  wire [7:0] p1_array_index_133949_comb;
  wire [7:0] p1_array_index_133950_comb;
  wire [7:0] p1_array_index_133951_comb;
  wire [7:0] p1_array_index_133952_comb;
  wire [7:0] p1_array_index_133953_comb;
  wire [7:0] p1_array_index_133954_comb;
  wire [7:0] p1_array_index_133955_comb;
  wire [7:0] p1_array_index_133956_comb;
  wire [7:0] p1_array_index_133957_comb;
  wire [7:0] p1_array_index_133958_comb;
  wire [7:0] p1_array_index_133959_comb;
  wire [7:0] p1_array_index_133960_comb;
  wire [7:0] p1_array_index_133961_comb;
  wire [7:0] p1_array_index_133962_comb;
  wire [7:0] p1_array_index_133975_comb;
  wire [7:0] p1_array_index_133976_comb;
  wire [7:0] p1_array_index_133977_comb;
  wire [7:0] p1_array_index_133978_comb;
  wire [7:0] p1_array_index_133979_comb;
  wire [7:0] p1_array_index_133980_comb;
  wire [7:0] p1_array_index_133981_comb;
  wire [7:0] p1_array_index_133982_comb;
  wire [7:0] p1_array_index_133983_comb;
  wire [7:0] p1_array_index_133984_comb;
  wire [7:0] p1_array_index_133985_comb;
  wire [7:0] p1_array_index_133986_comb;
  wire [7:0] p1_shifted__26_squeezed_comb;
  wire [7:0] p1_shifted__29_squeezed_comb;
  wire [7:0] p1_shifted__34_squeezed_comb;
  wire [7:0] p1_shifted__37_squeezed_comb;
  wire [7:0] p1_shifted__27_squeezed_comb;
  wire [7:0] p1_shifted__28_squeezed_comb;
  wire [7:0] p1_shifted__35_squeezed_comb;
  wire [7:0] p1_shifted__36_squeezed_comb;
  wire [7:0] p1_shifted__24_squeezed_comb;
  wire [7:0] p1_shifted__31_squeezed_comb;
  wire [7:0] p1_shifted__32_squeezed_comb;
  wire [7:0] p1_shifted__39_squeezed_comb;
  wire [7:0] p1_shifted__25_squeezed_comb;
  wire [7:0] p1_shifted__30_squeezed_comb;
  wire [7:0] p1_shifted__33_squeezed_comb;
  wire [7:0] p1_shifted__38_squeezed_comb;
  wire [7:0] p1_shifted__18_squeezed_comb;
  wire [7:0] p1_shifted__21_squeezed_comb;
  wire [7:0] p1_shifted__42_squeezed_comb;
  wire [7:0] p1_shifted__45_squeezed_comb;
  wire [7:0] p1_shifted__16_squeezed_comb;
  wire [7:0] p1_shifted__17_squeezed_comb;
  wire [7:0] p1_shifted__19_squeezed_comb;
  wire [7:0] p1_shifted__20_squeezed_comb;
  wire [7:0] p1_shifted__22_squeezed_comb;
  wire [7:0] p1_shifted__23_squeezed_comb;
  wire [7:0] p1_shifted__40_squeezed_comb;
  wire [7:0] p1_shifted__41_squeezed_comb;
  wire [7:0] p1_shifted__43_squeezed_comb;
  wire [7:0] p1_shifted__44_squeezed_comb;
  wire [7:0] p1_shifted__46_squeezed_comb;
  wire [7:0] p1_shifted__47_squeezed_comb;
  wire [7:0] p1_shifted__2_squeezed_comb;
  wire [7:0] p1_shifted__5_squeezed_comb;
  wire [7:0] p1_shifted__10_squeezed_comb;
  wire [7:0] p1_shifted__13_squeezed_comb;
  wire [7:0] p1_shifted__50_squeezed_comb;
  wire [7:0] p1_shifted__53_squeezed_comb;
  wire [7:0] p1_shifted__58_squeezed_comb;
  wire [7:0] p1_shifted__61_squeezed_comb;
  wire [7:0] p1_shifted_squeezed_comb;
  wire [7:0] p1_shifted__1_squeezed_comb;
  wire [7:0] p1_shifted__3_squeezed_comb;
  wire [7:0] p1_shifted__4_squeezed_comb;
  wire [7:0] p1_shifted__6_squeezed_comb;
  wire [7:0] p1_shifted__7_squeezed_comb;
  wire [7:0] p1_shifted__8_squeezed_comb;
  wire [7:0] p1_shifted__9_squeezed_comb;
  wire [7:0] p1_shifted__11_squeezed_comb;
  wire [7:0] p1_shifted__12_squeezed_comb;
  wire [7:0] p1_shifted__14_squeezed_comb;
  wire [7:0] p1_shifted__15_squeezed_comb;
  wire [7:0] p1_shifted__48_squeezed_comb;
  wire [7:0] p1_shifted__49_squeezed_comb;
  wire [7:0] p1_shifted__51_squeezed_comb;
  wire [7:0] p1_shifted__52_squeezed_comb;
  wire [7:0] p1_shifted__54_squeezed_comb;
  wire [7:0] p1_shifted__55_squeezed_comb;
  wire [7:0] p1_shifted__56_squeezed_comb;
  wire [7:0] p1_shifted__57_squeezed_comb;
  wire [7:0] p1_shifted__59_squeezed_comb;
  wire [7:0] p1_shifted__60_squeezed_comb;
  wire [7:0] p1_shifted__62_squeezed_comb;
  wire [7:0] p1_shifted__63_squeezed_comb;
  wire [15:0] p1_smul_57378_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___12_comb;
  wire [15:0] p1_smul_57384_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___15_comb;
  wire [15:0] p1_smul_57394_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___16_comb;
  wire [15:0] p1_smul_57400_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___19_comb;
  wire [15:0] p1_smul_57636_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___77_comb;
  wire [15:0] p1_smul_57638_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___78_comb;
  wire [15:0] p1_smul_57652_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___81_comb;
  wire [15:0] p1_smul_57654_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___82_comb;
  wire [15:0] p1_smul_57886_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___108_comb;
  wire [15:0] p1_smul_57900_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___111_comb;
  wire [15:0] p1_smul_57902_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___112_comb;
  wire [15:0] p1_smul_57916_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___115_comb;
  wire [15:0] p1_smul_58144_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___173_comb;
  wire [15:0] p1_smul_58154_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___174_comb;
  wire [15:0] p1_smul_58160_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___177_comb;
  wire [15:0] p1_smul_58170_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___178_comb;
  wire [7:0] p1_smul_57326_TrailingBits___144_comb;
  wire [7:0] p1_smul_57326_TrailingBits___145_comb;
  wire [7:0] p1_smul_57326_TrailingBits___146_comb;
  wire [7:0] p1_smul_57326_TrailingBits___147_comb;
  wire [7:0] p1_smul_57326_TrailingBits___148_comb;
  wire [7:0] p1_smul_57326_TrailingBits___149_comb;
  wire [7:0] p1_smul_57326_TrailingBits___150_comb;
  wire [7:0] p1_smul_57326_TrailingBits___151_comb;
  wire [7:0] p1_smul_57326_TrailingBits___168_comb;
  wire [7:0] p1_smul_57326_TrailingBits___169_comb;
  wire [7:0] p1_smul_57326_TrailingBits___170_comb;
  wire [7:0] p1_smul_57326_TrailingBits___171_comb;
  wire [7:0] p1_smul_57326_TrailingBits___172_comb;
  wire [7:0] p1_smul_57326_TrailingBits___173_comb;
  wire [7:0] p1_smul_57326_TrailingBits___174_comb;
  wire [7:0] p1_smul_57326_TrailingBits___175_comb;
  wire [7:0] p1_smul_57326_TrailingBits___128_comb;
  wire [7:0] p1_smul_57326_TrailingBits___129_comb;
  wire [7:0] p1_smul_57326_TrailingBits___130_comb;
  wire [7:0] p1_smul_57326_TrailingBits___131_comb;
  wire [7:0] p1_smul_57326_TrailingBits___132_comb;
  wire [7:0] p1_smul_57326_TrailingBits___133_comb;
  wire [7:0] p1_smul_57326_TrailingBits___134_comb;
  wire [7:0] p1_smul_57326_TrailingBits___135_comb;
  wire [7:0] p1_smul_57326_TrailingBits___136_comb;
  wire [7:0] p1_smul_57326_TrailingBits___137_comb;
  wire [7:0] p1_smul_57326_TrailingBits___138_comb;
  wire [7:0] p1_smul_57326_TrailingBits___139_comb;
  wire [7:0] p1_smul_57326_TrailingBits___140_comb;
  wire [7:0] p1_smul_57326_TrailingBits___141_comb;
  wire [7:0] p1_smul_57326_TrailingBits___142_comb;
  wire [7:0] p1_smul_57326_TrailingBits___143_comb;
  wire [7:0] p1_smul_57326_TrailingBits___152_comb;
  wire [7:0] p1_smul_57326_TrailingBits___153_comb;
  wire [7:0] p1_smul_57326_TrailingBits___154_comb;
  wire [7:0] p1_smul_57326_TrailingBits___155_comb;
  wire [7:0] p1_smul_57326_TrailingBits___156_comb;
  wire [7:0] p1_smul_57326_TrailingBits___157_comb;
  wire [7:0] p1_smul_57326_TrailingBits___158_comb;
  wire [7:0] p1_smul_57326_TrailingBits___159_comb;
  wire [7:0] p1_smul_57326_TrailingBits___160_comb;
  wire [7:0] p1_smul_57326_TrailingBits___161_comb;
  wire [7:0] p1_smul_57326_TrailingBits___162_comb;
  wire [7:0] p1_smul_57326_TrailingBits___163_comb;
  wire [7:0] p1_smul_57326_TrailingBits___164_comb;
  wire [7:0] p1_smul_57326_TrailingBits___165_comb;
  wire [7:0] p1_smul_57326_TrailingBits___166_comb;
  wire [7:0] p1_smul_57326_TrailingBits___167_comb;
  wire [7:0] p1_smul_57326_TrailingBits___176_comb;
  wire [7:0] p1_smul_57326_TrailingBits___177_comb;
  wire [7:0] p1_smul_57326_TrailingBits___178_comb;
  wire [7:0] p1_smul_57326_TrailingBits___179_comb;
  wire [7:0] p1_smul_57326_TrailingBits___180_comb;
  wire [7:0] p1_smul_57326_TrailingBits___181_comb;
  wire [7:0] p1_smul_57326_TrailingBits___182_comb;
  wire [7:0] p1_smul_57326_TrailingBits___183_comb;
  wire [7:0] p1_smul_57326_TrailingBits___184_comb;
  wire [7:0] p1_smul_57326_TrailingBits___185_comb;
  wire [7:0] p1_smul_57326_TrailingBits___186_comb;
  wire [7:0] p1_smul_57326_TrailingBits___187_comb;
  wire [7:0] p1_smul_57326_TrailingBits___188_comb;
  wire [7:0] p1_smul_57326_TrailingBits___189_comb;
  wire [7:0] p1_smul_57326_TrailingBits___190_comb;
  wire [7:0] p1_smul_57326_TrailingBits___191_comb;
  wire [15:0] p1_smul_57362_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___8_comb;
  wire [15:0] p1_smul_57368_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___11_comb;
  wire [15:0] p1_smul_57410_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___20_comb;
  wire [15:0] p1_smul_57416_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___23_comb;
  wire [14:0] p1_smul_57486_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___8_comb;
  wire [14:0] p1_smul_57488_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___40_comb;
  wire [14:0] p1_smul_57490_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___41_comb;
  wire [14:0] p1_smul_57492_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___9_comb;
  wire [14:0] p1_smul_57494_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___10_comb;
  wire [14:0] p1_smul_57496_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___42_comb;
  wire [14:0] p1_smul_57498_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___43_comb;
  wire [14:0] p1_smul_57500_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___11_comb;
  wire [14:0] p1_smul_57534_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___20_comb;
  wire [14:0] p1_smul_57536_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___52_comb;
  wire [14:0] p1_smul_57538_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___53_comb;
  wire [14:0] p1_smul_57540_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___21_comb;
  wire [14:0] p1_smul_57542_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___22_comb;
  wire [14:0] p1_smul_57544_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___54_comb;
  wire [14:0] p1_smul_57546_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___55_comb;
  wire [14:0] p1_smul_57548_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___23_comb;
  wire [15:0] p1_smul_57620_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___73_comb;
  wire [15:0] p1_smul_57622_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___74_comb;
  wire [15:0] p1_smul_57668_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___85_comb;
  wire [15:0] p1_smul_57670_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___86_comb;
  wire [15:0] p1_smul_57870_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___104_comb;
  wire [15:0] p1_smul_57884_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___107_comb;
  wire [15:0] p1_smul_57918_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___116_comb;
  wire [15:0] p1_smul_57932_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___119_comb;
  wire [14:0] p1_smul_57998_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___136_comb;
  wire [14:0] p1_smul_58000_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___40_comb;
  wire [14:0] p1_smul_58002_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___137_comb;
  wire [14:0] p1_smul_58004_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___41_comb;
  wire [14:0] p1_smul_58006_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___42_comb;
  wire [14:0] p1_smul_58008_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___138_comb;
  wire [14:0] p1_smul_58010_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___43_comb;
  wire [14:0] p1_smul_58012_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___139_comb;
  wire [14:0] p1_smul_58046_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___148_comb;
  wire [14:0] p1_smul_58048_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___52_comb;
  wire [14:0] p1_smul_58050_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___149_comb;
  wire [14:0] p1_smul_58052_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___53_comb;
  wire [14:0] p1_smul_58054_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___54_comb;
  wire [14:0] p1_smul_58056_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___150_comb;
  wire [14:0] p1_smul_58058_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___55_comb;
  wire [14:0] p1_smul_58060_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___151_comb;
  wire [15:0] p1_smul_58128_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___169_comb;
  wire [15:0] p1_smul_58138_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___170_comb;
  wire [15:0] p1_smul_58176_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___181_comb;
  wire [15:0] p1_smul_58186_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___182_comb;
  wire [15:0] p1_smul_57330_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits__comb;
  wire [15:0] p1_smul_57336_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___3_comb;
  wire [15:0] p1_smul_57346_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___4_comb;
  wire [15:0] p1_smul_57352_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___7_comb;
  wire [15:0] p1_smul_57426_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___24_comb;
  wire [15:0] p1_smul_57432_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___27_comb;
  wire [15:0] p1_smul_57442_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___28_comb;
  wire [15:0] p1_smul_57448_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___31_comb;
  wire [14:0] p1_smul_57454_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits__comb;
  wire [14:0] p1_smul_57456_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___32_comb;
  wire [14:0] p1_smul_57458_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___33_comb;
  wire [14:0] p1_smul_57460_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___1_comb;
  wire [14:0] p1_smul_57462_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___2_comb;
  wire [14:0] p1_smul_57464_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___34_comb;
  wire [14:0] p1_smul_57466_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___35_comb;
  wire [14:0] p1_smul_57468_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___3_comb;
  wire [14:0] p1_smul_57470_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___4_comb;
  wire [14:0] p1_smul_57472_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___36_comb;
  wire [14:0] p1_smul_57474_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___37_comb;
  wire [14:0] p1_smul_57476_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___5_comb;
  wire [14:0] p1_smul_57478_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___6_comb;
  wire [14:0] p1_smul_57480_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___38_comb;
  wire [14:0] p1_smul_57482_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___39_comb;
  wire [14:0] p1_smul_57484_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___7_comb;
  wire [14:0] p1_smul_57502_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___12_comb;
  wire [14:0] p1_smul_57504_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___44_comb;
  wire [14:0] p1_smul_57506_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___45_comb;
  wire [14:0] p1_smul_57508_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___13_comb;
  wire [14:0] p1_smul_57510_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___14_comb;
  wire [14:0] p1_smul_57512_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___46_comb;
  wire [14:0] p1_smul_57514_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___47_comb;
  wire [14:0] p1_smul_57516_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___15_comb;
  wire [14:0] p1_smul_57518_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___16_comb;
  wire [14:0] p1_smul_57520_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___48_comb;
  wire [14:0] p1_smul_57522_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___49_comb;
  wire [14:0] p1_smul_57524_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___17_comb;
  wire [14:0] p1_smul_57526_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___18_comb;
  wire [14:0] p1_smul_57528_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___50_comb;
  wire [14:0] p1_smul_57530_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___51_comb;
  wire [14:0] p1_smul_57532_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___19_comb;
  wire [14:0] p1_smul_57550_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___24_comb;
  wire [14:0] p1_smul_57552_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___56_comb;
  wire [14:0] p1_smul_57554_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___57_comb;
  wire [14:0] p1_smul_57556_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___25_comb;
  wire [14:0] p1_smul_57558_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___26_comb;
  wire [14:0] p1_smul_57560_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___58_comb;
  wire [14:0] p1_smul_57562_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___59_comb;
  wire [14:0] p1_smul_57564_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___27_comb;
  wire [14:0] p1_smul_57566_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___28_comb;
  wire [14:0] p1_smul_57568_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___60_comb;
  wire [14:0] p1_smul_57570_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___61_comb;
  wire [14:0] p1_smul_57572_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___29_comb;
  wire [14:0] p1_smul_57574_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___30_comb;
  wire [14:0] p1_smul_57576_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___62_comb;
  wire [14:0] p1_smul_57578_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___63_comb;
  wire [14:0] p1_smul_57580_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___31_comb;
  wire [15:0] p1_smul_57588_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___65_comb;
  wire [15:0] p1_smul_57590_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___66_comb;
  wire [15:0] p1_smul_57604_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___69_comb;
  wire [15:0] p1_smul_57606_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___70_comb;
  wire [15:0] p1_smul_57684_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___89_comb;
  wire [15:0] p1_smul_57686_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___90_comb;
  wire [15:0] p1_smul_57700_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___93_comb;
  wire [15:0] p1_smul_57702_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___94_comb;
  wire [15:0] p1_smul_57838_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___96_comb;
  wire [15:0] p1_smul_57852_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___99_comb;
  wire [15:0] p1_smul_57854_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___100_comb;
  wire [15:0] p1_smul_57868_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___103_comb;
  wire [15:0] p1_smul_57934_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___120_comb;
  wire [15:0] p1_smul_57948_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___123_comb;
  wire [15:0] p1_smul_57950_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___124_comb;
  wire [15:0] p1_smul_57964_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___127_comb;
  wire [14:0] p1_smul_57966_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___128_comb;
  wire [14:0] p1_smul_57968_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___32_comb;
  wire [14:0] p1_smul_57970_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___129_comb;
  wire [14:0] p1_smul_57972_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___33_comb;
  wire [14:0] p1_smul_57974_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___34_comb;
  wire [14:0] p1_smul_57976_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___130_comb;
  wire [14:0] p1_smul_57978_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___35_comb;
  wire [14:0] p1_smul_57980_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___131_comb;
  wire [14:0] p1_smul_57982_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___132_comb;
  wire [14:0] p1_smul_57984_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___36_comb;
  wire [14:0] p1_smul_57986_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___133_comb;
  wire [14:0] p1_smul_57988_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___37_comb;
  wire [14:0] p1_smul_57990_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___38_comb;
  wire [14:0] p1_smul_57992_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___134_comb;
  wire [14:0] p1_smul_57994_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___39_comb;
  wire [14:0] p1_smul_57996_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___135_comb;
  wire [14:0] p1_smul_58014_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___140_comb;
  wire [14:0] p1_smul_58016_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___44_comb;
  wire [14:0] p1_smul_58018_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___141_comb;
  wire [14:0] p1_smul_58020_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___45_comb;
  wire [14:0] p1_smul_58022_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___46_comb;
  wire [14:0] p1_smul_58024_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___142_comb;
  wire [14:0] p1_smul_58026_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___47_comb;
  wire [14:0] p1_smul_58028_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___143_comb;
  wire [14:0] p1_smul_58030_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___144_comb;
  wire [14:0] p1_smul_58032_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___48_comb;
  wire [14:0] p1_smul_58034_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___145_comb;
  wire [14:0] p1_smul_58036_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___49_comb;
  wire [14:0] p1_smul_58038_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___50_comb;
  wire [14:0] p1_smul_58040_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___146_comb;
  wire [14:0] p1_smul_58042_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___51_comb;
  wire [14:0] p1_smul_58044_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___147_comb;
  wire [14:0] p1_smul_58062_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___152_comb;
  wire [14:0] p1_smul_58064_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___56_comb;
  wire [14:0] p1_smul_58066_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___153_comb;
  wire [14:0] p1_smul_58068_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___57_comb;
  wire [14:0] p1_smul_58070_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___58_comb;
  wire [14:0] p1_smul_58072_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___154_comb;
  wire [14:0] p1_smul_58074_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___59_comb;
  wire [14:0] p1_smul_58076_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___155_comb;
  wire [14:0] p1_smul_58078_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___156_comb;
  wire [14:0] p1_smul_58080_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___60_comb;
  wire [14:0] p1_smul_58082_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___157_comb;
  wire [14:0] p1_smul_58084_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___61_comb;
  wire [14:0] p1_smul_58086_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___62_comb;
  wire [14:0] p1_smul_58088_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___158_comb;
  wire [14:0] p1_smul_58090_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___63_comb;
  wire [14:0] p1_smul_58092_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___159_comb;
  wire [15:0] p1_smul_58096_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___161_comb;
  wire [15:0] p1_smul_58106_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___162_comb;
  wire [15:0] p1_smul_58112_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___165_comb;
  wire [15:0] p1_smul_58122_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___166_comb;
  wire [15:0] p1_smul_58192_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___185_comb;
  wire [15:0] p1_smul_58202_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___186_comb;
  wire [15:0] p1_smul_58208_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___189_comb;
  wire [15:0] p1_smul_58218_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___190_comb;
  wire [24:0] p1_concat_135019_comb;
  wire [13:0] p1_smul_57380_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___13_comb;
  wire [13:0] p1_smul_57382_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___14_comb;
  wire [24:0] p1_concat_135024_comb;
  wire [24:0] p1_concat_135025_comb;
  wire [13:0] p1_smul_57396_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___17_comb;
  wire [13:0] p1_smul_57398_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___18_comb;
  wire [24:0] p1_concat_135030_comb;
  wire [13:0] p1_smul_57632_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___76_comb;
  wire [24:0] p1_concat_135097_comb;
  wire [24:0] p1_concat_135098_comb;
  wire [13:0] p1_smul_57642_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___79_comb;
  wire [13:0] p1_smul_57648_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___80_comb;
  wire [24:0] p1_concat_135103_comb;
  wire [24:0] p1_concat_135104_comb;
  wire [13:0] p1_smul_57658_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___83_comb;
  wire [24:0] p1_concat_135123_comb;
  wire [13:0] p1_smul_57890_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___109_comb;
  wire [13:0] p1_smul_57896_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___110_comb;
  wire [24:0] p1_concat_135128_comb;
  wire [24:0] p1_concat_135129_comb;
  wire [13:0] p1_smul_57906_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___113_comb;
  wire [13:0] p1_smul_57912_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___114_comb;
  wire [24:0] p1_concat_135134_comb;
  wire [13:0] p1_smul_58142_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___172_comb;
  wire [24:0] p1_concat_135201_comb;
  wire [24:0] p1_concat_135202_comb;
  wire [13:0] p1_smul_58156_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___175_comb;
  wire [13:0] p1_smul_58158_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___176_comb;
  wire [24:0] p1_concat_135207_comb;
  wire [24:0] p1_concat_135208_comb;
  wire [13:0] p1_smul_58172_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___179_comb;
  wire [15:0] p1_shifted__16_comb;
  wire [15:0] p1_shifted__17_comb;
  wire [15:0] p1_shifted__18_comb;
  wire [15:0] p1_shifted__19_comb;
  wire [15:0] p1_shifted__20_comb;
  wire [15:0] p1_shifted__21_comb;
  wire [15:0] p1_shifted__22_comb;
  wire [15:0] p1_shifted__23_comb;
  wire [15:0] p1_shifted__40_comb;
  wire [15:0] p1_shifted__41_comb;
  wire [15:0] p1_shifted__42_comb;
  wire [15:0] p1_shifted__43_comb;
  wire [15:0] p1_shifted__44_comb;
  wire [15:0] p1_shifted__45_comb;
  wire [15:0] p1_shifted__46_comb;
  wire [15:0] p1_shifted__47_comb;
  wire [15:0] p1_shifted_comb;
  wire [15:0] p1_shifted__1_comb;
  wire [15:0] p1_shifted__2_comb;
  wire [15:0] p1_shifted__3_comb;
  wire [15:0] p1_shifted__4_comb;
  wire [15:0] p1_shifted__5_comb;
  wire [15:0] p1_shifted__6_comb;
  wire [15:0] p1_shifted__7_comb;
  wire [15:0] p1_shifted__8_comb;
  wire [15:0] p1_shifted__9_comb;
  wire [15:0] p1_shifted__10_comb;
  wire [15:0] p1_shifted__11_comb;
  wire [15:0] p1_shifted__12_comb;
  wire [15:0] p1_shifted__13_comb;
  wire [15:0] p1_shifted__14_comb;
  wire [15:0] p1_shifted__15_comb;
  wire [15:0] p1_shifted__24_comb;
  wire [15:0] p1_shifted__25_comb;
  wire [15:0] p1_shifted__26_comb;
  wire [15:0] p1_shifted__27_comb;
  wire [15:0] p1_shifted__28_comb;
  wire [15:0] p1_shifted__29_comb;
  wire [15:0] p1_shifted__30_comb;
  wire [15:0] p1_shifted__31_comb;
  wire [15:0] p1_shifted__32_comb;
  wire [15:0] p1_shifted__33_comb;
  wire [15:0] p1_shifted__34_comb;
  wire [15:0] p1_shifted__35_comb;
  wire [15:0] p1_shifted__36_comb;
  wire [15:0] p1_shifted__37_comb;
  wire [15:0] p1_shifted__38_comb;
  wire [15:0] p1_shifted__39_comb;
  wire [15:0] p1_shifted__48_comb;
  wire [15:0] p1_shifted__49_comb;
  wire [15:0] p1_shifted__50_comb;
  wire [15:0] p1_shifted__51_comb;
  wire [15:0] p1_shifted__52_comb;
  wire [15:0] p1_shifted__53_comb;
  wire [15:0] p1_shifted__54_comb;
  wire [15:0] p1_shifted__55_comb;
  wire [15:0] p1_shifted__56_comb;
  wire [15:0] p1_shifted__57_comb;
  wire [15:0] p1_shifted__58_comb;
  wire [15:0] p1_shifted__59_comb;
  wire [15:0] p1_shifted__60_comb;
  wire [15:0] p1_shifted__61_comb;
  wire [15:0] p1_shifted__62_comb;
  wire [15:0] p1_shifted__63_comb;
  wire [24:0] p1_concat_134899_comb;
  wire [13:0] p1_smul_57364_NarrowedMult__comb;
  wire [13:0] p1_smul_57366_NarrowedMult__comb;
  wire [24:0] p1_concat_134902_comb;
  wire [24:0] p1_concat_134903_comb;
  wire [13:0] p1_smul_57412_NarrowedMult__comb;
  wire [13:0] p1_smul_57414_NarrowedMult__comb;
  wire [24:0] p1_concat_134906_comb;
  wire [24:0] p1_concat_134907_comb;
  wire [23:0] p1_concat_134908_comb;
  wire [23:0] p1_concat_134909_comb;
  wire [24:0] p1_concat_134910_comb;
  wire [24:0] p1_concat_134911_comb;
  wire [23:0] p1_concat_134912_comb;
  wire [23:0] p1_concat_134913_comb;
  wire [24:0] p1_concat_134914_comb;
  wire [24:0] p1_concat_134915_comb;
  wire [23:0] p1_concat_134916_comb;
  wire [23:0] p1_concat_134917_comb;
  wire [24:0] p1_concat_134918_comb;
  wire [24:0] p1_concat_134919_comb;
  wire [23:0] p1_concat_134920_comb;
  wire [23:0] p1_concat_134921_comb;
  wire [24:0] p1_concat_134922_comb;
  wire [13:0] p1_smul_57616_NarrowedMult__comb;
  wire [24:0] p1_concat_134924_comb;
  wire [24:0] p1_concat_134925_comb;
  wire [13:0] p1_smul_57626_NarrowedMult__comb;
  wire [13:0] p1_smul_57664_NarrowedMult__comb;
  wire [24:0] p1_concat_134928_comb;
  wire [24:0] p1_concat_134929_comb;
  wire [13:0] p1_smul_57674_NarrowedMult__comb;
  wire [24:0] p1_concat_134931_comb;
  wire [13:0] p1_smul_57874_NarrowedMult__comb;
  wire [13:0] p1_smul_57880_NarrowedMult__comb;
  wire [24:0] p1_concat_134934_comb;
  wire [24:0] p1_concat_134935_comb;
  wire [13:0] p1_smul_57922_NarrowedMult__comb;
  wire [13:0] p1_smul_57928_NarrowedMult__comb;
  wire [24:0] p1_concat_134938_comb;
  wire [23:0] p1_concat_134939_comb;
  wire [24:0] p1_concat_134940_comb;
  wire [23:0] p1_concat_134941_comb;
  wire [24:0] p1_concat_134942_comb;
  wire [24:0] p1_concat_134943_comb;
  wire [23:0] p1_concat_134944_comb;
  wire [24:0] p1_concat_134945_comb;
  wire [23:0] p1_concat_134946_comb;
  wire [23:0] p1_concat_134947_comb;
  wire [24:0] p1_concat_134948_comb;
  wire [23:0] p1_concat_134949_comb;
  wire [24:0] p1_concat_134950_comb;
  wire [24:0] p1_concat_134951_comb;
  wire [23:0] p1_concat_134952_comb;
  wire [24:0] p1_concat_134953_comb;
  wire [23:0] p1_concat_134954_comb;
  wire [13:0] p1_smul_58126_NarrowedMult__comb;
  wire [24:0] p1_concat_134956_comb;
  wire [24:0] p1_concat_134957_comb;
  wire [13:0] p1_smul_58140_NarrowedMult__comb;
  wire [13:0] p1_smul_58174_NarrowedMult__comb;
  wire [24:0] p1_concat_134960_comb;
  wire [24:0] p1_concat_134961_comb;
  wire [13:0] p1_smul_58188_NarrowedMult__comb;
  wire [24:0] p1_concat_135011_comb;
  wire [13:0] p1_smul_57332_NarrowedMult__comb;
  wire [13:0] p1_smul_57334_NarrowedMult__comb;
  wire [24:0] p1_concat_135014_comb;
  wire [24:0] p1_concat_135015_comb;
  wire [13:0] p1_smul_57348_NarrowedMult__comb;
  wire [13:0] p1_smul_57350_NarrowedMult__comb;
  wire [24:0] p1_concat_135018_comb;
  wire [24:0] p1_concat_135031_comb;
  wire [13:0] p1_smul_57428_NarrowedMult__comb;
  wire [13:0] p1_smul_57430_NarrowedMult__comb;
  wire [24:0] p1_concat_135034_comb;
  wire [24:0] p1_concat_135035_comb;
  wire [13:0] p1_smul_57444_NarrowedMult__comb;
  wire [13:0] p1_smul_57446_NarrowedMult__comb;
  wire [24:0] p1_concat_135038_comb;
  wire [24:0] p1_concat_135039_comb;
  wire [23:0] p1_concat_135040_comb;
  wire [23:0] p1_concat_135041_comb;
  wire [24:0] p1_concat_135042_comb;
  wire [24:0] p1_concat_135043_comb;
  wire [23:0] p1_concat_135044_comb;
  wire [23:0] p1_concat_135045_comb;
  wire [24:0] p1_concat_135046_comb;
  wire [24:0] p1_concat_135047_comb;
  wire [23:0] p1_concat_135048_comb;
  wire [23:0] p1_concat_135049_comb;
  wire [24:0] p1_concat_135050_comb;
  wire [24:0] p1_concat_135051_comb;
  wire [23:0] p1_concat_135052_comb;
  wire [23:0] p1_concat_135053_comb;
  wire [24:0] p1_concat_135054_comb;
  wire [24:0] p1_concat_135055_comb;
  wire [23:0] p1_concat_135056_comb;
  wire [23:0] p1_concat_135057_comb;
  wire [24:0] p1_concat_135058_comb;
  wire [24:0] p1_concat_135059_comb;
  wire [23:0] p1_concat_135060_comb;
  wire [23:0] p1_concat_135061_comb;
  wire [24:0] p1_concat_135062_comb;
  wire [24:0] p1_concat_135063_comb;
  wire [23:0] p1_concat_135064_comb;
  wire [23:0] p1_concat_135065_comb;
  wire [24:0] p1_concat_135066_comb;
  wire [24:0] p1_concat_135067_comb;
  wire [23:0] p1_concat_135068_comb;
  wire [23:0] p1_concat_135069_comb;
  wire [24:0] p1_concat_135070_comb;
  wire [24:0] p1_concat_135071_comb;
  wire [23:0] p1_concat_135072_comb;
  wire [23:0] p1_concat_135073_comb;
  wire [24:0] p1_concat_135074_comb;
  wire [24:0] p1_concat_135075_comb;
  wire [23:0] p1_concat_135076_comb;
  wire [23:0] p1_concat_135077_comb;
  wire [24:0] p1_concat_135078_comb;
  wire [24:0] p1_concat_135079_comb;
  wire [23:0] p1_concat_135080_comb;
  wire [23:0] p1_concat_135081_comb;
  wire [24:0] p1_concat_135082_comb;
  wire [24:0] p1_concat_135083_comb;
  wire [23:0] p1_concat_135084_comb;
  wire [23:0] p1_concat_135085_comb;
  wire [24:0] p1_concat_135086_comb;
  wire [13:0] p1_smul_57584_NarrowedMult__comb;
  wire [24:0] p1_concat_135088_comb;
  wire [24:0] p1_concat_135089_comb;
  wire [13:0] p1_smul_57594_NarrowedMult__comb;
  wire [13:0] p1_smul_57600_NarrowedMult__comb;
  wire [24:0] p1_concat_135092_comb;
  wire [24:0] p1_concat_135093_comb;
  wire [13:0] p1_smul_57610_NarrowedMult__comb;
  wire [13:0] p1_smul_57680_NarrowedMult__comb;
  wire [24:0] p1_concat_135108_comb;
  wire [24:0] p1_concat_135109_comb;
  wire [13:0] p1_smul_57690_NarrowedMult__comb;
  wire [13:0] p1_smul_57696_NarrowedMult__comb;
  wire [24:0] p1_concat_135112_comb;
  wire [24:0] p1_concat_135113_comb;
  wire [13:0] p1_smul_57706_NarrowedMult__comb;
  wire [24:0] p1_concat_135115_comb;
  wire [13:0] p1_smul_57842_NarrowedMult__comb;
  wire [13:0] p1_smul_57848_NarrowedMult__comb;
  wire [24:0] p1_concat_135118_comb;
  wire [24:0] p1_concat_135119_comb;
  wire [13:0] p1_smul_57858_NarrowedMult__comb;
  wire [13:0] p1_smul_57864_NarrowedMult__comb;
  wire [24:0] p1_concat_135122_comb;
  wire [24:0] p1_concat_135135_comb;
  wire [13:0] p1_smul_57938_NarrowedMult__comb;
  wire [13:0] p1_smul_57944_NarrowedMult__comb;
  wire [24:0] p1_concat_135138_comb;
  wire [24:0] p1_concat_135139_comb;
  wire [13:0] p1_smul_57954_NarrowedMult__comb;
  wire [13:0] p1_smul_57960_NarrowedMult__comb;
  wire [24:0] p1_concat_135142_comb;
  wire [23:0] p1_concat_135143_comb;
  wire [24:0] p1_concat_135144_comb;
  wire [23:0] p1_concat_135145_comb;
  wire [24:0] p1_concat_135146_comb;
  wire [24:0] p1_concat_135147_comb;
  wire [23:0] p1_concat_135148_comb;
  wire [24:0] p1_concat_135149_comb;
  wire [23:0] p1_concat_135150_comb;
  wire [23:0] p1_concat_135151_comb;
  wire [24:0] p1_concat_135152_comb;
  wire [23:0] p1_concat_135153_comb;
  wire [24:0] p1_concat_135154_comb;
  wire [24:0] p1_concat_135155_comb;
  wire [23:0] p1_concat_135156_comb;
  wire [24:0] p1_concat_135157_comb;
  wire [23:0] p1_concat_135158_comb;
  wire [23:0] p1_concat_135159_comb;
  wire [24:0] p1_concat_135160_comb;
  wire [23:0] p1_concat_135161_comb;
  wire [24:0] p1_concat_135162_comb;
  wire [24:0] p1_concat_135163_comb;
  wire [23:0] p1_concat_135164_comb;
  wire [24:0] p1_concat_135165_comb;
  wire [23:0] p1_concat_135166_comb;
  wire [23:0] p1_concat_135167_comb;
  wire [24:0] p1_concat_135168_comb;
  wire [23:0] p1_concat_135169_comb;
  wire [24:0] p1_concat_135170_comb;
  wire [24:0] p1_concat_135171_comb;
  wire [23:0] p1_concat_135172_comb;
  wire [24:0] p1_concat_135173_comb;
  wire [23:0] p1_concat_135174_comb;
  wire [23:0] p1_concat_135175_comb;
  wire [24:0] p1_concat_135176_comb;
  wire [23:0] p1_concat_135177_comb;
  wire [24:0] p1_concat_135178_comb;
  wire [24:0] p1_concat_135179_comb;
  wire [23:0] p1_concat_135180_comb;
  wire [24:0] p1_concat_135181_comb;
  wire [23:0] p1_concat_135182_comb;
  wire [23:0] p1_concat_135183_comb;
  wire [24:0] p1_concat_135184_comb;
  wire [23:0] p1_concat_135185_comb;
  wire [24:0] p1_concat_135186_comb;
  wire [24:0] p1_concat_135187_comb;
  wire [23:0] p1_concat_135188_comb;
  wire [24:0] p1_concat_135189_comb;
  wire [23:0] p1_concat_135190_comb;
  wire [13:0] p1_smul_58094_NarrowedMult__comb;
  wire [24:0] p1_concat_135192_comb;
  wire [24:0] p1_concat_135193_comb;
  wire [13:0] p1_smul_58108_NarrowedMult__comb;
  wire [13:0] p1_smul_58110_NarrowedMult__comb;
  wire [24:0] p1_concat_135196_comb;
  wire [24:0] p1_concat_135197_comb;
  wire [13:0] p1_smul_58124_NarrowedMult__comb;
  wire [13:0] p1_smul_58190_NarrowedMult__comb;
  wire [24:0] p1_concat_135212_comb;
  wire [24:0] p1_concat_135213_comb;
  wire [13:0] p1_smul_58204_NarrowedMult__comb;
  wire [13:0] p1_smul_58206_NarrowedMult__comb;
  wire [24:0] p1_concat_135216_comb;
  wire [24:0] p1_concat_135217_comb;
  wire [13:0] p1_smul_58220_NarrowedMult__comb;
  wire p1_slt_135220_comb;
  wire p1_slt_135222_comb;
  wire p1_slt_135224_comb;
  wire p1_slt_135226_comb;
  wire p1_slt_135228_comb;
  wire p1_slt_135230_comb;
  wire p1_slt_135232_comb;
  wire p1_slt_135234_comb;
  wire p1_slt_135236_comb;
  wire p1_slt_135238_comb;
  wire p1_slt_135240_comb;
  wire p1_slt_135242_comb;
  wire p1_slt_135244_comb;
  wire p1_slt_135246_comb;
  wire p1_slt_135248_comb;
  wire p1_slt_135250_comb;
  wire p1_slt_135252_comb;
  wire p1_slt_135254_comb;
  wire p1_slt_135256_comb;
  wire p1_slt_135258_comb;
  wire p1_slt_135260_comb;
  wire p1_slt_135262_comb;
  wire p1_slt_135264_comb;
  wire p1_slt_135266_comb;
  wire p1_slt_135268_comb;
  wire p1_slt_135270_comb;
  wire p1_slt_135272_comb;
  wire p1_slt_135274_comb;
  wire p1_slt_135276_comb;
  wire p1_slt_135278_comb;
  wire p1_slt_135280_comb;
  wire p1_slt_135282_comb;
  wire p1_slt_135284_comb;
  wire p1_slt_135286_comb;
  wire p1_slt_135288_comb;
  wire p1_slt_135290_comb;
  wire p1_slt_135292_comb;
  wire p1_slt_135294_comb;
  wire p1_slt_135296_comb;
  wire p1_slt_135298_comb;
  wire p1_slt_135300_comb;
  wire p1_slt_135302_comb;
  wire p1_slt_135304_comb;
  wire p1_slt_135306_comb;
  wire p1_slt_135308_comb;
  wire p1_slt_135310_comb;
  wire p1_slt_135312_comb;
  wire p1_slt_135314_comb;
  wire p1_slt_135316_comb;
  wire p1_slt_135318_comb;
  wire p1_slt_135320_comb;
  wire p1_slt_135322_comb;
  wire p1_slt_135324_comb;
  wire p1_slt_135326_comb;
  wire p1_slt_135328_comb;
  wire p1_slt_135330_comb;
  wire p1_slt_135332_comb;
  wire p1_slt_135334_comb;
  wire p1_slt_135336_comb;
  wire p1_slt_135338_comb;
  wire p1_slt_135340_comb;
  wire p1_slt_135342_comb;
  wire p1_slt_135344_comb;
  wire p1_slt_135346_comb;
  wire [31:0] p1_prod__199_comb;
  wire [22:0] p1_concat_135348_comb;
  wire [22:0] p1_concat_135349_comb;
  wire [31:0] p1_prod__214_comb;
  wire [31:0] p1_prod__263_comb;
  wire [22:0] p1_concat_135352_comb;
  wire [22:0] p1_concat_135353_comb;
  wire [31:0] p1_prod__278_comb;
  wire [22:0] p1_concat_135355_comb;
  wire [31:0] p1_prod__216_comb;
  wire [31:0] p1_prod__223_comb;
  wire [22:0] p1_concat_135358_comb;
  wire [22:0] p1_concat_135359_comb;
  wire [31:0] p1_prod__280_comb;
  wire [31:0] p1_prod__287_comb;
  wire [22:0] p1_concat_135362_comb;
  wire [31:0] p1_prod__212_comb;
  wire [22:0] p1_concat_135364_comb;
  wire [22:0] p1_concat_135365_comb;
  wire [31:0] p1_prod__250_comb;
  wire [31:0] p1_prod__276_comb;
  wire [22:0] p1_concat_135368_comb;
  wire [22:0] p1_concat_135369_comb;
  wire [31:0] p1_prod__314_comb;
  wire [22:0] p1_concat_135371_comb;
  wire [31:0] p1_prod__234_comb;
  wire [31:0] p1_prod__254_comb;
  wire [22:0] p1_concat_135374_comb;
  wire [22:0] p1_concat_135375_comb;
  wire [31:0] p1_prod__298_comb;
  wire [31:0] p1_prod__318_comb;
  wire [22:0] p1_concat_135378_comb;
  wire p1_sgt_135507_comb;
  wire p1_sgt_135508_comb;
  wire p1_sgt_135509_comb;
  wire p1_sgt_135510_comb;
  wire p1_sgt_135511_comb;
  wire p1_sgt_135512_comb;
  wire p1_sgt_135513_comb;
  wire p1_sgt_135514_comb;
  wire p1_sgt_135515_comb;
  wire p1_sgt_135516_comb;
  wire p1_sgt_135517_comb;
  wire p1_sgt_135518_comb;
  wire p1_sgt_135519_comb;
  wire p1_sgt_135520_comb;
  wire p1_sgt_135521_comb;
  wire p1_sgt_135522_comb;
  wire p1_sgt_135523_comb;
  wire p1_sgt_135524_comb;
  wire p1_sgt_135525_comb;
  wire p1_sgt_135526_comb;
  wire p1_sgt_135527_comb;
  wire p1_sgt_135528_comb;
  wire p1_sgt_135529_comb;
  wire p1_sgt_135530_comb;
  wire p1_sgt_135531_comb;
  wire p1_sgt_135532_comb;
  wire p1_sgt_135533_comb;
  wire p1_sgt_135534_comb;
  wire p1_sgt_135535_comb;
  wire p1_sgt_135536_comb;
  wire p1_sgt_135537_comb;
  wire p1_sgt_135538_comb;
  wire p1_sgt_135539_comb;
  wire p1_sgt_135540_comb;
  wire p1_sgt_135541_comb;
  wire p1_sgt_135542_comb;
  wire p1_sgt_135543_comb;
  wire p1_sgt_135544_comb;
  wire p1_sgt_135545_comb;
  wire p1_sgt_135546_comb;
  wire p1_sgt_135547_comb;
  wire p1_sgt_135548_comb;
  wire p1_sgt_135549_comb;
  wire p1_sgt_135550_comb;
  wire p1_sgt_135551_comb;
  wire p1_sgt_135552_comb;
  wire p1_sgt_135553_comb;
  wire p1_sgt_135554_comb;
  wire p1_sgt_135555_comb;
  wire p1_sgt_135556_comb;
  wire p1_sgt_135557_comb;
  wire p1_sgt_135558_comb;
  wire p1_sgt_135559_comb;
  wire p1_sgt_135560_comb;
  wire p1_sgt_135561_comb;
  wire p1_sgt_135562_comb;
  wire p1_sgt_135563_comb;
  wire p1_sgt_135564_comb;
  wire p1_sgt_135565_comb;
  wire p1_sgt_135566_comb;
  wire p1_sgt_135567_comb;
  wire p1_sgt_135568_comb;
  wire p1_sgt_135569_comb;
  wire p1_sgt_135570_comb;
  assign p1_array_index_133943_comb = p0_x[3'h3][3'h2];
  assign p1_array_index_133944_comb = p0_x[3'h3][3'h5];
  assign p1_array_index_133945_comb = p0_x[3'h4][3'h2];
  assign p1_array_index_133946_comb = p0_x[3'h4][3'h5];
  assign p1_array_index_133965_comb = p0_x[3'h3][3'h3];
  assign p1_array_index_133966_comb = p0_x[3'h3][3'h4];
  assign p1_array_index_133971_comb = p0_x[3'h4][3'h3];
  assign p1_array_index_133972_comb = p0_x[3'h4][3'h4];
  assign p1_array_index_133963_comb = p0_x[3'h3][3'h0];
  assign p1_array_index_133968_comb = p0_x[3'h3][3'h7];
  assign p1_array_index_133969_comb = p0_x[3'h4][3'h0];
  assign p1_array_index_133974_comb = p0_x[3'h4][3'h7];
  assign p1_array_index_133964_comb = p0_x[3'h3][3'h1];
  assign p1_array_index_133967_comb = p0_x[3'h3][3'h6];
  assign p1_array_index_133970_comb = p0_x[3'h4][3'h1];
  assign p1_array_index_133973_comb = p0_x[3'h4][3'h6];
  assign p1_array_index_133923_comb = p0_x[3'h2][3'h2];
  assign p1_array_index_133924_comb = p0_x[3'h2][3'h5];
  assign p1_array_index_133925_comb = p0_x[3'h5][3'h2];
  assign p1_array_index_133926_comb = p0_x[3'h5][3'h5];
  assign p1_array_index_133927_comb = p0_x[3'h2][3'h0];
  assign p1_array_index_133928_comb = p0_x[3'h2][3'h1];
  assign p1_array_index_133929_comb = p0_x[3'h2][3'h3];
  assign p1_array_index_133930_comb = p0_x[3'h2][3'h4];
  assign p1_array_index_133931_comb = p0_x[3'h2][3'h6];
  assign p1_array_index_133932_comb = p0_x[3'h2][3'h7];
  assign p1_array_index_133933_comb = p0_x[3'h5][3'h0];
  assign p1_array_index_133934_comb = p0_x[3'h5][3'h1];
  assign p1_array_index_133935_comb = p0_x[3'h5][3'h3];
  assign p1_array_index_133936_comb = p0_x[3'h5][3'h4];
  assign p1_array_index_133937_comb = p0_x[3'h5][3'h6];
  assign p1_array_index_133938_comb = p0_x[3'h5][3'h7];
  assign p1_array_index_133939_comb = p0_x[3'h0][3'h2];
  assign p1_array_index_133940_comb = p0_x[3'h0][3'h5];
  assign p1_array_index_133941_comb = p0_x[3'h1][3'h2];
  assign p1_array_index_133942_comb = p0_x[3'h1][3'h5];
  assign p1_array_index_133947_comb = p0_x[3'h6][3'h2];
  assign p1_array_index_133948_comb = p0_x[3'h6][3'h5];
  assign p1_array_index_133949_comb = p0_x[3'h7][3'h2];
  assign p1_array_index_133950_comb = p0_x[3'h7][3'h5];
  assign p1_array_index_133951_comb = p0_x[3'h0][3'h0];
  assign p1_array_index_133952_comb = p0_x[3'h0][3'h1];
  assign p1_array_index_133953_comb = p0_x[3'h0][3'h3];
  assign p1_array_index_133954_comb = p0_x[3'h0][3'h4];
  assign p1_array_index_133955_comb = p0_x[3'h0][3'h6];
  assign p1_array_index_133956_comb = p0_x[3'h0][3'h7];
  assign p1_array_index_133957_comb = p0_x[3'h1][3'h0];
  assign p1_array_index_133958_comb = p0_x[3'h1][3'h1];
  assign p1_array_index_133959_comb = p0_x[3'h1][3'h3];
  assign p1_array_index_133960_comb = p0_x[3'h1][3'h4];
  assign p1_array_index_133961_comb = p0_x[3'h1][3'h6];
  assign p1_array_index_133962_comb = p0_x[3'h1][3'h7];
  assign p1_array_index_133975_comb = p0_x[3'h6][3'h0];
  assign p1_array_index_133976_comb = p0_x[3'h6][3'h1];
  assign p1_array_index_133977_comb = p0_x[3'h6][3'h3];
  assign p1_array_index_133978_comb = p0_x[3'h6][3'h4];
  assign p1_array_index_133979_comb = p0_x[3'h6][3'h6];
  assign p1_array_index_133980_comb = p0_x[3'h6][3'h7];
  assign p1_array_index_133981_comb = p0_x[3'h7][3'h0];
  assign p1_array_index_133982_comb = p0_x[3'h7][3'h1];
  assign p1_array_index_133983_comb = p0_x[3'h7][3'h3];
  assign p1_array_index_133984_comb = p0_x[3'h7][3'h4];
  assign p1_array_index_133985_comb = p0_x[3'h7][3'h6];
  assign p1_array_index_133986_comb = p0_x[3'h7][3'h7];
  assign p1_shifted__26_squeezed_comb = {~p1_array_index_133943_comb[7], p1_array_index_133943_comb[6:0]};
  assign p1_shifted__29_squeezed_comb = {~p1_array_index_133944_comb[7], p1_array_index_133944_comb[6:0]};
  assign p1_shifted__34_squeezed_comb = {~p1_array_index_133945_comb[7], p1_array_index_133945_comb[6:0]};
  assign p1_shifted__37_squeezed_comb = {~p1_array_index_133946_comb[7], p1_array_index_133946_comb[6:0]};
  assign p1_shifted__27_squeezed_comb = {~p1_array_index_133965_comb[7], p1_array_index_133965_comb[6:0]};
  assign p1_shifted__28_squeezed_comb = {~p1_array_index_133966_comb[7], p1_array_index_133966_comb[6:0]};
  assign p1_shifted__35_squeezed_comb = {~p1_array_index_133971_comb[7], p1_array_index_133971_comb[6:0]};
  assign p1_shifted__36_squeezed_comb = {~p1_array_index_133972_comb[7], p1_array_index_133972_comb[6:0]};
  assign p1_shifted__24_squeezed_comb = {~p1_array_index_133963_comb[7], p1_array_index_133963_comb[6:0]};
  assign p1_shifted__31_squeezed_comb = {~p1_array_index_133968_comb[7], p1_array_index_133968_comb[6:0]};
  assign p1_shifted__32_squeezed_comb = {~p1_array_index_133969_comb[7], p1_array_index_133969_comb[6:0]};
  assign p1_shifted__39_squeezed_comb = {~p1_array_index_133974_comb[7], p1_array_index_133974_comb[6:0]};
  assign p1_shifted__25_squeezed_comb = {~p1_array_index_133964_comb[7], p1_array_index_133964_comb[6:0]};
  assign p1_shifted__30_squeezed_comb = {~p1_array_index_133967_comb[7], p1_array_index_133967_comb[6:0]};
  assign p1_shifted__33_squeezed_comb = {~p1_array_index_133970_comb[7], p1_array_index_133970_comb[6:0]};
  assign p1_shifted__38_squeezed_comb = {~p1_array_index_133973_comb[7], p1_array_index_133973_comb[6:0]};
  assign p1_shifted__18_squeezed_comb = {~p1_array_index_133923_comb[7], p1_array_index_133923_comb[6:0]};
  assign p1_shifted__21_squeezed_comb = {~p1_array_index_133924_comb[7], p1_array_index_133924_comb[6:0]};
  assign p1_shifted__42_squeezed_comb = {~p1_array_index_133925_comb[7], p1_array_index_133925_comb[6:0]};
  assign p1_shifted__45_squeezed_comb = {~p1_array_index_133926_comb[7], p1_array_index_133926_comb[6:0]};
  assign p1_shifted__16_squeezed_comb = {~p1_array_index_133927_comb[7], p1_array_index_133927_comb[6:0]};
  assign p1_shifted__17_squeezed_comb = {~p1_array_index_133928_comb[7], p1_array_index_133928_comb[6:0]};
  assign p1_shifted__19_squeezed_comb = {~p1_array_index_133929_comb[7], p1_array_index_133929_comb[6:0]};
  assign p1_shifted__20_squeezed_comb = {~p1_array_index_133930_comb[7], p1_array_index_133930_comb[6:0]};
  assign p1_shifted__22_squeezed_comb = {~p1_array_index_133931_comb[7], p1_array_index_133931_comb[6:0]};
  assign p1_shifted__23_squeezed_comb = {~p1_array_index_133932_comb[7], p1_array_index_133932_comb[6:0]};
  assign p1_shifted__40_squeezed_comb = {~p1_array_index_133933_comb[7], p1_array_index_133933_comb[6:0]};
  assign p1_shifted__41_squeezed_comb = {~p1_array_index_133934_comb[7], p1_array_index_133934_comb[6:0]};
  assign p1_shifted__43_squeezed_comb = {~p1_array_index_133935_comb[7], p1_array_index_133935_comb[6:0]};
  assign p1_shifted__44_squeezed_comb = {~p1_array_index_133936_comb[7], p1_array_index_133936_comb[6:0]};
  assign p1_shifted__46_squeezed_comb = {~p1_array_index_133937_comb[7], p1_array_index_133937_comb[6:0]};
  assign p1_shifted__47_squeezed_comb = {~p1_array_index_133938_comb[7], p1_array_index_133938_comb[6:0]};
  assign p1_shifted__2_squeezed_comb = {~p1_array_index_133939_comb[7], p1_array_index_133939_comb[6:0]};
  assign p1_shifted__5_squeezed_comb = {~p1_array_index_133940_comb[7], p1_array_index_133940_comb[6:0]};
  assign p1_shifted__10_squeezed_comb = {~p1_array_index_133941_comb[7], p1_array_index_133941_comb[6:0]};
  assign p1_shifted__13_squeezed_comb = {~p1_array_index_133942_comb[7], p1_array_index_133942_comb[6:0]};
  assign p1_shifted__50_squeezed_comb = {~p1_array_index_133947_comb[7], p1_array_index_133947_comb[6:0]};
  assign p1_shifted__53_squeezed_comb = {~p1_array_index_133948_comb[7], p1_array_index_133948_comb[6:0]};
  assign p1_shifted__58_squeezed_comb = {~p1_array_index_133949_comb[7], p1_array_index_133949_comb[6:0]};
  assign p1_shifted__61_squeezed_comb = {~p1_array_index_133950_comb[7], p1_array_index_133950_comb[6:0]};
  assign p1_shifted_squeezed_comb = {~p1_array_index_133951_comb[7], p1_array_index_133951_comb[6:0]};
  assign p1_shifted__1_squeezed_comb = {~p1_array_index_133952_comb[7], p1_array_index_133952_comb[6:0]};
  assign p1_shifted__3_squeezed_comb = {~p1_array_index_133953_comb[7], p1_array_index_133953_comb[6:0]};
  assign p1_shifted__4_squeezed_comb = {~p1_array_index_133954_comb[7], p1_array_index_133954_comb[6:0]};
  assign p1_shifted__6_squeezed_comb = {~p1_array_index_133955_comb[7], p1_array_index_133955_comb[6:0]};
  assign p1_shifted__7_squeezed_comb = {~p1_array_index_133956_comb[7], p1_array_index_133956_comb[6:0]};
  assign p1_shifted__8_squeezed_comb = {~p1_array_index_133957_comb[7], p1_array_index_133957_comb[6:0]};
  assign p1_shifted__9_squeezed_comb = {~p1_array_index_133958_comb[7], p1_array_index_133958_comb[6:0]};
  assign p1_shifted__11_squeezed_comb = {~p1_array_index_133959_comb[7], p1_array_index_133959_comb[6:0]};
  assign p1_shifted__12_squeezed_comb = {~p1_array_index_133960_comb[7], p1_array_index_133960_comb[6:0]};
  assign p1_shifted__14_squeezed_comb = {~p1_array_index_133961_comb[7], p1_array_index_133961_comb[6:0]};
  assign p1_shifted__15_squeezed_comb = {~p1_array_index_133962_comb[7], p1_array_index_133962_comb[6:0]};
  assign p1_shifted__48_squeezed_comb = {~p1_array_index_133975_comb[7], p1_array_index_133975_comb[6:0]};
  assign p1_shifted__49_squeezed_comb = {~p1_array_index_133976_comb[7], p1_array_index_133976_comb[6:0]};
  assign p1_shifted__51_squeezed_comb = {~p1_array_index_133977_comb[7], p1_array_index_133977_comb[6:0]};
  assign p1_shifted__52_squeezed_comb = {~p1_array_index_133978_comb[7], p1_array_index_133978_comb[6:0]};
  assign p1_shifted__54_squeezed_comb = {~p1_array_index_133979_comb[7], p1_array_index_133979_comb[6:0]};
  assign p1_shifted__55_squeezed_comb = {~p1_array_index_133980_comb[7], p1_array_index_133980_comb[6:0]};
  assign p1_shifted__56_squeezed_comb = {~p1_array_index_133981_comb[7], p1_array_index_133981_comb[6:0]};
  assign p1_shifted__57_squeezed_comb = {~p1_array_index_133982_comb[7], p1_array_index_133982_comb[6:0]};
  assign p1_shifted__59_squeezed_comb = {~p1_array_index_133983_comb[7], p1_array_index_133983_comb[6:0]};
  assign p1_shifted__60_squeezed_comb = {~p1_array_index_133984_comb[7], p1_array_index_133984_comb[6:0]};
  assign p1_shifted__62_squeezed_comb = {~p1_array_index_133985_comb[7], p1_array_index_133985_comb[6:0]};
  assign p1_shifted__63_squeezed_comb = {~p1_array_index_133986_comb[7], p1_array_index_133986_comb[6:0]};
  assign p1_smul_57378_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__26_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___12_comb = 9'h000;
  assign p1_smul_57384_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__29_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___15_comb = 9'h000;
  assign p1_smul_57394_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__34_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___16_comb = 9'h000;
  assign p1_smul_57400_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__37_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___19_comb = 9'h000;
  assign p1_smul_57636_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__27_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___77_comb = 9'h000;
  assign p1_smul_57638_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__28_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___78_comb = 9'h000;
  assign p1_smul_57652_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__35_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___81_comb = 9'h000;
  assign p1_smul_57654_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__36_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___82_comb = 9'h000;
  assign p1_smul_57886_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__24_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___108_comb = 9'h000;
  assign p1_smul_57900_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__31_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___111_comb = 9'h000;
  assign p1_smul_57902_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__32_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___112_comb = 9'h000;
  assign p1_smul_57916_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__39_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___115_comb = 9'h000;
  assign p1_smul_58144_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__25_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___173_comb = 9'h000;
  assign p1_smul_58154_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__30_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___174_comb = 9'h000;
  assign p1_smul_58160_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__33_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___177_comb = 9'h000;
  assign p1_smul_58170_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__38_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___178_comb = 9'h000;
  assign p1_smul_57326_TrailingBits___144_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___145_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___146_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___147_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___148_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___149_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___150_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___151_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___168_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___169_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___170_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___171_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___172_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___173_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___174_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___175_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___128_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___129_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___130_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___131_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___132_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___133_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___134_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___135_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___136_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___137_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___138_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___139_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___140_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___141_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___142_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___143_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___152_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___153_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___154_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___155_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___156_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___157_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___158_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___159_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___160_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___161_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___162_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___163_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___164_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___165_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___166_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___167_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___176_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___177_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___178_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___179_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___180_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___181_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___182_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___183_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___184_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___185_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___186_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___187_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___188_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___189_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___190_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___191_comb = 8'h00;
  assign p1_smul_57362_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__18_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___8_comb = 9'h000;
  assign p1_smul_57368_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__21_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___11_comb = 9'h000;
  assign p1_smul_57410_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__42_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___20_comb = 9'h000;
  assign p1_smul_57416_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__45_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___23_comb = 9'h000;
  assign p1_smul_57486_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__16_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___8_comb = 10'h000;
  assign p1_smul_57488_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__17_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___40_comb = 9'h000;
  assign p1_smul_57490_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__18_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___41_comb = 9'h000;
  assign p1_smul_57492_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__19_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___9_comb = 10'h000;
  assign p1_smul_57494_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__20_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___10_comb = 10'h000;
  assign p1_smul_57496_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__21_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___42_comb = 9'h000;
  assign p1_smul_57498_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__22_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___43_comb = 9'h000;
  assign p1_smul_57500_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__23_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___11_comb = 10'h000;
  assign p1_smul_57534_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__40_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___20_comb = 10'h000;
  assign p1_smul_57536_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__41_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___52_comb = 9'h000;
  assign p1_smul_57538_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__42_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___53_comb = 9'h000;
  assign p1_smul_57540_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__43_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___21_comb = 10'h000;
  assign p1_smul_57542_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__44_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___22_comb = 10'h000;
  assign p1_smul_57544_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__45_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___54_comb = 9'h000;
  assign p1_smul_57546_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__46_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___55_comb = 9'h000;
  assign p1_smul_57548_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__47_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___23_comb = 10'h000;
  assign p1_smul_57620_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__19_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___73_comb = 9'h000;
  assign p1_smul_57622_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__20_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___74_comb = 9'h000;
  assign p1_smul_57668_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__43_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___85_comb = 9'h000;
  assign p1_smul_57670_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__44_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___86_comb = 9'h000;
  assign p1_smul_57870_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__16_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___104_comb = 9'h000;
  assign p1_smul_57884_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__23_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___107_comb = 9'h000;
  assign p1_smul_57918_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__40_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___116_comb = 9'h000;
  assign p1_smul_57932_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__47_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___119_comb = 9'h000;
  assign p1_smul_57998_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__16_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___136_comb = 9'h000;
  assign p1_smul_58000_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__17_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___40_comb = 10'h000;
  assign p1_smul_58002_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__18_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___137_comb = 9'h000;
  assign p1_smul_58004_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__19_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___41_comb = 10'h000;
  assign p1_smul_58006_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__20_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___42_comb = 10'h000;
  assign p1_smul_58008_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__21_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___138_comb = 9'h000;
  assign p1_smul_58010_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__22_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___43_comb = 10'h000;
  assign p1_smul_58012_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__23_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___139_comb = 9'h000;
  assign p1_smul_58046_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__40_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___148_comb = 9'h000;
  assign p1_smul_58048_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__41_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___52_comb = 10'h000;
  assign p1_smul_58050_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__42_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___149_comb = 9'h000;
  assign p1_smul_58052_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__43_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___53_comb = 10'h000;
  assign p1_smul_58054_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__44_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___54_comb = 10'h000;
  assign p1_smul_58056_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__45_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___150_comb = 9'h000;
  assign p1_smul_58058_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__46_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___55_comb = 10'h000;
  assign p1_smul_58060_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__47_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___151_comb = 9'h000;
  assign p1_smul_58128_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__17_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___169_comb = 9'h000;
  assign p1_smul_58138_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__22_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___170_comb = 9'h000;
  assign p1_smul_58176_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__41_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___181_comb = 9'h000;
  assign p1_smul_58186_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__46_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___182_comb = 9'h000;
  assign p1_smul_57330_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__2_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits__comb = 9'h000;
  assign p1_smul_57336_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__5_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___3_comb = 9'h000;
  assign p1_smul_57346_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__10_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___4_comb = 9'h000;
  assign p1_smul_57352_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__13_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___7_comb = 9'h000;
  assign p1_smul_57426_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__50_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___24_comb = 9'h000;
  assign p1_smul_57432_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__53_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___27_comb = 9'h000;
  assign p1_smul_57442_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__58_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___28_comb = 9'h000;
  assign p1_smul_57448_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__61_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___31_comb = 9'h000;
  assign p1_smul_57454_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits__comb = 10'h000;
  assign p1_smul_57456_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__1_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___32_comb = 9'h000;
  assign p1_smul_57458_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__2_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___33_comb = 9'h000;
  assign p1_smul_57460_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__3_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___1_comb = 10'h000;
  assign p1_smul_57462_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__4_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___2_comb = 10'h000;
  assign p1_smul_57464_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__5_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___34_comb = 9'h000;
  assign p1_smul_57466_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__6_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___35_comb = 9'h000;
  assign p1_smul_57468_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__7_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___3_comb = 10'h000;
  assign p1_smul_57470_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__8_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___4_comb = 10'h000;
  assign p1_smul_57472_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__9_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___36_comb = 9'h000;
  assign p1_smul_57474_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__10_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___37_comb = 9'h000;
  assign p1_smul_57476_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__11_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___5_comb = 10'h000;
  assign p1_smul_57478_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__12_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___6_comb = 10'h000;
  assign p1_smul_57480_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__13_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___38_comb = 9'h000;
  assign p1_smul_57482_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__14_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___39_comb = 9'h000;
  assign p1_smul_57484_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__15_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___7_comb = 10'h000;
  assign p1_smul_57502_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__24_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___12_comb = 10'h000;
  assign p1_smul_57504_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__25_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___44_comb = 9'h000;
  assign p1_smul_57506_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__26_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___45_comb = 9'h000;
  assign p1_smul_57508_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__27_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___13_comb = 10'h000;
  assign p1_smul_57510_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__28_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___14_comb = 10'h000;
  assign p1_smul_57512_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__29_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___46_comb = 9'h000;
  assign p1_smul_57514_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__30_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___47_comb = 9'h000;
  assign p1_smul_57516_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__31_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___15_comb = 10'h000;
  assign p1_smul_57518_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__32_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___16_comb = 10'h000;
  assign p1_smul_57520_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__33_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___48_comb = 9'h000;
  assign p1_smul_57522_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__34_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___49_comb = 9'h000;
  assign p1_smul_57524_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__35_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___17_comb = 10'h000;
  assign p1_smul_57526_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__36_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___18_comb = 10'h000;
  assign p1_smul_57528_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__37_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___50_comb = 9'h000;
  assign p1_smul_57530_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__38_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___51_comb = 9'h000;
  assign p1_smul_57532_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__39_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___19_comb = 10'h000;
  assign p1_smul_57550_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__48_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___24_comb = 10'h000;
  assign p1_smul_57552_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__49_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___56_comb = 9'h000;
  assign p1_smul_57554_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__50_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___57_comb = 9'h000;
  assign p1_smul_57556_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__51_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___25_comb = 10'h000;
  assign p1_smul_57558_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__52_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___26_comb = 10'h000;
  assign p1_smul_57560_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__53_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___58_comb = 9'h000;
  assign p1_smul_57562_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__54_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___59_comb = 9'h000;
  assign p1_smul_57564_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__55_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___27_comb = 10'h000;
  assign p1_smul_57566_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__56_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___28_comb = 10'h000;
  assign p1_smul_57568_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__57_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___60_comb = 9'h000;
  assign p1_smul_57570_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__58_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___61_comb = 9'h000;
  assign p1_smul_57572_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__59_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___29_comb = 10'h000;
  assign p1_smul_57574_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__60_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___30_comb = 10'h000;
  assign p1_smul_57576_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__61_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___62_comb = 9'h000;
  assign p1_smul_57578_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__62_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___63_comb = 9'h000;
  assign p1_smul_57580_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__63_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___31_comb = 10'h000;
  assign p1_smul_57588_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__3_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___65_comb = 9'h000;
  assign p1_smul_57590_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__4_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___66_comb = 9'h000;
  assign p1_smul_57604_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__11_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___69_comb = 9'h000;
  assign p1_smul_57606_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__12_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___70_comb = 9'h000;
  assign p1_smul_57684_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__51_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___89_comb = 9'h000;
  assign p1_smul_57686_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__52_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___90_comb = 9'h000;
  assign p1_smul_57700_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__59_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___93_comb = 9'h000;
  assign p1_smul_57702_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__60_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___94_comb = 9'h000;
  assign p1_smul_57838_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___96_comb = 9'h000;
  assign p1_smul_57852_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__7_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___99_comb = 9'h000;
  assign p1_smul_57854_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__8_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___100_comb = 9'h000;
  assign p1_smul_57868_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__15_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___103_comb = 9'h000;
  assign p1_smul_57934_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__48_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___120_comb = 9'h000;
  assign p1_smul_57948_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__55_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___123_comb = 9'h000;
  assign p1_smul_57950_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__56_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___124_comb = 9'h000;
  assign p1_smul_57964_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__63_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___127_comb = 9'h000;
  assign p1_smul_57966_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___128_comb = 9'h000;
  assign p1_smul_57968_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__1_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___32_comb = 10'h000;
  assign p1_smul_57970_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__2_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___129_comb = 9'h000;
  assign p1_smul_57972_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__3_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___33_comb = 10'h000;
  assign p1_smul_57974_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__4_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___34_comb = 10'h000;
  assign p1_smul_57976_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__5_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___130_comb = 9'h000;
  assign p1_smul_57978_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__6_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___35_comb = 10'h000;
  assign p1_smul_57980_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__7_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___131_comb = 9'h000;
  assign p1_smul_57982_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__8_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___132_comb = 9'h000;
  assign p1_smul_57984_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__9_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___36_comb = 10'h000;
  assign p1_smul_57986_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__10_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___133_comb = 9'h000;
  assign p1_smul_57988_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__11_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___37_comb = 10'h000;
  assign p1_smul_57990_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__12_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___38_comb = 10'h000;
  assign p1_smul_57992_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__13_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___134_comb = 9'h000;
  assign p1_smul_57994_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__14_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___39_comb = 10'h000;
  assign p1_smul_57996_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__15_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___135_comb = 9'h000;
  assign p1_smul_58014_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__24_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___140_comb = 9'h000;
  assign p1_smul_58016_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__25_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___44_comb = 10'h000;
  assign p1_smul_58018_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__26_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___141_comb = 9'h000;
  assign p1_smul_58020_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__27_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___45_comb = 10'h000;
  assign p1_smul_58022_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__28_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___46_comb = 10'h000;
  assign p1_smul_58024_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__29_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___142_comb = 9'h000;
  assign p1_smul_58026_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__30_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___47_comb = 10'h000;
  assign p1_smul_58028_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__31_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___143_comb = 9'h000;
  assign p1_smul_58030_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__32_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___144_comb = 9'h000;
  assign p1_smul_58032_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__33_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___48_comb = 10'h000;
  assign p1_smul_58034_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__34_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___145_comb = 9'h000;
  assign p1_smul_58036_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__35_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___49_comb = 10'h000;
  assign p1_smul_58038_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__36_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___50_comb = 10'h000;
  assign p1_smul_58040_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__37_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___146_comb = 9'h000;
  assign p1_smul_58042_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__38_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___51_comb = 10'h000;
  assign p1_smul_58044_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__39_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___147_comb = 9'h000;
  assign p1_smul_58062_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__48_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___152_comb = 9'h000;
  assign p1_smul_58064_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__49_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___56_comb = 10'h000;
  assign p1_smul_58066_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__50_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___153_comb = 9'h000;
  assign p1_smul_58068_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__51_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___57_comb = 10'h000;
  assign p1_smul_58070_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__52_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___58_comb = 10'h000;
  assign p1_smul_58072_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__53_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___154_comb = 9'h000;
  assign p1_smul_58074_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__54_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___59_comb = 10'h000;
  assign p1_smul_58076_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__55_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___155_comb = 9'h000;
  assign p1_smul_58078_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__56_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___156_comb = 9'h000;
  assign p1_smul_58080_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__57_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___60_comb = 10'h000;
  assign p1_smul_58082_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__58_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___157_comb = 9'h000;
  assign p1_smul_58084_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__59_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___61_comb = 10'h000;
  assign p1_smul_58086_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__60_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___62_comb = 10'h000;
  assign p1_smul_58088_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__61_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___158_comb = 9'h000;
  assign p1_smul_58090_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__62_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___63_comb = 10'h000;
  assign p1_smul_58092_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__63_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___159_comb = 9'h000;
  assign p1_smul_58096_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__1_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___161_comb = 9'h000;
  assign p1_smul_58106_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__6_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___162_comb = 9'h000;
  assign p1_smul_58112_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__9_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___165_comb = 9'h000;
  assign p1_smul_58122_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__14_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___166_comb = 9'h000;
  assign p1_smul_58192_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__49_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___185_comb = 9'h000;
  assign p1_smul_58202_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__54_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___186_comb = 9'h000;
  assign p1_smul_58208_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__57_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___189_comb = 9'h000;
  assign p1_smul_58218_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__62_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___190_comb = 9'h000;
  assign p1_concat_135019_comb = {p1_smul_57378_NarrowedMult__comb, p1_smul_57330_TrailingBits___12_comb};
  assign p1_smul_57380_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__27_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___13_comb = 9'h000;
  assign p1_smul_57382_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__28_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___14_comb = 9'h000;
  assign p1_concat_135024_comb = {p1_smul_57384_NarrowedMult__comb, p1_smul_57330_TrailingBits___15_comb};
  assign p1_concat_135025_comb = {p1_smul_57394_NarrowedMult__comb, p1_smul_57330_TrailingBits___16_comb};
  assign p1_smul_57396_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__35_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___17_comb = 9'h000;
  assign p1_smul_57398_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__36_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___18_comb = 9'h000;
  assign p1_concat_135030_comb = {p1_smul_57400_NarrowedMult__comb, p1_smul_57330_TrailingBits___19_comb};
  assign p1_smul_57632_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__25_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___76_comb = 9'h000;
  assign p1_concat_135097_comb = {p1_smul_57636_NarrowedMult__comb, p1_smul_57330_TrailingBits___77_comb};
  assign p1_concat_135098_comb = {p1_smul_57638_NarrowedMult__comb, p1_smul_57330_TrailingBits___78_comb};
  assign p1_smul_57642_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__30_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___79_comb = 9'h000;
  assign p1_smul_57648_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__33_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___80_comb = 9'h000;
  assign p1_concat_135103_comb = {p1_smul_57652_NarrowedMult__comb, p1_smul_57330_TrailingBits___81_comb};
  assign p1_concat_135104_comb = {p1_smul_57654_NarrowedMult__comb, p1_smul_57330_TrailingBits___82_comb};
  assign p1_smul_57658_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__38_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___83_comb = 9'h000;
  assign p1_concat_135123_comb = {p1_smul_57886_NarrowedMult__comb, p1_smul_57330_TrailingBits___108_comb};
  assign p1_smul_57890_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__26_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___109_comb = 9'h000;
  assign p1_smul_57896_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__29_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___110_comb = 9'h000;
  assign p1_concat_135128_comb = {p1_smul_57900_NarrowedMult__comb, p1_smul_57330_TrailingBits___111_comb};
  assign p1_concat_135129_comb = {p1_smul_57902_NarrowedMult__comb, p1_smul_57330_TrailingBits___112_comb};
  assign p1_smul_57906_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__34_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___113_comb = 9'h000;
  assign p1_smul_57912_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__37_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___114_comb = 9'h000;
  assign p1_concat_135134_comb = {p1_smul_57916_NarrowedMult__comb, p1_smul_57330_TrailingBits___115_comb};
  assign p1_smul_58142_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__24_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___172_comb = 9'h000;
  assign p1_concat_135201_comb = {p1_smul_58144_NarrowedMult__comb, p1_smul_57330_TrailingBits___173_comb};
  assign p1_concat_135202_comb = {p1_smul_58154_NarrowedMult__comb, p1_smul_57330_TrailingBits___174_comb};
  assign p1_smul_58156_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__31_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___175_comb = 9'h000;
  assign p1_smul_58158_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__32_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___176_comb = 9'h000;
  assign p1_concat_135207_comb = {p1_smul_58160_NarrowedMult__comb, p1_smul_57330_TrailingBits___177_comb};
  assign p1_concat_135208_comb = {p1_smul_58170_NarrowedMult__comb, p1_smul_57330_TrailingBits___178_comb};
  assign p1_smul_58172_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__39_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___179_comb = 9'h000;
  assign p1_shifted__16_comb = {~p1_array_index_133927_comb[7], p1_array_index_133927_comb[6:0], p1_smul_57326_TrailingBits___144_comb};
  assign p1_shifted__17_comb = {~p1_array_index_133928_comb[7], p1_array_index_133928_comb[6:0], p1_smul_57326_TrailingBits___145_comb};
  assign p1_shifted__18_comb = {~p1_array_index_133923_comb[7], p1_array_index_133923_comb[6:0], p1_smul_57326_TrailingBits___146_comb};
  assign p1_shifted__19_comb = {~p1_array_index_133929_comb[7], p1_array_index_133929_comb[6:0], p1_smul_57326_TrailingBits___147_comb};
  assign p1_shifted__20_comb = {~p1_array_index_133930_comb[7], p1_array_index_133930_comb[6:0], p1_smul_57326_TrailingBits___148_comb};
  assign p1_shifted__21_comb = {~p1_array_index_133924_comb[7], p1_array_index_133924_comb[6:0], p1_smul_57326_TrailingBits___149_comb};
  assign p1_shifted__22_comb = {~p1_array_index_133931_comb[7], p1_array_index_133931_comb[6:0], p1_smul_57326_TrailingBits___150_comb};
  assign p1_shifted__23_comb = {~p1_array_index_133932_comb[7], p1_array_index_133932_comb[6:0], p1_smul_57326_TrailingBits___151_comb};
  assign p1_shifted__40_comb = {~p1_array_index_133933_comb[7], p1_array_index_133933_comb[6:0], p1_smul_57326_TrailingBits___168_comb};
  assign p1_shifted__41_comb = {~p1_array_index_133934_comb[7], p1_array_index_133934_comb[6:0], p1_smul_57326_TrailingBits___169_comb};
  assign p1_shifted__42_comb = {~p1_array_index_133925_comb[7], p1_array_index_133925_comb[6:0], p1_smul_57326_TrailingBits___170_comb};
  assign p1_shifted__43_comb = {~p1_array_index_133935_comb[7], p1_array_index_133935_comb[6:0], p1_smul_57326_TrailingBits___171_comb};
  assign p1_shifted__44_comb = {~p1_array_index_133936_comb[7], p1_array_index_133936_comb[6:0], p1_smul_57326_TrailingBits___172_comb};
  assign p1_shifted__45_comb = {~p1_array_index_133926_comb[7], p1_array_index_133926_comb[6:0], p1_smul_57326_TrailingBits___173_comb};
  assign p1_shifted__46_comb = {~p1_array_index_133937_comb[7], p1_array_index_133937_comb[6:0], p1_smul_57326_TrailingBits___174_comb};
  assign p1_shifted__47_comb = {~p1_array_index_133938_comb[7], p1_array_index_133938_comb[6:0], p1_smul_57326_TrailingBits___175_comb};
  assign p1_shifted_comb = {~p1_array_index_133951_comb[7], p1_array_index_133951_comb[6:0], p1_smul_57326_TrailingBits___128_comb};
  assign p1_shifted__1_comb = {~p1_array_index_133952_comb[7], p1_array_index_133952_comb[6:0], p1_smul_57326_TrailingBits___129_comb};
  assign p1_shifted__2_comb = {~p1_array_index_133939_comb[7], p1_array_index_133939_comb[6:0], p1_smul_57326_TrailingBits___130_comb};
  assign p1_shifted__3_comb = {~p1_array_index_133953_comb[7], p1_array_index_133953_comb[6:0], p1_smul_57326_TrailingBits___131_comb};
  assign p1_shifted__4_comb = {~p1_array_index_133954_comb[7], p1_array_index_133954_comb[6:0], p1_smul_57326_TrailingBits___132_comb};
  assign p1_shifted__5_comb = {~p1_array_index_133940_comb[7], p1_array_index_133940_comb[6:0], p1_smul_57326_TrailingBits___133_comb};
  assign p1_shifted__6_comb = {~p1_array_index_133955_comb[7], p1_array_index_133955_comb[6:0], p1_smul_57326_TrailingBits___134_comb};
  assign p1_shifted__7_comb = {~p1_array_index_133956_comb[7], p1_array_index_133956_comb[6:0], p1_smul_57326_TrailingBits___135_comb};
  assign p1_shifted__8_comb = {~p1_array_index_133957_comb[7], p1_array_index_133957_comb[6:0], p1_smul_57326_TrailingBits___136_comb};
  assign p1_shifted__9_comb = {~p1_array_index_133958_comb[7], p1_array_index_133958_comb[6:0], p1_smul_57326_TrailingBits___137_comb};
  assign p1_shifted__10_comb = {~p1_array_index_133941_comb[7], p1_array_index_133941_comb[6:0], p1_smul_57326_TrailingBits___138_comb};
  assign p1_shifted__11_comb = {~p1_array_index_133959_comb[7], p1_array_index_133959_comb[6:0], p1_smul_57326_TrailingBits___139_comb};
  assign p1_shifted__12_comb = {~p1_array_index_133960_comb[7], p1_array_index_133960_comb[6:0], p1_smul_57326_TrailingBits___140_comb};
  assign p1_shifted__13_comb = {~p1_array_index_133942_comb[7], p1_array_index_133942_comb[6:0], p1_smul_57326_TrailingBits___141_comb};
  assign p1_shifted__14_comb = {~p1_array_index_133961_comb[7], p1_array_index_133961_comb[6:0], p1_smul_57326_TrailingBits___142_comb};
  assign p1_shifted__15_comb = {~p1_array_index_133962_comb[7], p1_array_index_133962_comb[6:0], p1_smul_57326_TrailingBits___143_comb};
  assign p1_shifted__24_comb = {~p1_array_index_133963_comb[7], p1_array_index_133963_comb[6:0], p1_smul_57326_TrailingBits___152_comb};
  assign p1_shifted__25_comb = {~p1_array_index_133964_comb[7], p1_array_index_133964_comb[6:0], p1_smul_57326_TrailingBits___153_comb};
  assign p1_shifted__26_comb = {~p1_array_index_133943_comb[7], p1_array_index_133943_comb[6:0], p1_smul_57326_TrailingBits___154_comb};
  assign p1_shifted__27_comb = {~p1_array_index_133965_comb[7], p1_array_index_133965_comb[6:0], p1_smul_57326_TrailingBits___155_comb};
  assign p1_shifted__28_comb = {~p1_array_index_133966_comb[7], p1_array_index_133966_comb[6:0], p1_smul_57326_TrailingBits___156_comb};
  assign p1_shifted__29_comb = {~p1_array_index_133944_comb[7], p1_array_index_133944_comb[6:0], p1_smul_57326_TrailingBits___157_comb};
  assign p1_shifted__30_comb = {~p1_array_index_133967_comb[7], p1_array_index_133967_comb[6:0], p1_smul_57326_TrailingBits___158_comb};
  assign p1_shifted__31_comb = {~p1_array_index_133968_comb[7], p1_array_index_133968_comb[6:0], p1_smul_57326_TrailingBits___159_comb};
  assign p1_shifted__32_comb = {~p1_array_index_133969_comb[7], p1_array_index_133969_comb[6:0], p1_smul_57326_TrailingBits___160_comb};
  assign p1_shifted__33_comb = {~p1_array_index_133970_comb[7], p1_array_index_133970_comb[6:0], p1_smul_57326_TrailingBits___161_comb};
  assign p1_shifted__34_comb = {~p1_array_index_133945_comb[7], p1_array_index_133945_comb[6:0], p1_smul_57326_TrailingBits___162_comb};
  assign p1_shifted__35_comb = {~p1_array_index_133971_comb[7], p1_array_index_133971_comb[6:0], p1_smul_57326_TrailingBits___163_comb};
  assign p1_shifted__36_comb = {~p1_array_index_133972_comb[7], p1_array_index_133972_comb[6:0], p1_smul_57326_TrailingBits___164_comb};
  assign p1_shifted__37_comb = {~p1_array_index_133946_comb[7], p1_array_index_133946_comb[6:0], p1_smul_57326_TrailingBits___165_comb};
  assign p1_shifted__38_comb = {~p1_array_index_133973_comb[7], p1_array_index_133973_comb[6:0], p1_smul_57326_TrailingBits___166_comb};
  assign p1_shifted__39_comb = {~p1_array_index_133974_comb[7], p1_array_index_133974_comb[6:0], p1_smul_57326_TrailingBits___167_comb};
  assign p1_shifted__48_comb = {~p1_array_index_133975_comb[7], p1_array_index_133975_comb[6:0], p1_smul_57326_TrailingBits___176_comb};
  assign p1_shifted__49_comb = {~p1_array_index_133976_comb[7], p1_array_index_133976_comb[6:0], p1_smul_57326_TrailingBits___177_comb};
  assign p1_shifted__50_comb = {~p1_array_index_133947_comb[7], p1_array_index_133947_comb[6:0], p1_smul_57326_TrailingBits___178_comb};
  assign p1_shifted__51_comb = {~p1_array_index_133977_comb[7], p1_array_index_133977_comb[6:0], p1_smul_57326_TrailingBits___179_comb};
  assign p1_shifted__52_comb = {~p1_array_index_133978_comb[7], p1_array_index_133978_comb[6:0], p1_smul_57326_TrailingBits___180_comb};
  assign p1_shifted__53_comb = {~p1_array_index_133948_comb[7], p1_array_index_133948_comb[6:0], p1_smul_57326_TrailingBits___181_comb};
  assign p1_shifted__54_comb = {~p1_array_index_133979_comb[7], p1_array_index_133979_comb[6:0], p1_smul_57326_TrailingBits___182_comb};
  assign p1_shifted__55_comb = {~p1_array_index_133980_comb[7], p1_array_index_133980_comb[6:0], p1_smul_57326_TrailingBits___183_comb};
  assign p1_shifted__56_comb = {~p1_array_index_133981_comb[7], p1_array_index_133981_comb[6:0], p1_smul_57326_TrailingBits___184_comb};
  assign p1_shifted__57_comb = {~p1_array_index_133982_comb[7], p1_array_index_133982_comb[6:0], p1_smul_57326_TrailingBits___185_comb};
  assign p1_shifted__58_comb = {~p1_array_index_133949_comb[7], p1_array_index_133949_comb[6:0], p1_smul_57326_TrailingBits___186_comb};
  assign p1_shifted__59_comb = {~p1_array_index_133983_comb[7], p1_array_index_133983_comb[6:0], p1_smul_57326_TrailingBits___187_comb};
  assign p1_shifted__60_comb = {~p1_array_index_133984_comb[7], p1_array_index_133984_comb[6:0], p1_smul_57326_TrailingBits___188_comb};
  assign p1_shifted__61_comb = {~p1_array_index_133950_comb[7], p1_array_index_133950_comb[6:0], p1_smul_57326_TrailingBits___189_comb};
  assign p1_shifted__62_comb = {~p1_array_index_133985_comb[7], p1_array_index_133985_comb[6:0], p1_smul_57326_TrailingBits___190_comb};
  assign p1_shifted__63_comb = {~p1_array_index_133986_comb[7], p1_array_index_133986_comb[6:0], p1_smul_57326_TrailingBits___191_comb};
  assign p1_concat_134899_comb = {p1_smul_57362_NarrowedMult__comb, p1_smul_57330_TrailingBits___8_comb};
  assign p1_smul_57364_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__19_squeezed_comb, 6'h19);
  assign p1_smul_57366_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__20_squeezed_comb, 6'h27);
  assign p1_concat_134902_comb = {p1_smul_57368_NarrowedMult__comb, p1_smul_57330_TrailingBits___11_comb};
  assign p1_concat_134903_comb = {p1_smul_57410_NarrowedMult__comb, p1_smul_57330_TrailingBits___20_comb};
  assign p1_smul_57412_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__43_squeezed_comb, 6'h19);
  assign p1_smul_57414_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__44_squeezed_comb, 6'h27);
  assign p1_concat_134906_comb = {p1_smul_57416_NarrowedMult__comb, p1_smul_57330_TrailingBits___23_comb};
  assign p1_concat_134907_comb = {p1_smul_57486_NarrowedMult__comb, p1_smul_57454_TrailingBits___8_comb};
  assign p1_concat_134908_comb = {p1_smul_57488_NarrowedMult__comb, p1_smul_57330_TrailingBits___40_comb};
  assign p1_concat_134909_comb = {p1_smul_57490_NarrowedMult__comb, p1_smul_57330_TrailingBits___41_comb};
  assign p1_concat_134910_comb = {p1_smul_57492_NarrowedMult__comb, p1_smul_57454_TrailingBits___9_comb};
  assign p1_concat_134911_comb = {p1_smul_57494_NarrowedMult__comb, p1_smul_57454_TrailingBits___10_comb};
  assign p1_concat_134912_comb = {p1_smul_57496_NarrowedMult__comb, p1_smul_57330_TrailingBits___42_comb};
  assign p1_concat_134913_comb = {p1_smul_57498_NarrowedMult__comb, p1_smul_57330_TrailingBits___43_comb};
  assign p1_concat_134914_comb = {p1_smul_57500_NarrowedMult__comb, p1_smul_57454_TrailingBits___11_comb};
  assign p1_concat_134915_comb = {p1_smul_57534_NarrowedMult__comb, p1_smul_57454_TrailingBits___20_comb};
  assign p1_concat_134916_comb = {p1_smul_57536_NarrowedMult__comb, p1_smul_57330_TrailingBits___52_comb};
  assign p1_concat_134917_comb = {p1_smul_57538_NarrowedMult__comb, p1_smul_57330_TrailingBits___53_comb};
  assign p1_concat_134918_comb = {p1_smul_57540_NarrowedMult__comb, p1_smul_57454_TrailingBits___21_comb};
  assign p1_concat_134919_comb = {p1_smul_57542_NarrowedMult__comb, p1_smul_57454_TrailingBits___22_comb};
  assign p1_concat_134920_comb = {p1_smul_57544_NarrowedMult__comb, p1_smul_57330_TrailingBits___54_comb};
  assign p1_concat_134921_comb = {p1_smul_57546_NarrowedMult__comb, p1_smul_57330_TrailingBits___55_comb};
  assign p1_concat_134922_comb = {p1_smul_57548_NarrowedMult__comb, p1_smul_57454_TrailingBits___23_comb};
  assign p1_smul_57616_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__17_squeezed_comb, 6'h27);
  assign p1_concat_134924_comb = {p1_smul_57620_NarrowedMult__comb, p1_smul_57330_TrailingBits___73_comb};
  assign p1_concat_134925_comb = {p1_smul_57622_NarrowedMult__comb, p1_smul_57330_TrailingBits___74_comb};
  assign p1_smul_57626_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__22_squeezed_comb, 6'h19);
  assign p1_smul_57664_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__41_squeezed_comb, 6'h27);
  assign p1_concat_134928_comb = {p1_smul_57668_NarrowedMult__comb, p1_smul_57330_TrailingBits___85_comb};
  assign p1_concat_134929_comb = {p1_smul_57670_NarrowedMult__comb, p1_smul_57330_TrailingBits___86_comb};
  assign p1_smul_57674_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__46_squeezed_comb, 6'h19);
  assign p1_concat_134931_comb = {p1_smul_57870_NarrowedMult__comb, p1_smul_57330_TrailingBits___104_comb};
  assign p1_smul_57874_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__18_squeezed_comb, 6'h27);
  assign p1_smul_57880_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__21_squeezed_comb, 6'h27);
  assign p1_concat_134934_comb = {p1_smul_57884_NarrowedMult__comb, p1_smul_57330_TrailingBits___107_comb};
  assign p1_concat_134935_comb = {p1_smul_57918_NarrowedMult__comb, p1_smul_57330_TrailingBits___116_comb};
  assign p1_smul_57922_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__42_squeezed_comb, 6'h27);
  assign p1_smul_57928_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__45_squeezed_comb, 6'h27);
  assign p1_concat_134938_comb = {p1_smul_57932_NarrowedMult__comb, p1_smul_57330_TrailingBits___119_comb};
  assign p1_concat_134939_comb = {p1_smul_57998_NarrowedMult__comb, p1_smul_57330_TrailingBits___136_comb};
  assign p1_concat_134940_comb = {p1_smul_58000_NarrowedMult__comb, p1_smul_57454_TrailingBits___40_comb};
  assign p1_concat_134941_comb = {p1_smul_58002_NarrowedMult__comb, p1_smul_57330_TrailingBits___137_comb};
  assign p1_concat_134942_comb = {p1_smul_58004_NarrowedMult__comb, p1_smul_57454_TrailingBits___41_comb};
  assign p1_concat_134943_comb = {p1_smul_58006_NarrowedMult__comb, p1_smul_57454_TrailingBits___42_comb};
  assign p1_concat_134944_comb = {p1_smul_58008_NarrowedMult__comb, p1_smul_57330_TrailingBits___138_comb};
  assign p1_concat_134945_comb = {p1_smul_58010_NarrowedMult__comb, p1_smul_57454_TrailingBits___43_comb};
  assign p1_concat_134946_comb = {p1_smul_58012_NarrowedMult__comb, p1_smul_57330_TrailingBits___139_comb};
  assign p1_concat_134947_comb = {p1_smul_58046_NarrowedMult__comb, p1_smul_57330_TrailingBits___148_comb};
  assign p1_concat_134948_comb = {p1_smul_58048_NarrowedMult__comb, p1_smul_57454_TrailingBits___52_comb};
  assign p1_concat_134949_comb = {p1_smul_58050_NarrowedMult__comb, p1_smul_57330_TrailingBits___149_comb};
  assign p1_concat_134950_comb = {p1_smul_58052_NarrowedMult__comb, p1_smul_57454_TrailingBits___53_comb};
  assign p1_concat_134951_comb = {p1_smul_58054_NarrowedMult__comb, p1_smul_57454_TrailingBits___54_comb};
  assign p1_concat_134952_comb = {p1_smul_58056_NarrowedMult__comb, p1_smul_57330_TrailingBits___150_comb};
  assign p1_concat_134953_comb = {p1_smul_58058_NarrowedMult__comb, p1_smul_57454_TrailingBits___55_comb};
  assign p1_concat_134954_comb = {p1_smul_58060_NarrowedMult__comb, p1_smul_57330_TrailingBits___151_comb};
  assign p1_smul_58126_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__16_squeezed_comb, 6'h19);
  assign p1_concat_134956_comb = {p1_smul_58128_NarrowedMult__comb, p1_smul_57330_TrailingBits___169_comb};
  assign p1_concat_134957_comb = {p1_smul_58138_NarrowedMult__comb, p1_smul_57330_TrailingBits___170_comb};
  assign p1_smul_58140_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__23_squeezed_comb, 6'h19);
  assign p1_smul_58174_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__40_squeezed_comb, 6'h19);
  assign p1_concat_134960_comb = {p1_smul_58176_NarrowedMult__comb, p1_smul_57330_TrailingBits___181_comb};
  assign p1_concat_134961_comb = {p1_smul_58186_NarrowedMult__comb, p1_smul_57330_TrailingBits___182_comb};
  assign p1_smul_58188_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__47_squeezed_comb, 6'h19);
  assign p1_concat_135011_comb = {p1_smul_57330_NarrowedMult__comb, p1_smul_57330_TrailingBits__comb};
  assign p1_smul_57332_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__3_squeezed_comb, 6'h19);
  assign p1_smul_57334_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__4_squeezed_comb, 6'h27);
  assign p1_concat_135014_comb = {p1_smul_57336_NarrowedMult__comb, p1_smul_57330_TrailingBits___3_comb};
  assign p1_concat_135015_comb = {p1_smul_57346_NarrowedMult__comb, p1_smul_57330_TrailingBits___4_comb};
  assign p1_smul_57348_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__11_squeezed_comb, 6'h19);
  assign p1_smul_57350_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__12_squeezed_comb, 6'h27);
  assign p1_concat_135018_comb = {p1_smul_57352_NarrowedMult__comb, p1_smul_57330_TrailingBits___7_comb};
  assign p1_concat_135031_comb = {p1_smul_57426_NarrowedMult__comb, p1_smul_57330_TrailingBits___24_comb};
  assign p1_smul_57428_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__51_squeezed_comb, 6'h19);
  assign p1_smul_57430_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__52_squeezed_comb, 6'h27);
  assign p1_concat_135034_comb = {p1_smul_57432_NarrowedMult__comb, p1_smul_57330_TrailingBits___27_comb};
  assign p1_concat_135035_comb = {p1_smul_57442_NarrowedMult__comb, p1_smul_57330_TrailingBits___28_comb};
  assign p1_smul_57444_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__59_squeezed_comb, 6'h19);
  assign p1_smul_57446_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__60_squeezed_comb, 6'h27);
  assign p1_concat_135038_comb = {p1_smul_57448_NarrowedMult__comb, p1_smul_57330_TrailingBits___31_comb};
  assign p1_concat_135039_comb = {p1_smul_57454_NarrowedMult__comb, p1_smul_57454_TrailingBits__comb};
  assign p1_concat_135040_comb = {p1_smul_57456_NarrowedMult__comb, p1_smul_57330_TrailingBits___32_comb};
  assign p1_concat_135041_comb = {p1_smul_57458_NarrowedMult__comb, p1_smul_57330_TrailingBits___33_comb};
  assign p1_concat_135042_comb = {p1_smul_57460_NarrowedMult__comb, p1_smul_57454_TrailingBits___1_comb};
  assign p1_concat_135043_comb = {p1_smul_57462_NarrowedMult__comb, p1_smul_57454_TrailingBits___2_comb};
  assign p1_concat_135044_comb = {p1_smul_57464_NarrowedMult__comb, p1_smul_57330_TrailingBits___34_comb};
  assign p1_concat_135045_comb = {p1_smul_57466_NarrowedMult__comb, p1_smul_57330_TrailingBits___35_comb};
  assign p1_concat_135046_comb = {p1_smul_57468_NarrowedMult__comb, p1_smul_57454_TrailingBits___3_comb};
  assign p1_concat_135047_comb = {p1_smul_57470_NarrowedMult__comb, p1_smul_57454_TrailingBits___4_comb};
  assign p1_concat_135048_comb = {p1_smul_57472_NarrowedMult__comb, p1_smul_57330_TrailingBits___36_comb};
  assign p1_concat_135049_comb = {p1_smul_57474_NarrowedMult__comb, p1_smul_57330_TrailingBits___37_comb};
  assign p1_concat_135050_comb = {p1_smul_57476_NarrowedMult__comb, p1_smul_57454_TrailingBits___5_comb};
  assign p1_concat_135051_comb = {p1_smul_57478_NarrowedMult__comb, p1_smul_57454_TrailingBits___6_comb};
  assign p1_concat_135052_comb = {p1_smul_57480_NarrowedMult__comb, p1_smul_57330_TrailingBits___38_comb};
  assign p1_concat_135053_comb = {p1_smul_57482_NarrowedMult__comb, p1_smul_57330_TrailingBits___39_comb};
  assign p1_concat_135054_comb = {p1_smul_57484_NarrowedMult__comb, p1_smul_57454_TrailingBits___7_comb};
  assign p1_concat_135055_comb = {p1_smul_57502_NarrowedMult__comb, p1_smul_57454_TrailingBits___12_comb};
  assign p1_concat_135056_comb = {p1_smul_57504_NarrowedMult__comb, p1_smul_57330_TrailingBits___44_comb};
  assign p1_concat_135057_comb = {p1_smul_57506_NarrowedMult__comb, p1_smul_57330_TrailingBits___45_comb};
  assign p1_concat_135058_comb = {p1_smul_57508_NarrowedMult__comb, p1_smul_57454_TrailingBits___13_comb};
  assign p1_concat_135059_comb = {p1_smul_57510_NarrowedMult__comb, p1_smul_57454_TrailingBits___14_comb};
  assign p1_concat_135060_comb = {p1_smul_57512_NarrowedMult__comb, p1_smul_57330_TrailingBits___46_comb};
  assign p1_concat_135061_comb = {p1_smul_57514_NarrowedMult__comb, p1_smul_57330_TrailingBits___47_comb};
  assign p1_concat_135062_comb = {p1_smul_57516_NarrowedMult__comb, p1_smul_57454_TrailingBits___15_comb};
  assign p1_concat_135063_comb = {p1_smul_57518_NarrowedMult__comb, p1_smul_57454_TrailingBits___16_comb};
  assign p1_concat_135064_comb = {p1_smul_57520_NarrowedMult__comb, p1_smul_57330_TrailingBits___48_comb};
  assign p1_concat_135065_comb = {p1_smul_57522_NarrowedMult__comb, p1_smul_57330_TrailingBits___49_comb};
  assign p1_concat_135066_comb = {p1_smul_57524_NarrowedMult__comb, p1_smul_57454_TrailingBits___17_comb};
  assign p1_concat_135067_comb = {p1_smul_57526_NarrowedMult__comb, p1_smul_57454_TrailingBits___18_comb};
  assign p1_concat_135068_comb = {p1_smul_57528_NarrowedMult__comb, p1_smul_57330_TrailingBits___50_comb};
  assign p1_concat_135069_comb = {p1_smul_57530_NarrowedMult__comb, p1_smul_57330_TrailingBits___51_comb};
  assign p1_concat_135070_comb = {p1_smul_57532_NarrowedMult__comb, p1_smul_57454_TrailingBits___19_comb};
  assign p1_concat_135071_comb = {p1_smul_57550_NarrowedMult__comb, p1_smul_57454_TrailingBits___24_comb};
  assign p1_concat_135072_comb = {p1_smul_57552_NarrowedMult__comb, p1_smul_57330_TrailingBits___56_comb};
  assign p1_concat_135073_comb = {p1_smul_57554_NarrowedMult__comb, p1_smul_57330_TrailingBits___57_comb};
  assign p1_concat_135074_comb = {p1_smul_57556_NarrowedMult__comb, p1_smul_57454_TrailingBits___25_comb};
  assign p1_concat_135075_comb = {p1_smul_57558_NarrowedMult__comb, p1_smul_57454_TrailingBits___26_comb};
  assign p1_concat_135076_comb = {p1_smul_57560_NarrowedMult__comb, p1_smul_57330_TrailingBits___58_comb};
  assign p1_concat_135077_comb = {p1_smul_57562_NarrowedMult__comb, p1_smul_57330_TrailingBits___59_comb};
  assign p1_concat_135078_comb = {p1_smul_57564_NarrowedMult__comb, p1_smul_57454_TrailingBits___27_comb};
  assign p1_concat_135079_comb = {p1_smul_57566_NarrowedMult__comb, p1_smul_57454_TrailingBits___28_comb};
  assign p1_concat_135080_comb = {p1_smul_57568_NarrowedMult__comb, p1_smul_57330_TrailingBits___60_comb};
  assign p1_concat_135081_comb = {p1_smul_57570_NarrowedMult__comb, p1_smul_57330_TrailingBits___61_comb};
  assign p1_concat_135082_comb = {p1_smul_57572_NarrowedMult__comb, p1_smul_57454_TrailingBits___29_comb};
  assign p1_concat_135083_comb = {p1_smul_57574_NarrowedMult__comb, p1_smul_57454_TrailingBits___30_comb};
  assign p1_concat_135084_comb = {p1_smul_57576_NarrowedMult__comb, p1_smul_57330_TrailingBits___62_comb};
  assign p1_concat_135085_comb = {p1_smul_57578_NarrowedMult__comb, p1_smul_57330_TrailingBits___63_comb};
  assign p1_concat_135086_comb = {p1_smul_57580_NarrowedMult__comb, p1_smul_57454_TrailingBits___31_comb};
  assign p1_smul_57584_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__1_squeezed_comb, 6'h27);
  assign p1_concat_135088_comb = {p1_smul_57588_NarrowedMult__comb, p1_smul_57330_TrailingBits___65_comb};
  assign p1_concat_135089_comb = {p1_smul_57590_NarrowedMult__comb, p1_smul_57330_TrailingBits___66_comb};
  assign p1_smul_57594_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__6_squeezed_comb, 6'h19);
  assign p1_smul_57600_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__9_squeezed_comb, 6'h27);
  assign p1_concat_135092_comb = {p1_smul_57604_NarrowedMult__comb, p1_smul_57330_TrailingBits___69_comb};
  assign p1_concat_135093_comb = {p1_smul_57606_NarrowedMult__comb, p1_smul_57330_TrailingBits___70_comb};
  assign p1_smul_57610_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__14_squeezed_comb, 6'h19);
  assign p1_smul_57680_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__49_squeezed_comb, 6'h27);
  assign p1_concat_135108_comb = {p1_smul_57684_NarrowedMult__comb, p1_smul_57330_TrailingBits___89_comb};
  assign p1_concat_135109_comb = {p1_smul_57686_NarrowedMult__comb, p1_smul_57330_TrailingBits___90_comb};
  assign p1_smul_57690_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__54_squeezed_comb, 6'h19);
  assign p1_smul_57696_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__57_squeezed_comb, 6'h27);
  assign p1_concat_135112_comb = {p1_smul_57700_NarrowedMult__comb, p1_smul_57330_TrailingBits___93_comb};
  assign p1_concat_135113_comb = {p1_smul_57702_NarrowedMult__comb, p1_smul_57330_TrailingBits___94_comb};
  assign p1_smul_57706_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__62_squeezed_comb, 6'h19);
  assign p1_concat_135115_comb = {p1_smul_57838_NarrowedMult__comb, p1_smul_57330_TrailingBits___96_comb};
  assign p1_smul_57842_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__2_squeezed_comb, 6'h27);
  assign p1_smul_57848_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__5_squeezed_comb, 6'h27);
  assign p1_concat_135118_comb = {p1_smul_57852_NarrowedMult__comb, p1_smul_57330_TrailingBits___99_comb};
  assign p1_concat_135119_comb = {p1_smul_57854_NarrowedMult__comb, p1_smul_57330_TrailingBits___100_comb};
  assign p1_smul_57858_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__10_squeezed_comb, 6'h27);
  assign p1_smul_57864_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__13_squeezed_comb, 6'h27);
  assign p1_concat_135122_comb = {p1_smul_57868_NarrowedMult__comb, p1_smul_57330_TrailingBits___103_comb};
  assign p1_concat_135135_comb = {p1_smul_57934_NarrowedMult__comb, p1_smul_57330_TrailingBits___120_comb};
  assign p1_smul_57938_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__50_squeezed_comb, 6'h27);
  assign p1_smul_57944_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__53_squeezed_comb, 6'h27);
  assign p1_concat_135138_comb = {p1_smul_57948_NarrowedMult__comb, p1_smul_57330_TrailingBits___123_comb};
  assign p1_concat_135139_comb = {p1_smul_57950_NarrowedMult__comb, p1_smul_57330_TrailingBits___124_comb};
  assign p1_smul_57954_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__58_squeezed_comb, 6'h27);
  assign p1_smul_57960_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__61_squeezed_comb, 6'h27);
  assign p1_concat_135142_comb = {p1_smul_57964_NarrowedMult__comb, p1_smul_57330_TrailingBits___127_comb};
  assign p1_concat_135143_comb = {p1_smul_57966_NarrowedMult__comb, p1_smul_57330_TrailingBits___128_comb};
  assign p1_concat_135144_comb = {p1_smul_57968_NarrowedMult__comb, p1_smul_57454_TrailingBits___32_comb};
  assign p1_concat_135145_comb = {p1_smul_57970_NarrowedMult__comb, p1_smul_57330_TrailingBits___129_comb};
  assign p1_concat_135146_comb = {p1_smul_57972_NarrowedMult__comb, p1_smul_57454_TrailingBits___33_comb};
  assign p1_concat_135147_comb = {p1_smul_57974_NarrowedMult__comb, p1_smul_57454_TrailingBits___34_comb};
  assign p1_concat_135148_comb = {p1_smul_57976_NarrowedMult__comb, p1_smul_57330_TrailingBits___130_comb};
  assign p1_concat_135149_comb = {p1_smul_57978_NarrowedMult__comb, p1_smul_57454_TrailingBits___35_comb};
  assign p1_concat_135150_comb = {p1_smul_57980_NarrowedMult__comb, p1_smul_57330_TrailingBits___131_comb};
  assign p1_concat_135151_comb = {p1_smul_57982_NarrowedMult__comb, p1_smul_57330_TrailingBits___132_comb};
  assign p1_concat_135152_comb = {p1_smul_57984_NarrowedMult__comb, p1_smul_57454_TrailingBits___36_comb};
  assign p1_concat_135153_comb = {p1_smul_57986_NarrowedMult__comb, p1_smul_57330_TrailingBits___133_comb};
  assign p1_concat_135154_comb = {p1_smul_57988_NarrowedMult__comb, p1_smul_57454_TrailingBits___37_comb};
  assign p1_concat_135155_comb = {p1_smul_57990_NarrowedMult__comb, p1_smul_57454_TrailingBits___38_comb};
  assign p1_concat_135156_comb = {p1_smul_57992_NarrowedMult__comb, p1_smul_57330_TrailingBits___134_comb};
  assign p1_concat_135157_comb = {p1_smul_57994_NarrowedMult__comb, p1_smul_57454_TrailingBits___39_comb};
  assign p1_concat_135158_comb = {p1_smul_57996_NarrowedMult__comb, p1_smul_57330_TrailingBits___135_comb};
  assign p1_concat_135159_comb = {p1_smul_58014_NarrowedMult__comb, p1_smul_57330_TrailingBits___140_comb};
  assign p1_concat_135160_comb = {p1_smul_58016_NarrowedMult__comb, p1_smul_57454_TrailingBits___44_comb};
  assign p1_concat_135161_comb = {p1_smul_58018_NarrowedMult__comb, p1_smul_57330_TrailingBits___141_comb};
  assign p1_concat_135162_comb = {p1_smul_58020_NarrowedMult__comb, p1_smul_57454_TrailingBits___45_comb};
  assign p1_concat_135163_comb = {p1_smul_58022_NarrowedMult__comb, p1_smul_57454_TrailingBits___46_comb};
  assign p1_concat_135164_comb = {p1_smul_58024_NarrowedMult__comb, p1_smul_57330_TrailingBits___142_comb};
  assign p1_concat_135165_comb = {p1_smul_58026_NarrowedMult__comb, p1_smul_57454_TrailingBits___47_comb};
  assign p1_concat_135166_comb = {p1_smul_58028_NarrowedMult__comb, p1_smul_57330_TrailingBits___143_comb};
  assign p1_concat_135167_comb = {p1_smul_58030_NarrowedMult__comb, p1_smul_57330_TrailingBits___144_comb};
  assign p1_concat_135168_comb = {p1_smul_58032_NarrowedMult__comb, p1_smul_57454_TrailingBits___48_comb};
  assign p1_concat_135169_comb = {p1_smul_58034_NarrowedMult__comb, p1_smul_57330_TrailingBits___145_comb};
  assign p1_concat_135170_comb = {p1_smul_58036_NarrowedMult__comb, p1_smul_57454_TrailingBits___49_comb};
  assign p1_concat_135171_comb = {p1_smul_58038_NarrowedMult__comb, p1_smul_57454_TrailingBits___50_comb};
  assign p1_concat_135172_comb = {p1_smul_58040_NarrowedMult__comb, p1_smul_57330_TrailingBits___146_comb};
  assign p1_concat_135173_comb = {p1_smul_58042_NarrowedMult__comb, p1_smul_57454_TrailingBits___51_comb};
  assign p1_concat_135174_comb = {p1_smul_58044_NarrowedMult__comb, p1_smul_57330_TrailingBits___147_comb};
  assign p1_concat_135175_comb = {p1_smul_58062_NarrowedMult__comb, p1_smul_57330_TrailingBits___152_comb};
  assign p1_concat_135176_comb = {p1_smul_58064_NarrowedMult__comb, p1_smul_57454_TrailingBits___56_comb};
  assign p1_concat_135177_comb = {p1_smul_58066_NarrowedMult__comb, p1_smul_57330_TrailingBits___153_comb};
  assign p1_concat_135178_comb = {p1_smul_58068_NarrowedMult__comb, p1_smul_57454_TrailingBits___57_comb};
  assign p1_concat_135179_comb = {p1_smul_58070_NarrowedMult__comb, p1_smul_57454_TrailingBits___58_comb};
  assign p1_concat_135180_comb = {p1_smul_58072_NarrowedMult__comb, p1_smul_57330_TrailingBits___154_comb};
  assign p1_concat_135181_comb = {p1_smul_58074_NarrowedMult__comb, p1_smul_57454_TrailingBits___59_comb};
  assign p1_concat_135182_comb = {p1_smul_58076_NarrowedMult__comb, p1_smul_57330_TrailingBits___155_comb};
  assign p1_concat_135183_comb = {p1_smul_58078_NarrowedMult__comb, p1_smul_57330_TrailingBits___156_comb};
  assign p1_concat_135184_comb = {p1_smul_58080_NarrowedMult__comb, p1_smul_57454_TrailingBits___60_comb};
  assign p1_concat_135185_comb = {p1_smul_58082_NarrowedMult__comb, p1_smul_57330_TrailingBits___157_comb};
  assign p1_concat_135186_comb = {p1_smul_58084_NarrowedMult__comb, p1_smul_57454_TrailingBits___61_comb};
  assign p1_concat_135187_comb = {p1_smul_58086_NarrowedMult__comb, p1_smul_57454_TrailingBits___62_comb};
  assign p1_concat_135188_comb = {p1_smul_58088_NarrowedMult__comb, p1_smul_57330_TrailingBits___158_comb};
  assign p1_concat_135189_comb = {p1_smul_58090_NarrowedMult__comb, p1_smul_57454_TrailingBits___63_comb};
  assign p1_concat_135190_comb = {p1_smul_58092_NarrowedMult__comb, p1_smul_57330_TrailingBits___159_comb};
  assign p1_smul_58094_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted_squeezed_comb, 6'h19);
  assign p1_concat_135192_comb = {p1_smul_58096_NarrowedMult__comb, p1_smul_57330_TrailingBits___161_comb};
  assign p1_concat_135193_comb = {p1_smul_58106_NarrowedMult__comb, p1_smul_57330_TrailingBits___162_comb};
  assign p1_smul_58108_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__7_squeezed_comb, 6'h19);
  assign p1_smul_58110_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__8_squeezed_comb, 6'h19);
  assign p1_concat_135196_comb = {p1_smul_58112_NarrowedMult__comb, p1_smul_57330_TrailingBits___165_comb};
  assign p1_concat_135197_comb = {p1_smul_58122_NarrowedMult__comb, p1_smul_57330_TrailingBits___166_comb};
  assign p1_smul_58124_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__15_squeezed_comb, 6'h19);
  assign p1_smul_58190_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__48_squeezed_comb, 6'h19);
  assign p1_concat_135212_comb = {p1_smul_58192_NarrowedMult__comb, p1_smul_57330_TrailingBits___185_comb};
  assign p1_concat_135213_comb = {p1_smul_58202_NarrowedMult__comb, p1_smul_57330_TrailingBits___186_comb};
  assign p1_smul_58204_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__55_squeezed_comb, 6'h19);
  assign p1_smul_58206_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__56_squeezed_comb, 6'h19);
  assign p1_concat_135216_comb = {p1_smul_58208_NarrowedMult__comb, p1_smul_57330_TrailingBits___189_comb};
  assign p1_concat_135217_comb = {p1_smul_58218_NarrowedMult__comb, p1_smul_57330_TrailingBits___190_comb};
  assign p1_smul_58220_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__63_squeezed_comb, 6'h19);
  assign p1_slt_135220_comb = $signed(p1_shifted__16_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135222_comb = $signed(p1_shifted__17_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135224_comb = $signed(p1_shifted__18_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135226_comb = $signed(p1_shifted__19_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135228_comb = $signed(p1_shifted__20_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135230_comb = $signed(p1_shifted__21_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135232_comb = $signed(p1_shifted__22_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135234_comb = $signed(p1_shifted__23_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135236_comb = $signed(p1_shifted__40_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135238_comb = $signed(p1_shifted__41_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135240_comb = $signed(p1_shifted__42_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135242_comb = $signed(p1_shifted__43_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135244_comb = $signed(p1_shifted__44_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135246_comb = $signed(p1_shifted__45_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135248_comb = $signed(p1_shifted__46_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135250_comb = $signed(p1_shifted__47_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135252_comb = $signed(p1_shifted_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135254_comb = $signed(p1_shifted__1_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135256_comb = $signed(p1_shifted__2_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135258_comb = $signed(p1_shifted__3_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135260_comb = $signed(p1_shifted__4_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135262_comb = $signed(p1_shifted__5_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135264_comb = $signed(p1_shifted__6_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135266_comb = $signed(p1_shifted__7_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135268_comb = $signed(p1_shifted__8_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135270_comb = $signed(p1_shifted__9_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135272_comb = $signed(p1_shifted__10_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135274_comb = $signed(p1_shifted__11_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135276_comb = $signed(p1_shifted__12_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135278_comb = $signed(p1_shifted__13_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135280_comb = $signed(p1_shifted__14_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135282_comb = $signed(p1_shifted__15_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135284_comb = $signed(p1_shifted__24_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135286_comb = $signed(p1_shifted__25_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135288_comb = $signed(p1_shifted__26_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135290_comb = $signed(p1_shifted__27_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135292_comb = $signed(p1_shifted__28_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135294_comb = $signed(p1_shifted__29_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135296_comb = $signed(p1_shifted__30_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135298_comb = $signed(p1_shifted__31_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135300_comb = $signed(p1_shifted__32_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135302_comb = $signed(p1_shifted__33_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135304_comb = $signed(p1_shifted__34_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135306_comb = $signed(p1_shifted__35_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135308_comb = $signed(p1_shifted__36_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135310_comb = $signed(p1_shifted__37_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135312_comb = $signed(p1_shifted__38_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135314_comb = $signed(p1_shifted__39_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135316_comb = $signed(p1_shifted__48_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135318_comb = $signed(p1_shifted__49_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135320_comb = $signed(p1_shifted__50_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135322_comb = $signed(p1_shifted__51_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135324_comb = $signed(p1_shifted__52_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135326_comb = $signed(p1_shifted__53_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135328_comb = $signed(p1_shifted__54_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135330_comb = $signed(p1_shifted__55_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135332_comb = $signed(p1_shifted__56_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135334_comb = $signed(p1_shifted__57_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135336_comb = $signed(p1_shifted__58_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135338_comb = $signed(p1_shifted__59_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135340_comb = $signed(p1_shifted__60_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135342_comb = $signed(p1_shifted__61_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135344_comb = $signed(p1_shifted__62_squeezed_comb) < $signed(8'h80);
  assign p1_slt_135346_comb = $signed(p1_shifted__63_squeezed_comb) < $signed(8'h80);
  assign p1_prod__199_comb = {{7{p1_concat_135019_comb[24]}}, p1_concat_135019_comb};
  assign p1_concat_135348_comb = {p1_smul_57380_NarrowedMult__comb, p1_smul_57330_TrailingBits___13_comb};
  assign p1_concat_135349_comb = {p1_smul_57382_NarrowedMult__comb, p1_smul_57330_TrailingBits___14_comb};
  assign p1_prod__214_comb = {{7{p1_concat_135024_comb[24]}}, p1_concat_135024_comb};
  assign p1_prod__263_comb = {{7{p1_concat_135025_comb[24]}}, p1_concat_135025_comb};
  assign p1_concat_135352_comb = {p1_smul_57396_NarrowedMult__comb, p1_smul_57330_TrailingBits___17_comb};
  assign p1_concat_135353_comb = {p1_smul_57398_NarrowedMult__comb, p1_smul_57330_TrailingBits___18_comb};
  assign p1_prod__278_comb = {{7{p1_concat_135030_comb[24]}}, p1_concat_135030_comb};
  assign p1_concat_135355_comb = {p1_smul_57632_NarrowedMult__comb, p1_smul_57330_TrailingBits___76_comb};
  assign p1_prod__216_comb = {{7{p1_concat_135097_comb[24]}}, p1_concat_135097_comb};
  assign p1_prod__223_comb = {{7{p1_concat_135098_comb[24]}}, p1_concat_135098_comb};
  assign p1_concat_135358_comb = {p1_smul_57642_NarrowedMult__comb, p1_smul_57330_TrailingBits___79_comb};
  assign p1_concat_135359_comb = {p1_smul_57648_NarrowedMult__comb, p1_smul_57330_TrailingBits___80_comb};
  assign p1_prod__280_comb = {{7{p1_concat_135103_comb[24]}}, p1_concat_135103_comb};
  assign p1_prod__287_comb = {{7{p1_concat_135104_comb[24]}}, p1_concat_135104_comb};
  assign p1_concat_135362_comb = {p1_smul_57658_NarrowedMult__comb, p1_smul_57330_TrailingBits___83_comb};
  assign p1_prod__212_comb = {{7{p1_concat_135123_comb[24]}}, p1_concat_135123_comb};
  assign p1_concat_135364_comb = {p1_smul_57890_NarrowedMult__comb, p1_smul_57330_TrailingBits___109_comb};
  assign p1_concat_135365_comb = {p1_smul_57896_NarrowedMult__comb, p1_smul_57330_TrailingBits___110_comb};
  assign p1_prod__250_comb = {{7{p1_concat_135128_comb[24]}}, p1_concat_135128_comb};
  assign p1_prod__276_comb = {{7{p1_concat_135129_comb[24]}}, p1_concat_135129_comb};
  assign p1_concat_135368_comb = {p1_smul_57906_NarrowedMult__comb, p1_smul_57330_TrailingBits___113_comb};
  assign p1_concat_135369_comb = {p1_smul_57912_NarrowedMult__comb, p1_smul_57330_TrailingBits___114_comb};
  assign p1_prod__314_comb = {{7{p1_concat_135134_comb[24]}}, p1_concat_135134_comb};
  assign p1_concat_135371_comb = {p1_smul_58142_NarrowedMult__comb, p1_smul_57330_TrailingBits___172_comb};
  assign p1_prod__234_comb = {{7{p1_concat_135201_comb[24]}}, p1_concat_135201_comb};
  assign p1_prod__254_comb = {{7{p1_concat_135202_comb[24]}}, p1_concat_135202_comb};
  assign p1_concat_135374_comb = {p1_smul_58156_NarrowedMult__comb, p1_smul_57330_TrailingBits___175_comb};
  assign p1_concat_135375_comb = {p1_smul_58158_NarrowedMult__comb, p1_smul_57330_TrailingBits___176_comb};
  assign p1_prod__298_comb = {{7{p1_concat_135207_comb[24]}}, p1_concat_135207_comb};
  assign p1_prod__318_comb = {{7{p1_concat_135208_comb[24]}}, p1_concat_135208_comb};
  assign p1_concat_135378_comb = {p1_smul_58172_NarrowedMult__comb, p1_smul_57330_TrailingBits___179_comb};
  assign p1_sgt_135507_comb = $signed(p1_shifted__16_comb) > $signed(16'h7fff);
  assign p1_sgt_135508_comb = $signed(p1_shifted__17_comb) > $signed(16'h7fff);
  assign p1_sgt_135509_comb = $signed(p1_shifted__18_comb) > $signed(16'h7fff);
  assign p1_sgt_135510_comb = $signed(p1_shifted__19_comb) > $signed(16'h7fff);
  assign p1_sgt_135511_comb = $signed(p1_shifted__20_comb) > $signed(16'h7fff);
  assign p1_sgt_135512_comb = $signed(p1_shifted__21_comb) > $signed(16'h7fff);
  assign p1_sgt_135513_comb = $signed(p1_shifted__22_comb) > $signed(16'h7fff);
  assign p1_sgt_135514_comb = $signed(p1_shifted__23_comb) > $signed(16'h7fff);
  assign p1_sgt_135515_comb = $signed(p1_shifted__40_comb) > $signed(16'h7fff);
  assign p1_sgt_135516_comb = $signed(p1_shifted__41_comb) > $signed(16'h7fff);
  assign p1_sgt_135517_comb = $signed(p1_shifted__42_comb) > $signed(16'h7fff);
  assign p1_sgt_135518_comb = $signed(p1_shifted__43_comb) > $signed(16'h7fff);
  assign p1_sgt_135519_comb = $signed(p1_shifted__44_comb) > $signed(16'h7fff);
  assign p1_sgt_135520_comb = $signed(p1_shifted__45_comb) > $signed(16'h7fff);
  assign p1_sgt_135521_comb = $signed(p1_shifted__46_comb) > $signed(16'h7fff);
  assign p1_sgt_135522_comb = $signed(p1_shifted__47_comb) > $signed(16'h7fff);
  assign p1_sgt_135523_comb = $signed(p1_shifted_comb) > $signed(16'h7fff);
  assign p1_sgt_135524_comb = $signed(p1_shifted__1_comb) > $signed(16'h7fff);
  assign p1_sgt_135525_comb = $signed(p1_shifted__2_comb) > $signed(16'h7fff);
  assign p1_sgt_135526_comb = $signed(p1_shifted__3_comb) > $signed(16'h7fff);
  assign p1_sgt_135527_comb = $signed(p1_shifted__4_comb) > $signed(16'h7fff);
  assign p1_sgt_135528_comb = $signed(p1_shifted__5_comb) > $signed(16'h7fff);
  assign p1_sgt_135529_comb = $signed(p1_shifted__6_comb) > $signed(16'h7fff);
  assign p1_sgt_135530_comb = $signed(p1_shifted__7_comb) > $signed(16'h7fff);
  assign p1_sgt_135531_comb = $signed(p1_shifted__8_comb) > $signed(16'h7fff);
  assign p1_sgt_135532_comb = $signed(p1_shifted__9_comb) > $signed(16'h7fff);
  assign p1_sgt_135533_comb = $signed(p1_shifted__10_comb) > $signed(16'h7fff);
  assign p1_sgt_135534_comb = $signed(p1_shifted__11_comb) > $signed(16'h7fff);
  assign p1_sgt_135535_comb = $signed(p1_shifted__12_comb) > $signed(16'h7fff);
  assign p1_sgt_135536_comb = $signed(p1_shifted__13_comb) > $signed(16'h7fff);
  assign p1_sgt_135537_comb = $signed(p1_shifted__14_comb) > $signed(16'h7fff);
  assign p1_sgt_135538_comb = $signed(p1_shifted__15_comb) > $signed(16'h7fff);
  assign p1_sgt_135539_comb = $signed(p1_shifted__24_comb) > $signed(16'h7fff);
  assign p1_sgt_135540_comb = $signed(p1_shifted__25_comb) > $signed(16'h7fff);
  assign p1_sgt_135541_comb = $signed(p1_shifted__26_comb) > $signed(16'h7fff);
  assign p1_sgt_135542_comb = $signed(p1_shifted__27_comb) > $signed(16'h7fff);
  assign p1_sgt_135543_comb = $signed(p1_shifted__28_comb) > $signed(16'h7fff);
  assign p1_sgt_135544_comb = $signed(p1_shifted__29_comb) > $signed(16'h7fff);
  assign p1_sgt_135545_comb = $signed(p1_shifted__30_comb) > $signed(16'h7fff);
  assign p1_sgt_135546_comb = $signed(p1_shifted__31_comb) > $signed(16'h7fff);
  assign p1_sgt_135547_comb = $signed(p1_shifted__32_comb) > $signed(16'h7fff);
  assign p1_sgt_135548_comb = $signed(p1_shifted__33_comb) > $signed(16'h7fff);
  assign p1_sgt_135549_comb = $signed(p1_shifted__34_comb) > $signed(16'h7fff);
  assign p1_sgt_135550_comb = $signed(p1_shifted__35_comb) > $signed(16'h7fff);
  assign p1_sgt_135551_comb = $signed(p1_shifted__36_comb) > $signed(16'h7fff);
  assign p1_sgt_135552_comb = $signed(p1_shifted__37_comb) > $signed(16'h7fff);
  assign p1_sgt_135553_comb = $signed(p1_shifted__38_comb) > $signed(16'h7fff);
  assign p1_sgt_135554_comb = $signed(p1_shifted__39_comb) > $signed(16'h7fff);
  assign p1_sgt_135555_comb = $signed(p1_shifted__48_comb) > $signed(16'h7fff);
  assign p1_sgt_135556_comb = $signed(p1_shifted__49_comb) > $signed(16'h7fff);
  assign p1_sgt_135557_comb = $signed(p1_shifted__50_comb) > $signed(16'h7fff);
  assign p1_sgt_135558_comb = $signed(p1_shifted__51_comb) > $signed(16'h7fff);
  assign p1_sgt_135559_comb = $signed(p1_shifted__52_comb) > $signed(16'h7fff);
  assign p1_sgt_135560_comb = $signed(p1_shifted__53_comb) > $signed(16'h7fff);
  assign p1_sgt_135561_comb = $signed(p1_shifted__54_comb) > $signed(16'h7fff);
  assign p1_sgt_135562_comb = $signed(p1_shifted__55_comb) > $signed(16'h7fff);
  assign p1_sgt_135563_comb = $signed(p1_shifted__56_comb) > $signed(16'h7fff);
  assign p1_sgt_135564_comb = $signed(p1_shifted__57_comb) > $signed(16'h7fff);
  assign p1_sgt_135565_comb = $signed(p1_shifted__58_comb) > $signed(16'h7fff);
  assign p1_sgt_135566_comb = $signed(p1_shifted__59_comb) > $signed(16'h7fff);
  assign p1_sgt_135567_comb = $signed(p1_shifted__60_comb) > $signed(16'h7fff);
  assign p1_sgt_135568_comb = $signed(p1_shifted__61_comb) > $signed(16'h7fff);
  assign p1_sgt_135569_comb = $signed(p1_shifted__62_comb) > $signed(16'h7fff);
  assign p1_sgt_135570_comb = $signed(p1_shifted__63_comb) > $signed(16'h7fff);

  // Registers for pipe stage 1:
  reg [7:0] p1_shifted__18_squeezed;
  reg [7:0] p1_shifted__21_squeezed;
  reg [7:0] p1_shifted__42_squeezed;
  reg [7:0] p1_shifted__45_squeezed;
  reg [7:0] p1_shifted__16_squeezed;
  reg [7:0] p1_shifted__17_squeezed;
  reg [7:0] p1_shifted__19_squeezed;
  reg [7:0] p1_shifted__20_squeezed;
  reg [7:0] p1_shifted__22_squeezed;
  reg [7:0] p1_shifted__23_squeezed;
  reg [7:0] p1_shifted__40_squeezed;
  reg [7:0] p1_shifted__41_squeezed;
  reg [7:0] p1_shifted__43_squeezed;
  reg [7:0] p1_shifted__44_squeezed;
  reg [7:0] p1_shifted__46_squeezed;
  reg [7:0] p1_shifted__47_squeezed;
  reg [7:0] p1_shifted__2_squeezed;
  reg [7:0] p1_shifted__5_squeezed;
  reg [7:0] p1_shifted__10_squeezed;
  reg [7:0] p1_shifted__13_squeezed;
  reg [7:0] p1_shifted__26_squeezed;
  reg [7:0] p1_shifted__29_squeezed;
  reg [7:0] p1_shifted__34_squeezed;
  reg [7:0] p1_shifted__37_squeezed;
  reg [7:0] p1_shifted__50_squeezed;
  reg [7:0] p1_shifted__53_squeezed;
  reg [7:0] p1_shifted__58_squeezed;
  reg [7:0] p1_shifted__61_squeezed;
  reg [7:0] p1_shifted_squeezed;
  reg [7:0] p1_shifted__1_squeezed;
  reg [7:0] p1_shifted__3_squeezed;
  reg [7:0] p1_shifted__4_squeezed;
  reg [7:0] p1_shifted__6_squeezed;
  reg [7:0] p1_shifted__7_squeezed;
  reg [7:0] p1_shifted__8_squeezed;
  reg [7:0] p1_shifted__9_squeezed;
  reg [7:0] p1_shifted__11_squeezed;
  reg [7:0] p1_shifted__12_squeezed;
  reg [7:0] p1_shifted__14_squeezed;
  reg [7:0] p1_shifted__15_squeezed;
  reg [7:0] p1_shifted__24_squeezed;
  reg [7:0] p1_shifted__25_squeezed;
  reg [7:0] p1_shifted__27_squeezed;
  reg [7:0] p1_shifted__28_squeezed;
  reg [7:0] p1_shifted__30_squeezed;
  reg [7:0] p1_shifted__31_squeezed;
  reg [7:0] p1_shifted__32_squeezed;
  reg [7:0] p1_shifted__33_squeezed;
  reg [7:0] p1_shifted__35_squeezed;
  reg [7:0] p1_shifted__36_squeezed;
  reg [7:0] p1_shifted__38_squeezed;
  reg [7:0] p1_shifted__39_squeezed;
  reg [7:0] p1_shifted__48_squeezed;
  reg [7:0] p1_shifted__49_squeezed;
  reg [7:0] p1_shifted__51_squeezed;
  reg [7:0] p1_shifted__52_squeezed;
  reg [7:0] p1_shifted__54_squeezed;
  reg [7:0] p1_shifted__55_squeezed;
  reg [7:0] p1_shifted__56_squeezed;
  reg [7:0] p1_shifted__57_squeezed;
  reg [7:0] p1_shifted__59_squeezed;
  reg [7:0] p1_shifted__60_squeezed;
  reg [7:0] p1_shifted__62_squeezed;
  reg [7:0] p1_shifted__63_squeezed;
  reg [14:0] p1_smul_57488_NarrowedMult_;
  reg [14:0] p1_smul_57490_NarrowedMult_;
  reg [14:0] p1_smul_57496_NarrowedMult_;
  reg [14:0] p1_smul_57498_NarrowedMult_;
  reg [14:0] p1_smul_57536_NarrowedMult_;
  reg [14:0] p1_smul_57538_NarrowedMult_;
  reg [14:0] p1_smul_57544_NarrowedMult_;
  reg [14:0] p1_smul_57546_NarrowedMult_;
  reg [14:0] p1_smul_57998_NarrowedMult_;
  reg [14:0] p1_smul_58002_NarrowedMult_;
  reg [14:0] p1_smul_58008_NarrowedMult_;
  reg [14:0] p1_smul_58012_NarrowedMult_;
  reg [14:0] p1_smul_58046_NarrowedMult_;
  reg [14:0] p1_smul_58050_NarrowedMult_;
  reg [14:0] p1_smul_58056_NarrowedMult_;
  reg [14:0] p1_smul_58060_NarrowedMult_;
  reg [14:0] p1_smul_57456_NarrowedMult_;
  reg [14:0] p1_smul_57458_NarrowedMult_;
  reg [14:0] p1_smul_57464_NarrowedMult_;
  reg [14:0] p1_smul_57466_NarrowedMult_;
  reg [14:0] p1_smul_57472_NarrowedMult_;
  reg [14:0] p1_smul_57474_NarrowedMult_;
  reg [14:0] p1_smul_57480_NarrowedMult_;
  reg [14:0] p1_smul_57482_NarrowedMult_;
  reg [14:0] p1_smul_57504_NarrowedMult_;
  reg [14:0] p1_smul_57506_NarrowedMult_;
  reg [14:0] p1_smul_57512_NarrowedMult_;
  reg [14:0] p1_smul_57514_NarrowedMult_;
  reg [14:0] p1_smul_57520_NarrowedMult_;
  reg [14:0] p1_smul_57522_NarrowedMult_;
  reg [14:0] p1_smul_57528_NarrowedMult_;
  reg [14:0] p1_smul_57530_NarrowedMult_;
  reg [14:0] p1_smul_57552_NarrowedMult_;
  reg [14:0] p1_smul_57554_NarrowedMult_;
  reg [14:0] p1_smul_57560_NarrowedMult_;
  reg [14:0] p1_smul_57562_NarrowedMult_;
  reg [14:0] p1_smul_57568_NarrowedMult_;
  reg [14:0] p1_smul_57570_NarrowedMult_;
  reg [14:0] p1_smul_57576_NarrowedMult_;
  reg [14:0] p1_smul_57578_NarrowedMult_;
  reg [14:0] p1_smul_57966_NarrowedMult_;
  reg [14:0] p1_smul_57970_NarrowedMult_;
  reg [14:0] p1_smul_57976_NarrowedMult_;
  reg [14:0] p1_smul_57980_NarrowedMult_;
  reg [14:0] p1_smul_57982_NarrowedMult_;
  reg [14:0] p1_smul_57986_NarrowedMult_;
  reg [14:0] p1_smul_57992_NarrowedMult_;
  reg [14:0] p1_smul_57996_NarrowedMult_;
  reg [14:0] p1_smul_58014_NarrowedMult_;
  reg [14:0] p1_smul_58018_NarrowedMult_;
  reg [14:0] p1_smul_58024_NarrowedMult_;
  reg [14:0] p1_smul_58028_NarrowedMult_;
  reg [14:0] p1_smul_58030_NarrowedMult_;
  reg [14:0] p1_smul_58034_NarrowedMult_;
  reg [14:0] p1_smul_58040_NarrowedMult_;
  reg [14:0] p1_smul_58044_NarrowedMult_;
  reg [14:0] p1_smul_58062_NarrowedMult_;
  reg [14:0] p1_smul_58066_NarrowedMult_;
  reg [14:0] p1_smul_58072_NarrowedMult_;
  reg [14:0] p1_smul_58076_NarrowedMult_;
  reg [14:0] p1_smul_58078_NarrowedMult_;
  reg [14:0] p1_smul_58082_NarrowedMult_;
  reg [14:0] p1_smul_58088_NarrowedMult_;
  reg [14:0] p1_smul_58092_NarrowedMult_;
  reg [24:0] p1_concat_134899;
  reg [13:0] p1_smul_57364_NarrowedMult_;
  reg [13:0] p1_smul_57366_NarrowedMult_;
  reg [24:0] p1_concat_134902;
  reg [24:0] p1_concat_134903;
  reg [13:0] p1_smul_57412_NarrowedMult_;
  reg [13:0] p1_smul_57414_NarrowedMult_;
  reg [24:0] p1_concat_134906;
  reg [24:0] p1_concat_134907;
  reg [23:0] p1_concat_134908;
  reg [23:0] p1_concat_134909;
  reg [24:0] p1_concat_134910;
  reg [24:0] p1_concat_134911;
  reg [23:0] p1_concat_134912;
  reg [23:0] p1_concat_134913;
  reg [24:0] p1_concat_134914;
  reg [24:0] p1_concat_134915;
  reg [23:0] p1_concat_134916;
  reg [23:0] p1_concat_134917;
  reg [24:0] p1_concat_134918;
  reg [24:0] p1_concat_134919;
  reg [23:0] p1_concat_134920;
  reg [23:0] p1_concat_134921;
  reg [24:0] p1_concat_134922;
  reg [13:0] p1_smul_57616_NarrowedMult_;
  reg [24:0] p1_concat_134924;
  reg [24:0] p1_concat_134925;
  reg [13:0] p1_smul_57626_NarrowedMult_;
  reg [13:0] p1_smul_57664_NarrowedMult_;
  reg [24:0] p1_concat_134928;
  reg [24:0] p1_concat_134929;
  reg [13:0] p1_smul_57674_NarrowedMult_;
  reg [24:0] p1_concat_134931;
  reg [13:0] p1_smul_57874_NarrowedMult_;
  reg [13:0] p1_smul_57880_NarrowedMult_;
  reg [24:0] p1_concat_134934;
  reg [24:0] p1_concat_134935;
  reg [13:0] p1_smul_57922_NarrowedMult_;
  reg [13:0] p1_smul_57928_NarrowedMult_;
  reg [24:0] p1_concat_134938;
  reg [23:0] p1_concat_134939;
  reg [24:0] p1_concat_134940;
  reg [23:0] p1_concat_134941;
  reg [24:0] p1_concat_134942;
  reg [24:0] p1_concat_134943;
  reg [23:0] p1_concat_134944;
  reg [24:0] p1_concat_134945;
  reg [23:0] p1_concat_134946;
  reg [23:0] p1_concat_134947;
  reg [24:0] p1_concat_134948;
  reg [23:0] p1_concat_134949;
  reg [24:0] p1_concat_134950;
  reg [24:0] p1_concat_134951;
  reg [23:0] p1_concat_134952;
  reg [24:0] p1_concat_134953;
  reg [23:0] p1_concat_134954;
  reg [13:0] p1_smul_58126_NarrowedMult_;
  reg [24:0] p1_concat_134956;
  reg [24:0] p1_concat_134957;
  reg [13:0] p1_smul_58140_NarrowedMult_;
  reg [13:0] p1_smul_58174_NarrowedMult_;
  reg [24:0] p1_concat_134960;
  reg [24:0] p1_concat_134961;
  reg [13:0] p1_smul_58188_NarrowedMult_;
  reg [24:0] p1_concat_135011;
  reg [13:0] p1_smul_57332_NarrowedMult_;
  reg [13:0] p1_smul_57334_NarrowedMult_;
  reg [24:0] p1_concat_135014;
  reg [24:0] p1_concat_135015;
  reg [13:0] p1_smul_57348_NarrowedMult_;
  reg [13:0] p1_smul_57350_NarrowedMult_;
  reg [24:0] p1_concat_135018;
  reg [24:0] p1_concat_135031;
  reg [13:0] p1_smul_57428_NarrowedMult_;
  reg [13:0] p1_smul_57430_NarrowedMult_;
  reg [24:0] p1_concat_135034;
  reg [24:0] p1_concat_135035;
  reg [13:0] p1_smul_57444_NarrowedMult_;
  reg [13:0] p1_smul_57446_NarrowedMult_;
  reg [24:0] p1_concat_135038;
  reg [24:0] p1_concat_135039;
  reg [23:0] p1_concat_135040;
  reg [23:0] p1_concat_135041;
  reg [24:0] p1_concat_135042;
  reg [24:0] p1_concat_135043;
  reg [23:0] p1_concat_135044;
  reg [23:0] p1_concat_135045;
  reg [24:0] p1_concat_135046;
  reg [24:0] p1_concat_135047;
  reg [23:0] p1_concat_135048;
  reg [23:0] p1_concat_135049;
  reg [24:0] p1_concat_135050;
  reg [24:0] p1_concat_135051;
  reg [23:0] p1_concat_135052;
  reg [23:0] p1_concat_135053;
  reg [24:0] p1_concat_135054;
  reg [24:0] p1_concat_135055;
  reg [23:0] p1_concat_135056;
  reg [23:0] p1_concat_135057;
  reg [24:0] p1_concat_135058;
  reg [24:0] p1_concat_135059;
  reg [23:0] p1_concat_135060;
  reg [23:0] p1_concat_135061;
  reg [24:0] p1_concat_135062;
  reg [24:0] p1_concat_135063;
  reg [23:0] p1_concat_135064;
  reg [23:0] p1_concat_135065;
  reg [24:0] p1_concat_135066;
  reg [24:0] p1_concat_135067;
  reg [23:0] p1_concat_135068;
  reg [23:0] p1_concat_135069;
  reg [24:0] p1_concat_135070;
  reg [24:0] p1_concat_135071;
  reg [23:0] p1_concat_135072;
  reg [23:0] p1_concat_135073;
  reg [24:0] p1_concat_135074;
  reg [24:0] p1_concat_135075;
  reg [23:0] p1_concat_135076;
  reg [23:0] p1_concat_135077;
  reg [24:0] p1_concat_135078;
  reg [24:0] p1_concat_135079;
  reg [23:0] p1_concat_135080;
  reg [23:0] p1_concat_135081;
  reg [24:0] p1_concat_135082;
  reg [24:0] p1_concat_135083;
  reg [23:0] p1_concat_135084;
  reg [23:0] p1_concat_135085;
  reg [24:0] p1_concat_135086;
  reg [13:0] p1_smul_57584_NarrowedMult_;
  reg [24:0] p1_concat_135088;
  reg [24:0] p1_concat_135089;
  reg [13:0] p1_smul_57594_NarrowedMult_;
  reg [13:0] p1_smul_57600_NarrowedMult_;
  reg [24:0] p1_concat_135092;
  reg [24:0] p1_concat_135093;
  reg [13:0] p1_smul_57610_NarrowedMult_;
  reg [13:0] p1_smul_57680_NarrowedMult_;
  reg [24:0] p1_concat_135108;
  reg [24:0] p1_concat_135109;
  reg [13:0] p1_smul_57690_NarrowedMult_;
  reg [13:0] p1_smul_57696_NarrowedMult_;
  reg [24:0] p1_concat_135112;
  reg [24:0] p1_concat_135113;
  reg [13:0] p1_smul_57706_NarrowedMult_;
  reg [24:0] p1_concat_135115;
  reg [13:0] p1_smul_57842_NarrowedMult_;
  reg [13:0] p1_smul_57848_NarrowedMult_;
  reg [24:0] p1_concat_135118;
  reg [24:0] p1_concat_135119;
  reg [13:0] p1_smul_57858_NarrowedMult_;
  reg [13:0] p1_smul_57864_NarrowedMult_;
  reg [24:0] p1_concat_135122;
  reg [24:0] p1_concat_135135;
  reg [13:0] p1_smul_57938_NarrowedMult_;
  reg [13:0] p1_smul_57944_NarrowedMult_;
  reg [24:0] p1_concat_135138;
  reg [24:0] p1_concat_135139;
  reg [13:0] p1_smul_57954_NarrowedMult_;
  reg [13:0] p1_smul_57960_NarrowedMult_;
  reg [24:0] p1_concat_135142;
  reg [23:0] p1_concat_135143;
  reg [24:0] p1_concat_135144;
  reg [23:0] p1_concat_135145;
  reg [24:0] p1_concat_135146;
  reg [24:0] p1_concat_135147;
  reg [23:0] p1_concat_135148;
  reg [24:0] p1_concat_135149;
  reg [23:0] p1_concat_135150;
  reg [23:0] p1_concat_135151;
  reg [24:0] p1_concat_135152;
  reg [23:0] p1_concat_135153;
  reg [24:0] p1_concat_135154;
  reg [24:0] p1_concat_135155;
  reg [23:0] p1_concat_135156;
  reg [24:0] p1_concat_135157;
  reg [23:0] p1_concat_135158;
  reg [23:0] p1_concat_135159;
  reg [24:0] p1_concat_135160;
  reg [23:0] p1_concat_135161;
  reg [24:0] p1_concat_135162;
  reg [24:0] p1_concat_135163;
  reg [23:0] p1_concat_135164;
  reg [24:0] p1_concat_135165;
  reg [23:0] p1_concat_135166;
  reg [23:0] p1_concat_135167;
  reg [24:0] p1_concat_135168;
  reg [23:0] p1_concat_135169;
  reg [24:0] p1_concat_135170;
  reg [24:0] p1_concat_135171;
  reg [23:0] p1_concat_135172;
  reg [24:0] p1_concat_135173;
  reg [23:0] p1_concat_135174;
  reg [23:0] p1_concat_135175;
  reg [24:0] p1_concat_135176;
  reg [23:0] p1_concat_135177;
  reg [24:0] p1_concat_135178;
  reg [24:0] p1_concat_135179;
  reg [23:0] p1_concat_135180;
  reg [24:0] p1_concat_135181;
  reg [23:0] p1_concat_135182;
  reg [23:0] p1_concat_135183;
  reg [24:0] p1_concat_135184;
  reg [23:0] p1_concat_135185;
  reg [24:0] p1_concat_135186;
  reg [24:0] p1_concat_135187;
  reg [23:0] p1_concat_135188;
  reg [24:0] p1_concat_135189;
  reg [23:0] p1_concat_135190;
  reg [13:0] p1_smul_58094_NarrowedMult_;
  reg [24:0] p1_concat_135192;
  reg [24:0] p1_concat_135193;
  reg [13:0] p1_smul_58108_NarrowedMult_;
  reg [13:0] p1_smul_58110_NarrowedMult_;
  reg [24:0] p1_concat_135196;
  reg [24:0] p1_concat_135197;
  reg [13:0] p1_smul_58124_NarrowedMult_;
  reg [13:0] p1_smul_58190_NarrowedMult_;
  reg [24:0] p1_concat_135212;
  reg [24:0] p1_concat_135213;
  reg [13:0] p1_smul_58204_NarrowedMult_;
  reg [13:0] p1_smul_58206_NarrowedMult_;
  reg [24:0] p1_concat_135216;
  reg [24:0] p1_concat_135217;
  reg [13:0] p1_smul_58220_NarrowedMult_;
  reg p1_slt_135220;
  reg p1_slt_135222;
  reg p1_slt_135224;
  reg p1_slt_135226;
  reg p1_slt_135228;
  reg p1_slt_135230;
  reg p1_slt_135232;
  reg p1_slt_135234;
  reg p1_slt_135236;
  reg p1_slt_135238;
  reg p1_slt_135240;
  reg p1_slt_135242;
  reg p1_slt_135244;
  reg p1_slt_135246;
  reg p1_slt_135248;
  reg p1_slt_135250;
  reg p1_slt_135252;
  reg p1_slt_135254;
  reg p1_slt_135256;
  reg p1_slt_135258;
  reg p1_slt_135260;
  reg p1_slt_135262;
  reg p1_slt_135264;
  reg p1_slt_135266;
  reg p1_slt_135268;
  reg p1_slt_135270;
  reg p1_slt_135272;
  reg p1_slt_135274;
  reg p1_slt_135276;
  reg p1_slt_135278;
  reg p1_slt_135280;
  reg p1_slt_135282;
  reg p1_slt_135284;
  reg p1_slt_135286;
  reg p1_slt_135288;
  reg p1_slt_135290;
  reg p1_slt_135292;
  reg p1_slt_135294;
  reg p1_slt_135296;
  reg p1_slt_135298;
  reg p1_slt_135300;
  reg p1_slt_135302;
  reg p1_slt_135304;
  reg p1_slt_135306;
  reg p1_slt_135308;
  reg p1_slt_135310;
  reg p1_slt_135312;
  reg p1_slt_135314;
  reg p1_slt_135316;
  reg p1_slt_135318;
  reg p1_slt_135320;
  reg p1_slt_135322;
  reg p1_slt_135324;
  reg p1_slt_135326;
  reg p1_slt_135328;
  reg p1_slt_135330;
  reg p1_slt_135332;
  reg p1_slt_135334;
  reg p1_slt_135336;
  reg p1_slt_135338;
  reg p1_slt_135340;
  reg p1_slt_135342;
  reg p1_slt_135344;
  reg p1_slt_135346;
  reg [31:0] p1_prod__199;
  reg [22:0] p1_concat_135348;
  reg [22:0] p1_concat_135349;
  reg [31:0] p1_prod__214;
  reg [31:0] p1_prod__263;
  reg [22:0] p1_concat_135352;
  reg [22:0] p1_concat_135353;
  reg [31:0] p1_prod__278;
  reg [22:0] p1_concat_135355;
  reg [31:0] p1_prod__216;
  reg [31:0] p1_prod__223;
  reg [22:0] p1_concat_135358;
  reg [22:0] p1_concat_135359;
  reg [31:0] p1_prod__280;
  reg [31:0] p1_prod__287;
  reg [22:0] p1_concat_135362;
  reg [31:0] p1_prod__212;
  reg [22:0] p1_concat_135364;
  reg [22:0] p1_concat_135365;
  reg [31:0] p1_prod__250;
  reg [31:0] p1_prod__276;
  reg [22:0] p1_concat_135368;
  reg [22:0] p1_concat_135369;
  reg [31:0] p1_prod__314;
  reg [22:0] p1_concat_135371;
  reg [31:0] p1_prod__234;
  reg [31:0] p1_prod__254;
  reg [22:0] p1_concat_135374;
  reg [22:0] p1_concat_135375;
  reg [31:0] p1_prod__298;
  reg [31:0] p1_prod__318;
  reg [22:0] p1_concat_135378;
  reg p1_sgt_135507;
  reg p1_sgt_135508;
  reg p1_sgt_135509;
  reg p1_sgt_135510;
  reg p1_sgt_135511;
  reg p1_sgt_135512;
  reg p1_sgt_135513;
  reg p1_sgt_135514;
  reg p1_sgt_135515;
  reg p1_sgt_135516;
  reg p1_sgt_135517;
  reg p1_sgt_135518;
  reg p1_sgt_135519;
  reg p1_sgt_135520;
  reg p1_sgt_135521;
  reg p1_sgt_135522;
  reg p1_sgt_135523;
  reg p1_sgt_135524;
  reg p1_sgt_135525;
  reg p1_sgt_135526;
  reg p1_sgt_135527;
  reg p1_sgt_135528;
  reg p1_sgt_135529;
  reg p1_sgt_135530;
  reg p1_sgt_135531;
  reg p1_sgt_135532;
  reg p1_sgt_135533;
  reg p1_sgt_135534;
  reg p1_sgt_135535;
  reg p1_sgt_135536;
  reg p1_sgt_135537;
  reg p1_sgt_135538;
  reg p1_sgt_135539;
  reg p1_sgt_135540;
  reg p1_sgt_135541;
  reg p1_sgt_135542;
  reg p1_sgt_135543;
  reg p1_sgt_135544;
  reg p1_sgt_135545;
  reg p1_sgt_135546;
  reg p1_sgt_135547;
  reg p1_sgt_135548;
  reg p1_sgt_135549;
  reg p1_sgt_135550;
  reg p1_sgt_135551;
  reg p1_sgt_135552;
  reg p1_sgt_135553;
  reg p1_sgt_135554;
  reg p1_sgt_135555;
  reg p1_sgt_135556;
  reg p1_sgt_135557;
  reg p1_sgt_135558;
  reg p1_sgt_135559;
  reg p1_sgt_135560;
  reg p1_sgt_135561;
  reg p1_sgt_135562;
  reg p1_sgt_135563;
  reg p1_sgt_135564;
  reg p1_sgt_135565;
  reg p1_sgt_135566;
  reg p1_sgt_135567;
  reg p1_sgt_135568;
  reg p1_sgt_135569;
  reg p1_sgt_135570;
  always @ (posedge clk) begin
    p1_shifted__18_squeezed <= p1_shifted__18_squeezed_comb;
    p1_shifted__21_squeezed <= p1_shifted__21_squeezed_comb;
    p1_shifted__42_squeezed <= p1_shifted__42_squeezed_comb;
    p1_shifted__45_squeezed <= p1_shifted__45_squeezed_comb;
    p1_shifted__16_squeezed <= p1_shifted__16_squeezed_comb;
    p1_shifted__17_squeezed <= p1_shifted__17_squeezed_comb;
    p1_shifted__19_squeezed <= p1_shifted__19_squeezed_comb;
    p1_shifted__20_squeezed <= p1_shifted__20_squeezed_comb;
    p1_shifted__22_squeezed <= p1_shifted__22_squeezed_comb;
    p1_shifted__23_squeezed <= p1_shifted__23_squeezed_comb;
    p1_shifted__40_squeezed <= p1_shifted__40_squeezed_comb;
    p1_shifted__41_squeezed <= p1_shifted__41_squeezed_comb;
    p1_shifted__43_squeezed <= p1_shifted__43_squeezed_comb;
    p1_shifted__44_squeezed <= p1_shifted__44_squeezed_comb;
    p1_shifted__46_squeezed <= p1_shifted__46_squeezed_comb;
    p1_shifted__47_squeezed <= p1_shifted__47_squeezed_comb;
    p1_shifted__2_squeezed <= p1_shifted__2_squeezed_comb;
    p1_shifted__5_squeezed <= p1_shifted__5_squeezed_comb;
    p1_shifted__10_squeezed <= p1_shifted__10_squeezed_comb;
    p1_shifted__13_squeezed <= p1_shifted__13_squeezed_comb;
    p1_shifted__26_squeezed <= p1_shifted__26_squeezed_comb;
    p1_shifted__29_squeezed <= p1_shifted__29_squeezed_comb;
    p1_shifted__34_squeezed <= p1_shifted__34_squeezed_comb;
    p1_shifted__37_squeezed <= p1_shifted__37_squeezed_comb;
    p1_shifted__50_squeezed <= p1_shifted__50_squeezed_comb;
    p1_shifted__53_squeezed <= p1_shifted__53_squeezed_comb;
    p1_shifted__58_squeezed <= p1_shifted__58_squeezed_comb;
    p1_shifted__61_squeezed <= p1_shifted__61_squeezed_comb;
    p1_shifted_squeezed <= p1_shifted_squeezed_comb;
    p1_shifted__1_squeezed <= p1_shifted__1_squeezed_comb;
    p1_shifted__3_squeezed <= p1_shifted__3_squeezed_comb;
    p1_shifted__4_squeezed <= p1_shifted__4_squeezed_comb;
    p1_shifted__6_squeezed <= p1_shifted__6_squeezed_comb;
    p1_shifted__7_squeezed <= p1_shifted__7_squeezed_comb;
    p1_shifted__8_squeezed <= p1_shifted__8_squeezed_comb;
    p1_shifted__9_squeezed <= p1_shifted__9_squeezed_comb;
    p1_shifted__11_squeezed <= p1_shifted__11_squeezed_comb;
    p1_shifted__12_squeezed <= p1_shifted__12_squeezed_comb;
    p1_shifted__14_squeezed <= p1_shifted__14_squeezed_comb;
    p1_shifted__15_squeezed <= p1_shifted__15_squeezed_comb;
    p1_shifted__24_squeezed <= p1_shifted__24_squeezed_comb;
    p1_shifted__25_squeezed <= p1_shifted__25_squeezed_comb;
    p1_shifted__27_squeezed <= p1_shifted__27_squeezed_comb;
    p1_shifted__28_squeezed <= p1_shifted__28_squeezed_comb;
    p1_shifted__30_squeezed <= p1_shifted__30_squeezed_comb;
    p1_shifted__31_squeezed <= p1_shifted__31_squeezed_comb;
    p1_shifted__32_squeezed <= p1_shifted__32_squeezed_comb;
    p1_shifted__33_squeezed <= p1_shifted__33_squeezed_comb;
    p1_shifted__35_squeezed <= p1_shifted__35_squeezed_comb;
    p1_shifted__36_squeezed <= p1_shifted__36_squeezed_comb;
    p1_shifted__38_squeezed <= p1_shifted__38_squeezed_comb;
    p1_shifted__39_squeezed <= p1_shifted__39_squeezed_comb;
    p1_shifted__48_squeezed <= p1_shifted__48_squeezed_comb;
    p1_shifted__49_squeezed <= p1_shifted__49_squeezed_comb;
    p1_shifted__51_squeezed <= p1_shifted__51_squeezed_comb;
    p1_shifted__52_squeezed <= p1_shifted__52_squeezed_comb;
    p1_shifted__54_squeezed <= p1_shifted__54_squeezed_comb;
    p1_shifted__55_squeezed <= p1_shifted__55_squeezed_comb;
    p1_shifted__56_squeezed <= p1_shifted__56_squeezed_comb;
    p1_shifted__57_squeezed <= p1_shifted__57_squeezed_comb;
    p1_shifted__59_squeezed <= p1_shifted__59_squeezed_comb;
    p1_shifted__60_squeezed <= p1_shifted__60_squeezed_comb;
    p1_shifted__62_squeezed <= p1_shifted__62_squeezed_comb;
    p1_shifted__63_squeezed <= p1_shifted__63_squeezed_comb;
    p1_smul_57488_NarrowedMult_ <= p1_smul_57488_NarrowedMult__comb;
    p1_smul_57490_NarrowedMult_ <= p1_smul_57490_NarrowedMult__comb;
    p1_smul_57496_NarrowedMult_ <= p1_smul_57496_NarrowedMult__comb;
    p1_smul_57498_NarrowedMult_ <= p1_smul_57498_NarrowedMult__comb;
    p1_smul_57536_NarrowedMult_ <= p1_smul_57536_NarrowedMult__comb;
    p1_smul_57538_NarrowedMult_ <= p1_smul_57538_NarrowedMult__comb;
    p1_smul_57544_NarrowedMult_ <= p1_smul_57544_NarrowedMult__comb;
    p1_smul_57546_NarrowedMult_ <= p1_smul_57546_NarrowedMult__comb;
    p1_smul_57998_NarrowedMult_ <= p1_smul_57998_NarrowedMult__comb;
    p1_smul_58002_NarrowedMult_ <= p1_smul_58002_NarrowedMult__comb;
    p1_smul_58008_NarrowedMult_ <= p1_smul_58008_NarrowedMult__comb;
    p1_smul_58012_NarrowedMult_ <= p1_smul_58012_NarrowedMult__comb;
    p1_smul_58046_NarrowedMult_ <= p1_smul_58046_NarrowedMult__comb;
    p1_smul_58050_NarrowedMult_ <= p1_smul_58050_NarrowedMult__comb;
    p1_smul_58056_NarrowedMult_ <= p1_smul_58056_NarrowedMult__comb;
    p1_smul_58060_NarrowedMult_ <= p1_smul_58060_NarrowedMult__comb;
    p1_smul_57456_NarrowedMult_ <= p1_smul_57456_NarrowedMult__comb;
    p1_smul_57458_NarrowedMult_ <= p1_smul_57458_NarrowedMult__comb;
    p1_smul_57464_NarrowedMult_ <= p1_smul_57464_NarrowedMult__comb;
    p1_smul_57466_NarrowedMult_ <= p1_smul_57466_NarrowedMult__comb;
    p1_smul_57472_NarrowedMult_ <= p1_smul_57472_NarrowedMult__comb;
    p1_smul_57474_NarrowedMult_ <= p1_smul_57474_NarrowedMult__comb;
    p1_smul_57480_NarrowedMult_ <= p1_smul_57480_NarrowedMult__comb;
    p1_smul_57482_NarrowedMult_ <= p1_smul_57482_NarrowedMult__comb;
    p1_smul_57504_NarrowedMult_ <= p1_smul_57504_NarrowedMult__comb;
    p1_smul_57506_NarrowedMult_ <= p1_smul_57506_NarrowedMult__comb;
    p1_smul_57512_NarrowedMult_ <= p1_smul_57512_NarrowedMult__comb;
    p1_smul_57514_NarrowedMult_ <= p1_smul_57514_NarrowedMult__comb;
    p1_smul_57520_NarrowedMult_ <= p1_smul_57520_NarrowedMult__comb;
    p1_smul_57522_NarrowedMult_ <= p1_smul_57522_NarrowedMult__comb;
    p1_smul_57528_NarrowedMult_ <= p1_smul_57528_NarrowedMult__comb;
    p1_smul_57530_NarrowedMult_ <= p1_smul_57530_NarrowedMult__comb;
    p1_smul_57552_NarrowedMult_ <= p1_smul_57552_NarrowedMult__comb;
    p1_smul_57554_NarrowedMult_ <= p1_smul_57554_NarrowedMult__comb;
    p1_smul_57560_NarrowedMult_ <= p1_smul_57560_NarrowedMult__comb;
    p1_smul_57562_NarrowedMult_ <= p1_smul_57562_NarrowedMult__comb;
    p1_smul_57568_NarrowedMult_ <= p1_smul_57568_NarrowedMult__comb;
    p1_smul_57570_NarrowedMult_ <= p1_smul_57570_NarrowedMult__comb;
    p1_smul_57576_NarrowedMult_ <= p1_smul_57576_NarrowedMult__comb;
    p1_smul_57578_NarrowedMult_ <= p1_smul_57578_NarrowedMult__comb;
    p1_smul_57966_NarrowedMult_ <= p1_smul_57966_NarrowedMult__comb;
    p1_smul_57970_NarrowedMult_ <= p1_smul_57970_NarrowedMult__comb;
    p1_smul_57976_NarrowedMult_ <= p1_smul_57976_NarrowedMult__comb;
    p1_smul_57980_NarrowedMult_ <= p1_smul_57980_NarrowedMult__comb;
    p1_smul_57982_NarrowedMult_ <= p1_smul_57982_NarrowedMult__comb;
    p1_smul_57986_NarrowedMult_ <= p1_smul_57986_NarrowedMult__comb;
    p1_smul_57992_NarrowedMult_ <= p1_smul_57992_NarrowedMult__comb;
    p1_smul_57996_NarrowedMult_ <= p1_smul_57996_NarrowedMult__comb;
    p1_smul_58014_NarrowedMult_ <= p1_smul_58014_NarrowedMult__comb;
    p1_smul_58018_NarrowedMult_ <= p1_smul_58018_NarrowedMult__comb;
    p1_smul_58024_NarrowedMult_ <= p1_smul_58024_NarrowedMult__comb;
    p1_smul_58028_NarrowedMult_ <= p1_smul_58028_NarrowedMult__comb;
    p1_smul_58030_NarrowedMult_ <= p1_smul_58030_NarrowedMult__comb;
    p1_smul_58034_NarrowedMult_ <= p1_smul_58034_NarrowedMult__comb;
    p1_smul_58040_NarrowedMult_ <= p1_smul_58040_NarrowedMult__comb;
    p1_smul_58044_NarrowedMult_ <= p1_smul_58044_NarrowedMult__comb;
    p1_smul_58062_NarrowedMult_ <= p1_smul_58062_NarrowedMult__comb;
    p1_smul_58066_NarrowedMult_ <= p1_smul_58066_NarrowedMult__comb;
    p1_smul_58072_NarrowedMult_ <= p1_smul_58072_NarrowedMult__comb;
    p1_smul_58076_NarrowedMult_ <= p1_smul_58076_NarrowedMult__comb;
    p1_smul_58078_NarrowedMult_ <= p1_smul_58078_NarrowedMult__comb;
    p1_smul_58082_NarrowedMult_ <= p1_smul_58082_NarrowedMult__comb;
    p1_smul_58088_NarrowedMult_ <= p1_smul_58088_NarrowedMult__comb;
    p1_smul_58092_NarrowedMult_ <= p1_smul_58092_NarrowedMult__comb;
    p1_concat_134899 <= p1_concat_134899_comb;
    p1_smul_57364_NarrowedMult_ <= p1_smul_57364_NarrowedMult__comb;
    p1_smul_57366_NarrowedMult_ <= p1_smul_57366_NarrowedMult__comb;
    p1_concat_134902 <= p1_concat_134902_comb;
    p1_concat_134903 <= p1_concat_134903_comb;
    p1_smul_57412_NarrowedMult_ <= p1_smul_57412_NarrowedMult__comb;
    p1_smul_57414_NarrowedMult_ <= p1_smul_57414_NarrowedMult__comb;
    p1_concat_134906 <= p1_concat_134906_comb;
    p1_concat_134907 <= p1_concat_134907_comb;
    p1_concat_134908 <= p1_concat_134908_comb;
    p1_concat_134909 <= p1_concat_134909_comb;
    p1_concat_134910 <= p1_concat_134910_comb;
    p1_concat_134911 <= p1_concat_134911_comb;
    p1_concat_134912 <= p1_concat_134912_comb;
    p1_concat_134913 <= p1_concat_134913_comb;
    p1_concat_134914 <= p1_concat_134914_comb;
    p1_concat_134915 <= p1_concat_134915_comb;
    p1_concat_134916 <= p1_concat_134916_comb;
    p1_concat_134917 <= p1_concat_134917_comb;
    p1_concat_134918 <= p1_concat_134918_comb;
    p1_concat_134919 <= p1_concat_134919_comb;
    p1_concat_134920 <= p1_concat_134920_comb;
    p1_concat_134921 <= p1_concat_134921_comb;
    p1_concat_134922 <= p1_concat_134922_comb;
    p1_smul_57616_NarrowedMult_ <= p1_smul_57616_NarrowedMult__comb;
    p1_concat_134924 <= p1_concat_134924_comb;
    p1_concat_134925 <= p1_concat_134925_comb;
    p1_smul_57626_NarrowedMult_ <= p1_smul_57626_NarrowedMult__comb;
    p1_smul_57664_NarrowedMult_ <= p1_smul_57664_NarrowedMult__comb;
    p1_concat_134928 <= p1_concat_134928_comb;
    p1_concat_134929 <= p1_concat_134929_comb;
    p1_smul_57674_NarrowedMult_ <= p1_smul_57674_NarrowedMult__comb;
    p1_concat_134931 <= p1_concat_134931_comb;
    p1_smul_57874_NarrowedMult_ <= p1_smul_57874_NarrowedMult__comb;
    p1_smul_57880_NarrowedMult_ <= p1_smul_57880_NarrowedMult__comb;
    p1_concat_134934 <= p1_concat_134934_comb;
    p1_concat_134935 <= p1_concat_134935_comb;
    p1_smul_57922_NarrowedMult_ <= p1_smul_57922_NarrowedMult__comb;
    p1_smul_57928_NarrowedMult_ <= p1_smul_57928_NarrowedMult__comb;
    p1_concat_134938 <= p1_concat_134938_comb;
    p1_concat_134939 <= p1_concat_134939_comb;
    p1_concat_134940 <= p1_concat_134940_comb;
    p1_concat_134941 <= p1_concat_134941_comb;
    p1_concat_134942 <= p1_concat_134942_comb;
    p1_concat_134943 <= p1_concat_134943_comb;
    p1_concat_134944 <= p1_concat_134944_comb;
    p1_concat_134945 <= p1_concat_134945_comb;
    p1_concat_134946 <= p1_concat_134946_comb;
    p1_concat_134947 <= p1_concat_134947_comb;
    p1_concat_134948 <= p1_concat_134948_comb;
    p1_concat_134949 <= p1_concat_134949_comb;
    p1_concat_134950 <= p1_concat_134950_comb;
    p1_concat_134951 <= p1_concat_134951_comb;
    p1_concat_134952 <= p1_concat_134952_comb;
    p1_concat_134953 <= p1_concat_134953_comb;
    p1_concat_134954 <= p1_concat_134954_comb;
    p1_smul_58126_NarrowedMult_ <= p1_smul_58126_NarrowedMult__comb;
    p1_concat_134956 <= p1_concat_134956_comb;
    p1_concat_134957 <= p1_concat_134957_comb;
    p1_smul_58140_NarrowedMult_ <= p1_smul_58140_NarrowedMult__comb;
    p1_smul_58174_NarrowedMult_ <= p1_smul_58174_NarrowedMult__comb;
    p1_concat_134960 <= p1_concat_134960_comb;
    p1_concat_134961 <= p1_concat_134961_comb;
    p1_smul_58188_NarrowedMult_ <= p1_smul_58188_NarrowedMult__comb;
    p1_concat_135011 <= p1_concat_135011_comb;
    p1_smul_57332_NarrowedMult_ <= p1_smul_57332_NarrowedMult__comb;
    p1_smul_57334_NarrowedMult_ <= p1_smul_57334_NarrowedMult__comb;
    p1_concat_135014 <= p1_concat_135014_comb;
    p1_concat_135015 <= p1_concat_135015_comb;
    p1_smul_57348_NarrowedMult_ <= p1_smul_57348_NarrowedMult__comb;
    p1_smul_57350_NarrowedMult_ <= p1_smul_57350_NarrowedMult__comb;
    p1_concat_135018 <= p1_concat_135018_comb;
    p1_concat_135031 <= p1_concat_135031_comb;
    p1_smul_57428_NarrowedMult_ <= p1_smul_57428_NarrowedMult__comb;
    p1_smul_57430_NarrowedMult_ <= p1_smul_57430_NarrowedMult__comb;
    p1_concat_135034 <= p1_concat_135034_comb;
    p1_concat_135035 <= p1_concat_135035_comb;
    p1_smul_57444_NarrowedMult_ <= p1_smul_57444_NarrowedMult__comb;
    p1_smul_57446_NarrowedMult_ <= p1_smul_57446_NarrowedMult__comb;
    p1_concat_135038 <= p1_concat_135038_comb;
    p1_concat_135039 <= p1_concat_135039_comb;
    p1_concat_135040 <= p1_concat_135040_comb;
    p1_concat_135041 <= p1_concat_135041_comb;
    p1_concat_135042 <= p1_concat_135042_comb;
    p1_concat_135043 <= p1_concat_135043_comb;
    p1_concat_135044 <= p1_concat_135044_comb;
    p1_concat_135045 <= p1_concat_135045_comb;
    p1_concat_135046 <= p1_concat_135046_comb;
    p1_concat_135047 <= p1_concat_135047_comb;
    p1_concat_135048 <= p1_concat_135048_comb;
    p1_concat_135049 <= p1_concat_135049_comb;
    p1_concat_135050 <= p1_concat_135050_comb;
    p1_concat_135051 <= p1_concat_135051_comb;
    p1_concat_135052 <= p1_concat_135052_comb;
    p1_concat_135053 <= p1_concat_135053_comb;
    p1_concat_135054 <= p1_concat_135054_comb;
    p1_concat_135055 <= p1_concat_135055_comb;
    p1_concat_135056 <= p1_concat_135056_comb;
    p1_concat_135057 <= p1_concat_135057_comb;
    p1_concat_135058 <= p1_concat_135058_comb;
    p1_concat_135059 <= p1_concat_135059_comb;
    p1_concat_135060 <= p1_concat_135060_comb;
    p1_concat_135061 <= p1_concat_135061_comb;
    p1_concat_135062 <= p1_concat_135062_comb;
    p1_concat_135063 <= p1_concat_135063_comb;
    p1_concat_135064 <= p1_concat_135064_comb;
    p1_concat_135065 <= p1_concat_135065_comb;
    p1_concat_135066 <= p1_concat_135066_comb;
    p1_concat_135067 <= p1_concat_135067_comb;
    p1_concat_135068 <= p1_concat_135068_comb;
    p1_concat_135069 <= p1_concat_135069_comb;
    p1_concat_135070 <= p1_concat_135070_comb;
    p1_concat_135071 <= p1_concat_135071_comb;
    p1_concat_135072 <= p1_concat_135072_comb;
    p1_concat_135073 <= p1_concat_135073_comb;
    p1_concat_135074 <= p1_concat_135074_comb;
    p1_concat_135075 <= p1_concat_135075_comb;
    p1_concat_135076 <= p1_concat_135076_comb;
    p1_concat_135077 <= p1_concat_135077_comb;
    p1_concat_135078 <= p1_concat_135078_comb;
    p1_concat_135079 <= p1_concat_135079_comb;
    p1_concat_135080 <= p1_concat_135080_comb;
    p1_concat_135081 <= p1_concat_135081_comb;
    p1_concat_135082 <= p1_concat_135082_comb;
    p1_concat_135083 <= p1_concat_135083_comb;
    p1_concat_135084 <= p1_concat_135084_comb;
    p1_concat_135085 <= p1_concat_135085_comb;
    p1_concat_135086 <= p1_concat_135086_comb;
    p1_smul_57584_NarrowedMult_ <= p1_smul_57584_NarrowedMult__comb;
    p1_concat_135088 <= p1_concat_135088_comb;
    p1_concat_135089 <= p1_concat_135089_comb;
    p1_smul_57594_NarrowedMult_ <= p1_smul_57594_NarrowedMult__comb;
    p1_smul_57600_NarrowedMult_ <= p1_smul_57600_NarrowedMult__comb;
    p1_concat_135092 <= p1_concat_135092_comb;
    p1_concat_135093 <= p1_concat_135093_comb;
    p1_smul_57610_NarrowedMult_ <= p1_smul_57610_NarrowedMult__comb;
    p1_smul_57680_NarrowedMult_ <= p1_smul_57680_NarrowedMult__comb;
    p1_concat_135108 <= p1_concat_135108_comb;
    p1_concat_135109 <= p1_concat_135109_comb;
    p1_smul_57690_NarrowedMult_ <= p1_smul_57690_NarrowedMult__comb;
    p1_smul_57696_NarrowedMult_ <= p1_smul_57696_NarrowedMult__comb;
    p1_concat_135112 <= p1_concat_135112_comb;
    p1_concat_135113 <= p1_concat_135113_comb;
    p1_smul_57706_NarrowedMult_ <= p1_smul_57706_NarrowedMult__comb;
    p1_concat_135115 <= p1_concat_135115_comb;
    p1_smul_57842_NarrowedMult_ <= p1_smul_57842_NarrowedMult__comb;
    p1_smul_57848_NarrowedMult_ <= p1_smul_57848_NarrowedMult__comb;
    p1_concat_135118 <= p1_concat_135118_comb;
    p1_concat_135119 <= p1_concat_135119_comb;
    p1_smul_57858_NarrowedMult_ <= p1_smul_57858_NarrowedMult__comb;
    p1_smul_57864_NarrowedMult_ <= p1_smul_57864_NarrowedMult__comb;
    p1_concat_135122 <= p1_concat_135122_comb;
    p1_concat_135135 <= p1_concat_135135_comb;
    p1_smul_57938_NarrowedMult_ <= p1_smul_57938_NarrowedMult__comb;
    p1_smul_57944_NarrowedMult_ <= p1_smul_57944_NarrowedMult__comb;
    p1_concat_135138 <= p1_concat_135138_comb;
    p1_concat_135139 <= p1_concat_135139_comb;
    p1_smul_57954_NarrowedMult_ <= p1_smul_57954_NarrowedMult__comb;
    p1_smul_57960_NarrowedMult_ <= p1_smul_57960_NarrowedMult__comb;
    p1_concat_135142 <= p1_concat_135142_comb;
    p1_concat_135143 <= p1_concat_135143_comb;
    p1_concat_135144 <= p1_concat_135144_comb;
    p1_concat_135145 <= p1_concat_135145_comb;
    p1_concat_135146 <= p1_concat_135146_comb;
    p1_concat_135147 <= p1_concat_135147_comb;
    p1_concat_135148 <= p1_concat_135148_comb;
    p1_concat_135149 <= p1_concat_135149_comb;
    p1_concat_135150 <= p1_concat_135150_comb;
    p1_concat_135151 <= p1_concat_135151_comb;
    p1_concat_135152 <= p1_concat_135152_comb;
    p1_concat_135153 <= p1_concat_135153_comb;
    p1_concat_135154 <= p1_concat_135154_comb;
    p1_concat_135155 <= p1_concat_135155_comb;
    p1_concat_135156 <= p1_concat_135156_comb;
    p1_concat_135157 <= p1_concat_135157_comb;
    p1_concat_135158 <= p1_concat_135158_comb;
    p1_concat_135159 <= p1_concat_135159_comb;
    p1_concat_135160 <= p1_concat_135160_comb;
    p1_concat_135161 <= p1_concat_135161_comb;
    p1_concat_135162 <= p1_concat_135162_comb;
    p1_concat_135163 <= p1_concat_135163_comb;
    p1_concat_135164 <= p1_concat_135164_comb;
    p1_concat_135165 <= p1_concat_135165_comb;
    p1_concat_135166 <= p1_concat_135166_comb;
    p1_concat_135167 <= p1_concat_135167_comb;
    p1_concat_135168 <= p1_concat_135168_comb;
    p1_concat_135169 <= p1_concat_135169_comb;
    p1_concat_135170 <= p1_concat_135170_comb;
    p1_concat_135171 <= p1_concat_135171_comb;
    p1_concat_135172 <= p1_concat_135172_comb;
    p1_concat_135173 <= p1_concat_135173_comb;
    p1_concat_135174 <= p1_concat_135174_comb;
    p1_concat_135175 <= p1_concat_135175_comb;
    p1_concat_135176 <= p1_concat_135176_comb;
    p1_concat_135177 <= p1_concat_135177_comb;
    p1_concat_135178 <= p1_concat_135178_comb;
    p1_concat_135179 <= p1_concat_135179_comb;
    p1_concat_135180 <= p1_concat_135180_comb;
    p1_concat_135181 <= p1_concat_135181_comb;
    p1_concat_135182 <= p1_concat_135182_comb;
    p1_concat_135183 <= p1_concat_135183_comb;
    p1_concat_135184 <= p1_concat_135184_comb;
    p1_concat_135185 <= p1_concat_135185_comb;
    p1_concat_135186 <= p1_concat_135186_comb;
    p1_concat_135187 <= p1_concat_135187_comb;
    p1_concat_135188 <= p1_concat_135188_comb;
    p1_concat_135189 <= p1_concat_135189_comb;
    p1_concat_135190 <= p1_concat_135190_comb;
    p1_smul_58094_NarrowedMult_ <= p1_smul_58094_NarrowedMult__comb;
    p1_concat_135192 <= p1_concat_135192_comb;
    p1_concat_135193 <= p1_concat_135193_comb;
    p1_smul_58108_NarrowedMult_ <= p1_smul_58108_NarrowedMult__comb;
    p1_smul_58110_NarrowedMult_ <= p1_smul_58110_NarrowedMult__comb;
    p1_concat_135196 <= p1_concat_135196_comb;
    p1_concat_135197 <= p1_concat_135197_comb;
    p1_smul_58124_NarrowedMult_ <= p1_smul_58124_NarrowedMult__comb;
    p1_smul_58190_NarrowedMult_ <= p1_smul_58190_NarrowedMult__comb;
    p1_concat_135212 <= p1_concat_135212_comb;
    p1_concat_135213 <= p1_concat_135213_comb;
    p1_smul_58204_NarrowedMult_ <= p1_smul_58204_NarrowedMult__comb;
    p1_smul_58206_NarrowedMult_ <= p1_smul_58206_NarrowedMult__comb;
    p1_concat_135216 <= p1_concat_135216_comb;
    p1_concat_135217 <= p1_concat_135217_comb;
    p1_smul_58220_NarrowedMult_ <= p1_smul_58220_NarrowedMult__comb;
    p1_slt_135220 <= p1_slt_135220_comb;
    p1_slt_135222 <= p1_slt_135222_comb;
    p1_slt_135224 <= p1_slt_135224_comb;
    p1_slt_135226 <= p1_slt_135226_comb;
    p1_slt_135228 <= p1_slt_135228_comb;
    p1_slt_135230 <= p1_slt_135230_comb;
    p1_slt_135232 <= p1_slt_135232_comb;
    p1_slt_135234 <= p1_slt_135234_comb;
    p1_slt_135236 <= p1_slt_135236_comb;
    p1_slt_135238 <= p1_slt_135238_comb;
    p1_slt_135240 <= p1_slt_135240_comb;
    p1_slt_135242 <= p1_slt_135242_comb;
    p1_slt_135244 <= p1_slt_135244_comb;
    p1_slt_135246 <= p1_slt_135246_comb;
    p1_slt_135248 <= p1_slt_135248_comb;
    p1_slt_135250 <= p1_slt_135250_comb;
    p1_slt_135252 <= p1_slt_135252_comb;
    p1_slt_135254 <= p1_slt_135254_comb;
    p1_slt_135256 <= p1_slt_135256_comb;
    p1_slt_135258 <= p1_slt_135258_comb;
    p1_slt_135260 <= p1_slt_135260_comb;
    p1_slt_135262 <= p1_slt_135262_comb;
    p1_slt_135264 <= p1_slt_135264_comb;
    p1_slt_135266 <= p1_slt_135266_comb;
    p1_slt_135268 <= p1_slt_135268_comb;
    p1_slt_135270 <= p1_slt_135270_comb;
    p1_slt_135272 <= p1_slt_135272_comb;
    p1_slt_135274 <= p1_slt_135274_comb;
    p1_slt_135276 <= p1_slt_135276_comb;
    p1_slt_135278 <= p1_slt_135278_comb;
    p1_slt_135280 <= p1_slt_135280_comb;
    p1_slt_135282 <= p1_slt_135282_comb;
    p1_slt_135284 <= p1_slt_135284_comb;
    p1_slt_135286 <= p1_slt_135286_comb;
    p1_slt_135288 <= p1_slt_135288_comb;
    p1_slt_135290 <= p1_slt_135290_comb;
    p1_slt_135292 <= p1_slt_135292_comb;
    p1_slt_135294 <= p1_slt_135294_comb;
    p1_slt_135296 <= p1_slt_135296_comb;
    p1_slt_135298 <= p1_slt_135298_comb;
    p1_slt_135300 <= p1_slt_135300_comb;
    p1_slt_135302 <= p1_slt_135302_comb;
    p1_slt_135304 <= p1_slt_135304_comb;
    p1_slt_135306 <= p1_slt_135306_comb;
    p1_slt_135308 <= p1_slt_135308_comb;
    p1_slt_135310 <= p1_slt_135310_comb;
    p1_slt_135312 <= p1_slt_135312_comb;
    p1_slt_135314 <= p1_slt_135314_comb;
    p1_slt_135316 <= p1_slt_135316_comb;
    p1_slt_135318 <= p1_slt_135318_comb;
    p1_slt_135320 <= p1_slt_135320_comb;
    p1_slt_135322 <= p1_slt_135322_comb;
    p1_slt_135324 <= p1_slt_135324_comb;
    p1_slt_135326 <= p1_slt_135326_comb;
    p1_slt_135328 <= p1_slt_135328_comb;
    p1_slt_135330 <= p1_slt_135330_comb;
    p1_slt_135332 <= p1_slt_135332_comb;
    p1_slt_135334 <= p1_slt_135334_comb;
    p1_slt_135336 <= p1_slt_135336_comb;
    p1_slt_135338 <= p1_slt_135338_comb;
    p1_slt_135340 <= p1_slt_135340_comb;
    p1_slt_135342 <= p1_slt_135342_comb;
    p1_slt_135344 <= p1_slt_135344_comb;
    p1_slt_135346 <= p1_slt_135346_comb;
    p1_prod__199 <= p1_prod__199_comb;
    p1_concat_135348 <= p1_concat_135348_comb;
    p1_concat_135349 <= p1_concat_135349_comb;
    p1_prod__214 <= p1_prod__214_comb;
    p1_prod__263 <= p1_prod__263_comb;
    p1_concat_135352 <= p1_concat_135352_comb;
    p1_concat_135353 <= p1_concat_135353_comb;
    p1_prod__278 <= p1_prod__278_comb;
    p1_concat_135355 <= p1_concat_135355_comb;
    p1_prod__216 <= p1_prod__216_comb;
    p1_prod__223 <= p1_prod__223_comb;
    p1_concat_135358 <= p1_concat_135358_comb;
    p1_concat_135359 <= p1_concat_135359_comb;
    p1_prod__280 <= p1_prod__280_comb;
    p1_prod__287 <= p1_prod__287_comb;
    p1_concat_135362 <= p1_concat_135362_comb;
    p1_prod__212 <= p1_prod__212_comb;
    p1_concat_135364 <= p1_concat_135364_comb;
    p1_concat_135365 <= p1_concat_135365_comb;
    p1_prod__250 <= p1_prod__250_comb;
    p1_prod__276 <= p1_prod__276_comb;
    p1_concat_135368 <= p1_concat_135368_comb;
    p1_concat_135369 <= p1_concat_135369_comb;
    p1_prod__314 <= p1_prod__314_comb;
    p1_concat_135371 <= p1_concat_135371_comb;
    p1_prod__234 <= p1_prod__234_comb;
    p1_prod__254 <= p1_prod__254_comb;
    p1_concat_135374 <= p1_concat_135374_comb;
    p1_concat_135375 <= p1_concat_135375_comb;
    p1_prod__298 <= p1_prod__298_comb;
    p1_prod__318 <= p1_prod__318_comb;
    p1_concat_135378 <= p1_concat_135378_comb;
    p1_sgt_135507 <= p1_sgt_135507_comb;
    p1_sgt_135508 <= p1_sgt_135508_comb;
    p1_sgt_135509 <= p1_sgt_135509_comb;
    p1_sgt_135510 <= p1_sgt_135510_comb;
    p1_sgt_135511 <= p1_sgt_135511_comb;
    p1_sgt_135512 <= p1_sgt_135512_comb;
    p1_sgt_135513 <= p1_sgt_135513_comb;
    p1_sgt_135514 <= p1_sgt_135514_comb;
    p1_sgt_135515 <= p1_sgt_135515_comb;
    p1_sgt_135516 <= p1_sgt_135516_comb;
    p1_sgt_135517 <= p1_sgt_135517_comb;
    p1_sgt_135518 <= p1_sgt_135518_comb;
    p1_sgt_135519 <= p1_sgt_135519_comb;
    p1_sgt_135520 <= p1_sgt_135520_comb;
    p1_sgt_135521 <= p1_sgt_135521_comb;
    p1_sgt_135522 <= p1_sgt_135522_comb;
    p1_sgt_135523 <= p1_sgt_135523_comb;
    p1_sgt_135524 <= p1_sgt_135524_comb;
    p1_sgt_135525 <= p1_sgt_135525_comb;
    p1_sgt_135526 <= p1_sgt_135526_comb;
    p1_sgt_135527 <= p1_sgt_135527_comb;
    p1_sgt_135528 <= p1_sgt_135528_comb;
    p1_sgt_135529 <= p1_sgt_135529_comb;
    p1_sgt_135530 <= p1_sgt_135530_comb;
    p1_sgt_135531 <= p1_sgt_135531_comb;
    p1_sgt_135532 <= p1_sgt_135532_comb;
    p1_sgt_135533 <= p1_sgt_135533_comb;
    p1_sgt_135534 <= p1_sgt_135534_comb;
    p1_sgt_135535 <= p1_sgt_135535_comb;
    p1_sgt_135536 <= p1_sgt_135536_comb;
    p1_sgt_135537 <= p1_sgt_135537_comb;
    p1_sgt_135538 <= p1_sgt_135538_comb;
    p1_sgt_135539 <= p1_sgt_135539_comb;
    p1_sgt_135540 <= p1_sgt_135540_comb;
    p1_sgt_135541 <= p1_sgt_135541_comb;
    p1_sgt_135542 <= p1_sgt_135542_comb;
    p1_sgt_135543 <= p1_sgt_135543_comb;
    p1_sgt_135544 <= p1_sgt_135544_comb;
    p1_sgt_135545 <= p1_sgt_135545_comb;
    p1_sgt_135546 <= p1_sgt_135546_comb;
    p1_sgt_135547 <= p1_sgt_135547_comb;
    p1_sgt_135548 <= p1_sgt_135548_comb;
    p1_sgt_135549 <= p1_sgt_135549_comb;
    p1_sgt_135550 <= p1_sgt_135550_comb;
    p1_sgt_135551 <= p1_sgt_135551_comb;
    p1_sgt_135552 <= p1_sgt_135552_comb;
    p1_sgt_135553 <= p1_sgt_135553_comb;
    p1_sgt_135554 <= p1_sgt_135554_comb;
    p1_sgt_135555 <= p1_sgt_135555_comb;
    p1_sgt_135556 <= p1_sgt_135556_comb;
    p1_sgt_135557 <= p1_sgt_135557_comb;
    p1_sgt_135558 <= p1_sgt_135558_comb;
    p1_sgt_135559 <= p1_sgt_135559_comb;
    p1_sgt_135560 <= p1_sgt_135560_comb;
    p1_sgt_135561 <= p1_sgt_135561_comb;
    p1_sgt_135562 <= p1_sgt_135562_comb;
    p1_sgt_135563 <= p1_sgt_135563_comb;
    p1_sgt_135564 <= p1_sgt_135564_comb;
    p1_sgt_135565 <= p1_sgt_135565_comb;
    p1_sgt_135566 <= p1_sgt_135566_comb;
    p1_sgt_135567 <= p1_sgt_135567_comb;
    p1_sgt_135568 <= p1_sgt_135568_comb;
    p1_sgt_135569 <= p1_sgt_135569_comb;
    p1_sgt_135570 <= p1_sgt_135570_comb;
  end

  // ===== Pipe stage 2:
  wire [8:0] p2_smul_57330_TrailingBits___9_comb;
  wire [8:0] p2_smul_57330_TrailingBits___10_comb;
  wire [8:0] p2_smul_57330_TrailingBits___21_comb;
  wire [8:0] p2_smul_57330_TrailingBits___22_comb;
  wire [8:0] p2_smul_57330_TrailingBits___72_comb;
  wire [8:0] p2_smul_57330_TrailingBits___75_comb;
  wire [8:0] p2_smul_57330_TrailingBits___84_comb;
  wire [8:0] p2_smul_57330_TrailingBits___87_comb;
  wire [8:0] p2_smul_57330_TrailingBits___105_comb;
  wire [8:0] p2_smul_57330_TrailingBits___106_comb;
  wire [8:0] p2_smul_57330_TrailingBits___117_comb;
  wire [8:0] p2_smul_57330_TrailingBits___118_comb;
  wire [8:0] p2_smul_57330_TrailingBits___168_comb;
  wire [8:0] p2_smul_57330_TrailingBits___171_comb;
  wire [8:0] p2_smul_57330_TrailingBits___180_comb;
  wire [8:0] p2_smul_57330_TrailingBits___183_comb;
  wire [8:0] p2_smul_57330_TrailingBits___1_comb;
  wire [8:0] p2_smul_57330_TrailingBits___2_comb;
  wire [8:0] p2_smul_57330_TrailingBits___5_comb;
  wire [8:0] p2_smul_57330_TrailingBits___6_comb;
  wire [8:0] p2_smul_57330_TrailingBits___25_comb;
  wire [8:0] p2_smul_57330_TrailingBits___26_comb;
  wire [8:0] p2_smul_57330_TrailingBits___29_comb;
  wire [8:0] p2_smul_57330_TrailingBits___30_comb;
  wire [8:0] p2_smul_57330_TrailingBits___64_comb;
  wire [8:0] p2_smul_57330_TrailingBits___67_comb;
  wire [8:0] p2_smul_57330_TrailingBits___68_comb;
  wire [8:0] p2_smul_57330_TrailingBits___71_comb;
  wire [8:0] p2_smul_57330_TrailingBits___88_comb;
  wire [8:0] p2_smul_57330_TrailingBits___91_comb;
  wire [8:0] p2_smul_57330_TrailingBits___92_comb;
  wire [8:0] p2_smul_57330_TrailingBits___95_comb;
  wire [8:0] p2_smul_57330_TrailingBits___97_comb;
  wire [8:0] p2_smul_57330_TrailingBits___98_comb;
  wire [8:0] p2_smul_57330_TrailingBits___101_comb;
  wire [8:0] p2_smul_57330_TrailingBits___102_comb;
  wire [8:0] p2_smul_57330_TrailingBits___121_comb;
  wire [8:0] p2_smul_57330_TrailingBits___122_comb;
  wire [8:0] p2_smul_57330_TrailingBits___125_comb;
  wire [8:0] p2_smul_57330_TrailingBits___126_comb;
  wire [8:0] p2_smul_57330_TrailingBits___160_comb;
  wire [8:0] p2_smul_57330_TrailingBits___163_comb;
  wire [8:0] p2_smul_57330_TrailingBits___164_comb;
  wire [8:0] p2_smul_57330_TrailingBits___167_comb;
  wire [8:0] p2_smul_57330_TrailingBits___184_comb;
  wire [8:0] p2_smul_57330_TrailingBits___187_comb;
  wire [8:0] p2_smul_57330_TrailingBits___188_comb;
  wire [8:0] p2_smul_57330_TrailingBits___191_comb;
  wire [31:0] p2_prod__135_comb;
  wire [22:0] p2_concat_136661_comb;
  wire [22:0] p2_concat_136662_comb;
  wire [31:0] p2_prod__150_comb;
  wire [31:0] p2_prod__327_comb;
  wire [22:0] p2_concat_136667_comb;
  wire [22:0] p2_concat_136668_comb;
  wire [31:0] p2_prod__342_comb;
  wire [31:0] p2_prod__133_comb;
  wire [31:0] p2_prod__136_comb;
  wire [31:0] p2_prod__140_comb;
  wire [31:0] p2_prod__145_comb;
  wire [31:0] p2_prod__151_comb;
  wire [31:0] p2_prod__158_comb;
  wire [31:0] p2_prod__165_comb;
  wire [31:0] p2_prod__171_comb;
  wire [31:0] p2_prod__325_comb;
  wire [31:0] p2_prod__328_comb;
  wire [31:0] p2_prod__332_comb;
  wire [31:0] p2_prod__337_comb;
  wire [31:0] p2_prod__343_comb;
  wire [31:0] p2_prod__350_comb;
  wire [31:0] p2_prod__357_comb;
  wire [31:0] p2_prod__363_comb;
  wire [22:0] p2_concat_136695_comb;
  wire [31:0] p2_prod__152_comb;
  wire [31:0] p2_prod__159_comb;
  wire [22:0] p2_concat_136700_comb;
  wire [22:0] p2_concat_136701_comb;
  wire [31:0] p2_prod__344_comb;
  wire [31:0] p2_prod__351_comb;
  wire [22:0] p2_concat_136706_comb;
  wire [31:0] p2_prod__148_comb;
  wire [22:0] p2_concat_136709_comb;
  wire [22:0] p2_concat_136710_comb;
  wire [31:0] p2_prod__186_comb;
  wire [31:0] p2_prod__340_comb;
  wire [22:0] p2_concat_136715_comb;
  wire [22:0] p2_concat_136716_comb;
  wire [31:0] p2_prod__378_comb;
  wire [31:0] p2_prod__155_comb;
  wire [31:0] p2_prod__162_comb;
  wire [31:0] p2_prod__169_comb;
  wire [31:0] p2_prod__175_comb;
  wire [31:0] p2_prod__180_comb;
  wire [31:0] p2_prod__184_comb;
  wire [31:0] p2_prod__187_comb;
  wire [31:0] p2_prod__189_comb;
  wire [31:0] p2_prod__347_comb;
  wire [31:0] p2_prod__354_comb;
  wire [31:0] p2_prod__361_comb;
  wire [31:0] p2_prod__367_comb;
  wire [31:0] p2_prod__372_comb;
  wire [31:0] p2_prod__376_comb;
  wire [31:0] p2_prod__379_comb;
  wire [31:0] p2_prod__381_comb;
  wire [22:0] p2_concat_136743_comb;
  wire [31:0] p2_prod__170_comb;
  wire [31:0] p2_prod__190_comb;
  wire [22:0] p2_concat_136748_comb;
  wire [22:0] p2_concat_136749_comb;
  wire [31:0] p2_prod__362_comb;
  wire [31:0] p2_prod__382_comb;
  wire [22:0] p2_concat_136754_comb;
  wire [31:0] p2_prod__10_comb;
  wire [22:0] p2_concat_136805_comb;
  wire [22:0] p2_concat_136806_comb;
  wire [31:0] p2_prod__13_comb;
  wire [31:0] p2_prod__71_comb;
  wire [22:0] p2_concat_136811_comb;
  wire [22:0] p2_concat_136812_comb;
  wire [31:0] p2_prod__86_comb;
  wire [31:0] p2_prod__391_comb;
  wire [22:0] p2_concat_136821_comb;
  wire [22:0] p2_concat_136822_comb;
  wire [31:0] p2_prod__406_comb;
  wire [31:0] p2_prod__455_comb;
  wire [22:0] p2_concat_136827_comb;
  wire [22:0] p2_concat_136828_comb;
  wire [31:0] p2_prod__470_comb;
  wire [31:0] p2_prod__16_comb;
  wire [31:0] p2_prod__17_comb;
  wire [31:0] p2_prod__18_comb;
  wire [31:0] p2_prod__19_comb;
  wire [31:0] p2_prod__20_comb;
  wire [31:0] p2_prod__21_comb;
  wire [31:0] p2_prod__22_comb;
  wire [31:0] p2_prod__23_comb;
  wire [31:0] p2_prod__69_comb;
  wire [31:0] p2_prod__72_comb;
  wire [31:0] p2_prod__76_comb;
  wire [31:0] p2_prod__81_comb;
  wire [31:0] p2_prod__87_comb;
  wire [31:0] p2_prod__94_comb;
  wire [31:0] p2_prod__101_comb;
  wire [31:0] p2_prod__107_comb;
  wire [31:0] p2_prod__197_comb;
  wire [31:0] p2_prod__200_comb;
  wire [31:0] p2_prod__204_comb;
  wire [31:0] p2_prod__209_comb;
  wire [31:0] p2_prod__215_comb;
  wire [31:0] p2_prod__222_comb;
  wire [31:0] p2_prod__229_comb;
  wire [31:0] p2_prod__235_comb;
  wire [31:0] p2_prod__261_comb;
  wire [31:0] p2_prod__264_comb;
  wire [31:0] p2_prod__268_comb;
  wire [31:0] p2_prod__273_comb;
  wire [31:0] p2_prod__279_comb;
  wire [31:0] p2_prod__286_comb;
  wire [31:0] p2_prod__293_comb;
  wire [31:0] p2_prod__299_comb;
  wire [31:0] p2_prod__389_comb;
  wire [31:0] p2_prod__392_comb;
  wire [31:0] p2_prod__396_comb;
  wire [31:0] p2_prod__401_comb;
  wire [31:0] p2_prod__407_comb;
  wire [31:0] p2_prod__414_comb;
  wire [31:0] p2_prod__421_comb;
  wire [31:0] p2_prod__427_comb;
  wire [31:0] p2_prod__453_comb;
  wire [31:0] p2_prod__456_comb;
  wire [31:0] p2_prod__460_comb;
  wire [31:0] p2_prod__465_comb;
  wire [31:0] p2_prod__471_comb;
  wire [31:0] p2_prod__478_comb;
  wire [31:0] p2_prod__485_comb;
  wire [31:0] p2_prod__491_comb;
  wire [22:0] p2_concat_136903_comb;
  wire [31:0] p2_prod__27_comb;
  wire [31:0] p2_prod__28_comb;
  wire [22:0] p2_concat_136908_comb;
  wire [22:0] p2_concat_136909_comb;
  wire [31:0] p2_prod__88_comb;
  wire [31:0] p2_prod__95_comb;
  wire [22:0] p2_concat_136914_comb;
  wire [22:0] p2_concat_136919_comb;
  wire [31:0] p2_prod__408_comb;
  wire [31:0] p2_prod__415_comb;
  wire [22:0] p2_concat_136924_comb;
  wire [22:0] p2_concat_136925_comb;
  wire [31:0] p2_prod__472_comb;
  wire [31:0] p2_prod__479_comb;
  wire [22:0] p2_concat_136930_comb;
  wire [31:0] p2_prod__40_comb;
  wire [22:0] p2_concat_136933_comb;
  wire [22:0] p2_concat_136934_comb;
  wire [31:0] p2_prod__47_comb;
  wire [31:0] p2_prod__84_comb;
  wire [22:0] p2_concat_136939_comb;
  wire [22:0] p2_concat_136940_comb;
  wire [31:0] p2_prod__122_comb;
  wire [31:0] p2_prod__404_comb;
  wire [22:0] p2_concat_136949_comb;
  wire [22:0] p2_concat_136950_comb;
  wire [31:0] p2_prod__442_comb;
  wire [31:0] p2_prod__468_comb;
  wire [22:0] p2_concat_136955_comb;
  wire [22:0] p2_concat_136956_comb;
  wire [31:0] p2_prod__506_comb;
  wire [31:0] p2_prod__48_comb;
  wire [31:0] p2_prod__49_comb;
  wire [31:0] p2_prod__50_comb;
  wire [31:0] p2_prod__51_comb;
  wire [31:0] p2_prod__52_comb;
  wire [31:0] p2_prod__53_comb;
  wire [31:0] p2_prod__54_comb;
  wire [31:0] p2_prod__55_comb;
  wire [31:0] p2_prod__91_comb;
  wire [31:0] p2_prod__98_comb;
  wire [31:0] p2_prod__105_comb;
  wire [31:0] p2_prod__111_comb;
  wire [31:0] p2_prod__116_comb;
  wire [31:0] p2_prod__120_comb;
  wire [31:0] p2_prod__123_comb;
  wire [31:0] p2_prod__125_comb;
  wire [31:0] p2_prod__219_comb;
  wire [31:0] p2_prod__226_comb;
  wire [31:0] p2_prod__233_comb;
  wire [31:0] p2_prod__239_comb;
  wire [31:0] p2_prod__244_comb;
  wire [31:0] p2_prod__248_comb;
  wire [31:0] p2_prod__251_comb;
  wire [31:0] p2_prod__253_comb;
  wire [31:0] p2_prod__283_comb;
  wire [31:0] p2_prod__290_comb;
  wire [31:0] p2_prod__297_comb;
  wire [31:0] p2_prod__303_comb;
  wire [31:0] p2_prod__308_comb;
  wire [31:0] p2_prod__312_comb;
  wire [31:0] p2_prod__315_comb;
  wire [31:0] p2_prod__317_comb;
  wire [31:0] p2_prod__411_comb;
  wire [31:0] p2_prod__418_comb;
  wire [31:0] p2_prod__425_comb;
  wire [31:0] p2_prod__431_comb;
  wire [31:0] p2_prod__436_comb;
  wire [31:0] p2_prod__440_comb;
  wire [31:0] p2_prod__443_comb;
  wire [31:0] p2_prod__445_comb;
  wire [31:0] p2_prod__475_comb;
  wire [31:0] p2_prod__482_comb;
  wire [31:0] p2_prod__489_comb;
  wire [31:0] p2_prod__495_comb;
  wire [31:0] p2_prod__500_comb;
  wire [31:0] p2_prod__504_comb;
  wire [31:0] p2_prod__507_comb;
  wire [31:0] p2_prod__509_comb;
  wire [22:0] p2_concat_137031_comb;
  wire [31:0] p2_prod__57_comb;
  wire [31:0] p2_prod__62_comb;
  wire [22:0] p2_concat_137036_comb;
  wire [22:0] p2_concat_137037_comb;
  wire [31:0] p2_prod__106_comb;
  wire [31:0] p2_prod__126_comb;
  wire [22:0] p2_concat_137042_comb;
  wire [22:0] p2_concat_137047_comb;
  wire [31:0] p2_prod__426_comb;
  wire [31:0] p2_prod__446_comb;
  wire [22:0] p2_concat_137052_comb;
  wire [22:0] p2_concat_137053_comb;
  wire [31:0] p2_prod__490_comb;
  wire [31:0] p2_prod__510_comb;
  wire [22:0] p2_concat_137058_comb;
  wire [7:0] p2_smul_57326_TrailingBits___16_comb;
  wire [7:0] p2_smul_57326_TrailingBits___17_comb;
  wire [7:0] p2_smul_57326_TrailingBits___18_comb;
  wire [7:0] p2_smul_57326_TrailingBits___19_comb;
  wire [7:0] p2_smul_57326_TrailingBits___20_comb;
  wire [7:0] p2_smul_57326_TrailingBits___21_comb;
  wire [7:0] p2_smul_57326_TrailingBits___22_comb;
  wire [7:0] p2_smul_57326_TrailingBits___23_comb;
  wire [7:0] p2_smul_57326_TrailingBits___40_comb;
  wire [7:0] p2_smul_57326_TrailingBits___41_comb;
  wire [7:0] p2_smul_57326_TrailingBits___42_comb;
  wire [7:0] p2_smul_57326_TrailingBits___43_comb;
  wire [7:0] p2_smul_57326_TrailingBits___44_comb;
  wire [7:0] p2_smul_57326_TrailingBits___45_comb;
  wire [7:0] p2_smul_57326_TrailingBits___46_comb;
  wire [7:0] p2_smul_57326_TrailingBits___47_comb;
  wire [7:0] p2_smul_57326_TrailingBits__comb;
  wire [7:0] p2_smul_57326_TrailingBits___1_comb;
  wire [7:0] p2_smul_57326_TrailingBits___2_comb;
  wire [7:0] p2_smul_57326_TrailingBits___3_comb;
  wire [7:0] p2_smul_57326_TrailingBits___4_comb;
  wire [7:0] p2_smul_57326_TrailingBits___5_comb;
  wire [7:0] p2_smul_57326_TrailingBits___6_comb;
  wire [7:0] p2_smul_57326_TrailingBits___7_comb;
  wire [7:0] p2_smul_57326_TrailingBits___8_comb;
  wire [7:0] p2_smul_57326_TrailingBits___9_comb;
  wire [7:0] p2_smul_57326_TrailingBits___10_comb;
  wire [7:0] p2_smul_57326_TrailingBits___11_comb;
  wire [7:0] p2_smul_57326_TrailingBits___12_comb;
  wire [7:0] p2_smul_57326_TrailingBits___13_comb;
  wire [7:0] p2_smul_57326_TrailingBits___14_comb;
  wire [7:0] p2_smul_57326_TrailingBits___15_comb;
  wire [7:0] p2_smul_57326_TrailingBits___24_comb;
  wire [7:0] p2_smul_57326_TrailingBits___25_comb;
  wire [7:0] p2_smul_57326_TrailingBits___26_comb;
  wire [7:0] p2_smul_57326_TrailingBits___27_comb;
  wire [7:0] p2_smul_57326_TrailingBits___28_comb;
  wire [7:0] p2_smul_57326_TrailingBits___29_comb;
  wire [7:0] p2_smul_57326_TrailingBits___30_comb;
  wire [7:0] p2_smul_57326_TrailingBits___31_comb;
  wire [7:0] p2_smul_57326_TrailingBits___32_comb;
  wire [7:0] p2_smul_57326_TrailingBits___33_comb;
  wire [7:0] p2_smul_57326_TrailingBits___34_comb;
  wire [7:0] p2_smul_57326_TrailingBits___35_comb;
  wire [7:0] p2_smul_57326_TrailingBits___36_comb;
  wire [7:0] p2_smul_57326_TrailingBits___37_comb;
  wire [7:0] p2_smul_57326_TrailingBits___38_comb;
  wire [7:0] p2_smul_57326_TrailingBits___39_comb;
  wire [7:0] p2_smul_57326_TrailingBits___48_comb;
  wire [7:0] p2_smul_57326_TrailingBits___49_comb;
  wire [7:0] p2_smul_57326_TrailingBits___50_comb;
  wire [7:0] p2_smul_57326_TrailingBits___51_comb;
  wire [7:0] p2_smul_57326_TrailingBits___52_comb;
  wire [7:0] p2_smul_57326_TrailingBits___53_comb;
  wire [7:0] p2_smul_57326_TrailingBits___54_comb;
  wire [7:0] p2_smul_57326_TrailingBits___55_comb;
  wire [7:0] p2_smul_57326_TrailingBits___56_comb;
  wire [7:0] p2_smul_57326_TrailingBits___57_comb;
  wire [7:0] p2_smul_57326_TrailingBits___58_comb;
  wire [7:0] p2_smul_57326_TrailingBits___59_comb;
  wire [7:0] p2_smul_57326_TrailingBits___60_comb;
  wire [7:0] p2_smul_57326_TrailingBits___61_comb;
  wire [7:0] p2_smul_57326_TrailingBits___62_comb;
  wire [7:0] p2_smul_57326_TrailingBits___63_comb;
  wire [31:0] p2_or_137427_comb;
  wire [31:0] p2_prod__203_comb;
  wire [31:0] p2_prod__208_comb;
  wire [31:0] p2_or_137434_comb;
  wire [31:0] p2_or_137441_comb;
  wire [31:0] p2_prod__267_comb;
  wire [31:0] p2_prod__272_comb;
  wire [31:0] p2_or_137448_comb;
  wire [31:0] p2_prod__205_comb;
  wire [31:0] p2_or_137633_comb;
  wire [31:0] p2_or_137636_comb;
  wire [31:0] p2_prod__236_comb;
  wire [31:0] p2_prod__269_comb;
  wire [31:0] p2_or_137647_comb;
  wire [31:0] p2_or_137650_comb;
  wire [31:0] p2_prod__300_comb;
  wire [31:0] p2_or_137761_comb;
  wire [31:0] p2_prod__225_comb;
  wire [31:0] p2_prod__243_comb;
  wire [31:0] p2_or_137772_comb;
  wire [31:0] p2_or_137775_comb;
  wire [31:0] p2_prod__289_comb;
  wire [31:0] p2_prod__307_comb;
  wire [31:0] p2_or_137786_comb;
  wire [31:0] p2_prod__227_comb;
  wire [31:0] p2_or_137967_comb;
  wire [31:0] p2_or_137974_comb;
  wire [31:0] p2_prod__255_comb;
  wire [31:0] p2_prod__291_comb;
  wire [31:0] p2_or_137981_comb;
  wire [31:0] p2_or_137988_comb;
  wire [31:0] p2_prod__319_comb;
  wire [16:0] p2_smul_57742_NarrowedMult__comb;
  wire [16:0] p2_smul_57744_NarrowedMult__comb;
  wire [16:0] p2_smul_57746_NarrowedMult__comb;
  wire [16:0] p2_smul_57748_NarrowedMult__comb;
  wire [16:0] p2_smul_57750_NarrowedMult__comb;
  wire [16:0] p2_smul_57752_NarrowedMult__comb;
  wire [16:0] p2_smul_57754_NarrowedMult__comb;
  wire [16:0] p2_smul_57756_NarrowedMult__comb;
  wire [16:0] p2_smul_57790_NarrowedMult__comb;
  wire [16:0] p2_smul_57792_NarrowedMult__comb;
  wire [16:0] p2_smul_57794_NarrowedMult__comb;
  wire [16:0] p2_smul_57796_NarrowedMult__comb;
  wire [16:0] p2_smul_57798_NarrowedMult__comb;
  wire [16:0] p2_smul_57800_NarrowedMult__comb;
  wire [16:0] p2_smul_57802_NarrowedMult__comb;
  wire [16:0] p2_smul_57804_NarrowedMult__comb;
  wire [16:0] p2_smul_57710_NarrowedMult__comb;
  wire [16:0] p2_smul_57712_NarrowedMult__comb;
  wire [16:0] p2_smul_57714_NarrowedMult__comb;
  wire [16:0] p2_smul_57716_NarrowedMult__comb;
  wire [16:0] p2_smul_57718_NarrowedMult__comb;
  wire [16:0] p2_smul_57720_NarrowedMult__comb;
  wire [16:0] p2_smul_57722_NarrowedMult__comb;
  wire [16:0] p2_smul_57724_NarrowedMult__comb;
  wire [16:0] p2_smul_57726_NarrowedMult__comb;
  wire [16:0] p2_smul_57728_NarrowedMult__comb;
  wire [16:0] p2_smul_57730_NarrowedMult__comb;
  wire [16:0] p2_smul_57732_NarrowedMult__comb;
  wire [16:0] p2_smul_57734_NarrowedMult__comb;
  wire [16:0] p2_smul_57736_NarrowedMult__comb;
  wire [16:0] p2_smul_57738_NarrowedMult__comb;
  wire [16:0] p2_smul_57740_NarrowedMult__comb;
  wire [16:0] p2_smul_57758_NarrowedMult__comb;
  wire [16:0] p2_smul_57760_NarrowedMult__comb;
  wire [16:0] p2_smul_57762_NarrowedMult__comb;
  wire [16:0] p2_smul_57764_NarrowedMult__comb;
  wire [16:0] p2_smul_57766_NarrowedMult__comb;
  wire [16:0] p2_smul_57768_NarrowedMult__comb;
  wire [16:0] p2_smul_57770_NarrowedMult__comb;
  wire [16:0] p2_smul_57772_NarrowedMult__comb;
  wire [16:0] p2_smul_57774_NarrowedMult__comb;
  wire [16:0] p2_smul_57776_NarrowedMult__comb;
  wire [16:0] p2_smul_57778_NarrowedMult__comb;
  wire [16:0] p2_smul_57780_NarrowedMult__comb;
  wire [16:0] p2_smul_57782_NarrowedMult__comb;
  wire [16:0] p2_smul_57784_NarrowedMult__comb;
  wire [16:0] p2_smul_57786_NarrowedMult__comb;
  wire [16:0] p2_smul_57788_NarrowedMult__comb;
  wire [16:0] p2_smul_57806_NarrowedMult__comb;
  wire [16:0] p2_smul_57808_NarrowedMult__comb;
  wire [16:0] p2_smul_57810_NarrowedMult__comb;
  wire [16:0] p2_smul_57812_NarrowedMult__comb;
  wire [16:0] p2_smul_57814_NarrowedMult__comb;
  wire [16:0] p2_smul_57816_NarrowedMult__comb;
  wire [16:0] p2_smul_57818_NarrowedMult__comb;
  wire [16:0] p2_smul_57820_NarrowedMult__comb;
  wire [16:0] p2_smul_57822_NarrowedMult__comb;
  wire [16:0] p2_smul_57824_NarrowedMult__comb;
  wire [16:0] p2_smul_57826_NarrowedMult__comb;
  wire [16:0] p2_smul_57828_NarrowedMult__comb;
  wire [16:0] p2_smul_57830_NarrowedMult__comb;
  wire [16:0] p2_smul_57832_NarrowedMult__comb;
  wire [16:0] p2_smul_57834_NarrowedMult__comb;
  wire [16:0] p2_smul_57836_NarrowedMult__comb;
  wire [31:0] p2_or_137095_comb;
  wire [31:0] p2_prod__139_comb;
  wire [31:0] p2_prod__144_comb;
  wire [31:0] p2_or_137102_comb;
  wire [31:0] p2_or_137109_comb;
  wire [31:0] p2_prod__331_comb;
  wire [31:0] p2_prod__336_comb;
  wire [31:0] p2_or_137116_comb;
  wire [31:0] p2_or_137121_comb;
  wire [31:0] p2_or_137128_comb;
  wire [31:0] p2_or_137131_comb;
  wire [31:0] p2_or_137138_comb;
  wire [31:0] p2_or_137141_comb;
  wire [31:0] p2_or_137148_comb;
  wire [31:0] p2_or_137151_comb;
  wire [31:0] p2_or_137158_comb;
  wire [31:0] p2_prod__141_comb;
  wire [31:0] p2_or_137165_comb;
  wire [31:0] p2_or_137168_comb;
  wire [31:0] p2_prod__172_comb;
  wire [31:0] p2_prod__333_comb;
  wire [31:0] p2_or_137179_comb;
  wire [31:0] p2_or_137182_comb;
  wire [31:0] p2_prod__364_comb;
  wire [31:0] p2_or_137205_comb;
  wire [31:0] p2_prod__161_comb;
  wire [31:0] p2_prod__179_comb;
  wire [31:0] p2_or_137216_comb;
  wire [31:0] p2_or_137219_comb;
  wire [31:0] p2_prod__353_comb;
  wire [31:0] p2_prod__371_comb;
  wire [31:0] p2_or_137230_comb;
  wire [31:0] p2_or_137235_comb;
  wire [31:0] p2_or_137240_comb;
  wire [31:0] p2_or_137243_comb;
  wire [31:0] p2_or_137248_comb;
  wire [31:0] p2_or_137255_comb;
  wire [31:0] p2_or_137260_comb;
  wire [31:0] p2_or_137263_comb;
  wire [31:0] p2_or_137268_comb;
  wire [31:0] p2_prod__163_comb;
  wire [31:0] p2_or_137275_comb;
  wire [31:0] p2_or_137282_comb;
  wire [31:0] p2_prod__191_comb;
  wire [31:0] p2_prod__355_comb;
  wire [31:0] p2_or_137289_comb;
  wire [31:0] p2_or_137296_comb;
  wire [31:0] p2_prod__383_comb;
  wire [31:0] p2_or_137399_comb;
  wire [31:0] p2_prod__11_comb;
  wire [31:0] p2_prod__12_comb;
  wire [31:0] p2_or_137406_comb;
  wire [31:0] p2_or_137413_comb;
  wire [31:0] p2_prod__75_comb;
  wire [31:0] p2_prod__80_comb;
  wire [31:0] p2_or_137420_comb;
  wire [31:0] p2_or_137455_comb;
  wire [31:0] p2_prod__395_comb;
  wire [31:0] p2_prod__400_comb;
  wire [31:0] p2_or_137462_comb;
  wire [31:0] p2_or_137469_comb;
  wire [31:0] p2_prod__459_comb;
  wire [31:0] p2_prod__464_comb;
  wire [31:0] p2_or_137476_comb;
  wire [31:0] p2_or_137481_comb;
  wire [31:0] p2_or_137488_comb;
  wire [31:0] p2_or_137491_comb;
  wire [31:0] p2_or_137498_comb;
  wire [31:0] p2_or_137501_comb;
  wire [31:0] p2_or_137508_comb;
  wire [31:0] p2_or_137511_comb;
  wire [31:0] p2_or_137518_comb;
  wire [31:0] p2_or_137521_comb;
  wire [31:0] p2_or_137528_comb;
  wire [31:0] p2_or_137531_comb;
  wire [31:0] p2_or_137538_comb;
  wire [31:0] p2_or_137541_comb;
  wire [31:0] p2_or_137548_comb;
  wire [31:0] p2_or_137551_comb;
  wire [31:0] p2_or_137558_comb;
  wire [31:0] p2_or_137561_comb;
  wire [31:0] p2_or_137568_comb;
  wire [31:0] p2_or_137571_comb;
  wire [31:0] p2_or_137578_comb;
  wire [31:0] p2_or_137581_comb;
  wire [31:0] p2_or_137588_comb;
  wire [31:0] p2_or_137591_comb;
  wire [31:0] p2_or_137598_comb;
  wire [31:0] p2_prod__25_comb;
  wire [31:0] p2_or_137605_comb;
  wire [31:0] p2_or_137608_comb;
  wire [31:0] p2_prod__30_comb;
  wire [31:0] p2_prod__77_comb;
  wire [31:0] p2_or_137619_comb;
  wire [31:0] p2_or_137622_comb;
  wire [31:0] p2_prod__108_comb;
  wire [31:0] p2_prod__397_comb;
  wire [31:0] p2_or_137661_comb;
  wire [31:0] p2_or_137664_comb;
  wire [31:0] p2_prod__428_comb;
  wire [31:0] p2_prod__461_comb;
  wire [31:0] p2_or_137675_comb;
  wire [31:0] p2_or_137678_comb;
  wire [31:0] p2_prod__492_comb;
  wire [31:0] p2_or_137733_comb;
  wire [31:0] p2_prod__42_comb;
  wire [31:0] p2_prod__45_comb;
  wire [31:0] p2_or_137744_comb;
  wire [31:0] p2_or_137747_comb;
  wire [31:0] p2_prod__97_comb;
  wire [31:0] p2_prod__115_comb;
  wire [31:0] p2_or_137758_comb;
  wire [31:0] p2_or_137789_comb;
  wire [31:0] p2_prod__417_comb;
  wire [31:0] p2_prod__435_comb;
  wire [31:0] p2_or_137800_comb;
  wire [31:0] p2_or_137803_comb;
  wire [31:0] p2_prod__481_comb;
  wire [31:0] p2_prod__499_comb;
  wire [31:0] p2_or_137814_comb;
  wire [31:0] p2_or_137819_comb;
  wire [31:0] p2_or_137824_comb;
  wire [31:0] p2_or_137827_comb;
  wire [31:0] p2_or_137832_comb;
  wire [31:0] p2_or_137839_comb;
  wire [31:0] p2_or_137844_comb;
  wire [31:0] p2_or_137847_comb;
  wire [31:0] p2_or_137852_comb;
  wire [31:0] p2_or_137859_comb;
  wire [31:0] p2_or_137864_comb;
  wire [31:0] p2_or_137867_comb;
  wire [31:0] p2_or_137872_comb;
  wire [31:0] p2_or_137879_comb;
  wire [31:0] p2_or_137884_comb;
  wire [31:0] p2_or_137887_comb;
  wire [31:0] p2_or_137892_comb;
  wire [31:0] p2_or_137899_comb;
  wire [31:0] p2_or_137904_comb;
  wire [31:0] p2_or_137907_comb;
  wire [31:0] p2_or_137912_comb;
  wire [31:0] p2_or_137919_comb;
  wire [31:0] p2_or_137924_comb;
  wire [31:0] p2_or_137927_comb;
  wire [31:0] p2_or_137932_comb;
  wire [31:0] p2_prod__56_comb;
  wire [31:0] p2_or_137939_comb;
  wire [31:0] p2_or_137946_comb;
  wire [31:0] p2_prod__63_comb;
  wire [31:0] p2_prod__99_comb;
  wire [31:0] p2_or_137953_comb;
  wire [31:0] p2_or_137960_comb;
  wire [31:0] p2_prod__127_comb;
  wire [31:0] p2_prod__419_comb;
  wire [31:0] p2_or_137995_comb;
  wire [31:0] p2_or_138002_comb;
  wire [31:0] p2_prod__447_comb;
  wire [31:0] p2_prod__483_comb;
  wire [31:0] p2_or_138009_comb;
  wire [31:0] p2_or_138016_comb;
  wire [31:0] p2_prod__511_comb;
  wire [16:0] p2_smul_57374_NarrowedMult__comb;
  wire [16:0] p2_smul_57376_NarrowedMult__comb;
  wire [31:0] p2_or_138426_comb;
  wire [31:0] p2_or_138427_comb;
  wire [16:0] p2_smul_57386_NarrowedMult__comb;
  wire [16:0] p2_smul_57388_NarrowedMult__comb;
  wire [16:0] p2_smul_57390_NarrowedMult__comb;
  wire [16:0] p2_smul_57392_NarrowedMult__comb;
  wire [31:0] p2_or_138442_comb;
  wire [31:0] p2_or_138443_comb;
  wire [16:0] p2_smul_57402_NarrowedMult__comb;
  wire [16:0] p2_smul_57404_NarrowedMult__comb;
  wire [16:0] p2_smul_57630_NarrowedMult__comb;
  wire [31:0] p2_or_138637_comb;
  wire [16:0] p2_smul_57634_NarrowedMult__comb;
  wire [16:0] p2_smul_57640_NarrowedMult__comb;
  wire [31:0] p2_or_138648_comb;
  wire [16:0] p2_smul_57644_NarrowedMult__comb;
  wire [16:0] p2_smul_57646_NarrowedMult__comb;
  wire [31:0] p2_or_138653_comb;
  wire [16:0] p2_smul_57650_NarrowedMult__comb;
  wire [16:0] p2_smul_57656_NarrowedMult__comb;
  wire [31:0] p2_or_138664_comb;
  wire [16:0] p2_smul_57660_NarrowedMult__comb;
  wire [16:0] p2_smul_57888_NarrowedMult__comb;
  wire [31:0] p2_or_138832_comb;
  wire [16:0] p2_smul_57892_NarrowedMult__comb;
  wire [16:0] p2_smul_57894_NarrowedMult__comb;
  wire [31:0] p2_or_138837_comb;
  wire [16:0] p2_smul_57898_NarrowedMult__comb;
  wire [16:0] p2_smul_57904_NarrowedMult__comb;
  wire [31:0] p2_or_138848_comb;
  wire [16:0] p2_smul_57908_NarrowedMult__comb;
  wire [16:0] p2_smul_57910_NarrowedMult__comb;
  wire [31:0] p2_or_138853_comb;
  wire [16:0] p2_smul_57914_NarrowedMult__comb;
  wire [31:0] p2_or_139043_comb;
  wire [16:0] p2_smul_58146_NarrowedMult__comb;
  wire [16:0] p2_smul_58148_NarrowedMult__comb;
  wire [16:0] p2_smul_58150_NarrowedMult__comb;
  wire [16:0] p2_smul_58152_NarrowedMult__comb;
  wire [31:0] p2_or_139058_comb;
  wire [31:0] p2_or_139059_comb;
  wire [16:0] p2_smul_58162_NarrowedMult__comb;
  wire [16:0] p2_smul_58164_NarrowedMult__comb;
  wire [16:0] p2_smul_58166_NarrowedMult__comb;
  wire [16:0] p2_smul_58168_NarrowedMult__comb;
  wire [31:0] p2_or_139074_comb;
  wire [16:0] p2_smul_57358_NarrowedMult__comb;
  wire [16:0] p2_smul_57360_NarrowedMult__comb;
  wire [31:0] p2_or_138058_comb;
  wire [31:0] p2_or_138059_comb;
  wire [16:0] p2_smul_57370_NarrowedMult__comb;
  wire [16:0] p2_smul_57372_NarrowedMult__comb;
  wire [16:0] p2_smul_57406_NarrowedMult__comb;
  wire [16:0] p2_smul_57408_NarrowedMult__comb;
  wire [31:0] p2_or_138074_comb;
  wire [31:0] p2_or_138075_comb;
  wire [16:0] p2_smul_57418_NarrowedMult__comb;
  wire [16:0] p2_smul_57420_NarrowedMult__comb;
  wire [16:0] p2_smul_57614_NarrowedMult__comb;
  wire [31:0] p2_or_138125_comb;
  wire [16:0] p2_smul_57618_NarrowedMult__comb;
  wire [16:0] p2_smul_57624_NarrowedMult__comb;
  wire [31:0] p2_or_138136_comb;
  wire [16:0] p2_smul_57628_NarrowedMult__comb;
  wire [16:0] p2_smul_57662_NarrowedMult__comb;
  wire [31:0] p2_or_138141_comb;
  wire [16:0] p2_smul_57666_NarrowedMult__comb;
  wire [16:0] p2_smul_57672_NarrowedMult__comb;
  wire [31:0] p2_or_138152_comb;
  wire [16:0] p2_smul_57676_NarrowedMult__comb;
  wire [16:0] p2_smul_57872_NarrowedMult__comb;
  wire [31:0] p2_or_138192_comb;
  wire [16:0] p2_smul_57876_NarrowedMult__comb;
  wire [16:0] p2_smul_57878_NarrowedMult__comb;
  wire [31:0] p2_or_138197_comb;
  wire [16:0] p2_smul_57882_NarrowedMult__comb;
  wire [16:0] p2_smul_57920_NarrowedMult__comb;
  wire [31:0] p2_or_138208_comb;
  wire [16:0] p2_smul_57924_NarrowedMult__comb;
  wire [16:0] p2_smul_57926_NarrowedMult__comb;
  wire [31:0] p2_or_138213_comb;
  wire [16:0] p2_smul_57930_NarrowedMult__comb;
  wire [31:0] p2_or_138259_comb;
  wire [16:0] p2_smul_58130_NarrowedMult__comb;
  wire [16:0] p2_smul_58132_NarrowedMult__comb;
  wire [16:0] p2_smul_58134_NarrowedMult__comb;
  wire [16:0] p2_smul_58136_NarrowedMult__comb;
  wire [31:0] p2_or_138274_comb;
  wire [31:0] p2_or_138275_comb;
  wire [16:0] p2_smul_58178_NarrowedMult__comb;
  wire [16:0] p2_smul_58180_NarrowedMult__comb;
  wire [16:0] p2_smul_58182_NarrowedMult__comb;
  wire [16:0] p2_smul_58184_NarrowedMult__comb;
  wire [31:0] p2_or_138290_comb;
  wire [16:0] p2_smul_57326_NarrowedMult__comb;
  wire [16:0] p2_smul_57328_NarrowedMult__comb;
  wire [31:0] p2_or_138394_comb;
  wire [31:0] p2_or_138395_comb;
  wire [16:0] p2_smul_57338_NarrowedMult__comb;
  wire [16:0] p2_smul_57340_NarrowedMult__comb;
  wire [16:0] p2_smul_57342_NarrowedMult__comb;
  wire [16:0] p2_smul_57344_NarrowedMult__comb;
  wire [31:0] p2_or_138410_comb;
  wire [31:0] p2_or_138411_comb;
  wire [16:0] p2_smul_57354_NarrowedMult__comb;
  wire [16:0] p2_smul_57356_NarrowedMult__comb;
  wire [16:0] p2_smul_57422_NarrowedMult__comb;
  wire [16:0] p2_smul_57424_NarrowedMult__comb;
  wire [31:0] p2_or_138458_comb;
  wire [31:0] p2_or_138459_comb;
  wire [16:0] p2_smul_57434_NarrowedMult__comb;
  wire [16:0] p2_smul_57436_NarrowedMult__comb;
  wire [16:0] p2_smul_57438_NarrowedMult__comb;
  wire [16:0] p2_smul_57440_NarrowedMult__comb;
  wire [31:0] p2_or_138474_comb;
  wire [31:0] p2_or_138475_comb;
  wire [16:0] p2_smul_57450_NarrowedMult__comb;
  wire [16:0] p2_smul_57452_NarrowedMult__comb;
  wire [16:0] p2_smul_57582_NarrowedMult__comb;
  wire [31:0] p2_or_138605_comb;
  wire [16:0] p2_smul_57586_NarrowedMult__comb;
  wire [16:0] p2_smul_57592_NarrowedMult__comb;
  wire [31:0] p2_or_138616_comb;
  wire [16:0] p2_smul_57596_NarrowedMult__comb;
  wire [16:0] p2_smul_57598_NarrowedMult__comb;
  wire [31:0] p2_or_138621_comb;
  wire [16:0] p2_smul_57602_NarrowedMult__comb;
  wire [16:0] p2_smul_57608_NarrowedMult__comb;
  wire [31:0] p2_or_138632_comb;
  wire [16:0] p2_smul_57612_NarrowedMult__comb;
  wire [16:0] p2_smul_57678_NarrowedMult__comb;
  wire [31:0] p2_or_138669_comb;
  wire [16:0] p2_smul_57682_NarrowedMult__comb;
  wire [16:0] p2_smul_57688_NarrowedMult__comb;
  wire [31:0] p2_or_138680_comb;
  wire [16:0] p2_smul_57692_NarrowedMult__comb;
  wire [16:0] p2_smul_57694_NarrowedMult__comb;
  wire [31:0] p2_or_138685_comb;
  wire [16:0] p2_smul_57698_NarrowedMult__comb;
  wire [16:0] p2_smul_57704_NarrowedMult__comb;
  wire [31:0] p2_or_138696_comb;
  wire [16:0] p2_smul_57708_NarrowedMult__comb;
  wire [16:0] p2_smul_57840_NarrowedMult__comb;
  wire [31:0] p2_or_138800_comb;
  wire [16:0] p2_smul_57844_NarrowedMult__comb;
  wire [16:0] p2_smul_57846_NarrowedMult__comb;
  wire [31:0] p2_or_138805_comb;
  wire [16:0] p2_smul_57850_NarrowedMult__comb;
  wire [16:0] p2_smul_57856_NarrowedMult__comb;
  wire [31:0] p2_or_138816_comb;
  wire [16:0] p2_smul_57860_NarrowedMult__comb;
  wire [16:0] p2_smul_57862_NarrowedMult__comb;
  wire [31:0] p2_or_138821_comb;
  wire [16:0] p2_smul_57866_NarrowedMult__comb;
  wire [16:0] p2_smul_57936_NarrowedMult__comb;
  wire [31:0] p2_or_138864_comb;
  wire [16:0] p2_smul_57940_NarrowedMult__comb;
  wire [16:0] p2_smul_57942_NarrowedMult__comb;
  wire [31:0] p2_or_138869_comb;
  wire [16:0] p2_smul_57946_NarrowedMult__comb;
  wire [16:0] p2_smul_57952_NarrowedMult__comb;
  wire [31:0] p2_or_138880_comb;
  wire [16:0] p2_smul_57956_NarrowedMult__comb;
  wire [16:0] p2_smul_57958_NarrowedMult__comb;
  wire [31:0] p2_or_138885_comb;
  wire [16:0] p2_smul_57962_NarrowedMult__comb;
  wire [31:0] p2_or_139011_comb;
  wire [16:0] p2_smul_58098_NarrowedMult__comb;
  wire [16:0] p2_smul_58100_NarrowedMult__comb;
  wire [16:0] p2_smul_58102_NarrowedMult__comb;
  wire [16:0] p2_smul_58104_NarrowedMult__comb;
  wire [31:0] p2_or_139026_comb;
  wire [31:0] p2_or_139027_comb;
  wire [16:0] p2_smul_58114_NarrowedMult__comb;
  wire [16:0] p2_smul_58116_NarrowedMult__comb;
  wire [16:0] p2_smul_58118_NarrowedMult__comb;
  wire [16:0] p2_smul_58120_NarrowedMult__comb;
  wire [31:0] p2_or_139042_comb;
  wire [31:0] p2_or_139075_comb;
  wire [16:0] p2_smul_58194_NarrowedMult__comb;
  wire [16:0] p2_smul_58196_NarrowedMult__comb;
  wire [16:0] p2_smul_58198_NarrowedMult__comb;
  wire [16:0] p2_smul_58200_NarrowedMult__comb;
  wire [31:0] p2_or_139090_comb;
  wire [31:0] p2_or_139091_comb;
  wire [16:0] p2_smul_58210_NarrowedMult__comb;
  wire [16:0] p2_smul_58212_NarrowedMult__comb;
  wire [16:0] p2_smul_58214_NarrowedMult__comb;
  wire [16:0] p2_smul_58216_NarrowedMult__comb;
  wire [31:0] p2_or_139106_comb;
  wire [15:0] p2_sel_139107_comb;
  wire [15:0] p2_sel_139108_comb;
  wire [15:0] p2_sel_139109_comb;
  wire [15:0] p2_sel_139110_comb;
  wire [15:0] p2_sel_139111_comb;
  wire [15:0] p2_sel_139112_comb;
  wire [15:0] p2_sel_139113_comb;
  wire [15:0] p2_sel_139114_comb;
  wire [15:0] p2_sel_139115_comb;
  wire [15:0] p2_sel_139116_comb;
  wire [15:0] p2_sel_139117_comb;
  wire [15:0] p2_sel_139118_comb;
  wire [15:0] p2_sel_139119_comb;
  wire [15:0] p2_sel_139120_comb;
  wire [15:0] p2_sel_139121_comb;
  wire [15:0] p2_sel_139122_comb;
  wire [15:0] p2_sel_139571_comb;
  wire [15:0] p2_sel_139572_comb;
  wire [15:0] p2_sel_139573_comb;
  wire [15:0] p2_sel_139574_comb;
  wire [15:0] p2_sel_139575_comb;
  wire [15:0] p2_sel_139576_comb;
  wire [15:0] p2_sel_139577_comb;
  wire [15:0] p2_sel_139578_comb;
  wire [15:0] p2_sel_139579_comb;
  wire [15:0] p2_sel_139580_comb;
  wire [15:0] p2_sel_139581_comb;
  wire [15:0] p2_sel_139582_comb;
  wire [15:0] p2_sel_139583_comb;
  wire [15:0] p2_sel_139584_comb;
  wire [15:0] p2_sel_139585_comb;
  wire [15:0] p2_sel_139586_comb;
  wire [15:0] p2_sel_139587_comb;
  wire [15:0] p2_sel_139588_comb;
  wire [15:0] p2_sel_139589_comb;
  wire [15:0] p2_sel_139590_comb;
  wire [15:0] p2_sel_139591_comb;
  wire [15:0] p2_sel_139592_comb;
  wire [15:0] p2_sel_139593_comb;
  wire [15:0] p2_sel_139594_comb;
  wire [15:0] p2_sel_139595_comb;
  wire [15:0] p2_sel_139596_comb;
  wire [15:0] p2_sel_139597_comb;
  wire [15:0] p2_sel_139598_comb;
  wire [15:0] p2_sel_139599_comb;
  wire [15:0] p2_sel_139600_comb;
  wire [15:0] p2_sel_139601_comb;
  wire [15:0] p2_sel_139602_comb;
  wire [15:0] p2_sel_139603_comb;
  wire [15:0] p2_sel_139604_comb;
  wire [15:0] p2_sel_139605_comb;
  wire [15:0] p2_sel_139606_comb;
  wire [15:0] p2_sel_139607_comb;
  wire [15:0] p2_sel_139608_comb;
  wire [15:0] p2_sel_139609_comb;
  wire [15:0] p2_sel_139610_comb;
  wire [15:0] p2_sel_139611_comb;
  wire [15:0] p2_sel_139612_comb;
  wire [15:0] p2_sel_139613_comb;
  wire [15:0] p2_sel_139614_comb;
  wire [15:0] p2_sel_139615_comb;
  wire [15:0] p2_sel_139616_comb;
  wire [15:0] p2_sel_139617_comb;
  wire [15:0] p2_sel_139618_comb;
  wire [15:0] p2_sel_142427_comb;
  wire [15:0] p2_sel_142428_comb;
  wire [15:0] p2_sel_142429_comb;
  wire [15:0] p2_sel_142430_comb;
  wire [15:0] p2_sel_142431_comb;
  wire [15:0] p2_sel_142432_comb;
  wire [15:0] p2_sel_142433_comb;
  wire [15:0] p2_sel_142434_comb;
  wire [15:0] p2_sel_142435_comb;
  wire [15:0] p2_sel_142436_comb;
  wire [15:0] p2_sel_142437_comb;
  wire [15:0] p2_sel_142438_comb;
  wire [15:0] p2_sel_142439_comb;
  wire [15:0] p2_sel_142440_comb;
  wire [15:0] p2_sel_142441_comb;
  wire [15:0] p2_sel_142442_comb;
  wire [15:0] p2_sel_142659_comb;
  wire [15:0] p2_sel_142660_comb;
  wire [15:0] p2_sel_142661_comb;
  wire [15:0] p2_sel_142662_comb;
  wire [15:0] p2_sel_142663_comb;
  wire [15:0] p2_sel_142664_comb;
  wire [15:0] p2_sel_142665_comb;
  wire [15:0] p2_sel_142666_comb;
  wire [15:0] p2_sel_142667_comb;
  wire [15:0] p2_sel_142668_comb;
  wire [15:0] p2_sel_142669_comb;
  wire [15:0] p2_sel_142670_comb;
  wire [15:0] p2_sel_142671_comb;
  wire [15:0] p2_sel_142672_comb;
  wire [15:0] p2_sel_142673_comb;
  wire [15:0] p2_sel_142674_comb;
  wire [15:0] p2_sel_142675_comb;
  wire [15:0] p2_sel_142676_comb;
  wire [15:0] p2_sel_142677_comb;
  wire [15:0] p2_sel_142678_comb;
  wire [15:0] p2_sel_142679_comb;
  wire [15:0] p2_sel_142680_comb;
  wire [15:0] p2_sel_142681_comb;
  wire [15:0] p2_sel_142682_comb;
  wire [15:0] p2_sel_142683_comb;
  wire [15:0] p2_sel_142684_comb;
  wire [15:0] p2_sel_142685_comb;
  wire [15:0] p2_sel_142686_comb;
  wire [15:0] p2_sel_142687_comb;
  wire [15:0] p2_sel_142688_comb;
  wire [15:0] p2_sel_142689_comb;
  wire [15:0] p2_sel_142690_comb;
  wire [15:0] p2_sel_142691_comb;
  wire [15:0] p2_sel_142692_comb;
  wire [15:0] p2_sel_142693_comb;
  wire [15:0] p2_sel_142694_comb;
  wire [15:0] p2_sel_142695_comb;
  wire [15:0] p2_sel_142696_comb;
  wire [15:0] p2_sel_142697_comb;
  wire [15:0] p2_sel_142698_comb;
  wire [15:0] p2_sel_142699_comb;
  wire [15:0] p2_sel_142700_comb;
  wire [15:0] p2_sel_142701_comb;
  wire [15:0] p2_sel_142702_comb;
  wire [15:0] p2_sel_142703_comb;
  wire [15:0] p2_sel_142704_comb;
  wire [15:0] p2_sel_142705_comb;
  wire [15:0] p2_sel_142706_comb;
  wire [16:0] p2_add_142371_comb;
  wire [16:0] p2_add_142372_comb;
  wire [16:0] p2_add_142373_comb;
  wire [16:0] p2_add_142374_comb;
  wire [16:0] p2_add_142375_comb;
  wire [16:0] p2_add_142376_comb;
  wire [16:0] p2_add_142377_comb;
  wire [16:0] p2_add_142378_comb;
  wire [16:0] p2_add_142491_comb;
  wire [16:0] p2_add_142492_comb;
  wire [16:0] p2_add_142493_comb;
  wire [16:0] p2_add_142494_comb;
  wire [16:0] p2_add_142495_comb;
  wire [16:0] p2_add_142496_comb;
  wire [16:0] p2_add_142497_comb;
  wire [16:0] p2_add_142498_comb;
  wire [16:0] p2_add_142499_comb;
  wire [16:0] p2_add_142500_comb;
  wire [16:0] p2_add_142501_comb;
  wire [16:0] p2_add_142502_comb;
  wire [16:0] p2_add_142503_comb;
  wire [16:0] p2_add_142504_comb;
  wire [16:0] p2_add_142505_comb;
  wire [16:0] p2_add_142506_comb;
  wire [16:0] p2_add_142507_comb;
  wire [16:0] p2_add_142508_comb;
  wire [16:0] p2_add_142509_comb;
  wire [16:0] p2_add_142510_comb;
  wire [16:0] p2_add_142511_comb;
  wire [16:0] p2_add_142512_comb;
  wire [16:0] p2_add_142513_comb;
  wire [16:0] p2_add_142514_comb;
  wire [15:0] p2_sel_142531_comb;
  wire [15:0] p2_sel_142532_comb;
  wire [15:0] p2_sel_142533_comb;
  wire [15:0] p2_sel_142534_comb;
  wire [15:0] p2_sel_142535_comb;
  wire [15:0] p2_sel_142536_comb;
  wire [15:0] p2_sel_142537_comb;
  wire [15:0] p2_sel_142538_comb;
  wire [15:0] p2_sel_142539_comb;
  wire [15:0] p2_sel_142540_comb;
  wire [15:0] p2_sel_142541_comb;
  wire [15:0] p2_sel_142542_comb;
  wire [15:0] p2_sel_142543_comb;
  wire [15:0] p2_sel_142544_comb;
  wire [15:0] p2_sel_142545_comb;
  wire [15:0] p2_sel_142546_comb;
  wire [15:0] p2_sel_142627_comb;
  wire [15:0] p2_sel_142628_comb;
  wire [15:0] p2_sel_142629_comb;
  wire [15:0] p2_sel_142630_comb;
  wire [15:0] p2_sel_142631_comb;
  wire [15:0] p2_sel_142632_comb;
  wire [15:0] p2_sel_142633_comb;
  wire [15:0] p2_sel_142634_comb;
  wire [15:0] p2_sel_142635_comb;
  wire [15:0] p2_sel_142636_comb;
  wire [15:0] p2_sel_142637_comb;
  wire [15:0] p2_sel_142638_comb;
  wire [15:0] p2_sel_142639_comb;
  wire [15:0] p2_sel_142640_comb;
  wire [15:0] p2_sel_142641_comb;
  wire [15:0] p2_sel_142642_comb;
  wire [15:0] p2_sel_142723_comb;
  wire [15:0] p2_sel_142724_comb;
  wire [15:0] p2_sel_142725_comb;
  wire [15:0] p2_sel_142726_comb;
  wire [15:0] p2_sel_142727_comb;
  wire [15:0] p2_sel_142728_comb;
  wire [15:0] p2_sel_142729_comb;
  wire [15:0] p2_sel_142730_comb;
  wire [15:0] p2_sel_142731_comb;
  wire [15:0] p2_sel_142732_comb;
  wire [15:0] p2_sel_142733_comb;
  wire [15:0] p2_sel_142734_comb;
  wire [15:0] p2_sel_142735_comb;
  wire [15:0] p2_sel_142736_comb;
  wire [15:0] p2_sel_142737_comb;
  wire [15:0] p2_sel_142738_comb;
  wire [15:0] p2_sel_142819_comb;
  wire [15:0] p2_sel_142820_comb;
  wire [15:0] p2_sel_142821_comb;
  wire [15:0] p2_sel_142822_comb;
  wire [15:0] p2_sel_142823_comb;
  wire [15:0] p2_sel_142824_comb;
  wire [15:0] p2_sel_142825_comb;
  wire [15:0] p2_sel_142826_comb;
  wire [15:0] p2_sel_142827_comb;
  wire [15:0] p2_sel_142828_comb;
  wire [15:0] p2_sel_142829_comb;
  wire [15:0] p2_sel_142830_comb;
  wire [15:0] p2_sel_142831_comb;
  wire [15:0] p2_sel_142832_comb;
  wire [15:0] p2_sel_142833_comb;
  wire [15:0] p2_sel_142834_comb;
  wire [15:0] p2_sel_142379_comb;
  wire [15:0] p2_sel_142380_comb;
  wire [15:0] p2_sel_142381_comb;
  wire [15:0] p2_sel_142382_comb;
  wire [15:0] p2_sel_142383_comb;
  wire [15:0] p2_sel_142384_comb;
  wire [15:0] p2_sel_142385_comb;
  wire [15:0] p2_sel_142386_comb;
  wire [15:0] p2_sel_142387_comb;
  wire [15:0] p2_sel_142388_comb;
  wire [15:0] p2_sel_142389_comb;
  wire [15:0] p2_sel_142390_comb;
  wire [15:0] p2_sel_142391_comb;
  wire [15:0] p2_sel_142392_comb;
  wire [15:0] p2_sel_142393_comb;
  wire [15:0] p2_sel_142394_comb;
  wire [15:0] p2_sel_142395_comb;
  wire [15:0] p2_sel_142396_comb;
  wire [15:0] p2_sel_142397_comb;
  wire [15:0] p2_sel_142398_comb;
  wire [15:0] p2_sel_142399_comb;
  wire [15:0] p2_sel_142400_comb;
  wire [15:0] p2_sel_142401_comb;
  wire [15:0] p2_sel_142402_comb;
  wire [15:0] p2_sel_142403_comb;
  wire [15:0] p2_sel_142404_comb;
  wire [15:0] p2_sel_142405_comb;
  wire [15:0] p2_sel_142406_comb;
  wire [15:0] p2_sel_142407_comb;
  wire [15:0] p2_sel_142408_comb;
  wire [15:0] p2_sel_142409_comb;
  wire [15:0] p2_sel_142410_comb;
  wire [15:0] p2_sel_142411_comb;
  wire [15:0] p2_sel_142412_comb;
  wire [15:0] p2_sel_142413_comb;
  wire [15:0] p2_sel_142414_comb;
  wire [15:0] p2_sel_142415_comb;
  wire [15:0] p2_sel_142416_comb;
  wire [15:0] p2_sel_142417_comb;
  wire [15:0] p2_sel_142418_comb;
  wire [15:0] p2_sel_142419_comb;
  wire [15:0] p2_sel_142420_comb;
  wire [15:0] p2_sel_142421_comb;
  wire [15:0] p2_sel_142422_comb;
  wire [15:0] p2_sel_142423_comb;
  wire [15:0] p2_sel_142424_comb;
  wire [15:0] p2_sel_142425_comb;
  wire [15:0] p2_sel_142426_comb;
  wire [15:0] p2_sel_142443_comb;
  wire [15:0] p2_sel_142444_comb;
  wire [15:0] p2_sel_142445_comb;
  wire [15:0] p2_sel_142446_comb;
  wire [15:0] p2_sel_142447_comb;
  wire [15:0] p2_sel_142448_comb;
  wire [15:0] p2_sel_142449_comb;
  wire [15:0] p2_sel_142450_comb;
  wire [15:0] p2_sel_142451_comb;
  wire [15:0] p2_sel_142452_comb;
  wire [15:0] p2_sel_142453_comb;
  wire [15:0] p2_sel_142454_comb;
  wire [15:0] p2_sel_142455_comb;
  wire [15:0] p2_sel_142456_comb;
  wire [15:0] p2_sel_142457_comb;
  wire [15:0] p2_sel_142458_comb;
  wire [15:0] p2_sel_142459_comb;
  wire [15:0] p2_sel_142460_comb;
  wire [15:0] p2_sel_142461_comb;
  wire [15:0] p2_sel_142462_comb;
  wire [15:0] p2_sel_142463_comb;
  wire [15:0] p2_sel_142464_comb;
  wire [15:0] p2_sel_142465_comb;
  wire [15:0] p2_sel_142466_comb;
  wire [15:0] p2_sel_142467_comb;
  wire [15:0] p2_sel_142468_comb;
  wire [15:0] p2_sel_142469_comb;
  wire [15:0] p2_sel_142470_comb;
  wire [15:0] p2_sel_142471_comb;
  wire [15:0] p2_sel_142472_comb;
  wire [15:0] p2_sel_142473_comb;
  wire [15:0] p2_sel_142474_comb;
  wire [15:0] p2_sel_142475_comb;
  wire [15:0] p2_sel_142476_comb;
  wire [15:0] p2_sel_142477_comb;
  wire [15:0] p2_sel_142478_comb;
  wire [15:0] p2_sel_142479_comb;
  wire [15:0] p2_sel_142480_comb;
  wire [15:0] p2_sel_142481_comb;
  wire [15:0] p2_sel_142482_comb;
  wire [15:0] p2_sel_142483_comb;
  wire [15:0] p2_sel_142484_comb;
  wire [15:0] p2_sel_142485_comb;
  wire [15:0] p2_sel_142486_comb;
  wire [15:0] p2_sel_142487_comb;
  wire [15:0] p2_sel_142488_comb;
  wire [15:0] p2_sel_142489_comb;
  wire [15:0] p2_sel_142490_comb;
  wire [15:0] p2_sel_142515_comb;
  wire [15:0] p2_sel_142516_comb;
  wire [15:0] p2_sel_142517_comb;
  wire [15:0] p2_sel_142518_comb;
  wire [15:0] p2_sel_142519_comb;
  wire [15:0] p2_sel_142520_comb;
  wire [15:0] p2_sel_142521_comb;
  wire [15:0] p2_sel_142522_comb;
  wire [15:0] p2_sel_142523_comb;
  wire [15:0] p2_sel_142524_comb;
  wire [15:0] p2_sel_142525_comb;
  wire [15:0] p2_sel_142526_comb;
  wire [15:0] p2_sel_142527_comb;
  wire [15:0] p2_sel_142528_comb;
  wire [15:0] p2_sel_142529_comb;
  wire [15:0] p2_sel_142530_comb;
  wire [15:0] p2_sel_142547_comb;
  wire [15:0] p2_sel_142548_comb;
  wire [15:0] p2_sel_142549_comb;
  wire [15:0] p2_sel_142550_comb;
  wire [15:0] p2_sel_142551_comb;
  wire [15:0] p2_sel_142552_comb;
  wire [15:0] p2_sel_142553_comb;
  wire [15:0] p2_sel_142554_comb;
  wire [15:0] p2_sel_142555_comb;
  wire [15:0] p2_sel_142556_comb;
  wire [15:0] p2_sel_142557_comb;
  wire [15:0] p2_sel_142558_comb;
  wire [15:0] p2_sel_142559_comb;
  wire [15:0] p2_sel_142560_comb;
  wire [15:0] p2_sel_142561_comb;
  wire [15:0] p2_sel_142562_comb;
  wire [15:0] p2_sel_142563_comb;
  wire [15:0] p2_sel_142564_comb;
  wire [15:0] p2_sel_142565_comb;
  wire [15:0] p2_sel_142566_comb;
  wire [15:0] p2_sel_142567_comb;
  wire [15:0] p2_sel_142568_comb;
  wire [15:0] p2_sel_142569_comb;
  wire [15:0] p2_sel_142570_comb;
  wire [15:0] p2_sel_142571_comb;
  wire [15:0] p2_sel_142572_comb;
  wire [15:0] p2_sel_142573_comb;
  wire [15:0] p2_sel_142574_comb;
  wire [15:0] p2_sel_142575_comb;
  wire [15:0] p2_sel_142576_comb;
  wire [15:0] p2_sel_142577_comb;
  wire [15:0] p2_sel_142578_comb;
  wire [15:0] p2_sel_142579_comb;
  wire [15:0] p2_sel_142580_comb;
  wire [15:0] p2_sel_142581_comb;
  wire [15:0] p2_sel_142582_comb;
  wire [15:0] p2_sel_142583_comb;
  wire [15:0] p2_sel_142584_comb;
  wire [15:0] p2_sel_142585_comb;
  wire [15:0] p2_sel_142586_comb;
  wire [15:0] p2_sel_142587_comb;
  wire [15:0] p2_sel_142588_comb;
  wire [15:0] p2_sel_142589_comb;
  wire [15:0] p2_sel_142590_comb;
  wire [15:0] p2_sel_142591_comb;
  wire [15:0] p2_sel_142592_comb;
  wire [15:0] p2_sel_142593_comb;
  wire [15:0] p2_sel_142594_comb;
  wire [15:0] p2_sel_142595_comb;
  wire [15:0] p2_sel_142596_comb;
  wire [15:0] p2_sel_142597_comb;
  wire [15:0] p2_sel_142598_comb;
  wire [15:0] p2_sel_142599_comb;
  wire [15:0] p2_sel_142600_comb;
  wire [15:0] p2_sel_142601_comb;
  wire [15:0] p2_sel_142602_comb;
  wire [15:0] p2_sel_142603_comb;
  wire [15:0] p2_sel_142604_comb;
  wire [15:0] p2_sel_142605_comb;
  wire [15:0] p2_sel_142606_comb;
  wire [15:0] p2_sel_142607_comb;
  wire [15:0] p2_sel_142608_comb;
  wire [15:0] p2_sel_142609_comb;
  wire [15:0] p2_sel_142610_comb;
  wire [15:0] p2_sel_142611_comb;
  wire [15:0] p2_sel_142612_comb;
  wire [15:0] p2_sel_142613_comb;
  wire [15:0] p2_sel_142614_comb;
  wire [15:0] p2_sel_142615_comb;
  wire [15:0] p2_sel_142616_comb;
  wire [15:0] p2_sel_142617_comb;
  wire [15:0] p2_sel_142618_comb;
  wire [15:0] p2_sel_142619_comb;
  wire [15:0] p2_sel_142620_comb;
  wire [15:0] p2_sel_142621_comb;
  wire [15:0] p2_sel_142622_comb;
  wire [15:0] p2_sel_142623_comb;
  wire [15:0] p2_sel_142624_comb;
  wire [15:0] p2_sel_142625_comb;
  wire [15:0] p2_sel_142626_comb;
  wire [15:0] p2_sel_142643_comb;
  wire [15:0] p2_sel_142644_comb;
  wire [15:0] p2_sel_142645_comb;
  wire [15:0] p2_sel_142646_comb;
  wire [15:0] p2_sel_142647_comb;
  wire [15:0] p2_sel_142648_comb;
  wire [15:0] p2_sel_142649_comb;
  wire [15:0] p2_sel_142650_comb;
  wire [15:0] p2_sel_142651_comb;
  wire [15:0] p2_sel_142652_comb;
  wire [15:0] p2_sel_142653_comb;
  wire [15:0] p2_sel_142654_comb;
  wire [15:0] p2_sel_142655_comb;
  wire [15:0] p2_sel_142656_comb;
  wire [15:0] p2_sel_142657_comb;
  wire [15:0] p2_sel_142658_comb;
  wire [15:0] p2_sel_142707_comb;
  wire [15:0] p2_sel_142708_comb;
  wire [15:0] p2_sel_142709_comb;
  wire [15:0] p2_sel_142710_comb;
  wire [15:0] p2_sel_142711_comb;
  wire [15:0] p2_sel_142712_comb;
  wire [15:0] p2_sel_142713_comb;
  wire [15:0] p2_sel_142714_comb;
  wire [15:0] p2_sel_142715_comb;
  wire [15:0] p2_sel_142716_comb;
  wire [15:0] p2_sel_142717_comb;
  wire [15:0] p2_sel_142718_comb;
  wire [15:0] p2_sel_142719_comb;
  wire [15:0] p2_sel_142720_comb;
  wire [15:0] p2_sel_142721_comb;
  wire [15:0] p2_sel_142722_comb;
  wire [15:0] p2_sel_142739_comb;
  wire [15:0] p2_sel_142740_comb;
  wire [15:0] p2_sel_142741_comb;
  wire [15:0] p2_sel_142742_comb;
  wire [15:0] p2_sel_142743_comb;
  wire [15:0] p2_sel_142744_comb;
  wire [15:0] p2_sel_142745_comb;
  wire [15:0] p2_sel_142746_comb;
  wire [15:0] p2_sel_142747_comb;
  wire [15:0] p2_sel_142748_comb;
  wire [15:0] p2_sel_142749_comb;
  wire [15:0] p2_sel_142750_comb;
  wire [15:0] p2_sel_142751_comb;
  wire [15:0] p2_sel_142752_comb;
  wire [15:0] p2_sel_142753_comb;
  wire [15:0] p2_sel_142754_comb;
  wire [15:0] p2_sel_142755_comb;
  wire [15:0] p2_sel_142756_comb;
  wire [15:0] p2_sel_142757_comb;
  wire [15:0] p2_sel_142758_comb;
  wire [15:0] p2_sel_142759_comb;
  wire [15:0] p2_sel_142760_comb;
  wire [15:0] p2_sel_142761_comb;
  wire [15:0] p2_sel_142762_comb;
  wire [15:0] p2_sel_142763_comb;
  wire [15:0] p2_sel_142764_comb;
  wire [15:0] p2_sel_142765_comb;
  wire [15:0] p2_sel_142766_comb;
  wire [15:0] p2_sel_142767_comb;
  wire [15:0] p2_sel_142768_comb;
  wire [15:0] p2_sel_142769_comb;
  wire [15:0] p2_sel_142770_comb;
  wire [15:0] p2_sel_142771_comb;
  wire [15:0] p2_sel_142772_comb;
  wire [15:0] p2_sel_142773_comb;
  wire [15:0] p2_sel_142774_comb;
  wire [15:0] p2_sel_142775_comb;
  wire [15:0] p2_sel_142776_comb;
  wire [15:0] p2_sel_142777_comb;
  wire [15:0] p2_sel_142778_comb;
  wire [15:0] p2_sel_142779_comb;
  wire [15:0] p2_sel_142780_comb;
  wire [15:0] p2_sel_142781_comb;
  wire [15:0] p2_sel_142782_comb;
  wire [15:0] p2_sel_142783_comb;
  wire [15:0] p2_sel_142784_comb;
  wire [15:0] p2_sel_142785_comb;
  wire [15:0] p2_sel_142786_comb;
  wire [15:0] p2_sel_142787_comb;
  wire [15:0] p2_sel_142788_comb;
  wire [15:0] p2_sel_142789_comb;
  wire [15:0] p2_sel_142790_comb;
  wire [15:0] p2_sel_142791_comb;
  wire [15:0] p2_sel_142792_comb;
  wire [15:0] p2_sel_142793_comb;
  wire [15:0] p2_sel_142794_comb;
  wire [15:0] p2_sel_142795_comb;
  wire [15:0] p2_sel_142796_comb;
  wire [15:0] p2_sel_142797_comb;
  wire [15:0] p2_sel_142798_comb;
  wire [15:0] p2_sel_142799_comb;
  wire [15:0] p2_sel_142800_comb;
  wire [15:0] p2_sel_142801_comb;
  wire [15:0] p2_sel_142802_comb;
  wire [15:0] p2_sel_142803_comb;
  wire [15:0] p2_sel_142804_comb;
  wire [15:0] p2_sel_142805_comb;
  wire [15:0] p2_sel_142806_comb;
  wire [15:0] p2_sel_142807_comb;
  wire [15:0] p2_sel_142808_comb;
  wire [15:0] p2_sel_142809_comb;
  wire [15:0] p2_sel_142810_comb;
  wire [15:0] p2_sel_142811_comb;
  wire [15:0] p2_sel_142812_comb;
  wire [15:0] p2_sel_142813_comb;
  wire [15:0] p2_sel_142814_comb;
  wire [15:0] p2_sel_142815_comb;
  wire [15:0] p2_sel_142816_comb;
  wire [15:0] p2_sel_142817_comb;
  wire [15:0] p2_sel_142818_comb;
  wire [15:0] p2_sel_142835_comb;
  wire [15:0] p2_sel_142836_comb;
  wire [15:0] p2_sel_142837_comb;
  wire [15:0] p2_sel_142838_comb;
  wire [15:0] p2_sel_142839_comb;
  wire [15:0] p2_sel_142840_comb;
  wire [15:0] p2_sel_142841_comb;
  wire [15:0] p2_sel_142842_comb;
  wire [15:0] p2_sel_142843_comb;
  wire [15:0] p2_sel_142844_comb;
  wire [15:0] p2_sel_142845_comb;
  wire [15:0] p2_sel_142846_comb;
  wire [15:0] p2_sel_142847_comb;
  wire [15:0] p2_sel_142848_comb;
  wire [15:0] p2_sel_142849_comb;
  wire [15:0] p2_sel_142850_comb;
  wire [31:0] p2_sum__989_comb;
  wire [31:0] p2_sum__990_comb;
  wire [31:0] p2_sum__991_comb;
  wire [31:0] p2_sum__992_comb;
  wire [31:0] p2_sum__884_comb;
  wire [31:0] p2_sum__885_comb;
  wire [31:0] p2_sum__886_comb;
  wire [31:0] p2_sum__887_comb;
  wire [31:0] p2_sum__1017_comb;
  wire [31:0] p2_sum__1018_comb;
  wire [31:0] p2_sum__1019_comb;
  wire [31:0] p2_sum__1020_comb;
  wire [31:0] p2_sum__1010_comb;
  wire [31:0] p2_sum__1011_comb;
  wire [31:0] p2_sum__1012_comb;
  wire [31:0] p2_sum__1013_comb;
  wire [31:0] p2_sum__961_comb;
  wire [31:0] p2_sum__962_comb;
  wire [31:0] p2_sum__963_comb;
  wire [31:0] p2_sum__964_comb;
  wire [31:0] p2_sum__926_comb;
  wire [31:0] p2_sum__927_comb;
  wire [31:0] p2_sum__928_comb;
  wire [31:0] p2_sum__929_comb;
  wire [31:0] p2_sum__835_comb;
  wire [31:0] p2_sum__836_comb;
  wire [31:0] p2_sum__837_comb;
  wire [31:0] p2_sum__838_comb;
  wire [31:0] p2_sum__779_comb;
  wire [31:0] p2_sum__780_comb;
  wire [31:0] p2_sum__781_comb;
  wire [31:0] p2_sum__782_comb;
  wire [16:0] p2_add_143359_comb;
  wire [16:0] p2_add_143360_comb;
  wire [16:0] p2_add_143361_comb;
  wire [16:0] p2_add_143362_comb;
  wire [16:0] p2_add_143363_comb;
  wire [16:0] p2_add_143364_comb;
  wire [16:0] p2_add_143365_comb;
  wire [16:0] p2_add_143366_comb;
  wire [16:0] p2_add_143475_comb;
  wire [16:0] p2_add_143476_comb;
  wire [16:0] p2_add_143477_comb;
  wire [16:0] p2_add_143478_comb;
  wire [16:0] p2_add_143479_comb;
  wire [16:0] p2_add_143480_comb;
  wire [16:0] p2_add_143481_comb;
  wire [16:0] p2_add_143482_comb;
  wire [16:0] p2_add_143483_comb;
  wire [16:0] p2_add_143484_comb;
  wire [16:0] p2_add_143485_comb;
  wire [16:0] p2_add_143486_comb;
  wire [16:0] p2_add_143487_comb;
  wire [16:0] p2_add_143488_comb;
  wire [16:0] p2_add_143489_comb;
  wire [16:0] p2_add_143490_comb;
  wire [16:0] p2_add_143491_comb;
  wire [16:0] p2_add_143492_comb;
  wire [16:0] p2_add_143493_comb;
  wire [16:0] p2_add_143494_comb;
  wire [16:0] p2_add_143495_comb;
  wire [16:0] p2_add_143496_comb;
  wire [16:0] p2_add_143497_comb;
  wire [16:0] p2_add_143498_comb;
  wire [31:0] p2_sum__993_comb;
  wire [31:0] p2_sum__994_comb;
  wire [31:0] p2_sum__888_comb;
  wire [31:0] p2_sum__889_comb;
  wire [31:0] p2_sum__1021_comb;
  wire [31:0] p2_sum__1022_comb;
  wire [31:0] p2_sum__1014_comb;
  wire [31:0] p2_sum__1015_comb;
  wire [31:0] p2_sum__965_comb;
  wire [31:0] p2_sum__966_comb;
  wire [31:0] p2_sum__930_comb;
  wire [31:0] p2_sum__931_comb;
  wire [31:0] p2_sum__839_comb;
  wire [31:0] p2_sum__840_comb;
  wire [31:0] p2_sum__783_comb;
  wire [31:0] p2_sum__784_comb;
  wire [16:0] p2_add_143411_comb;
  wire [16:0] p2_add_143412_comb;
  wire [16:0] p2_add_143413_comb;
  wire [16:0] p2_add_143414_comb;
  wire [16:0] p2_add_143415_comb;
  wire [16:0] p2_add_143416_comb;
  wire [16:0] p2_add_143417_comb;
  wire [16:0] p2_add_143418_comb;
  wire [16:0] p2_add_143459_comb;
  wire [16:0] p2_add_143460_comb;
  wire [16:0] p2_add_143461_comb;
  wire [16:0] p2_add_143462_comb;
  wire [16:0] p2_add_143463_comb;
  wire [16:0] p2_add_143464_comb;
  wire [16:0] p2_add_143465_comb;
  wire [16:0] p2_add_143466_comb;
  wire [16:0] p2_add_143507_comb;
  wire [16:0] p2_add_143508_comb;
  wire [16:0] p2_add_143509_comb;
  wire [16:0] p2_add_143510_comb;
  wire [16:0] p2_add_143511_comb;
  wire [16:0] p2_add_143512_comb;
  wire [16:0] p2_add_143513_comb;
  wire [16:0] p2_add_143514_comb;
  wire [16:0] p2_add_143555_comb;
  wire [16:0] p2_add_143556_comb;
  wire [16:0] p2_add_143557_comb;
  wire [16:0] p2_add_143558_comb;
  wire [16:0] p2_add_143559_comb;
  wire [16:0] p2_add_143560_comb;
  wire [16:0] p2_add_143561_comb;
  wire [16:0] p2_add_143562_comb;
  wire [24:0] p2_sum__1736_comb;
  wire [24:0] p2_sum__1737_comb;
  wire [24:0] p2_sum__1738_comb;
  wire [24:0] p2_sum__1739_comb;
  wire [24:0] p2_sum__1652_comb;
  wire [24:0] p2_sum__1653_comb;
  wire [24:0] p2_sum__1654_comb;
  wire [24:0] p2_sum__1655_comb;
  wire [24:0] p2_sum__1780_comb;
  wire [24:0] p2_sum__1781_comb;
  wire [24:0] p2_sum__1782_comb;
  wire [24:0] p2_sum__1783_comb;
  wire [24:0] p2_sum__1760_comb;
  wire [24:0] p2_sum__1761_comb;
  wire [24:0] p2_sum__1762_comb;
  wire [24:0] p2_sum__1763_comb;
  wire [24:0] p2_sum__1708_comb;
  wire [24:0] p2_sum__1709_comb;
  wire [24:0] p2_sum__1710_comb;
  wire [24:0] p2_sum__1711_comb;
  wire [24:0] p2_sum__1680_comb;
  wire [24:0] p2_sum__1681_comb;
  wire [24:0] p2_sum__1682_comb;
  wire [24:0] p2_sum__1683_comb;
  wire [24:0] p2_sum__1628_comb;
  wire [24:0] p2_sum__1629_comb;
  wire [24:0] p2_sum__1630_comb;
  wire [24:0] p2_sum__1631_comb;
  wire [24:0] p2_sum__1608_comb;
  wire [24:0] p2_sum__1609_comb;
  wire [24:0] p2_sum__1610_comb;
  wire [24:0] p2_sum__1611_comb;
  wire [16:0] p2_add_143335_comb;
  wire [16:0] p2_add_143336_comb;
  wire [16:0] p2_add_143337_comb;
  wire [16:0] p2_add_143338_comb;
  wire [16:0] p2_add_143339_comb;
  wire [16:0] p2_add_143340_comb;
  wire [16:0] p2_add_143341_comb;
  wire [16:0] p2_add_143342_comb;
  wire [16:0] p2_add_143343_comb;
  wire [16:0] p2_add_143344_comb;
  wire [16:0] p2_add_143345_comb;
  wire [16:0] p2_add_143346_comb;
  wire [16:0] p2_add_143347_comb;
  wire [16:0] p2_add_143348_comb;
  wire [16:0] p2_add_143349_comb;
  wire [16:0] p2_add_143350_comb;
  wire [16:0] p2_add_143351_comb;
  wire [16:0] p2_add_143352_comb;
  wire [16:0] p2_add_143353_comb;
  wire [16:0] p2_add_143354_comb;
  wire [16:0] p2_add_143355_comb;
  wire [16:0] p2_add_143356_comb;
  wire [16:0] p2_add_143357_comb;
  wire [16:0] p2_add_143358_comb;
  wire [16:0] p2_add_143367_comb;
  wire [16:0] p2_add_143368_comb;
  wire [16:0] p2_add_143369_comb;
  wire [16:0] p2_add_143370_comb;
  wire [16:0] p2_add_143371_comb;
  wire [16:0] p2_add_143372_comb;
  wire [16:0] p2_add_143373_comb;
  wire [16:0] p2_add_143374_comb;
  wire [16:0] p2_add_143375_comb;
  wire [16:0] p2_add_143376_comb;
  wire [16:0] p2_add_143377_comb;
  wire [16:0] p2_add_143378_comb;
  wire [16:0] p2_add_143379_comb;
  wire [16:0] p2_add_143380_comb;
  wire [16:0] p2_add_143381_comb;
  wire [16:0] p2_add_143382_comb;
  wire [16:0] p2_add_143383_comb;
  wire [16:0] p2_add_143384_comb;
  wire [16:0] p2_add_143385_comb;
  wire [16:0] p2_add_143386_comb;
  wire [16:0] p2_add_143387_comb;
  wire [16:0] p2_add_143388_comb;
  wire [16:0] p2_add_143389_comb;
  wire [16:0] p2_add_143390_comb;
  wire [16:0] p2_add_143403_comb;
  wire [16:0] p2_add_143404_comb;
  wire [16:0] p2_add_143405_comb;
  wire [16:0] p2_add_143406_comb;
  wire [16:0] p2_add_143407_comb;
  wire [16:0] p2_add_143408_comb;
  wire [16:0] p2_add_143409_comb;
  wire [16:0] p2_add_143410_comb;
  wire [16:0] p2_add_143419_comb;
  wire [16:0] p2_add_143420_comb;
  wire [16:0] p2_add_143421_comb;
  wire [16:0] p2_add_143422_comb;
  wire [16:0] p2_add_143423_comb;
  wire [16:0] p2_add_143424_comb;
  wire [16:0] p2_add_143425_comb;
  wire [16:0] p2_add_143426_comb;
  wire [16:0] p2_add_143427_comb;
  wire [16:0] p2_add_143428_comb;
  wire [16:0] p2_add_143429_comb;
  wire [16:0] p2_add_143430_comb;
  wire [16:0] p2_add_143431_comb;
  wire [16:0] p2_add_143432_comb;
  wire [16:0] p2_add_143433_comb;
  wire [16:0] p2_add_143434_comb;
  wire [16:0] p2_add_143435_comb;
  wire [16:0] p2_add_143436_comb;
  wire [16:0] p2_add_143437_comb;
  wire [16:0] p2_add_143438_comb;
  wire [16:0] p2_add_143439_comb;
  wire [16:0] p2_add_143440_comb;
  wire [16:0] p2_add_143441_comb;
  wire [16:0] p2_add_143442_comb;
  wire [16:0] p2_add_143443_comb;
  wire [16:0] p2_add_143444_comb;
  wire [16:0] p2_add_143445_comb;
  wire [16:0] p2_add_143446_comb;
  wire [16:0] p2_add_143447_comb;
  wire [16:0] p2_add_143448_comb;
  wire [16:0] p2_add_143449_comb;
  wire [16:0] p2_add_143450_comb;
  wire [16:0] p2_add_143451_comb;
  wire [16:0] p2_add_143452_comb;
  wire [16:0] p2_add_143453_comb;
  wire [16:0] p2_add_143454_comb;
  wire [16:0] p2_add_143455_comb;
  wire [16:0] p2_add_143456_comb;
  wire [16:0] p2_add_143457_comb;
  wire [16:0] p2_add_143458_comb;
  wire [16:0] p2_add_143467_comb;
  wire [16:0] p2_add_143468_comb;
  wire [16:0] p2_add_143469_comb;
  wire [16:0] p2_add_143470_comb;
  wire [16:0] p2_add_143471_comb;
  wire [16:0] p2_add_143472_comb;
  wire [16:0] p2_add_143473_comb;
  wire [16:0] p2_add_143474_comb;
  wire [16:0] p2_add_143499_comb;
  wire [16:0] p2_add_143500_comb;
  wire [16:0] p2_add_143501_comb;
  wire [16:0] p2_add_143502_comb;
  wire [16:0] p2_add_143503_comb;
  wire [16:0] p2_add_143504_comb;
  wire [16:0] p2_add_143505_comb;
  wire [16:0] p2_add_143506_comb;
  wire [16:0] p2_add_143515_comb;
  wire [16:0] p2_add_143516_comb;
  wire [16:0] p2_add_143517_comb;
  wire [16:0] p2_add_143518_comb;
  wire [16:0] p2_add_143519_comb;
  wire [16:0] p2_add_143520_comb;
  wire [16:0] p2_add_143521_comb;
  wire [16:0] p2_add_143522_comb;
  wire [16:0] p2_add_143523_comb;
  wire [16:0] p2_add_143524_comb;
  wire [16:0] p2_add_143525_comb;
  wire [16:0] p2_add_143526_comb;
  wire [16:0] p2_add_143527_comb;
  wire [16:0] p2_add_143528_comb;
  wire [16:0] p2_add_143529_comb;
  wire [16:0] p2_add_143530_comb;
  wire [16:0] p2_add_143531_comb;
  wire [16:0] p2_add_143532_comb;
  wire [16:0] p2_add_143533_comb;
  wire [16:0] p2_add_143534_comb;
  wire [16:0] p2_add_143535_comb;
  wire [16:0] p2_add_143536_comb;
  wire [16:0] p2_add_143537_comb;
  wire [16:0] p2_add_143538_comb;
  wire [16:0] p2_add_143539_comb;
  wire [16:0] p2_add_143540_comb;
  wire [16:0] p2_add_143541_comb;
  wire [16:0] p2_add_143542_comb;
  wire [16:0] p2_add_143543_comb;
  wire [16:0] p2_add_143544_comb;
  wire [16:0] p2_add_143545_comb;
  wire [16:0] p2_add_143546_comb;
  wire [16:0] p2_add_143547_comb;
  wire [16:0] p2_add_143548_comb;
  wire [16:0] p2_add_143549_comb;
  wire [16:0] p2_add_143550_comb;
  wire [16:0] p2_add_143551_comb;
  wire [16:0] p2_add_143552_comb;
  wire [16:0] p2_add_143553_comb;
  wire [16:0] p2_add_143554_comb;
  wire [16:0] p2_add_143563_comb;
  wire [16:0] p2_add_143564_comb;
  wire [16:0] p2_add_143565_comb;
  wire [16:0] p2_add_143566_comb;
  wire [16:0] p2_add_143567_comb;
  wire [16:0] p2_add_143568_comb;
  wire [16:0] p2_add_143569_comb;
  wire [16:0] p2_add_143570_comb;
  wire [31:0] p2_sum__995_comb;
  wire [31:0] p2_sum__890_comb;
  wire [31:0] p2_sum__1023_comb;
  wire [31:0] p2_sum__1016_comb;
  wire [31:0] p2_sum__967_comb;
  wire [31:0] p2_sum__932_comb;
  wire [31:0] p2_sum__841_comb;
  wire [31:0] p2_sum__785_comb;
  wire [24:0] p2_sum__1768_comb;
  wire [24:0] p2_sum__1769_comb;
  wire [24:0] p2_sum__1770_comb;
  wire [24:0] p2_sum__1771_comb;
  wire [24:0] p2_sum__1748_comb;
  wire [24:0] p2_sum__1749_comb;
  wire [24:0] p2_sum__1750_comb;
  wire [24:0] p2_sum__1751_comb;
  wire [24:0] p2_sum__1732_comb;
  wire [24:0] p2_sum__1733_comb;
  wire [24:0] p2_sum__1734_comb;
  wire [24:0] p2_sum__1735_comb;
  wire [24:0] p2_sum__1704_comb;
  wire [24:0] p2_sum__1705_comb;
  wire [24:0] p2_sum__1706_comb;
  wire [24:0] p2_sum__1707_comb;
  wire [24:0] p2_sum__1684_comb;
  wire [24:0] p2_sum__1685_comb;
  wire [24:0] p2_sum__1686_comb;
  wire [24:0] p2_sum__1687_comb;
  wire [24:0] p2_sum__1656_comb;
  wire [24:0] p2_sum__1657_comb;
  wire [24:0] p2_sum__1658_comb;
  wire [24:0] p2_sum__1659_comb;
  wire [24:0] p2_sum__1640_comb;
  wire [24:0] p2_sum__1641_comb;
  wire [24:0] p2_sum__1642_comb;
  wire [24:0] p2_sum__1643_comb;
  wire [24:0] p2_sum__1620_comb;
  wire [24:0] p2_sum__1621_comb;
  wire [24:0] p2_sum__1622_comb;
  wire [24:0] p2_sum__1623_comb;
  wire [24:0] p2_sum__1324_comb;
  wire [24:0] p2_sum__1325_comb;
  wire [24:0] p2_sum__1282_comb;
  wire [24:0] p2_sum__1283_comb;
  wire [24:0] p2_sum__1346_comb;
  wire [24:0] p2_sum__1347_comb;
  wire [24:0] p2_sum__1336_comb;
  wire [24:0] p2_sum__1337_comb;
  wire [24:0] p2_sum__1310_comb;
  wire [24:0] p2_sum__1311_comb;
  wire [24:0] p2_sum__1296_comb;
  wire [24:0] p2_sum__1297_comb;
  wire [24:0] p2_sum__1270_comb;
  wire [24:0] p2_sum__1271_comb;
  wire [24:0] p2_sum__1260_comb;
  wire [24:0] p2_sum__1261_comb;
  assign p2_smul_57330_TrailingBits___9_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___10_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___21_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___22_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___72_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___75_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___84_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___87_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___105_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___106_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___117_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___118_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___168_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___171_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___180_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___183_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___1_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___2_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___5_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___6_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___25_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___26_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___29_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___30_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___64_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___67_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___68_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___71_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___88_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___91_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___92_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___95_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___97_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___98_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___101_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___102_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___121_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___122_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___125_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___126_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___160_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___163_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___164_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___167_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___184_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___187_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___188_comb = 9'h000;
  assign p2_smul_57330_TrailingBits___191_comb = 9'h000;
  assign p2_prod__135_comb = {{7{p1_concat_134899[24]}}, p1_concat_134899};
  assign p2_concat_136661_comb = {p1_smul_57364_NarrowedMult_, p2_smul_57330_TrailingBits___9_comb};
  assign p2_concat_136662_comb = {p1_smul_57366_NarrowedMult_, p2_smul_57330_TrailingBits___10_comb};
  assign p2_prod__150_comb = {{7{p1_concat_134902[24]}}, p1_concat_134902};
  assign p2_prod__327_comb = {{7{p1_concat_134903[24]}}, p1_concat_134903};
  assign p2_concat_136667_comb = {p1_smul_57412_NarrowedMult_, p2_smul_57330_TrailingBits___21_comb};
  assign p2_concat_136668_comb = {p1_smul_57414_NarrowedMult_, p2_smul_57330_TrailingBits___22_comb};
  assign p2_prod__342_comb = {{7{p1_concat_134906[24]}}, p1_concat_134906};
  assign p2_prod__133_comb = {{7{p1_concat_134907[24]}}, p1_concat_134907};
  assign p2_prod__136_comb = {{8{p1_concat_134908[23]}}, p1_concat_134908};
  assign p2_prod__140_comb = {{8{p1_concat_134909[23]}}, p1_concat_134909};
  assign p2_prod__145_comb = {{7{p1_concat_134910[24]}}, p1_concat_134910};
  assign p2_prod__151_comb = {{7{p1_concat_134911[24]}}, p1_concat_134911};
  assign p2_prod__158_comb = {{8{p1_concat_134912[23]}}, p1_concat_134912};
  assign p2_prod__165_comb = {{8{p1_concat_134913[23]}}, p1_concat_134913};
  assign p2_prod__171_comb = {{7{p1_concat_134914[24]}}, p1_concat_134914};
  assign p2_prod__325_comb = {{7{p1_concat_134915[24]}}, p1_concat_134915};
  assign p2_prod__328_comb = {{8{p1_concat_134916[23]}}, p1_concat_134916};
  assign p2_prod__332_comb = {{8{p1_concat_134917[23]}}, p1_concat_134917};
  assign p2_prod__337_comb = {{7{p1_concat_134918[24]}}, p1_concat_134918};
  assign p2_prod__343_comb = {{7{p1_concat_134919[24]}}, p1_concat_134919};
  assign p2_prod__350_comb = {{8{p1_concat_134920[23]}}, p1_concat_134920};
  assign p2_prod__357_comb = {{8{p1_concat_134921[23]}}, p1_concat_134921};
  assign p2_prod__363_comb = {{7{p1_concat_134922[24]}}, p1_concat_134922};
  assign p2_concat_136695_comb = {p1_smul_57616_NarrowedMult_, p2_smul_57330_TrailingBits___72_comb};
  assign p2_prod__152_comb = {{7{p1_concat_134924[24]}}, p1_concat_134924};
  assign p2_prod__159_comb = {{7{p1_concat_134925[24]}}, p1_concat_134925};
  assign p2_concat_136700_comb = {p1_smul_57626_NarrowedMult_, p2_smul_57330_TrailingBits___75_comb};
  assign p2_concat_136701_comb = {p1_smul_57664_NarrowedMult_, p2_smul_57330_TrailingBits___84_comb};
  assign p2_prod__344_comb = {{7{p1_concat_134928[24]}}, p1_concat_134928};
  assign p2_prod__351_comb = {{7{p1_concat_134929[24]}}, p1_concat_134929};
  assign p2_concat_136706_comb = {p1_smul_57674_NarrowedMult_, p2_smul_57330_TrailingBits___87_comb};
  assign p2_prod__148_comb = {{7{p1_concat_134931[24]}}, p1_concat_134931};
  assign p2_concat_136709_comb = {p1_smul_57874_NarrowedMult_, p2_smul_57330_TrailingBits___105_comb};
  assign p2_concat_136710_comb = {p1_smul_57880_NarrowedMult_, p2_smul_57330_TrailingBits___106_comb};
  assign p2_prod__186_comb = {{7{p1_concat_134934[24]}}, p1_concat_134934};
  assign p2_prod__340_comb = {{7{p1_concat_134935[24]}}, p1_concat_134935};
  assign p2_concat_136715_comb = {p1_smul_57922_NarrowedMult_, p2_smul_57330_TrailingBits___117_comb};
  assign p2_concat_136716_comb = {p1_smul_57928_NarrowedMult_, p2_smul_57330_TrailingBits___118_comb};
  assign p2_prod__378_comb = {{7{p1_concat_134938[24]}}, p1_concat_134938};
  assign p2_prod__155_comb = {{8{p1_concat_134939[23]}}, p1_concat_134939};
  assign p2_prod__162_comb = {{7{p1_concat_134940[24]}}, p1_concat_134940};
  assign p2_prod__169_comb = {{8{p1_concat_134941[23]}}, p1_concat_134941};
  assign p2_prod__175_comb = {{7{p1_concat_134942[24]}}, p1_concat_134942};
  assign p2_prod__180_comb = {{7{p1_concat_134943[24]}}, p1_concat_134943};
  assign p2_prod__184_comb = {{8{p1_concat_134944[23]}}, p1_concat_134944};
  assign p2_prod__187_comb = {{7{p1_concat_134945[24]}}, p1_concat_134945};
  assign p2_prod__189_comb = {{8{p1_concat_134946[23]}}, p1_concat_134946};
  assign p2_prod__347_comb = {{8{p1_concat_134947[23]}}, p1_concat_134947};
  assign p2_prod__354_comb = {{7{p1_concat_134948[24]}}, p1_concat_134948};
  assign p2_prod__361_comb = {{8{p1_concat_134949[23]}}, p1_concat_134949};
  assign p2_prod__367_comb = {{7{p1_concat_134950[24]}}, p1_concat_134950};
  assign p2_prod__372_comb = {{7{p1_concat_134951[24]}}, p1_concat_134951};
  assign p2_prod__376_comb = {{8{p1_concat_134952[23]}}, p1_concat_134952};
  assign p2_prod__379_comb = {{7{p1_concat_134953[24]}}, p1_concat_134953};
  assign p2_prod__381_comb = {{8{p1_concat_134954[23]}}, p1_concat_134954};
  assign p2_concat_136743_comb = {p1_smul_58126_NarrowedMult_, p2_smul_57330_TrailingBits___168_comb};
  assign p2_prod__170_comb = {{7{p1_concat_134956[24]}}, p1_concat_134956};
  assign p2_prod__190_comb = {{7{p1_concat_134957[24]}}, p1_concat_134957};
  assign p2_concat_136748_comb = {p1_smul_58140_NarrowedMult_, p2_smul_57330_TrailingBits___171_comb};
  assign p2_concat_136749_comb = {p1_smul_58174_NarrowedMult_, p2_smul_57330_TrailingBits___180_comb};
  assign p2_prod__362_comb = {{7{p1_concat_134960[24]}}, p1_concat_134960};
  assign p2_prod__382_comb = {{7{p1_concat_134961[24]}}, p1_concat_134961};
  assign p2_concat_136754_comb = {p1_smul_58188_NarrowedMult_, p2_smul_57330_TrailingBits___183_comb};
  assign p2_prod__10_comb = {{7{p1_concat_135011[24]}}, p1_concat_135011};
  assign p2_concat_136805_comb = {p1_smul_57332_NarrowedMult_, p2_smul_57330_TrailingBits___1_comb};
  assign p2_concat_136806_comb = {p1_smul_57334_NarrowedMult_, p2_smul_57330_TrailingBits___2_comb};
  assign p2_prod__13_comb = {{7{p1_concat_135014[24]}}, p1_concat_135014};
  assign p2_prod__71_comb = {{7{p1_concat_135015[24]}}, p1_concat_135015};
  assign p2_concat_136811_comb = {p1_smul_57348_NarrowedMult_, p2_smul_57330_TrailingBits___5_comb};
  assign p2_concat_136812_comb = {p1_smul_57350_NarrowedMult_, p2_smul_57330_TrailingBits___6_comb};
  assign p2_prod__86_comb = {{7{p1_concat_135018[24]}}, p1_concat_135018};
  assign p2_prod__391_comb = {{7{p1_concat_135031[24]}}, p1_concat_135031};
  assign p2_concat_136821_comb = {p1_smul_57428_NarrowedMult_, p2_smul_57330_TrailingBits___25_comb};
  assign p2_concat_136822_comb = {p1_smul_57430_NarrowedMult_, p2_smul_57330_TrailingBits___26_comb};
  assign p2_prod__406_comb = {{7{p1_concat_135034[24]}}, p1_concat_135034};
  assign p2_prod__455_comb = {{7{p1_concat_135035[24]}}, p1_concat_135035};
  assign p2_concat_136827_comb = {p1_smul_57444_NarrowedMult_, p2_smul_57330_TrailingBits___29_comb};
  assign p2_concat_136828_comb = {p1_smul_57446_NarrowedMult_, p2_smul_57330_TrailingBits___30_comb};
  assign p2_prod__470_comb = {{7{p1_concat_135038[24]}}, p1_concat_135038};
  assign p2_prod__16_comb = {{7{p1_concat_135039[24]}}, p1_concat_135039};
  assign p2_prod__17_comb = {{8{p1_concat_135040[23]}}, p1_concat_135040};
  assign p2_prod__18_comb = {{8{p1_concat_135041[23]}}, p1_concat_135041};
  assign p2_prod__19_comb = {{7{p1_concat_135042[24]}}, p1_concat_135042};
  assign p2_prod__20_comb = {{7{p1_concat_135043[24]}}, p1_concat_135043};
  assign p2_prod__21_comb = {{8{p1_concat_135044[23]}}, p1_concat_135044};
  assign p2_prod__22_comb = {{8{p1_concat_135045[23]}}, p1_concat_135045};
  assign p2_prod__23_comb = {{7{p1_concat_135046[24]}}, p1_concat_135046};
  assign p2_prod__69_comb = {{7{p1_concat_135047[24]}}, p1_concat_135047};
  assign p2_prod__72_comb = {{8{p1_concat_135048[23]}}, p1_concat_135048};
  assign p2_prod__76_comb = {{8{p1_concat_135049[23]}}, p1_concat_135049};
  assign p2_prod__81_comb = {{7{p1_concat_135050[24]}}, p1_concat_135050};
  assign p2_prod__87_comb = {{7{p1_concat_135051[24]}}, p1_concat_135051};
  assign p2_prod__94_comb = {{8{p1_concat_135052[23]}}, p1_concat_135052};
  assign p2_prod__101_comb = {{8{p1_concat_135053[23]}}, p1_concat_135053};
  assign p2_prod__107_comb = {{7{p1_concat_135054[24]}}, p1_concat_135054};
  assign p2_prod__197_comb = {{7{p1_concat_135055[24]}}, p1_concat_135055};
  assign p2_prod__200_comb = {{8{p1_concat_135056[23]}}, p1_concat_135056};
  assign p2_prod__204_comb = {{8{p1_concat_135057[23]}}, p1_concat_135057};
  assign p2_prod__209_comb = {{7{p1_concat_135058[24]}}, p1_concat_135058};
  assign p2_prod__215_comb = {{7{p1_concat_135059[24]}}, p1_concat_135059};
  assign p2_prod__222_comb = {{8{p1_concat_135060[23]}}, p1_concat_135060};
  assign p2_prod__229_comb = {{8{p1_concat_135061[23]}}, p1_concat_135061};
  assign p2_prod__235_comb = {{7{p1_concat_135062[24]}}, p1_concat_135062};
  assign p2_prod__261_comb = {{7{p1_concat_135063[24]}}, p1_concat_135063};
  assign p2_prod__264_comb = {{8{p1_concat_135064[23]}}, p1_concat_135064};
  assign p2_prod__268_comb = {{8{p1_concat_135065[23]}}, p1_concat_135065};
  assign p2_prod__273_comb = {{7{p1_concat_135066[24]}}, p1_concat_135066};
  assign p2_prod__279_comb = {{7{p1_concat_135067[24]}}, p1_concat_135067};
  assign p2_prod__286_comb = {{8{p1_concat_135068[23]}}, p1_concat_135068};
  assign p2_prod__293_comb = {{8{p1_concat_135069[23]}}, p1_concat_135069};
  assign p2_prod__299_comb = {{7{p1_concat_135070[24]}}, p1_concat_135070};
  assign p2_prod__389_comb = {{7{p1_concat_135071[24]}}, p1_concat_135071};
  assign p2_prod__392_comb = {{8{p1_concat_135072[23]}}, p1_concat_135072};
  assign p2_prod__396_comb = {{8{p1_concat_135073[23]}}, p1_concat_135073};
  assign p2_prod__401_comb = {{7{p1_concat_135074[24]}}, p1_concat_135074};
  assign p2_prod__407_comb = {{7{p1_concat_135075[24]}}, p1_concat_135075};
  assign p2_prod__414_comb = {{8{p1_concat_135076[23]}}, p1_concat_135076};
  assign p2_prod__421_comb = {{8{p1_concat_135077[23]}}, p1_concat_135077};
  assign p2_prod__427_comb = {{7{p1_concat_135078[24]}}, p1_concat_135078};
  assign p2_prod__453_comb = {{7{p1_concat_135079[24]}}, p1_concat_135079};
  assign p2_prod__456_comb = {{8{p1_concat_135080[23]}}, p1_concat_135080};
  assign p2_prod__460_comb = {{8{p1_concat_135081[23]}}, p1_concat_135081};
  assign p2_prod__465_comb = {{7{p1_concat_135082[24]}}, p1_concat_135082};
  assign p2_prod__471_comb = {{7{p1_concat_135083[24]}}, p1_concat_135083};
  assign p2_prod__478_comb = {{8{p1_concat_135084[23]}}, p1_concat_135084};
  assign p2_prod__485_comb = {{8{p1_concat_135085[23]}}, p1_concat_135085};
  assign p2_prod__491_comb = {{7{p1_concat_135086[24]}}, p1_concat_135086};
  assign p2_concat_136903_comb = {p1_smul_57584_NarrowedMult_, p2_smul_57330_TrailingBits___64_comb};
  assign p2_prod__27_comb = {{7{p1_concat_135088[24]}}, p1_concat_135088};
  assign p2_prod__28_comb = {{7{p1_concat_135089[24]}}, p1_concat_135089};
  assign p2_concat_136908_comb = {p1_smul_57594_NarrowedMult_, p2_smul_57330_TrailingBits___67_comb};
  assign p2_concat_136909_comb = {p1_smul_57600_NarrowedMult_, p2_smul_57330_TrailingBits___68_comb};
  assign p2_prod__88_comb = {{7{p1_concat_135092[24]}}, p1_concat_135092};
  assign p2_prod__95_comb = {{7{p1_concat_135093[24]}}, p1_concat_135093};
  assign p2_concat_136914_comb = {p1_smul_57610_NarrowedMult_, p2_smul_57330_TrailingBits___71_comb};
  assign p2_concat_136919_comb = {p1_smul_57680_NarrowedMult_, p2_smul_57330_TrailingBits___88_comb};
  assign p2_prod__408_comb = {{7{p1_concat_135108[24]}}, p1_concat_135108};
  assign p2_prod__415_comb = {{7{p1_concat_135109[24]}}, p1_concat_135109};
  assign p2_concat_136924_comb = {p1_smul_57690_NarrowedMult_, p2_smul_57330_TrailingBits___91_comb};
  assign p2_concat_136925_comb = {p1_smul_57696_NarrowedMult_, p2_smul_57330_TrailingBits___92_comb};
  assign p2_prod__472_comb = {{7{p1_concat_135112[24]}}, p1_concat_135112};
  assign p2_prod__479_comb = {{7{p1_concat_135113[24]}}, p1_concat_135113};
  assign p2_concat_136930_comb = {p1_smul_57706_NarrowedMult_, p2_smul_57330_TrailingBits___95_comb};
  assign p2_prod__40_comb = {{7{p1_concat_135115[24]}}, p1_concat_135115};
  assign p2_concat_136933_comb = {p1_smul_57842_NarrowedMult_, p2_smul_57330_TrailingBits___97_comb};
  assign p2_concat_136934_comb = {p1_smul_57848_NarrowedMult_, p2_smul_57330_TrailingBits___98_comb};
  assign p2_prod__47_comb = {{7{p1_concat_135118[24]}}, p1_concat_135118};
  assign p2_prod__84_comb = {{7{p1_concat_135119[24]}}, p1_concat_135119};
  assign p2_concat_136939_comb = {p1_smul_57858_NarrowedMult_, p2_smul_57330_TrailingBits___101_comb};
  assign p2_concat_136940_comb = {p1_smul_57864_NarrowedMult_, p2_smul_57330_TrailingBits___102_comb};
  assign p2_prod__122_comb = {{7{p1_concat_135122[24]}}, p1_concat_135122};
  assign p2_prod__404_comb = {{7{p1_concat_135135[24]}}, p1_concat_135135};
  assign p2_concat_136949_comb = {p1_smul_57938_NarrowedMult_, p2_smul_57330_TrailingBits___121_comb};
  assign p2_concat_136950_comb = {p1_smul_57944_NarrowedMult_, p2_smul_57330_TrailingBits___122_comb};
  assign p2_prod__442_comb = {{7{p1_concat_135138[24]}}, p1_concat_135138};
  assign p2_prod__468_comb = {{7{p1_concat_135139[24]}}, p1_concat_135139};
  assign p2_concat_136955_comb = {p1_smul_57954_NarrowedMult_, p2_smul_57330_TrailingBits___125_comb};
  assign p2_concat_136956_comb = {p1_smul_57960_NarrowedMult_, p2_smul_57330_TrailingBits___126_comb};
  assign p2_prod__506_comb = {{7{p1_concat_135142[24]}}, p1_concat_135142};
  assign p2_prod__48_comb = {{8{p1_concat_135143[23]}}, p1_concat_135143};
  assign p2_prod__49_comb = {{7{p1_concat_135144[24]}}, p1_concat_135144};
  assign p2_prod__50_comb = {{8{p1_concat_135145[23]}}, p1_concat_135145};
  assign p2_prod__51_comb = {{7{p1_concat_135146[24]}}, p1_concat_135146};
  assign p2_prod__52_comb = {{7{p1_concat_135147[24]}}, p1_concat_135147};
  assign p2_prod__53_comb = {{8{p1_concat_135148[23]}}, p1_concat_135148};
  assign p2_prod__54_comb = {{7{p1_concat_135149[24]}}, p1_concat_135149};
  assign p2_prod__55_comb = {{8{p1_concat_135150[23]}}, p1_concat_135150};
  assign p2_prod__91_comb = {{8{p1_concat_135151[23]}}, p1_concat_135151};
  assign p2_prod__98_comb = {{7{p1_concat_135152[24]}}, p1_concat_135152};
  assign p2_prod__105_comb = {{8{p1_concat_135153[23]}}, p1_concat_135153};
  assign p2_prod__111_comb = {{7{p1_concat_135154[24]}}, p1_concat_135154};
  assign p2_prod__116_comb = {{7{p1_concat_135155[24]}}, p1_concat_135155};
  assign p2_prod__120_comb = {{8{p1_concat_135156[23]}}, p1_concat_135156};
  assign p2_prod__123_comb = {{7{p1_concat_135157[24]}}, p1_concat_135157};
  assign p2_prod__125_comb = {{8{p1_concat_135158[23]}}, p1_concat_135158};
  assign p2_prod__219_comb = {{8{p1_concat_135159[23]}}, p1_concat_135159};
  assign p2_prod__226_comb = {{7{p1_concat_135160[24]}}, p1_concat_135160};
  assign p2_prod__233_comb = {{8{p1_concat_135161[23]}}, p1_concat_135161};
  assign p2_prod__239_comb = {{7{p1_concat_135162[24]}}, p1_concat_135162};
  assign p2_prod__244_comb = {{7{p1_concat_135163[24]}}, p1_concat_135163};
  assign p2_prod__248_comb = {{8{p1_concat_135164[23]}}, p1_concat_135164};
  assign p2_prod__251_comb = {{7{p1_concat_135165[24]}}, p1_concat_135165};
  assign p2_prod__253_comb = {{8{p1_concat_135166[23]}}, p1_concat_135166};
  assign p2_prod__283_comb = {{8{p1_concat_135167[23]}}, p1_concat_135167};
  assign p2_prod__290_comb = {{7{p1_concat_135168[24]}}, p1_concat_135168};
  assign p2_prod__297_comb = {{8{p1_concat_135169[23]}}, p1_concat_135169};
  assign p2_prod__303_comb = {{7{p1_concat_135170[24]}}, p1_concat_135170};
  assign p2_prod__308_comb = {{7{p1_concat_135171[24]}}, p1_concat_135171};
  assign p2_prod__312_comb = {{8{p1_concat_135172[23]}}, p1_concat_135172};
  assign p2_prod__315_comb = {{7{p1_concat_135173[24]}}, p1_concat_135173};
  assign p2_prod__317_comb = {{8{p1_concat_135174[23]}}, p1_concat_135174};
  assign p2_prod__411_comb = {{8{p1_concat_135175[23]}}, p1_concat_135175};
  assign p2_prod__418_comb = {{7{p1_concat_135176[24]}}, p1_concat_135176};
  assign p2_prod__425_comb = {{8{p1_concat_135177[23]}}, p1_concat_135177};
  assign p2_prod__431_comb = {{7{p1_concat_135178[24]}}, p1_concat_135178};
  assign p2_prod__436_comb = {{7{p1_concat_135179[24]}}, p1_concat_135179};
  assign p2_prod__440_comb = {{8{p1_concat_135180[23]}}, p1_concat_135180};
  assign p2_prod__443_comb = {{7{p1_concat_135181[24]}}, p1_concat_135181};
  assign p2_prod__445_comb = {{8{p1_concat_135182[23]}}, p1_concat_135182};
  assign p2_prod__475_comb = {{8{p1_concat_135183[23]}}, p1_concat_135183};
  assign p2_prod__482_comb = {{7{p1_concat_135184[24]}}, p1_concat_135184};
  assign p2_prod__489_comb = {{8{p1_concat_135185[23]}}, p1_concat_135185};
  assign p2_prod__495_comb = {{7{p1_concat_135186[24]}}, p1_concat_135186};
  assign p2_prod__500_comb = {{7{p1_concat_135187[24]}}, p1_concat_135187};
  assign p2_prod__504_comb = {{8{p1_concat_135188[23]}}, p1_concat_135188};
  assign p2_prod__507_comb = {{7{p1_concat_135189[24]}}, p1_concat_135189};
  assign p2_prod__509_comb = {{8{p1_concat_135190[23]}}, p1_concat_135190};
  assign p2_concat_137031_comb = {p1_smul_58094_NarrowedMult_, p2_smul_57330_TrailingBits___160_comb};
  assign p2_prod__57_comb = {{7{p1_concat_135192[24]}}, p1_concat_135192};
  assign p2_prod__62_comb = {{7{p1_concat_135193[24]}}, p1_concat_135193};
  assign p2_concat_137036_comb = {p1_smul_58108_NarrowedMult_, p2_smul_57330_TrailingBits___163_comb};
  assign p2_concat_137037_comb = {p1_smul_58110_NarrowedMult_, p2_smul_57330_TrailingBits___164_comb};
  assign p2_prod__106_comb = {{7{p1_concat_135196[24]}}, p1_concat_135196};
  assign p2_prod__126_comb = {{7{p1_concat_135197[24]}}, p1_concat_135197};
  assign p2_concat_137042_comb = {p1_smul_58124_NarrowedMult_, p2_smul_57330_TrailingBits___167_comb};
  assign p2_concat_137047_comb = {p1_smul_58190_NarrowedMult_, p2_smul_57330_TrailingBits___184_comb};
  assign p2_prod__426_comb = {{7{p1_concat_135212[24]}}, p1_concat_135212};
  assign p2_prod__446_comb = {{7{p1_concat_135213[24]}}, p1_concat_135213};
  assign p2_concat_137052_comb = {p1_smul_58204_NarrowedMult_, p2_smul_57330_TrailingBits___187_comb};
  assign p2_concat_137053_comb = {p1_smul_58206_NarrowedMult_, p2_smul_57330_TrailingBits___188_comb};
  assign p2_prod__490_comb = {{7{p1_concat_135216[24]}}, p1_concat_135216};
  assign p2_prod__510_comb = {{7{p1_concat_135217[24]}}, p1_concat_135217};
  assign p2_concat_137058_comb = {p1_smul_58220_NarrowedMult_, p2_smul_57330_TrailingBits___191_comb};
  assign p2_smul_57326_TrailingBits___16_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___17_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___18_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___19_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___20_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___21_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___22_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___23_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___40_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___41_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___42_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___43_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___44_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___45_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___46_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___47_comb = 8'h00;
  assign p2_smul_57326_TrailingBits__comb = 8'h00;
  assign p2_smul_57326_TrailingBits___1_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___2_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___3_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___4_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___5_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___6_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___7_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___8_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___9_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___10_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___11_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___12_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___13_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___14_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___15_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___24_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___25_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___26_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___27_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___28_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___29_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___30_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___31_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___32_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___33_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___34_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___35_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___36_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___37_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___38_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___39_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___48_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___49_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___50_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___51_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___52_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___53_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___54_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___55_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___56_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___57_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___58_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___59_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___60_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___61_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___62_comb = 8'h00;
  assign p2_smul_57326_TrailingBits___63_comb = 8'h00;
  assign p2_or_137427_comb = p1_prod__199 | 32'h0000_0080;
  assign p2_prod__203_comb = {{9{p1_concat_135348[22]}}, p1_concat_135348};
  assign p2_prod__208_comb = {{9{p1_concat_135349[22]}}, p1_concat_135349};
  assign p2_or_137434_comb = p1_prod__214 | 32'h0000_0080;
  assign p2_or_137441_comb = p1_prod__263 | 32'h0000_0080;
  assign p2_prod__267_comb = {{9{p1_concat_135352[22]}}, p1_concat_135352};
  assign p2_prod__272_comb = {{9{p1_concat_135353[22]}}, p1_concat_135353};
  assign p2_or_137448_comb = p1_prod__278 | 32'h0000_0080;
  assign p2_prod__205_comb = {{9{p1_concat_135355[22]}}, p1_concat_135355};
  assign p2_or_137633_comb = p1_prod__216 | 32'h0000_0080;
  assign p2_or_137636_comb = p1_prod__223 | 32'h0000_0080;
  assign p2_prod__236_comb = {{9{p1_concat_135358[22]}}, p1_concat_135358};
  assign p2_prod__269_comb = {{9{p1_concat_135359[22]}}, p1_concat_135359};
  assign p2_or_137647_comb = p1_prod__280 | 32'h0000_0080;
  assign p2_or_137650_comb = p1_prod__287 | 32'h0000_0080;
  assign p2_prod__300_comb = {{9{p1_concat_135362[22]}}, p1_concat_135362};
  assign p2_or_137761_comb = p1_prod__212 | 32'h0000_0080;
  assign p2_prod__225_comb = {{9{p1_concat_135364[22]}}, p1_concat_135364};
  assign p2_prod__243_comb = {{9{p1_concat_135365[22]}}, p1_concat_135365};
  assign p2_or_137772_comb = p1_prod__250 | 32'h0000_0080;
  assign p2_or_137775_comb = p1_prod__276 | 32'h0000_0080;
  assign p2_prod__289_comb = {{9{p1_concat_135368[22]}}, p1_concat_135368};
  assign p2_prod__307_comb = {{9{p1_concat_135369[22]}}, p1_concat_135369};
  assign p2_or_137786_comb = p1_prod__314 | 32'h0000_0080;
  assign p2_prod__227_comb = {{9{p1_concat_135371[22]}}, p1_concat_135371};
  assign p2_or_137967_comb = p1_prod__234 | 32'h0000_0080;
  assign p2_or_137974_comb = p1_prod__254 | 32'h0000_0080;
  assign p2_prod__255_comb = {{9{p1_concat_135374[22]}}, p1_concat_135374};
  assign p2_prod__291_comb = {{9{p1_concat_135375[22]}}, p1_concat_135375};
  assign p2_or_137981_comb = p1_prod__298 | 32'h0000_0080;
  assign p2_or_137988_comb = p1_prod__318 | 32'h0000_0080;
  assign p2_prod__319_comb = {{9{p1_concat_135378[22]}}, p1_concat_135378};
  assign p2_smul_57742_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__16_squeezed, 9'h0b5);
  assign p2_smul_57744_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__17_squeezed, 9'h14b);
  assign p2_smul_57746_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__18_squeezed, 9'h14b);
  assign p2_smul_57748_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__19_squeezed, 9'h0b5);
  assign p2_smul_57750_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__20_squeezed, 9'h0b5);
  assign p2_smul_57752_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__21_squeezed, 9'h14b);
  assign p2_smul_57754_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__22_squeezed, 9'h14b);
  assign p2_smul_57756_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__23_squeezed, 9'h0b5);
  assign p2_smul_57790_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__40_squeezed, 9'h0b5);
  assign p2_smul_57792_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__41_squeezed, 9'h14b);
  assign p2_smul_57794_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__42_squeezed, 9'h14b);
  assign p2_smul_57796_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__43_squeezed, 9'h0b5);
  assign p2_smul_57798_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__44_squeezed, 9'h0b5);
  assign p2_smul_57800_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__45_squeezed, 9'h14b);
  assign p2_smul_57802_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__46_squeezed, 9'h14b);
  assign p2_smul_57804_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__47_squeezed, 9'h0b5);
  assign p2_smul_57710_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted_squeezed, 9'h0b5);
  assign p2_smul_57712_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__1_squeezed, 9'h14b);
  assign p2_smul_57714_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__2_squeezed, 9'h14b);
  assign p2_smul_57716_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__3_squeezed, 9'h0b5);
  assign p2_smul_57718_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__4_squeezed, 9'h0b5);
  assign p2_smul_57720_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__5_squeezed, 9'h14b);
  assign p2_smul_57722_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__6_squeezed, 9'h14b);
  assign p2_smul_57724_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__7_squeezed, 9'h0b5);
  assign p2_smul_57726_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__8_squeezed, 9'h0b5);
  assign p2_smul_57728_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__9_squeezed, 9'h14b);
  assign p2_smul_57730_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__10_squeezed, 9'h14b);
  assign p2_smul_57732_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__11_squeezed, 9'h0b5);
  assign p2_smul_57734_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__12_squeezed, 9'h0b5);
  assign p2_smul_57736_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__13_squeezed, 9'h14b);
  assign p2_smul_57738_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__14_squeezed, 9'h14b);
  assign p2_smul_57740_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__15_squeezed, 9'h0b5);
  assign p2_smul_57758_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__24_squeezed, 9'h0b5);
  assign p2_smul_57760_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__25_squeezed, 9'h14b);
  assign p2_smul_57762_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__26_squeezed, 9'h14b);
  assign p2_smul_57764_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__27_squeezed, 9'h0b5);
  assign p2_smul_57766_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__28_squeezed, 9'h0b5);
  assign p2_smul_57768_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__29_squeezed, 9'h14b);
  assign p2_smul_57770_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__30_squeezed, 9'h14b);
  assign p2_smul_57772_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__31_squeezed, 9'h0b5);
  assign p2_smul_57774_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__32_squeezed, 9'h0b5);
  assign p2_smul_57776_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__33_squeezed, 9'h14b);
  assign p2_smul_57778_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__34_squeezed, 9'h14b);
  assign p2_smul_57780_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__35_squeezed, 9'h0b5);
  assign p2_smul_57782_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__36_squeezed, 9'h0b5);
  assign p2_smul_57784_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__37_squeezed, 9'h14b);
  assign p2_smul_57786_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__38_squeezed, 9'h14b);
  assign p2_smul_57788_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__39_squeezed, 9'h0b5);
  assign p2_smul_57806_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__48_squeezed, 9'h0b5);
  assign p2_smul_57808_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__49_squeezed, 9'h14b);
  assign p2_smul_57810_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__50_squeezed, 9'h14b);
  assign p2_smul_57812_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__51_squeezed, 9'h0b5);
  assign p2_smul_57814_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__52_squeezed, 9'h0b5);
  assign p2_smul_57816_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__53_squeezed, 9'h14b);
  assign p2_smul_57818_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__54_squeezed, 9'h14b);
  assign p2_smul_57820_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__55_squeezed, 9'h0b5);
  assign p2_smul_57822_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__56_squeezed, 9'h0b5);
  assign p2_smul_57824_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__57_squeezed, 9'h14b);
  assign p2_smul_57826_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__58_squeezed, 9'h14b);
  assign p2_smul_57828_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__59_squeezed, 9'h0b5);
  assign p2_smul_57830_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__60_squeezed, 9'h0b5);
  assign p2_smul_57832_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__61_squeezed, 9'h14b);
  assign p2_smul_57834_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__62_squeezed, 9'h14b);
  assign p2_smul_57836_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__63_squeezed, 9'h0b5);
  assign p2_or_137095_comb = p2_prod__135_comb | 32'h0000_0080;
  assign p2_prod__139_comb = {{9{p2_concat_136661_comb[22]}}, p2_concat_136661_comb};
  assign p2_prod__144_comb = {{9{p2_concat_136662_comb[22]}}, p2_concat_136662_comb};
  assign p2_or_137102_comb = p2_prod__150_comb | 32'h0000_0080;
  assign p2_or_137109_comb = p2_prod__327_comb | 32'h0000_0080;
  assign p2_prod__331_comb = {{9{p2_concat_136667_comb[22]}}, p2_concat_136667_comb};
  assign p2_prod__336_comb = {{9{p2_concat_136668_comb[22]}}, p2_concat_136668_comb};
  assign p2_or_137116_comb = p2_prod__342_comb | 32'h0000_0080;
  assign p2_or_137121_comb = p2_prod__133_comb | 32'h0000_0080;
  assign p2_or_137128_comb = p2_prod__145_comb | 32'h0000_0080;
  assign p2_or_137131_comb = p2_prod__151_comb | 32'h0000_0080;
  assign p2_or_137138_comb = p2_prod__171_comb | 32'h0000_0080;
  assign p2_or_137141_comb = p2_prod__325_comb | 32'h0000_0080;
  assign p2_or_137148_comb = p2_prod__337_comb | 32'h0000_0080;
  assign p2_or_137151_comb = p2_prod__343_comb | 32'h0000_0080;
  assign p2_or_137158_comb = p2_prod__363_comb | 32'h0000_0080;
  assign p2_prod__141_comb = {{9{p2_concat_136695_comb[22]}}, p2_concat_136695_comb};
  assign p2_or_137165_comb = p2_prod__152_comb | 32'h0000_0080;
  assign p2_or_137168_comb = p2_prod__159_comb | 32'h0000_0080;
  assign p2_prod__172_comb = {{9{p2_concat_136700_comb[22]}}, p2_concat_136700_comb};
  assign p2_prod__333_comb = {{9{p2_concat_136701_comb[22]}}, p2_concat_136701_comb};
  assign p2_or_137179_comb = p2_prod__344_comb | 32'h0000_0080;
  assign p2_or_137182_comb = p2_prod__351_comb | 32'h0000_0080;
  assign p2_prod__364_comb = {{9{p2_concat_136706_comb[22]}}, p2_concat_136706_comb};
  assign p2_or_137205_comb = p2_prod__148_comb | 32'h0000_0080;
  assign p2_prod__161_comb = {{9{p2_concat_136709_comb[22]}}, p2_concat_136709_comb};
  assign p2_prod__179_comb = {{9{p2_concat_136710_comb[22]}}, p2_concat_136710_comb};
  assign p2_or_137216_comb = p2_prod__186_comb | 32'h0000_0080;
  assign p2_or_137219_comb = p2_prod__340_comb | 32'h0000_0080;
  assign p2_prod__353_comb = {{9{p2_concat_136715_comb[22]}}, p2_concat_136715_comb};
  assign p2_prod__371_comb = {{9{p2_concat_136716_comb[22]}}, p2_concat_136716_comb};
  assign p2_or_137230_comb = p2_prod__378_comb | 32'h0000_0080;
  assign p2_or_137235_comb = p2_prod__162_comb | 32'h0000_0080;
  assign p2_or_137240_comb = p2_prod__175_comb | 32'h0000_0080;
  assign p2_or_137243_comb = p2_prod__180_comb | 32'h0000_0080;
  assign p2_or_137248_comb = p2_prod__187_comb | 32'h0000_0080;
  assign p2_or_137255_comb = p2_prod__354_comb | 32'h0000_0080;
  assign p2_or_137260_comb = p2_prod__367_comb | 32'h0000_0080;
  assign p2_or_137263_comb = p2_prod__372_comb | 32'h0000_0080;
  assign p2_or_137268_comb = p2_prod__379_comb | 32'h0000_0080;
  assign p2_prod__163_comb = {{9{p2_concat_136743_comb[22]}}, p2_concat_136743_comb};
  assign p2_or_137275_comb = p2_prod__170_comb | 32'h0000_0080;
  assign p2_or_137282_comb = p2_prod__190_comb | 32'h0000_0080;
  assign p2_prod__191_comb = {{9{p2_concat_136748_comb[22]}}, p2_concat_136748_comb};
  assign p2_prod__355_comb = {{9{p2_concat_136749_comb[22]}}, p2_concat_136749_comb};
  assign p2_or_137289_comb = p2_prod__362_comb | 32'h0000_0080;
  assign p2_or_137296_comb = p2_prod__382_comb | 32'h0000_0080;
  assign p2_prod__383_comb = {{9{p2_concat_136754_comb[22]}}, p2_concat_136754_comb};
  assign p2_or_137399_comb = p2_prod__10_comb | 32'h0000_0080;
  assign p2_prod__11_comb = {{9{p2_concat_136805_comb[22]}}, p2_concat_136805_comb};
  assign p2_prod__12_comb = {{9{p2_concat_136806_comb[22]}}, p2_concat_136806_comb};
  assign p2_or_137406_comb = p2_prod__13_comb | 32'h0000_0080;
  assign p2_or_137413_comb = p2_prod__71_comb | 32'h0000_0080;
  assign p2_prod__75_comb = {{9{p2_concat_136811_comb[22]}}, p2_concat_136811_comb};
  assign p2_prod__80_comb = {{9{p2_concat_136812_comb[22]}}, p2_concat_136812_comb};
  assign p2_or_137420_comb = p2_prod__86_comb | 32'h0000_0080;
  assign p2_or_137455_comb = p2_prod__391_comb | 32'h0000_0080;
  assign p2_prod__395_comb = {{9{p2_concat_136821_comb[22]}}, p2_concat_136821_comb};
  assign p2_prod__400_comb = {{9{p2_concat_136822_comb[22]}}, p2_concat_136822_comb};
  assign p2_or_137462_comb = p2_prod__406_comb | 32'h0000_0080;
  assign p2_or_137469_comb = p2_prod__455_comb | 32'h0000_0080;
  assign p2_prod__459_comb = {{9{p2_concat_136827_comb[22]}}, p2_concat_136827_comb};
  assign p2_prod__464_comb = {{9{p2_concat_136828_comb[22]}}, p2_concat_136828_comb};
  assign p2_or_137476_comb = p2_prod__470_comb | 32'h0000_0080;
  assign p2_or_137481_comb = p2_prod__16_comb | 32'h0000_0080;
  assign p2_or_137488_comb = p2_prod__19_comb | 32'h0000_0080;
  assign p2_or_137491_comb = p2_prod__20_comb | 32'h0000_0080;
  assign p2_or_137498_comb = p2_prod__23_comb | 32'h0000_0080;
  assign p2_or_137501_comb = p2_prod__69_comb | 32'h0000_0080;
  assign p2_or_137508_comb = p2_prod__81_comb | 32'h0000_0080;
  assign p2_or_137511_comb = p2_prod__87_comb | 32'h0000_0080;
  assign p2_or_137518_comb = p2_prod__107_comb | 32'h0000_0080;
  assign p2_or_137521_comb = p2_prod__197_comb | 32'h0000_0080;
  assign p2_or_137528_comb = p2_prod__209_comb | 32'h0000_0080;
  assign p2_or_137531_comb = p2_prod__215_comb | 32'h0000_0080;
  assign p2_or_137538_comb = p2_prod__235_comb | 32'h0000_0080;
  assign p2_or_137541_comb = p2_prod__261_comb | 32'h0000_0080;
  assign p2_or_137548_comb = p2_prod__273_comb | 32'h0000_0080;
  assign p2_or_137551_comb = p2_prod__279_comb | 32'h0000_0080;
  assign p2_or_137558_comb = p2_prod__299_comb | 32'h0000_0080;
  assign p2_or_137561_comb = p2_prod__389_comb | 32'h0000_0080;
  assign p2_or_137568_comb = p2_prod__401_comb | 32'h0000_0080;
  assign p2_or_137571_comb = p2_prod__407_comb | 32'h0000_0080;
  assign p2_or_137578_comb = p2_prod__427_comb | 32'h0000_0080;
  assign p2_or_137581_comb = p2_prod__453_comb | 32'h0000_0080;
  assign p2_or_137588_comb = p2_prod__465_comb | 32'h0000_0080;
  assign p2_or_137591_comb = p2_prod__471_comb | 32'h0000_0080;
  assign p2_or_137598_comb = p2_prod__491_comb | 32'h0000_0080;
  assign p2_prod__25_comb = {{9{p2_concat_136903_comb[22]}}, p2_concat_136903_comb};
  assign p2_or_137605_comb = p2_prod__27_comb | 32'h0000_0080;
  assign p2_or_137608_comb = p2_prod__28_comb | 32'h0000_0080;
  assign p2_prod__30_comb = {{9{p2_concat_136908_comb[22]}}, p2_concat_136908_comb};
  assign p2_prod__77_comb = {{9{p2_concat_136909_comb[22]}}, p2_concat_136909_comb};
  assign p2_or_137619_comb = p2_prod__88_comb | 32'h0000_0080;
  assign p2_or_137622_comb = p2_prod__95_comb | 32'h0000_0080;
  assign p2_prod__108_comb = {{9{p2_concat_136914_comb[22]}}, p2_concat_136914_comb};
  assign p2_prod__397_comb = {{9{p2_concat_136919_comb[22]}}, p2_concat_136919_comb};
  assign p2_or_137661_comb = p2_prod__408_comb | 32'h0000_0080;
  assign p2_or_137664_comb = p2_prod__415_comb | 32'h0000_0080;
  assign p2_prod__428_comb = {{9{p2_concat_136924_comb[22]}}, p2_concat_136924_comb};
  assign p2_prod__461_comb = {{9{p2_concat_136925_comb[22]}}, p2_concat_136925_comb};
  assign p2_or_137675_comb = p2_prod__472_comb | 32'h0000_0080;
  assign p2_or_137678_comb = p2_prod__479_comb | 32'h0000_0080;
  assign p2_prod__492_comb = {{9{p2_concat_136930_comb[22]}}, p2_concat_136930_comb};
  assign p2_or_137733_comb = p2_prod__40_comb | 32'h0000_0080;
  assign p2_prod__42_comb = {{9{p2_concat_136933_comb[22]}}, p2_concat_136933_comb};
  assign p2_prod__45_comb = {{9{p2_concat_136934_comb[22]}}, p2_concat_136934_comb};
  assign p2_or_137744_comb = p2_prod__47_comb | 32'h0000_0080;
  assign p2_or_137747_comb = p2_prod__84_comb | 32'h0000_0080;
  assign p2_prod__97_comb = {{9{p2_concat_136939_comb[22]}}, p2_concat_136939_comb};
  assign p2_prod__115_comb = {{9{p2_concat_136940_comb[22]}}, p2_concat_136940_comb};
  assign p2_or_137758_comb = p2_prod__122_comb | 32'h0000_0080;
  assign p2_or_137789_comb = p2_prod__404_comb | 32'h0000_0080;
  assign p2_prod__417_comb = {{9{p2_concat_136949_comb[22]}}, p2_concat_136949_comb};
  assign p2_prod__435_comb = {{9{p2_concat_136950_comb[22]}}, p2_concat_136950_comb};
  assign p2_or_137800_comb = p2_prod__442_comb | 32'h0000_0080;
  assign p2_or_137803_comb = p2_prod__468_comb | 32'h0000_0080;
  assign p2_prod__481_comb = {{9{p2_concat_136955_comb[22]}}, p2_concat_136955_comb};
  assign p2_prod__499_comb = {{9{p2_concat_136956_comb[22]}}, p2_concat_136956_comb};
  assign p2_or_137814_comb = p2_prod__506_comb | 32'h0000_0080;
  assign p2_or_137819_comb = p2_prod__49_comb | 32'h0000_0080;
  assign p2_or_137824_comb = p2_prod__51_comb | 32'h0000_0080;
  assign p2_or_137827_comb = p2_prod__52_comb | 32'h0000_0080;
  assign p2_or_137832_comb = p2_prod__54_comb | 32'h0000_0080;
  assign p2_or_137839_comb = p2_prod__98_comb | 32'h0000_0080;
  assign p2_or_137844_comb = p2_prod__111_comb | 32'h0000_0080;
  assign p2_or_137847_comb = p2_prod__116_comb | 32'h0000_0080;
  assign p2_or_137852_comb = p2_prod__123_comb | 32'h0000_0080;
  assign p2_or_137859_comb = p2_prod__226_comb | 32'h0000_0080;
  assign p2_or_137864_comb = p2_prod__239_comb | 32'h0000_0080;
  assign p2_or_137867_comb = p2_prod__244_comb | 32'h0000_0080;
  assign p2_or_137872_comb = p2_prod__251_comb | 32'h0000_0080;
  assign p2_or_137879_comb = p2_prod__290_comb | 32'h0000_0080;
  assign p2_or_137884_comb = p2_prod__303_comb | 32'h0000_0080;
  assign p2_or_137887_comb = p2_prod__308_comb | 32'h0000_0080;
  assign p2_or_137892_comb = p2_prod__315_comb | 32'h0000_0080;
  assign p2_or_137899_comb = p2_prod__418_comb | 32'h0000_0080;
  assign p2_or_137904_comb = p2_prod__431_comb | 32'h0000_0080;
  assign p2_or_137907_comb = p2_prod__436_comb | 32'h0000_0080;
  assign p2_or_137912_comb = p2_prod__443_comb | 32'h0000_0080;
  assign p2_or_137919_comb = p2_prod__482_comb | 32'h0000_0080;
  assign p2_or_137924_comb = p2_prod__495_comb | 32'h0000_0080;
  assign p2_or_137927_comb = p2_prod__500_comb | 32'h0000_0080;
  assign p2_or_137932_comb = p2_prod__507_comb | 32'h0000_0080;
  assign p2_prod__56_comb = {{9{p2_concat_137031_comb[22]}}, p2_concat_137031_comb};
  assign p2_or_137939_comb = p2_prod__57_comb | 32'h0000_0080;
  assign p2_or_137946_comb = p2_prod__62_comb | 32'h0000_0080;
  assign p2_prod__63_comb = {{9{p2_concat_137036_comb[22]}}, p2_concat_137036_comb};
  assign p2_prod__99_comb = {{9{p2_concat_137037_comb[22]}}, p2_concat_137037_comb};
  assign p2_or_137953_comb = p2_prod__106_comb | 32'h0000_0080;
  assign p2_or_137960_comb = p2_prod__126_comb | 32'h0000_0080;
  assign p2_prod__127_comb = {{9{p2_concat_137042_comb[22]}}, p2_concat_137042_comb};
  assign p2_prod__419_comb = {{9{p2_concat_137047_comb[22]}}, p2_concat_137047_comb};
  assign p2_or_137995_comb = p2_prod__426_comb | 32'h0000_0080;
  assign p2_or_138002_comb = p2_prod__446_comb | 32'h0000_0080;
  assign p2_prod__447_comb = {{9{p2_concat_137052_comb[22]}}, p2_concat_137052_comb};
  assign p2_prod__483_comb = {{9{p2_concat_137053_comb[22]}}, p2_concat_137053_comb};
  assign p2_or_138009_comb = p2_prod__490_comb | 32'h0000_0080;
  assign p2_or_138016_comb = p2_prod__510_comb | 32'h0000_0080;
  assign p2_prod__511_comb = {{9{p2_concat_137058_comb[22]}}, p2_concat_137058_comb};
  assign p2_smul_57374_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__24_squeezed, 9'h0fb);
  assign p2_smul_57376_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__25_squeezed, 9'h0d5);
  assign p2_or_138426_comb = p2_prod__203_comb | 32'h0000_0080;
  assign p2_or_138427_comb = p2_prod__208_comb | 32'h0000_0080;
  assign p2_smul_57386_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__30_squeezed, 9'h12b);
  assign p2_smul_57388_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__31_squeezed, 9'h105);
  assign p2_smul_57390_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__32_squeezed, 9'h0fb);
  assign p2_smul_57392_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__33_squeezed, 9'h0d5);
  assign p2_or_138442_comb = p2_prod__267_comb | 32'h0000_0080;
  assign p2_or_138443_comb = p2_prod__272_comb | 32'h0000_0080;
  assign p2_smul_57402_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__38_squeezed, 9'h12b);
  assign p2_smul_57404_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__39_squeezed, 9'h105);
  assign p2_smul_57630_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__24_squeezed, 9'h0d5);
  assign p2_or_138637_comb = p2_prod__205_comb | 32'h0000_0080;
  assign p2_smul_57634_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__26_squeezed, 9'h105);
  assign p2_smul_57640_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__29_squeezed, 9'h0fb);
  assign p2_or_138648_comb = p2_prod__236_comb | 32'h0000_0080;
  assign p2_smul_57644_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__31_squeezed, 9'h12b);
  assign p2_smul_57646_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__32_squeezed, 9'h0d5);
  assign p2_or_138653_comb = p2_prod__269_comb | 32'h0000_0080;
  assign p2_smul_57650_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__34_squeezed, 9'h105);
  assign p2_smul_57656_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__37_squeezed, 9'h0fb);
  assign p2_or_138664_comb = p2_prod__300_comb | 32'h0000_0080;
  assign p2_smul_57660_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__39_squeezed, 9'h12b);
  assign p2_smul_57888_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__25_squeezed, 9'h105);
  assign p2_or_138832_comb = p2_prod__225_comb | 32'h0000_0080;
  assign p2_smul_57892_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__27_squeezed, 9'h0d5);
  assign p2_smul_57894_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__28_squeezed, 9'h0d5);
  assign p2_or_138837_comb = p2_prod__243_comb | 32'h0000_0080;
  assign p2_smul_57898_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__30_squeezed, 9'h105);
  assign p2_smul_57904_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__33_squeezed, 9'h105);
  assign p2_or_138848_comb = p2_prod__289_comb | 32'h0000_0080;
  assign p2_smul_57908_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__35_squeezed, 9'h0d5);
  assign p2_smul_57910_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__36_squeezed, 9'h0d5);
  assign p2_or_138853_comb = p2_prod__307_comb | 32'h0000_0080;
  assign p2_smul_57914_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__38_squeezed, 9'h105);
  assign p2_or_139043_comb = p2_prod__227_comb | 32'h0000_0080;
  assign p2_smul_58146_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__26_squeezed, 9'h0d5);
  assign p2_smul_58148_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__27_squeezed, 9'h105);
  assign p2_smul_58150_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__28_squeezed, 9'h105);
  assign p2_smul_58152_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__29_squeezed, 9'h0d5);
  assign p2_or_139058_comb = p2_prod__255_comb | 32'h0000_0080;
  assign p2_or_139059_comb = p2_prod__291_comb | 32'h0000_0080;
  assign p2_smul_58162_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__34_squeezed, 9'h0d5);
  assign p2_smul_58164_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__35_squeezed, 9'h105);
  assign p2_smul_58166_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__36_squeezed, 9'h105);
  assign p2_smul_58168_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__37_squeezed, 9'h0d5);
  assign p2_or_139074_comb = p2_prod__319_comb | 32'h0000_0080;
  assign p2_smul_57358_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__16_squeezed, 9'h0fb);
  assign p2_smul_57360_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__17_squeezed, 9'h0d5);
  assign p2_or_138058_comb = p2_prod__139_comb | 32'h0000_0080;
  assign p2_or_138059_comb = p2_prod__144_comb | 32'h0000_0080;
  assign p2_smul_57370_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__22_squeezed, 9'h12b);
  assign p2_smul_57372_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__23_squeezed, 9'h105);
  assign p2_smul_57406_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__40_squeezed, 9'h0fb);
  assign p2_smul_57408_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__41_squeezed, 9'h0d5);
  assign p2_or_138074_comb = p2_prod__331_comb | 32'h0000_0080;
  assign p2_or_138075_comb = p2_prod__336_comb | 32'h0000_0080;
  assign p2_smul_57418_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__46_squeezed, 9'h12b);
  assign p2_smul_57420_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__47_squeezed, 9'h105);
  assign p2_smul_57614_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__16_squeezed, 9'h0d5);
  assign p2_or_138125_comb = p2_prod__141_comb | 32'h0000_0080;
  assign p2_smul_57618_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__18_squeezed, 9'h105);
  assign p2_smul_57624_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__21_squeezed, 9'h0fb);
  assign p2_or_138136_comb = p2_prod__172_comb | 32'h0000_0080;
  assign p2_smul_57628_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__23_squeezed, 9'h12b);
  assign p2_smul_57662_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__40_squeezed, 9'h0d5);
  assign p2_or_138141_comb = p2_prod__333_comb | 32'h0000_0080;
  assign p2_smul_57666_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__42_squeezed, 9'h105);
  assign p2_smul_57672_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__45_squeezed, 9'h0fb);
  assign p2_or_138152_comb = p2_prod__364_comb | 32'h0000_0080;
  assign p2_smul_57676_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__47_squeezed, 9'h12b);
  assign p2_smul_57872_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__17_squeezed, 9'h105);
  assign p2_or_138192_comb = p2_prod__161_comb | 32'h0000_0080;
  assign p2_smul_57876_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__19_squeezed, 9'h0d5);
  assign p2_smul_57878_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__20_squeezed, 9'h0d5);
  assign p2_or_138197_comb = p2_prod__179_comb | 32'h0000_0080;
  assign p2_smul_57882_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__22_squeezed, 9'h105);
  assign p2_smul_57920_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__41_squeezed, 9'h105);
  assign p2_or_138208_comb = p2_prod__353_comb | 32'h0000_0080;
  assign p2_smul_57924_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__43_squeezed, 9'h0d5);
  assign p2_smul_57926_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__44_squeezed, 9'h0d5);
  assign p2_or_138213_comb = p2_prod__371_comb | 32'h0000_0080;
  assign p2_smul_57930_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__46_squeezed, 9'h105);
  assign p2_or_138259_comb = p2_prod__163_comb | 32'h0000_0080;
  assign p2_smul_58130_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__18_squeezed, 9'h0d5);
  assign p2_smul_58132_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__19_squeezed, 9'h105);
  assign p2_smul_58134_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__20_squeezed, 9'h105);
  assign p2_smul_58136_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__21_squeezed, 9'h0d5);
  assign p2_or_138274_comb = p2_prod__191_comb | 32'h0000_0080;
  assign p2_or_138275_comb = p2_prod__355_comb | 32'h0000_0080;
  assign p2_smul_58178_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__42_squeezed, 9'h0d5);
  assign p2_smul_58180_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__43_squeezed, 9'h105);
  assign p2_smul_58182_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__44_squeezed, 9'h105);
  assign p2_smul_58184_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__45_squeezed, 9'h0d5);
  assign p2_or_138290_comb = p2_prod__383_comb | 32'h0000_0080;
  assign p2_smul_57326_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted_squeezed, 9'h0fb);
  assign p2_smul_57328_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__1_squeezed, 9'h0d5);
  assign p2_or_138394_comb = p2_prod__11_comb | 32'h0000_0080;
  assign p2_or_138395_comb = p2_prod__12_comb | 32'h0000_0080;
  assign p2_smul_57338_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__6_squeezed, 9'h12b);
  assign p2_smul_57340_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__7_squeezed, 9'h105);
  assign p2_smul_57342_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__8_squeezed, 9'h0fb);
  assign p2_smul_57344_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__9_squeezed, 9'h0d5);
  assign p2_or_138410_comb = p2_prod__75_comb | 32'h0000_0080;
  assign p2_or_138411_comb = p2_prod__80_comb | 32'h0000_0080;
  assign p2_smul_57354_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__14_squeezed, 9'h12b);
  assign p2_smul_57356_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__15_squeezed, 9'h105);
  assign p2_smul_57422_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__48_squeezed, 9'h0fb);
  assign p2_smul_57424_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__49_squeezed, 9'h0d5);
  assign p2_or_138458_comb = p2_prod__395_comb | 32'h0000_0080;
  assign p2_or_138459_comb = p2_prod__400_comb | 32'h0000_0080;
  assign p2_smul_57434_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__54_squeezed, 9'h12b);
  assign p2_smul_57436_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__55_squeezed, 9'h105);
  assign p2_smul_57438_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__56_squeezed, 9'h0fb);
  assign p2_smul_57440_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__57_squeezed, 9'h0d5);
  assign p2_or_138474_comb = p2_prod__459_comb | 32'h0000_0080;
  assign p2_or_138475_comb = p2_prod__464_comb | 32'h0000_0080;
  assign p2_smul_57450_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__62_squeezed, 9'h12b);
  assign p2_smul_57452_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__63_squeezed, 9'h105);
  assign p2_smul_57582_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted_squeezed, 9'h0d5);
  assign p2_or_138605_comb = p2_prod__25_comb | 32'h0000_0080;
  assign p2_smul_57586_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__2_squeezed, 9'h105);
  assign p2_smul_57592_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__5_squeezed, 9'h0fb);
  assign p2_or_138616_comb = p2_prod__30_comb | 32'h0000_0080;
  assign p2_smul_57596_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__7_squeezed, 9'h12b);
  assign p2_smul_57598_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__8_squeezed, 9'h0d5);
  assign p2_or_138621_comb = p2_prod__77_comb | 32'h0000_0080;
  assign p2_smul_57602_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__10_squeezed, 9'h105);
  assign p2_smul_57608_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__13_squeezed, 9'h0fb);
  assign p2_or_138632_comb = p2_prod__108_comb | 32'h0000_0080;
  assign p2_smul_57612_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__15_squeezed, 9'h12b);
  assign p2_smul_57678_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__48_squeezed, 9'h0d5);
  assign p2_or_138669_comb = p2_prod__397_comb | 32'h0000_0080;
  assign p2_smul_57682_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__50_squeezed, 9'h105);
  assign p2_smul_57688_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__53_squeezed, 9'h0fb);
  assign p2_or_138680_comb = p2_prod__428_comb | 32'h0000_0080;
  assign p2_smul_57692_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__55_squeezed, 9'h12b);
  assign p2_smul_57694_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__56_squeezed, 9'h0d5);
  assign p2_or_138685_comb = p2_prod__461_comb | 32'h0000_0080;
  assign p2_smul_57698_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__58_squeezed, 9'h105);
  assign p2_smul_57704_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__61_squeezed, 9'h0fb);
  assign p2_or_138696_comb = p2_prod__492_comb | 32'h0000_0080;
  assign p2_smul_57708_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__63_squeezed, 9'h12b);
  assign p2_smul_57840_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__1_squeezed, 9'h105);
  assign p2_or_138800_comb = p2_prod__42_comb | 32'h0000_0080;
  assign p2_smul_57844_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__3_squeezed, 9'h0d5);
  assign p2_smul_57846_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__4_squeezed, 9'h0d5);
  assign p2_or_138805_comb = p2_prod__45_comb | 32'h0000_0080;
  assign p2_smul_57850_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__6_squeezed, 9'h105);
  assign p2_smul_57856_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__9_squeezed, 9'h105);
  assign p2_or_138816_comb = p2_prod__97_comb | 32'h0000_0080;
  assign p2_smul_57860_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__11_squeezed, 9'h0d5);
  assign p2_smul_57862_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__12_squeezed, 9'h0d5);
  assign p2_or_138821_comb = p2_prod__115_comb | 32'h0000_0080;
  assign p2_smul_57866_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__14_squeezed, 9'h105);
  assign p2_smul_57936_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__49_squeezed, 9'h105);
  assign p2_or_138864_comb = p2_prod__417_comb | 32'h0000_0080;
  assign p2_smul_57940_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__51_squeezed, 9'h0d5);
  assign p2_smul_57942_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__52_squeezed, 9'h0d5);
  assign p2_or_138869_comb = p2_prod__435_comb | 32'h0000_0080;
  assign p2_smul_57946_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__54_squeezed, 9'h105);
  assign p2_smul_57952_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__57_squeezed, 9'h105);
  assign p2_or_138880_comb = p2_prod__481_comb | 32'h0000_0080;
  assign p2_smul_57956_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__59_squeezed, 9'h0d5);
  assign p2_smul_57958_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__60_squeezed, 9'h0d5);
  assign p2_or_138885_comb = p2_prod__499_comb | 32'h0000_0080;
  assign p2_smul_57962_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__62_squeezed, 9'h105);
  assign p2_or_139011_comb = p2_prod__56_comb | 32'h0000_0080;
  assign p2_smul_58098_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__2_squeezed, 9'h0d5);
  assign p2_smul_58100_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__3_squeezed, 9'h105);
  assign p2_smul_58102_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__4_squeezed, 9'h105);
  assign p2_smul_58104_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__5_squeezed, 9'h0d5);
  assign p2_or_139026_comb = p2_prod__63_comb | 32'h0000_0080;
  assign p2_or_139027_comb = p2_prod__99_comb | 32'h0000_0080;
  assign p2_smul_58114_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__10_squeezed, 9'h0d5);
  assign p2_smul_58116_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__11_squeezed, 9'h105);
  assign p2_smul_58118_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__12_squeezed, 9'h105);
  assign p2_smul_58120_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__13_squeezed, 9'h0d5);
  assign p2_or_139042_comb = p2_prod__127_comb | 32'h0000_0080;
  assign p2_or_139075_comb = p2_prod__419_comb | 32'h0000_0080;
  assign p2_smul_58194_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__50_squeezed, 9'h0d5);
  assign p2_smul_58196_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__51_squeezed, 9'h105);
  assign p2_smul_58198_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__52_squeezed, 9'h105);
  assign p2_smul_58200_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__53_squeezed, 9'h0d5);
  assign p2_or_139090_comb = p2_prod__447_comb | 32'h0000_0080;
  assign p2_or_139091_comb = p2_prod__483_comb | 32'h0000_0080;
  assign p2_smul_58210_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__58_squeezed, 9'h0d5);
  assign p2_smul_58212_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__59_squeezed, 9'h105);
  assign p2_smul_58214_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__60_squeezed, 9'h105);
  assign p2_smul_58216_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__61_squeezed, 9'h0d5);
  assign p2_or_139106_comb = p2_prod__511_comb | 32'h0000_0080;
  assign p2_sel_139107_comb = p1_sgt_135507 ? 16'h7fff : {p1_slt_135220 ? 8'h80 : p1_shifted__16_squeezed, p2_smul_57326_TrailingBits___16_comb};
  assign p2_sel_139108_comb = p1_sgt_135508 ? 16'h7fff : {p1_slt_135222 ? 8'h80 : p1_shifted__17_squeezed, p2_smul_57326_TrailingBits___17_comb};
  assign p2_sel_139109_comb = p1_sgt_135509 ? 16'h7fff : {p1_slt_135224 ? 8'h80 : p1_shifted__18_squeezed, p2_smul_57326_TrailingBits___18_comb};
  assign p2_sel_139110_comb = p1_sgt_135510 ? 16'h7fff : {p1_slt_135226 ? 8'h80 : p1_shifted__19_squeezed, p2_smul_57326_TrailingBits___19_comb};
  assign p2_sel_139111_comb = p1_sgt_135511 ? 16'h7fff : {p1_slt_135228 ? 8'h80 : p1_shifted__20_squeezed, p2_smul_57326_TrailingBits___20_comb};
  assign p2_sel_139112_comb = p1_sgt_135512 ? 16'h7fff : {p1_slt_135230 ? 8'h80 : p1_shifted__21_squeezed, p2_smul_57326_TrailingBits___21_comb};
  assign p2_sel_139113_comb = p1_sgt_135513 ? 16'h7fff : {p1_slt_135232 ? 8'h80 : p1_shifted__22_squeezed, p2_smul_57326_TrailingBits___22_comb};
  assign p2_sel_139114_comb = p1_sgt_135514 ? 16'h7fff : {p1_slt_135234 ? 8'h80 : p1_shifted__23_squeezed, p2_smul_57326_TrailingBits___23_comb};
  assign p2_sel_139115_comb = p1_sgt_135515 ? 16'h7fff : {p1_slt_135236 ? 8'h80 : p1_shifted__40_squeezed, p2_smul_57326_TrailingBits___40_comb};
  assign p2_sel_139116_comb = p1_sgt_135516 ? 16'h7fff : {p1_slt_135238 ? 8'h80 : p1_shifted__41_squeezed, p2_smul_57326_TrailingBits___41_comb};
  assign p2_sel_139117_comb = p1_sgt_135517 ? 16'h7fff : {p1_slt_135240 ? 8'h80 : p1_shifted__42_squeezed, p2_smul_57326_TrailingBits___42_comb};
  assign p2_sel_139118_comb = p1_sgt_135518 ? 16'h7fff : {p1_slt_135242 ? 8'h80 : p1_shifted__43_squeezed, p2_smul_57326_TrailingBits___43_comb};
  assign p2_sel_139119_comb = p1_sgt_135519 ? 16'h7fff : {p1_slt_135244 ? 8'h80 : p1_shifted__44_squeezed, p2_smul_57326_TrailingBits___44_comb};
  assign p2_sel_139120_comb = p1_sgt_135520 ? 16'h7fff : {p1_slt_135246 ? 8'h80 : p1_shifted__45_squeezed, p2_smul_57326_TrailingBits___45_comb};
  assign p2_sel_139121_comb = p1_sgt_135521 ? 16'h7fff : {p1_slt_135248 ? 8'h80 : p1_shifted__46_squeezed, p2_smul_57326_TrailingBits___46_comb};
  assign p2_sel_139122_comb = p1_sgt_135522 ? 16'h7fff : {p1_slt_135250 ? 8'h80 : p1_shifted__47_squeezed, p2_smul_57326_TrailingBits___47_comb};
  assign p2_sel_139571_comb = p1_sgt_135523 ? 16'h7fff : {p1_slt_135252 ? 8'h80 : p1_shifted_squeezed, p2_smul_57326_TrailingBits__comb};
  assign p2_sel_139572_comb = p1_sgt_135524 ? 16'h7fff : {p1_slt_135254 ? 8'h80 : p1_shifted__1_squeezed, p2_smul_57326_TrailingBits___1_comb};
  assign p2_sel_139573_comb = p1_sgt_135525 ? 16'h7fff : {p1_slt_135256 ? 8'h80 : p1_shifted__2_squeezed, p2_smul_57326_TrailingBits___2_comb};
  assign p2_sel_139574_comb = p1_sgt_135526 ? 16'h7fff : {p1_slt_135258 ? 8'h80 : p1_shifted__3_squeezed, p2_smul_57326_TrailingBits___3_comb};
  assign p2_sel_139575_comb = p1_sgt_135527 ? 16'h7fff : {p1_slt_135260 ? 8'h80 : p1_shifted__4_squeezed, p2_smul_57326_TrailingBits___4_comb};
  assign p2_sel_139576_comb = p1_sgt_135528 ? 16'h7fff : {p1_slt_135262 ? 8'h80 : p1_shifted__5_squeezed, p2_smul_57326_TrailingBits___5_comb};
  assign p2_sel_139577_comb = p1_sgt_135529 ? 16'h7fff : {p1_slt_135264 ? 8'h80 : p1_shifted__6_squeezed, p2_smul_57326_TrailingBits___6_comb};
  assign p2_sel_139578_comb = p1_sgt_135530 ? 16'h7fff : {p1_slt_135266 ? 8'h80 : p1_shifted__7_squeezed, p2_smul_57326_TrailingBits___7_comb};
  assign p2_sel_139579_comb = p1_sgt_135531 ? 16'h7fff : {p1_slt_135268 ? 8'h80 : p1_shifted__8_squeezed, p2_smul_57326_TrailingBits___8_comb};
  assign p2_sel_139580_comb = p1_sgt_135532 ? 16'h7fff : {p1_slt_135270 ? 8'h80 : p1_shifted__9_squeezed, p2_smul_57326_TrailingBits___9_comb};
  assign p2_sel_139581_comb = p1_sgt_135533 ? 16'h7fff : {p1_slt_135272 ? 8'h80 : p1_shifted__10_squeezed, p2_smul_57326_TrailingBits___10_comb};
  assign p2_sel_139582_comb = p1_sgt_135534 ? 16'h7fff : {p1_slt_135274 ? 8'h80 : p1_shifted__11_squeezed, p2_smul_57326_TrailingBits___11_comb};
  assign p2_sel_139583_comb = p1_sgt_135535 ? 16'h7fff : {p1_slt_135276 ? 8'h80 : p1_shifted__12_squeezed, p2_smul_57326_TrailingBits___12_comb};
  assign p2_sel_139584_comb = p1_sgt_135536 ? 16'h7fff : {p1_slt_135278 ? 8'h80 : p1_shifted__13_squeezed, p2_smul_57326_TrailingBits___13_comb};
  assign p2_sel_139585_comb = p1_sgt_135537 ? 16'h7fff : {p1_slt_135280 ? 8'h80 : p1_shifted__14_squeezed, p2_smul_57326_TrailingBits___14_comb};
  assign p2_sel_139586_comb = p1_sgt_135538 ? 16'h7fff : {p1_slt_135282 ? 8'h80 : p1_shifted__15_squeezed, p2_smul_57326_TrailingBits___15_comb};
  assign p2_sel_139587_comb = p1_sgt_135539 ? 16'h7fff : {p1_slt_135284 ? 8'h80 : p1_shifted__24_squeezed, p2_smul_57326_TrailingBits___24_comb};
  assign p2_sel_139588_comb = p1_sgt_135540 ? 16'h7fff : {p1_slt_135286 ? 8'h80 : p1_shifted__25_squeezed, p2_smul_57326_TrailingBits___25_comb};
  assign p2_sel_139589_comb = p1_sgt_135541 ? 16'h7fff : {p1_slt_135288 ? 8'h80 : p1_shifted__26_squeezed, p2_smul_57326_TrailingBits___26_comb};
  assign p2_sel_139590_comb = p1_sgt_135542 ? 16'h7fff : {p1_slt_135290 ? 8'h80 : p1_shifted__27_squeezed, p2_smul_57326_TrailingBits___27_comb};
  assign p2_sel_139591_comb = p1_sgt_135543 ? 16'h7fff : {p1_slt_135292 ? 8'h80 : p1_shifted__28_squeezed, p2_smul_57326_TrailingBits___28_comb};
  assign p2_sel_139592_comb = p1_sgt_135544 ? 16'h7fff : {p1_slt_135294 ? 8'h80 : p1_shifted__29_squeezed, p2_smul_57326_TrailingBits___29_comb};
  assign p2_sel_139593_comb = p1_sgt_135545 ? 16'h7fff : {p1_slt_135296 ? 8'h80 : p1_shifted__30_squeezed, p2_smul_57326_TrailingBits___30_comb};
  assign p2_sel_139594_comb = p1_sgt_135546 ? 16'h7fff : {p1_slt_135298 ? 8'h80 : p1_shifted__31_squeezed, p2_smul_57326_TrailingBits___31_comb};
  assign p2_sel_139595_comb = p1_sgt_135547 ? 16'h7fff : {p1_slt_135300 ? 8'h80 : p1_shifted__32_squeezed, p2_smul_57326_TrailingBits___32_comb};
  assign p2_sel_139596_comb = p1_sgt_135548 ? 16'h7fff : {p1_slt_135302 ? 8'h80 : p1_shifted__33_squeezed, p2_smul_57326_TrailingBits___33_comb};
  assign p2_sel_139597_comb = p1_sgt_135549 ? 16'h7fff : {p1_slt_135304 ? 8'h80 : p1_shifted__34_squeezed, p2_smul_57326_TrailingBits___34_comb};
  assign p2_sel_139598_comb = p1_sgt_135550 ? 16'h7fff : {p1_slt_135306 ? 8'h80 : p1_shifted__35_squeezed, p2_smul_57326_TrailingBits___35_comb};
  assign p2_sel_139599_comb = p1_sgt_135551 ? 16'h7fff : {p1_slt_135308 ? 8'h80 : p1_shifted__36_squeezed, p2_smul_57326_TrailingBits___36_comb};
  assign p2_sel_139600_comb = p1_sgt_135552 ? 16'h7fff : {p1_slt_135310 ? 8'h80 : p1_shifted__37_squeezed, p2_smul_57326_TrailingBits___37_comb};
  assign p2_sel_139601_comb = p1_sgt_135553 ? 16'h7fff : {p1_slt_135312 ? 8'h80 : p1_shifted__38_squeezed, p2_smul_57326_TrailingBits___38_comb};
  assign p2_sel_139602_comb = p1_sgt_135554 ? 16'h7fff : {p1_slt_135314 ? 8'h80 : p1_shifted__39_squeezed, p2_smul_57326_TrailingBits___39_comb};
  assign p2_sel_139603_comb = p1_sgt_135555 ? 16'h7fff : {p1_slt_135316 ? 8'h80 : p1_shifted__48_squeezed, p2_smul_57326_TrailingBits___48_comb};
  assign p2_sel_139604_comb = p1_sgt_135556 ? 16'h7fff : {p1_slt_135318 ? 8'h80 : p1_shifted__49_squeezed, p2_smul_57326_TrailingBits___49_comb};
  assign p2_sel_139605_comb = p1_sgt_135557 ? 16'h7fff : {p1_slt_135320 ? 8'h80 : p1_shifted__50_squeezed, p2_smul_57326_TrailingBits___50_comb};
  assign p2_sel_139606_comb = p1_sgt_135558 ? 16'h7fff : {p1_slt_135322 ? 8'h80 : p1_shifted__51_squeezed, p2_smul_57326_TrailingBits___51_comb};
  assign p2_sel_139607_comb = p1_sgt_135559 ? 16'h7fff : {p1_slt_135324 ? 8'h80 : p1_shifted__52_squeezed, p2_smul_57326_TrailingBits___52_comb};
  assign p2_sel_139608_comb = p1_sgt_135560 ? 16'h7fff : {p1_slt_135326 ? 8'h80 : p1_shifted__53_squeezed, p2_smul_57326_TrailingBits___53_comb};
  assign p2_sel_139609_comb = p1_sgt_135561 ? 16'h7fff : {p1_slt_135328 ? 8'h80 : p1_shifted__54_squeezed, p2_smul_57326_TrailingBits___54_comb};
  assign p2_sel_139610_comb = p1_sgt_135562 ? 16'h7fff : {p1_slt_135330 ? 8'h80 : p1_shifted__55_squeezed, p2_smul_57326_TrailingBits___55_comb};
  assign p2_sel_139611_comb = p1_sgt_135563 ? 16'h7fff : {p1_slt_135332 ? 8'h80 : p1_shifted__56_squeezed, p2_smul_57326_TrailingBits___56_comb};
  assign p2_sel_139612_comb = p1_sgt_135564 ? 16'h7fff : {p1_slt_135334 ? 8'h80 : p1_shifted__57_squeezed, p2_smul_57326_TrailingBits___57_comb};
  assign p2_sel_139613_comb = p1_sgt_135565 ? 16'h7fff : {p1_slt_135336 ? 8'h80 : p1_shifted__58_squeezed, p2_smul_57326_TrailingBits___58_comb};
  assign p2_sel_139614_comb = p1_sgt_135566 ? 16'h7fff : {p1_slt_135338 ? 8'h80 : p1_shifted__59_squeezed, p2_smul_57326_TrailingBits___59_comb};
  assign p2_sel_139615_comb = p1_sgt_135567 ? 16'h7fff : {p1_slt_135340 ? 8'h80 : p1_shifted__60_squeezed, p2_smul_57326_TrailingBits___60_comb};
  assign p2_sel_139616_comb = p1_sgt_135568 ? 16'h7fff : {p1_slt_135342 ? 8'h80 : p1_shifted__61_squeezed, p2_smul_57326_TrailingBits___61_comb};
  assign p2_sel_139617_comb = p1_sgt_135569 ? 16'h7fff : {p1_slt_135344 ? 8'h80 : p1_shifted__62_squeezed, p2_smul_57326_TrailingBits___62_comb};
  assign p2_sel_139618_comb = p1_sgt_135570 ? 16'h7fff : {p1_slt_135346 ? 8'h80 : p1_shifted__63_squeezed, p2_smul_57326_TrailingBits___63_comb};
  assign p2_sel_142427_comb = $signed(p2_smul_57742_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57742_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57742_NarrowedMult__comb[15:0]);
  assign p2_sel_142428_comb = $signed(p2_smul_57744_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57744_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57744_NarrowedMult__comb[15:0]);
  assign p2_sel_142429_comb = $signed(p2_smul_57746_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57746_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57746_NarrowedMult__comb[15:0]);
  assign p2_sel_142430_comb = $signed(p2_smul_57748_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57748_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57748_NarrowedMult__comb[15:0]);
  assign p2_sel_142431_comb = $signed(p2_smul_57750_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57750_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57750_NarrowedMult__comb[15:0]);
  assign p2_sel_142432_comb = $signed(p2_smul_57752_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57752_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57752_NarrowedMult__comb[15:0]);
  assign p2_sel_142433_comb = $signed(p2_smul_57754_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57754_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57754_NarrowedMult__comb[15:0]);
  assign p2_sel_142434_comb = $signed(p2_smul_57756_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57756_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57756_NarrowedMult__comb[15:0]);
  assign p2_sel_142435_comb = $signed(p2_smul_57790_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57790_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57790_NarrowedMult__comb[15:0]);
  assign p2_sel_142436_comb = $signed(p2_smul_57792_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57792_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57792_NarrowedMult__comb[15:0]);
  assign p2_sel_142437_comb = $signed(p2_smul_57794_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57794_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57794_NarrowedMult__comb[15:0]);
  assign p2_sel_142438_comb = $signed(p2_smul_57796_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57796_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57796_NarrowedMult__comb[15:0]);
  assign p2_sel_142439_comb = $signed(p2_smul_57798_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57798_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57798_NarrowedMult__comb[15:0]);
  assign p2_sel_142440_comb = $signed(p2_smul_57800_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57800_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57800_NarrowedMult__comb[15:0]);
  assign p2_sel_142441_comb = $signed(p2_smul_57802_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57802_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57802_NarrowedMult__comb[15:0]);
  assign p2_sel_142442_comb = $signed(p2_smul_57804_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57804_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57804_NarrowedMult__comb[15:0]);
  assign p2_sel_142659_comb = $signed(p2_smul_57710_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57710_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57710_NarrowedMult__comb[15:0]);
  assign p2_sel_142660_comb = $signed(p2_smul_57712_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57712_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57712_NarrowedMult__comb[15:0]);
  assign p2_sel_142661_comb = $signed(p2_smul_57714_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57714_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57714_NarrowedMult__comb[15:0]);
  assign p2_sel_142662_comb = $signed(p2_smul_57716_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57716_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57716_NarrowedMult__comb[15:0]);
  assign p2_sel_142663_comb = $signed(p2_smul_57718_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57718_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57718_NarrowedMult__comb[15:0]);
  assign p2_sel_142664_comb = $signed(p2_smul_57720_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57720_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57720_NarrowedMult__comb[15:0]);
  assign p2_sel_142665_comb = $signed(p2_smul_57722_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57722_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57722_NarrowedMult__comb[15:0]);
  assign p2_sel_142666_comb = $signed(p2_smul_57724_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57724_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57724_NarrowedMult__comb[15:0]);
  assign p2_sel_142667_comb = $signed(p2_smul_57726_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57726_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57726_NarrowedMult__comb[15:0]);
  assign p2_sel_142668_comb = $signed(p2_smul_57728_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57728_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57728_NarrowedMult__comb[15:0]);
  assign p2_sel_142669_comb = $signed(p2_smul_57730_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57730_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57730_NarrowedMult__comb[15:0]);
  assign p2_sel_142670_comb = $signed(p2_smul_57732_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57732_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57732_NarrowedMult__comb[15:0]);
  assign p2_sel_142671_comb = $signed(p2_smul_57734_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57734_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57734_NarrowedMult__comb[15:0]);
  assign p2_sel_142672_comb = $signed(p2_smul_57736_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57736_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57736_NarrowedMult__comb[15:0]);
  assign p2_sel_142673_comb = $signed(p2_smul_57738_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57738_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57738_NarrowedMult__comb[15:0]);
  assign p2_sel_142674_comb = $signed(p2_smul_57740_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57740_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57740_NarrowedMult__comb[15:0]);
  assign p2_sel_142675_comb = $signed(p2_smul_57758_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57758_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57758_NarrowedMult__comb[15:0]);
  assign p2_sel_142676_comb = $signed(p2_smul_57760_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57760_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57760_NarrowedMult__comb[15:0]);
  assign p2_sel_142677_comb = $signed(p2_smul_57762_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57762_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57762_NarrowedMult__comb[15:0]);
  assign p2_sel_142678_comb = $signed(p2_smul_57764_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57764_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57764_NarrowedMult__comb[15:0]);
  assign p2_sel_142679_comb = $signed(p2_smul_57766_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57766_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57766_NarrowedMult__comb[15:0]);
  assign p2_sel_142680_comb = $signed(p2_smul_57768_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57768_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57768_NarrowedMult__comb[15:0]);
  assign p2_sel_142681_comb = $signed(p2_smul_57770_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57770_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57770_NarrowedMult__comb[15:0]);
  assign p2_sel_142682_comb = $signed(p2_smul_57772_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57772_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57772_NarrowedMult__comb[15:0]);
  assign p2_sel_142683_comb = $signed(p2_smul_57774_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57774_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57774_NarrowedMult__comb[15:0]);
  assign p2_sel_142684_comb = $signed(p2_smul_57776_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57776_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57776_NarrowedMult__comb[15:0]);
  assign p2_sel_142685_comb = $signed(p2_smul_57778_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57778_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57778_NarrowedMult__comb[15:0]);
  assign p2_sel_142686_comb = $signed(p2_smul_57780_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57780_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57780_NarrowedMult__comb[15:0]);
  assign p2_sel_142687_comb = $signed(p2_smul_57782_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57782_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57782_NarrowedMult__comb[15:0]);
  assign p2_sel_142688_comb = $signed(p2_smul_57784_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57784_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57784_NarrowedMult__comb[15:0]);
  assign p2_sel_142689_comb = $signed(p2_smul_57786_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57786_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57786_NarrowedMult__comb[15:0]);
  assign p2_sel_142690_comb = $signed(p2_smul_57788_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57788_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57788_NarrowedMult__comb[15:0]);
  assign p2_sel_142691_comb = $signed(p2_smul_57806_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57806_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57806_NarrowedMult__comb[15:0]);
  assign p2_sel_142692_comb = $signed(p2_smul_57808_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57808_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57808_NarrowedMult__comb[15:0]);
  assign p2_sel_142693_comb = $signed(p2_smul_57810_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57810_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57810_NarrowedMult__comb[15:0]);
  assign p2_sel_142694_comb = $signed(p2_smul_57812_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57812_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57812_NarrowedMult__comb[15:0]);
  assign p2_sel_142695_comb = $signed(p2_smul_57814_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57814_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57814_NarrowedMult__comb[15:0]);
  assign p2_sel_142696_comb = $signed(p2_smul_57816_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57816_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57816_NarrowedMult__comb[15:0]);
  assign p2_sel_142697_comb = $signed(p2_smul_57818_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57818_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57818_NarrowedMult__comb[15:0]);
  assign p2_sel_142698_comb = $signed(p2_smul_57820_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57820_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57820_NarrowedMult__comb[15:0]);
  assign p2_sel_142699_comb = $signed(p2_smul_57822_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57822_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57822_NarrowedMult__comb[15:0]);
  assign p2_sel_142700_comb = $signed(p2_smul_57824_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57824_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57824_NarrowedMult__comb[15:0]);
  assign p2_sel_142701_comb = $signed(p2_smul_57826_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57826_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57826_NarrowedMult__comb[15:0]);
  assign p2_sel_142702_comb = $signed(p2_smul_57828_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57828_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57828_NarrowedMult__comb[15:0]);
  assign p2_sel_142703_comb = $signed(p2_smul_57830_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57830_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57830_NarrowedMult__comb[15:0]);
  assign p2_sel_142704_comb = $signed(p2_smul_57832_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57832_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57832_NarrowedMult__comb[15:0]);
  assign p2_sel_142705_comb = $signed(p2_smul_57834_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57834_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57834_NarrowedMult__comb[15:0]);
  assign p2_sel_142706_comb = $signed(p2_smul_57836_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57836_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57836_NarrowedMult__comb[15:0]);
  assign p2_add_142371_comb = {{1{p2_sel_139107_comb[15]}}, p2_sel_139107_comb} + {{1{p2_sel_139108_comb[15]}}, p2_sel_139108_comb};
  assign p2_add_142372_comb = {{1{p2_sel_139109_comb[15]}}, p2_sel_139109_comb} + {{1{p2_sel_139110_comb[15]}}, p2_sel_139110_comb};
  assign p2_add_142373_comb = {{1{p2_sel_139111_comb[15]}}, p2_sel_139111_comb} + {{1{p2_sel_139112_comb[15]}}, p2_sel_139112_comb};
  assign p2_add_142374_comb = {{1{p2_sel_139113_comb[15]}}, p2_sel_139113_comb} + {{1{p2_sel_139114_comb[15]}}, p2_sel_139114_comb};
  assign p2_add_142375_comb = {{1{p2_sel_139115_comb[15]}}, p2_sel_139115_comb} + {{1{p2_sel_139116_comb[15]}}, p2_sel_139116_comb};
  assign p2_add_142376_comb = {{1{p2_sel_139117_comb[15]}}, p2_sel_139117_comb} + {{1{p2_sel_139118_comb[15]}}, p2_sel_139118_comb};
  assign p2_add_142377_comb = {{1{p2_sel_139119_comb[15]}}, p2_sel_139119_comb} + {{1{p2_sel_139120_comb[15]}}, p2_sel_139120_comb};
  assign p2_add_142378_comb = {{1{p2_sel_139121_comb[15]}}, p2_sel_139121_comb} + {{1{p2_sel_139122_comb[15]}}, p2_sel_139122_comb};
  assign p2_add_142491_comb = {{1{p2_sel_139571_comb[15]}}, p2_sel_139571_comb} + {{1{p2_sel_139572_comb[15]}}, p2_sel_139572_comb};
  assign p2_add_142492_comb = {{1{p2_sel_139573_comb[15]}}, p2_sel_139573_comb} + {{1{p2_sel_139574_comb[15]}}, p2_sel_139574_comb};
  assign p2_add_142493_comb = {{1{p2_sel_139575_comb[15]}}, p2_sel_139575_comb} + {{1{p2_sel_139576_comb[15]}}, p2_sel_139576_comb};
  assign p2_add_142494_comb = {{1{p2_sel_139577_comb[15]}}, p2_sel_139577_comb} + {{1{p2_sel_139578_comb[15]}}, p2_sel_139578_comb};
  assign p2_add_142495_comb = {{1{p2_sel_139579_comb[15]}}, p2_sel_139579_comb} + {{1{p2_sel_139580_comb[15]}}, p2_sel_139580_comb};
  assign p2_add_142496_comb = {{1{p2_sel_139581_comb[15]}}, p2_sel_139581_comb} + {{1{p2_sel_139582_comb[15]}}, p2_sel_139582_comb};
  assign p2_add_142497_comb = {{1{p2_sel_139583_comb[15]}}, p2_sel_139583_comb} + {{1{p2_sel_139584_comb[15]}}, p2_sel_139584_comb};
  assign p2_add_142498_comb = {{1{p2_sel_139585_comb[15]}}, p2_sel_139585_comb} + {{1{p2_sel_139586_comb[15]}}, p2_sel_139586_comb};
  assign p2_add_142499_comb = {{1{p2_sel_139587_comb[15]}}, p2_sel_139587_comb} + {{1{p2_sel_139588_comb[15]}}, p2_sel_139588_comb};
  assign p2_add_142500_comb = {{1{p2_sel_139589_comb[15]}}, p2_sel_139589_comb} + {{1{p2_sel_139590_comb[15]}}, p2_sel_139590_comb};
  assign p2_add_142501_comb = {{1{p2_sel_139591_comb[15]}}, p2_sel_139591_comb} + {{1{p2_sel_139592_comb[15]}}, p2_sel_139592_comb};
  assign p2_add_142502_comb = {{1{p2_sel_139593_comb[15]}}, p2_sel_139593_comb} + {{1{p2_sel_139594_comb[15]}}, p2_sel_139594_comb};
  assign p2_add_142503_comb = {{1{p2_sel_139595_comb[15]}}, p2_sel_139595_comb} + {{1{p2_sel_139596_comb[15]}}, p2_sel_139596_comb};
  assign p2_add_142504_comb = {{1{p2_sel_139597_comb[15]}}, p2_sel_139597_comb} + {{1{p2_sel_139598_comb[15]}}, p2_sel_139598_comb};
  assign p2_add_142505_comb = {{1{p2_sel_139599_comb[15]}}, p2_sel_139599_comb} + {{1{p2_sel_139600_comb[15]}}, p2_sel_139600_comb};
  assign p2_add_142506_comb = {{1{p2_sel_139601_comb[15]}}, p2_sel_139601_comb} + {{1{p2_sel_139602_comb[15]}}, p2_sel_139602_comb};
  assign p2_add_142507_comb = {{1{p2_sel_139603_comb[15]}}, p2_sel_139603_comb} + {{1{p2_sel_139604_comb[15]}}, p2_sel_139604_comb};
  assign p2_add_142508_comb = {{1{p2_sel_139605_comb[15]}}, p2_sel_139605_comb} + {{1{p2_sel_139606_comb[15]}}, p2_sel_139606_comb};
  assign p2_add_142509_comb = {{1{p2_sel_139607_comb[15]}}, p2_sel_139607_comb} + {{1{p2_sel_139608_comb[15]}}, p2_sel_139608_comb};
  assign p2_add_142510_comb = {{1{p2_sel_139609_comb[15]}}, p2_sel_139609_comb} + {{1{p2_sel_139610_comb[15]}}, p2_sel_139610_comb};
  assign p2_add_142511_comb = {{1{p2_sel_139611_comb[15]}}, p2_sel_139611_comb} + {{1{p2_sel_139612_comb[15]}}, p2_sel_139612_comb};
  assign p2_add_142512_comb = {{1{p2_sel_139613_comb[15]}}, p2_sel_139613_comb} + {{1{p2_sel_139614_comb[15]}}, p2_sel_139614_comb};
  assign p2_add_142513_comb = {{1{p2_sel_139615_comb[15]}}, p2_sel_139615_comb} + {{1{p2_sel_139616_comb[15]}}, p2_sel_139616_comb};
  assign p2_add_142514_comb = {{1{p2_sel_139617_comb[15]}}, p2_sel_139617_comb} + {{1{p2_sel_139618_comb[15]}}, p2_sel_139618_comb};
  assign p2_sel_142531_comb = $signed(p2_smul_57374_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57374_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57374_NarrowedMult__comb[15:0]);
  assign p2_sel_142532_comb = $signed(p2_smul_57376_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57376_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57376_NarrowedMult__comb[15:0]);
  assign p2_sel_142533_comb = $signed(p2_or_137427_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__199[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137427_comb[23:9], 1'h0};
  assign p2_sel_142534_comb = $signed(p2_or_138426_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138426_comb[23:9], 1'h0};
  assign p2_sel_142535_comb = $signed(p2_or_138427_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138427_comb[23:9], 1'h0};
  assign p2_sel_142536_comb = $signed(p2_or_137434_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__214[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137434_comb[23:9], 1'h0};
  assign p2_sel_142537_comb = $signed(p2_smul_57386_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57386_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57386_NarrowedMult__comb[15:0]);
  assign p2_sel_142538_comb = $signed(p2_smul_57388_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57388_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57388_NarrowedMult__comb[15:0]);
  assign p2_sel_142539_comb = $signed(p2_smul_57390_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57390_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57390_NarrowedMult__comb[15:0]);
  assign p2_sel_142540_comb = $signed(p2_smul_57392_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57392_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57392_NarrowedMult__comb[15:0]);
  assign p2_sel_142541_comb = $signed(p2_or_137441_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__263[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137441_comb[23:9], 1'h0};
  assign p2_sel_142542_comb = $signed(p2_or_138442_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138442_comb[23:9], 1'h0};
  assign p2_sel_142543_comb = $signed(p2_or_138443_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138443_comb[23:9], 1'h0};
  assign p2_sel_142544_comb = $signed(p2_or_137448_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__278[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137448_comb[23:9], 1'h0};
  assign p2_sel_142545_comb = $signed(p2_smul_57402_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57402_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57402_NarrowedMult__comb[15:0]);
  assign p2_sel_142546_comb = $signed(p2_smul_57404_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57404_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57404_NarrowedMult__comb[15:0]);
  assign p2_sel_142627_comb = $signed(p2_smul_57630_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57630_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57630_NarrowedMult__comb[15:0]);
  assign p2_sel_142628_comb = $signed(p2_or_138637_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138637_comb[23:9], 1'h0};
  assign p2_sel_142629_comb = $signed(p2_smul_57634_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57634_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57634_NarrowedMult__comb[15:0]);
  assign p2_sel_142630_comb = $signed(p2_or_137633_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__216[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137633_comb[23:9], 1'h0};
  assign p2_sel_142631_comb = $signed(p2_or_137636_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__223[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137636_comb[23:9], 1'h0};
  assign p2_sel_142632_comb = $signed(p2_smul_57640_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57640_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57640_NarrowedMult__comb[15:0]);
  assign p2_sel_142633_comb = $signed(p2_or_138648_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138648_comb[23:9], 1'h0};
  assign p2_sel_142634_comb = $signed(p2_smul_57644_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57644_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57644_NarrowedMult__comb[15:0]);
  assign p2_sel_142635_comb = $signed(p2_smul_57646_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57646_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57646_NarrowedMult__comb[15:0]);
  assign p2_sel_142636_comb = $signed(p2_or_138653_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138653_comb[23:9], 1'h0};
  assign p2_sel_142637_comb = $signed(p2_smul_57650_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57650_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57650_NarrowedMult__comb[15:0]);
  assign p2_sel_142638_comb = $signed(p2_or_137647_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__280[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137647_comb[23:9], 1'h0};
  assign p2_sel_142639_comb = $signed(p2_or_137650_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__287[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137650_comb[23:9], 1'h0};
  assign p2_sel_142640_comb = $signed(p2_smul_57656_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57656_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57656_NarrowedMult__comb[15:0]);
  assign p2_sel_142641_comb = $signed(p2_or_138664_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138664_comb[23:9], 1'h0};
  assign p2_sel_142642_comb = $signed(p2_smul_57660_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57660_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57660_NarrowedMult__comb[15:0]);
  assign p2_sel_142723_comb = $signed(p2_or_137761_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__212[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137761_comb[23:9], 1'h0};
  assign p2_sel_142724_comb = $signed(p2_smul_57888_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57888_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57888_NarrowedMult__comb[15:0]);
  assign p2_sel_142725_comb = $signed(p2_or_138832_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138832_comb[23:9], 1'h0};
  assign p2_sel_142726_comb = $signed(p2_smul_57892_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57892_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57892_NarrowedMult__comb[15:0]);
  assign p2_sel_142727_comb = $signed(p2_smul_57894_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57894_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57894_NarrowedMult__comb[15:0]);
  assign p2_sel_142728_comb = $signed(p2_or_138837_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138837_comb[23:9], 1'h0};
  assign p2_sel_142729_comb = $signed(p2_smul_57898_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57898_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57898_NarrowedMult__comb[15:0]);
  assign p2_sel_142730_comb = $signed(p2_or_137772_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__250[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137772_comb[23:9], 1'h0};
  assign p2_sel_142731_comb = $signed(p2_or_137775_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__276[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137775_comb[23:9], 1'h0};
  assign p2_sel_142732_comb = $signed(p2_smul_57904_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57904_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57904_NarrowedMult__comb[15:0]);
  assign p2_sel_142733_comb = $signed(p2_or_138848_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138848_comb[23:9], 1'h0};
  assign p2_sel_142734_comb = $signed(p2_smul_57908_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57908_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57908_NarrowedMult__comb[15:0]);
  assign p2_sel_142735_comb = $signed(p2_smul_57910_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57910_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57910_NarrowedMult__comb[15:0]);
  assign p2_sel_142736_comb = $signed(p2_or_138853_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138853_comb[23:9], 1'h0};
  assign p2_sel_142737_comb = $signed(p2_smul_57914_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57914_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57914_NarrowedMult__comb[15:0]);
  assign p2_sel_142738_comb = $signed(p2_or_137786_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__314[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137786_comb[23:9], 1'h0};
  assign p2_sel_142819_comb = $signed(p2_or_139043_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139043_comb[23:9], 1'h0};
  assign p2_sel_142820_comb = $signed(p2_or_137967_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__234[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137967_comb[23:9], 1'h0};
  assign p2_sel_142821_comb = $signed(p2_smul_58146_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58146_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58146_NarrowedMult__comb[15:0]);
  assign p2_sel_142822_comb = $signed(p2_smul_58148_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58148_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58148_NarrowedMult__comb[15:0]);
  assign p2_sel_142823_comb = $signed(p2_smul_58150_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58150_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58150_NarrowedMult__comb[15:0]);
  assign p2_sel_142824_comb = $signed(p2_smul_58152_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58152_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58152_NarrowedMult__comb[15:0]);
  assign p2_sel_142825_comb = $signed(p2_or_137974_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__254[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137974_comb[23:9], 1'h0};
  assign p2_sel_142826_comb = $signed(p2_or_139058_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139058_comb[23:9], 1'h0};
  assign p2_sel_142827_comb = $signed(p2_or_139059_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139059_comb[23:9], 1'h0};
  assign p2_sel_142828_comb = $signed(p2_or_137981_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__298[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137981_comb[23:9], 1'h0};
  assign p2_sel_142829_comb = $signed(p2_smul_58162_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58162_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58162_NarrowedMult__comb[15:0]);
  assign p2_sel_142830_comb = $signed(p2_smul_58164_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58164_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58164_NarrowedMult__comb[15:0]);
  assign p2_sel_142831_comb = $signed(p2_smul_58166_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58166_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58166_NarrowedMult__comb[15:0]);
  assign p2_sel_142832_comb = $signed(p2_smul_58168_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58168_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58168_NarrowedMult__comb[15:0]);
  assign p2_sel_142833_comb = $signed(p2_or_137988_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__318[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137988_comb[23:9], 1'h0};
  assign p2_sel_142834_comb = $signed(p2_or_139074_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139074_comb[23:9], 1'h0};
  assign p2_sel_142379_comb = $signed(p2_smul_57358_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57358_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57358_NarrowedMult__comb[15:0]);
  assign p2_sel_142380_comb = $signed(p2_smul_57360_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57360_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57360_NarrowedMult__comb[15:0]);
  assign p2_sel_142381_comb = $signed(p2_or_137095_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__135_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137095_comb[23:9], 1'h0};
  assign p2_sel_142382_comb = $signed(p2_or_138058_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138058_comb[23:9], 1'h0};
  assign p2_sel_142383_comb = $signed(p2_or_138059_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138059_comb[23:9], 1'h0};
  assign p2_sel_142384_comb = $signed(p2_or_137102_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__150_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137102_comb[23:9], 1'h0};
  assign p2_sel_142385_comb = $signed(p2_smul_57370_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57370_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57370_NarrowedMult__comb[15:0]);
  assign p2_sel_142386_comb = $signed(p2_smul_57372_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57372_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57372_NarrowedMult__comb[15:0]);
  assign p2_sel_142387_comb = $signed(p2_smul_57406_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57406_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57406_NarrowedMult__comb[15:0]);
  assign p2_sel_142388_comb = $signed(p2_smul_57408_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57408_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57408_NarrowedMult__comb[15:0]);
  assign p2_sel_142389_comb = $signed(p2_or_137109_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__327_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137109_comb[23:9], 1'h0};
  assign p2_sel_142390_comb = $signed(p2_or_138074_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138074_comb[23:9], 1'h0};
  assign p2_sel_142391_comb = $signed(p2_or_138075_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138075_comb[23:9], 1'h0};
  assign p2_sel_142392_comb = $signed(p2_or_137116_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__342_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137116_comb[23:9], 1'h0};
  assign p2_sel_142393_comb = $signed(p2_smul_57418_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57418_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57418_NarrowedMult__comb[15:0]);
  assign p2_sel_142394_comb = $signed(p2_smul_57420_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57420_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57420_NarrowedMult__comb[15:0]);
  assign p2_sel_142395_comb = $signed(p2_or_137121_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__133_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137121_comb[23:10], 2'h0};
  assign p2_sel_142396_comb = $signed(p2_prod__136_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__136_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57488_NarrowedMult_, 1'h0};
  assign p2_sel_142397_comb = $signed(p2_prod__140_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__140_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57490_NarrowedMult_, 1'h0};
  assign p2_sel_142398_comb = $signed(p2_or_137128_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__145_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137128_comb[23:10], 2'h0};
  assign p2_sel_142399_comb = $signed(p2_or_137131_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__151_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137131_comb[23:10], 2'h0};
  assign p2_sel_142400_comb = $signed(p2_prod__158_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__158_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57496_NarrowedMult_, 1'h0};
  assign p2_sel_142401_comb = $signed(p2_prod__165_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__165_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57498_NarrowedMult_, 1'h0};
  assign p2_sel_142402_comb = $signed(p2_or_137138_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__171_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137138_comb[23:10], 2'h0};
  assign p2_sel_142403_comb = $signed(p2_or_137141_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__325_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137141_comb[23:10], 2'h0};
  assign p2_sel_142404_comb = $signed(p2_prod__328_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__328_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57536_NarrowedMult_, 1'h0};
  assign p2_sel_142405_comb = $signed(p2_prod__332_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__332_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57538_NarrowedMult_, 1'h0};
  assign p2_sel_142406_comb = $signed(p2_or_137148_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__337_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137148_comb[23:10], 2'h0};
  assign p2_sel_142407_comb = $signed(p2_or_137151_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__343_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137151_comb[23:10], 2'h0};
  assign p2_sel_142408_comb = $signed(p2_prod__350_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__350_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57544_NarrowedMult_, 1'h0};
  assign p2_sel_142409_comb = $signed(p2_prod__357_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__357_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57546_NarrowedMult_, 1'h0};
  assign p2_sel_142410_comb = $signed(p2_or_137158_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__363_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137158_comb[23:10], 2'h0};
  assign p2_sel_142411_comb = $signed(p2_smul_57614_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57614_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57614_NarrowedMult__comb[15:0]);
  assign p2_sel_142412_comb = $signed(p2_or_138125_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138125_comb[23:9], 1'h0};
  assign p2_sel_142413_comb = $signed(p2_smul_57618_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57618_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57618_NarrowedMult__comb[15:0]);
  assign p2_sel_142414_comb = $signed(p2_or_137165_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__152_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137165_comb[23:9], 1'h0};
  assign p2_sel_142415_comb = $signed(p2_or_137168_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__159_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137168_comb[23:9], 1'h0};
  assign p2_sel_142416_comb = $signed(p2_smul_57624_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57624_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57624_NarrowedMult__comb[15:0]);
  assign p2_sel_142417_comb = $signed(p2_or_138136_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138136_comb[23:9], 1'h0};
  assign p2_sel_142418_comb = $signed(p2_smul_57628_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57628_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57628_NarrowedMult__comb[15:0]);
  assign p2_sel_142419_comb = $signed(p2_smul_57662_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57662_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57662_NarrowedMult__comb[15:0]);
  assign p2_sel_142420_comb = $signed(p2_or_138141_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138141_comb[23:9], 1'h0};
  assign p2_sel_142421_comb = $signed(p2_smul_57666_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57666_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57666_NarrowedMult__comb[15:0]);
  assign p2_sel_142422_comb = $signed(p2_or_137179_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__344_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137179_comb[23:9], 1'h0};
  assign p2_sel_142423_comb = $signed(p2_or_137182_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__351_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137182_comb[23:9], 1'h0};
  assign p2_sel_142424_comb = $signed(p2_smul_57672_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57672_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57672_NarrowedMult__comb[15:0]);
  assign p2_sel_142425_comb = $signed(p2_or_138152_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138152_comb[23:9], 1'h0};
  assign p2_sel_142426_comb = $signed(p2_smul_57676_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57676_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57676_NarrowedMult__comb[15:0]);
  assign p2_sel_142443_comb = $signed(p2_or_137205_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__148_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137205_comb[23:9], 1'h0};
  assign p2_sel_142444_comb = $signed(p2_smul_57872_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57872_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57872_NarrowedMult__comb[15:0]);
  assign p2_sel_142445_comb = $signed(p2_or_138192_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138192_comb[23:9], 1'h0};
  assign p2_sel_142446_comb = $signed(p2_smul_57876_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57876_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57876_NarrowedMult__comb[15:0]);
  assign p2_sel_142447_comb = $signed(p2_smul_57878_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57878_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57878_NarrowedMult__comb[15:0]);
  assign p2_sel_142448_comb = $signed(p2_or_138197_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138197_comb[23:9], 1'h0};
  assign p2_sel_142449_comb = $signed(p2_smul_57882_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57882_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57882_NarrowedMult__comb[15:0]);
  assign p2_sel_142450_comb = $signed(p2_or_137216_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__186_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137216_comb[23:9], 1'h0};
  assign p2_sel_142451_comb = $signed(p2_or_137219_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__340_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137219_comb[23:9], 1'h0};
  assign p2_sel_142452_comb = $signed(p2_smul_57920_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57920_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57920_NarrowedMult__comb[15:0]);
  assign p2_sel_142453_comb = $signed(p2_or_138208_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138208_comb[23:9], 1'h0};
  assign p2_sel_142454_comb = $signed(p2_smul_57924_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57924_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57924_NarrowedMult__comb[15:0]);
  assign p2_sel_142455_comb = $signed(p2_smul_57926_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57926_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57926_NarrowedMult__comb[15:0]);
  assign p2_sel_142456_comb = $signed(p2_or_138213_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138213_comb[23:9], 1'h0};
  assign p2_sel_142457_comb = $signed(p2_smul_57930_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57930_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57930_NarrowedMult__comb[15:0]);
  assign p2_sel_142458_comb = $signed(p2_or_137230_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__378_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137230_comb[23:9], 1'h0};
  assign p2_sel_142459_comb = $signed(p2_prod__155_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__155_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57998_NarrowedMult_, 1'h0};
  assign p2_sel_142460_comb = $signed(p2_or_137235_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__162_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137235_comb[23:10], 2'h0};
  assign p2_sel_142461_comb = $signed(p2_prod__169_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__169_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58002_NarrowedMult_, 1'h0};
  assign p2_sel_142462_comb = $signed(p2_or_137240_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__175_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137240_comb[23:10], 2'h0};
  assign p2_sel_142463_comb = $signed(p2_or_137243_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__180_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137243_comb[23:10], 2'h0};
  assign p2_sel_142464_comb = $signed(p2_prod__184_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__184_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58008_NarrowedMult_, 1'h0};
  assign p2_sel_142465_comb = $signed(p2_or_137248_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__187_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137248_comb[23:10], 2'h0};
  assign p2_sel_142466_comb = $signed(p2_prod__189_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__189_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58012_NarrowedMult_, 1'h0};
  assign p2_sel_142467_comb = $signed(p2_prod__347_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__347_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58046_NarrowedMult_, 1'h0};
  assign p2_sel_142468_comb = $signed(p2_or_137255_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__354_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137255_comb[23:10], 2'h0};
  assign p2_sel_142469_comb = $signed(p2_prod__361_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__361_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58050_NarrowedMult_, 1'h0};
  assign p2_sel_142470_comb = $signed(p2_or_137260_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__367_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137260_comb[23:10], 2'h0};
  assign p2_sel_142471_comb = $signed(p2_or_137263_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__372_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137263_comb[23:10], 2'h0};
  assign p2_sel_142472_comb = $signed(p2_prod__376_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__376_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58056_NarrowedMult_, 1'h0};
  assign p2_sel_142473_comb = $signed(p2_or_137268_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__379_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137268_comb[23:10], 2'h0};
  assign p2_sel_142474_comb = $signed(p2_prod__381_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__381_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58060_NarrowedMult_, 1'h0};
  assign p2_sel_142475_comb = $signed(p2_or_138259_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138259_comb[23:9], 1'h0};
  assign p2_sel_142476_comb = $signed(p2_or_137275_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__170_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137275_comb[23:9], 1'h0};
  assign p2_sel_142477_comb = $signed(p2_smul_58130_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58130_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58130_NarrowedMult__comb[15:0]);
  assign p2_sel_142478_comb = $signed(p2_smul_58132_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58132_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58132_NarrowedMult__comb[15:0]);
  assign p2_sel_142479_comb = $signed(p2_smul_58134_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58134_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58134_NarrowedMult__comb[15:0]);
  assign p2_sel_142480_comb = $signed(p2_smul_58136_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58136_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58136_NarrowedMult__comb[15:0]);
  assign p2_sel_142481_comb = $signed(p2_or_137282_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__190_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137282_comb[23:9], 1'h0};
  assign p2_sel_142482_comb = $signed(p2_or_138274_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138274_comb[23:9], 1'h0};
  assign p2_sel_142483_comb = $signed(p2_or_138275_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138275_comb[23:9], 1'h0};
  assign p2_sel_142484_comb = $signed(p2_or_137289_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__362_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137289_comb[23:9], 1'h0};
  assign p2_sel_142485_comb = $signed(p2_smul_58178_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58178_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58178_NarrowedMult__comb[15:0]);
  assign p2_sel_142486_comb = $signed(p2_smul_58180_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58180_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58180_NarrowedMult__comb[15:0]);
  assign p2_sel_142487_comb = $signed(p2_smul_58182_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58182_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58182_NarrowedMult__comb[15:0]);
  assign p2_sel_142488_comb = $signed(p2_smul_58184_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58184_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58184_NarrowedMult__comb[15:0]);
  assign p2_sel_142489_comb = $signed(p2_or_137296_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__382_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137296_comb[23:9], 1'h0};
  assign p2_sel_142490_comb = $signed(p2_or_138290_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138290_comb[23:9], 1'h0};
  assign p2_sel_142515_comb = $signed(p2_smul_57326_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57326_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57326_NarrowedMult__comb[15:0]);
  assign p2_sel_142516_comb = $signed(p2_smul_57328_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57328_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57328_NarrowedMult__comb[15:0]);
  assign p2_sel_142517_comb = $signed(p2_or_137399_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__10_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137399_comb[23:9], 1'h0};
  assign p2_sel_142518_comb = $signed(p2_or_138394_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138394_comb[23:9], 1'h0};
  assign p2_sel_142519_comb = $signed(p2_or_138395_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138395_comb[23:9], 1'h0};
  assign p2_sel_142520_comb = $signed(p2_or_137406_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__13_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137406_comb[23:9], 1'h0};
  assign p2_sel_142521_comb = $signed(p2_smul_57338_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57338_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57338_NarrowedMult__comb[15:0]);
  assign p2_sel_142522_comb = $signed(p2_smul_57340_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57340_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57340_NarrowedMult__comb[15:0]);
  assign p2_sel_142523_comb = $signed(p2_smul_57342_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57342_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57342_NarrowedMult__comb[15:0]);
  assign p2_sel_142524_comb = $signed(p2_smul_57344_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57344_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57344_NarrowedMult__comb[15:0]);
  assign p2_sel_142525_comb = $signed(p2_or_137413_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__71_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137413_comb[23:9], 1'h0};
  assign p2_sel_142526_comb = $signed(p2_or_138410_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138410_comb[23:9], 1'h0};
  assign p2_sel_142527_comb = $signed(p2_or_138411_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138411_comb[23:9], 1'h0};
  assign p2_sel_142528_comb = $signed(p2_or_137420_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__86_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137420_comb[23:9], 1'h0};
  assign p2_sel_142529_comb = $signed(p2_smul_57354_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57354_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57354_NarrowedMult__comb[15:0]);
  assign p2_sel_142530_comb = $signed(p2_smul_57356_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57356_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57356_NarrowedMult__comb[15:0]);
  assign p2_sel_142547_comb = $signed(p2_smul_57422_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57422_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57422_NarrowedMult__comb[15:0]);
  assign p2_sel_142548_comb = $signed(p2_smul_57424_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57424_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57424_NarrowedMult__comb[15:0]);
  assign p2_sel_142549_comb = $signed(p2_or_137455_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__391_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137455_comb[23:9], 1'h0};
  assign p2_sel_142550_comb = $signed(p2_or_138458_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138458_comb[23:9], 1'h0};
  assign p2_sel_142551_comb = $signed(p2_or_138459_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138459_comb[23:9], 1'h0};
  assign p2_sel_142552_comb = $signed(p2_or_137462_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__406_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137462_comb[23:9], 1'h0};
  assign p2_sel_142553_comb = $signed(p2_smul_57434_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57434_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57434_NarrowedMult__comb[15:0]);
  assign p2_sel_142554_comb = $signed(p2_smul_57436_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57436_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57436_NarrowedMult__comb[15:0]);
  assign p2_sel_142555_comb = $signed(p2_smul_57438_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57438_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57438_NarrowedMult__comb[15:0]);
  assign p2_sel_142556_comb = $signed(p2_smul_57440_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57440_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57440_NarrowedMult__comb[15:0]);
  assign p2_sel_142557_comb = $signed(p2_or_137469_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__455_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137469_comb[23:9], 1'h0};
  assign p2_sel_142558_comb = $signed(p2_or_138474_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138474_comb[23:9], 1'h0};
  assign p2_sel_142559_comb = $signed(p2_or_138475_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138475_comb[23:9], 1'h0};
  assign p2_sel_142560_comb = $signed(p2_or_137476_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__470_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137476_comb[23:9], 1'h0};
  assign p2_sel_142561_comb = $signed(p2_smul_57450_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57450_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57450_NarrowedMult__comb[15:0]);
  assign p2_sel_142562_comb = $signed(p2_smul_57452_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57452_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57452_NarrowedMult__comb[15:0]);
  assign p2_sel_142563_comb = $signed(p2_or_137481_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__16_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137481_comb[23:10], 2'h0};
  assign p2_sel_142564_comb = $signed(p2_prod__17_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__17_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57456_NarrowedMult_, 1'h0};
  assign p2_sel_142565_comb = $signed(p2_prod__18_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__18_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57458_NarrowedMult_, 1'h0};
  assign p2_sel_142566_comb = $signed(p2_or_137488_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__19_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137488_comb[23:10], 2'h0};
  assign p2_sel_142567_comb = $signed(p2_or_137491_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__20_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137491_comb[23:10], 2'h0};
  assign p2_sel_142568_comb = $signed(p2_prod__21_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__21_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57464_NarrowedMult_, 1'h0};
  assign p2_sel_142569_comb = $signed(p2_prod__22_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__22_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57466_NarrowedMult_, 1'h0};
  assign p2_sel_142570_comb = $signed(p2_or_137498_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__23_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137498_comb[23:10], 2'h0};
  assign p2_sel_142571_comb = $signed(p2_or_137501_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__69_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137501_comb[23:10], 2'h0};
  assign p2_sel_142572_comb = $signed(p2_prod__72_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__72_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57472_NarrowedMult_, 1'h0};
  assign p2_sel_142573_comb = $signed(p2_prod__76_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__76_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57474_NarrowedMult_, 1'h0};
  assign p2_sel_142574_comb = $signed(p2_or_137508_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__81_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137508_comb[23:10], 2'h0};
  assign p2_sel_142575_comb = $signed(p2_or_137511_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__87_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137511_comb[23:10], 2'h0};
  assign p2_sel_142576_comb = $signed(p2_prod__94_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__94_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57480_NarrowedMult_, 1'h0};
  assign p2_sel_142577_comb = $signed(p2_prod__101_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__101_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57482_NarrowedMult_, 1'h0};
  assign p2_sel_142578_comb = $signed(p2_or_137518_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__107_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137518_comb[23:10], 2'h0};
  assign p2_sel_142579_comb = $signed(p2_or_137521_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__197_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137521_comb[23:10], 2'h0};
  assign p2_sel_142580_comb = $signed(p2_prod__200_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__200_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57504_NarrowedMult_, 1'h0};
  assign p2_sel_142581_comb = $signed(p2_prod__204_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__204_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57506_NarrowedMult_, 1'h0};
  assign p2_sel_142582_comb = $signed(p2_or_137528_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__209_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137528_comb[23:10], 2'h0};
  assign p2_sel_142583_comb = $signed(p2_or_137531_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__215_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137531_comb[23:10], 2'h0};
  assign p2_sel_142584_comb = $signed(p2_prod__222_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__222_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57512_NarrowedMult_, 1'h0};
  assign p2_sel_142585_comb = $signed(p2_prod__229_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__229_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57514_NarrowedMult_, 1'h0};
  assign p2_sel_142586_comb = $signed(p2_or_137538_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__235_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137538_comb[23:10], 2'h0};
  assign p2_sel_142587_comb = $signed(p2_or_137541_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__261_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137541_comb[23:10], 2'h0};
  assign p2_sel_142588_comb = $signed(p2_prod__264_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__264_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57520_NarrowedMult_, 1'h0};
  assign p2_sel_142589_comb = $signed(p2_prod__268_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__268_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57522_NarrowedMult_, 1'h0};
  assign p2_sel_142590_comb = $signed(p2_or_137548_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__273_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137548_comb[23:10], 2'h0};
  assign p2_sel_142591_comb = $signed(p2_or_137551_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__279_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137551_comb[23:10], 2'h0};
  assign p2_sel_142592_comb = $signed(p2_prod__286_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__286_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57528_NarrowedMult_, 1'h0};
  assign p2_sel_142593_comb = $signed(p2_prod__293_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__293_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57530_NarrowedMult_, 1'h0};
  assign p2_sel_142594_comb = $signed(p2_or_137558_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__299_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137558_comb[23:10], 2'h0};
  assign p2_sel_142595_comb = $signed(p2_or_137561_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__389_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137561_comb[23:10], 2'h0};
  assign p2_sel_142596_comb = $signed(p2_prod__392_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__392_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57552_NarrowedMult_, 1'h0};
  assign p2_sel_142597_comb = $signed(p2_prod__396_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__396_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57554_NarrowedMult_, 1'h0};
  assign p2_sel_142598_comb = $signed(p2_or_137568_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__401_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137568_comb[23:10], 2'h0};
  assign p2_sel_142599_comb = $signed(p2_or_137571_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__407_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137571_comb[23:10], 2'h0};
  assign p2_sel_142600_comb = $signed(p2_prod__414_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__414_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57560_NarrowedMult_, 1'h0};
  assign p2_sel_142601_comb = $signed(p2_prod__421_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__421_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57562_NarrowedMult_, 1'h0};
  assign p2_sel_142602_comb = $signed(p2_or_137578_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__427_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137578_comb[23:10], 2'h0};
  assign p2_sel_142603_comb = $signed(p2_or_137581_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__453_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137581_comb[23:10], 2'h0};
  assign p2_sel_142604_comb = $signed(p2_prod__456_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__456_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57568_NarrowedMult_, 1'h0};
  assign p2_sel_142605_comb = $signed(p2_prod__460_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__460_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57570_NarrowedMult_, 1'h0};
  assign p2_sel_142606_comb = $signed(p2_or_137588_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__465_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137588_comb[23:10], 2'h0};
  assign p2_sel_142607_comb = $signed(p2_or_137591_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__471_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137591_comb[23:10], 2'h0};
  assign p2_sel_142608_comb = $signed(p2_prod__478_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__478_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57576_NarrowedMult_, 1'h0};
  assign p2_sel_142609_comb = $signed(p2_prod__485_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__485_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57578_NarrowedMult_, 1'h0};
  assign p2_sel_142610_comb = $signed(p2_or_137598_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__491_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137598_comb[23:10], 2'h0};
  assign p2_sel_142611_comb = $signed(p2_smul_57582_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57582_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57582_NarrowedMult__comb[15:0]);
  assign p2_sel_142612_comb = $signed(p2_or_138605_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138605_comb[23:9], 1'h0};
  assign p2_sel_142613_comb = $signed(p2_smul_57586_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57586_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57586_NarrowedMult__comb[15:0]);
  assign p2_sel_142614_comb = $signed(p2_or_137605_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__27_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137605_comb[23:9], 1'h0};
  assign p2_sel_142615_comb = $signed(p2_or_137608_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__28_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137608_comb[23:9], 1'h0};
  assign p2_sel_142616_comb = $signed(p2_smul_57592_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57592_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57592_NarrowedMult__comb[15:0]);
  assign p2_sel_142617_comb = $signed(p2_or_138616_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138616_comb[23:9], 1'h0};
  assign p2_sel_142618_comb = $signed(p2_smul_57596_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57596_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57596_NarrowedMult__comb[15:0]);
  assign p2_sel_142619_comb = $signed(p2_smul_57598_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57598_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57598_NarrowedMult__comb[15:0]);
  assign p2_sel_142620_comb = $signed(p2_or_138621_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138621_comb[23:9], 1'h0};
  assign p2_sel_142621_comb = $signed(p2_smul_57602_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57602_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57602_NarrowedMult__comb[15:0]);
  assign p2_sel_142622_comb = $signed(p2_or_137619_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__88_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137619_comb[23:9], 1'h0};
  assign p2_sel_142623_comb = $signed(p2_or_137622_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__95_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137622_comb[23:9], 1'h0};
  assign p2_sel_142624_comb = $signed(p2_smul_57608_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57608_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57608_NarrowedMult__comb[15:0]);
  assign p2_sel_142625_comb = $signed(p2_or_138632_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138632_comb[23:9], 1'h0};
  assign p2_sel_142626_comb = $signed(p2_smul_57612_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57612_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57612_NarrowedMult__comb[15:0]);
  assign p2_sel_142643_comb = $signed(p2_smul_57678_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57678_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57678_NarrowedMult__comb[15:0]);
  assign p2_sel_142644_comb = $signed(p2_or_138669_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138669_comb[23:9], 1'h0};
  assign p2_sel_142645_comb = $signed(p2_smul_57682_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57682_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57682_NarrowedMult__comb[15:0]);
  assign p2_sel_142646_comb = $signed(p2_or_137661_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__408_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137661_comb[23:9], 1'h0};
  assign p2_sel_142647_comb = $signed(p2_or_137664_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__415_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137664_comb[23:9], 1'h0};
  assign p2_sel_142648_comb = $signed(p2_smul_57688_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57688_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57688_NarrowedMult__comb[15:0]);
  assign p2_sel_142649_comb = $signed(p2_or_138680_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138680_comb[23:9], 1'h0};
  assign p2_sel_142650_comb = $signed(p2_smul_57692_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57692_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57692_NarrowedMult__comb[15:0]);
  assign p2_sel_142651_comb = $signed(p2_smul_57694_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57694_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57694_NarrowedMult__comb[15:0]);
  assign p2_sel_142652_comb = $signed(p2_or_138685_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138685_comb[23:9], 1'h0};
  assign p2_sel_142653_comb = $signed(p2_smul_57698_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57698_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57698_NarrowedMult__comb[15:0]);
  assign p2_sel_142654_comb = $signed(p2_or_137675_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__472_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137675_comb[23:9], 1'h0};
  assign p2_sel_142655_comb = $signed(p2_or_137678_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__479_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137678_comb[23:9], 1'h0};
  assign p2_sel_142656_comb = $signed(p2_smul_57704_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57704_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57704_NarrowedMult__comb[15:0]);
  assign p2_sel_142657_comb = $signed(p2_or_138696_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138696_comb[23:9], 1'h0};
  assign p2_sel_142658_comb = $signed(p2_smul_57708_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57708_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57708_NarrowedMult__comb[15:0]);
  assign p2_sel_142707_comb = $signed(p2_or_137733_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__40_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137733_comb[23:9], 1'h0};
  assign p2_sel_142708_comb = $signed(p2_smul_57840_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57840_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57840_NarrowedMult__comb[15:0]);
  assign p2_sel_142709_comb = $signed(p2_or_138800_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138800_comb[23:9], 1'h0};
  assign p2_sel_142710_comb = $signed(p2_smul_57844_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57844_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57844_NarrowedMult__comb[15:0]);
  assign p2_sel_142711_comb = $signed(p2_smul_57846_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57846_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57846_NarrowedMult__comb[15:0]);
  assign p2_sel_142712_comb = $signed(p2_or_138805_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138805_comb[23:9], 1'h0};
  assign p2_sel_142713_comb = $signed(p2_smul_57850_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57850_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57850_NarrowedMult__comb[15:0]);
  assign p2_sel_142714_comb = $signed(p2_or_137744_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__47_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137744_comb[23:9], 1'h0};
  assign p2_sel_142715_comb = $signed(p2_or_137747_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__84_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137747_comb[23:9], 1'h0};
  assign p2_sel_142716_comb = $signed(p2_smul_57856_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57856_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57856_NarrowedMult__comb[15:0]);
  assign p2_sel_142717_comb = $signed(p2_or_138816_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138816_comb[23:9], 1'h0};
  assign p2_sel_142718_comb = $signed(p2_smul_57860_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57860_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57860_NarrowedMult__comb[15:0]);
  assign p2_sel_142719_comb = $signed(p2_smul_57862_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57862_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57862_NarrowedMult__comb[15:0]);
  assign p2_sel_142720_comb = $signed(p2_or_138821_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138821_comb[23:9], 1'h0};
  assign p2_sel_142721_comb = $signed(p2_smul_57866_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57866_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57866_NarrowedMult__comb[15:0]);
  assign p2_sel_142722_comb = $signed(p2_or_137758_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__122_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137758_comb[23:9], 1'h0};
  assign p2_sel_142739_comb = $signed(p2_or_137789_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__404_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137789_comb[23:9], 1'h0};
  assign p2_sel_142740_comb = $signed(p2_smul_57936_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57936_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57936_NarrowedMult__comb[15:0]);
  assign p2_sel_142741_comb = $signed(p2_or_138864_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138864_comb[23:9], 1'h0};
  assign p2_sel_142742_comb = $signed(p2_smul_57940_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57940_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57940_NarrowedMult__comb[15:0]);
  assign p2_sel_142743_comb = $signed(p2_smul_57942_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57942_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57942_NarrowedMult__comb[15:0]);
  assign p2_sel_142744_comb = $signed(p2_or_138869_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138869_comb[23:9], 1'h0};
  assign p2_sel_142745_comb = $signed(p2_smul_57946_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57946_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57946_NarrowedMult__comb[15:0]);
  assign p2_sel_142746_comb = $signed(p2_or_137800_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__442_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137800_comb[23:9], 1'h0};
  assign p2_sel_142747_comb = $signed(p2_or_137803_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__468_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137803_comb[23:9], 1'h0};
  assign p2_sel_142748_comb = $signed(p2_smul_57952_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57952_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57952_NarrowedMult__comb[15:0]);
  assign p2_sel_142749_comb = $signed(p2_or_138880_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138880_comb[23:9], 1'h0};
  assign p2_sel_142750_comb = $signed(p2_smul_57956_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57956_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57956_NarrowedMult__comb[15:0]);
  assign p2_sel_142751_comb = $signed(p2_smul_57958_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57958_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57958_NarrowedMult__comb[15:0]);
  assign p2_sel_142752_comb = $signed(p2_or_138885_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_138885_comb[23:9], 1'h0};
  assign p2_sel_142753_comb = $signed(p2_smul_57962_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_57962_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_57962_NarrowedMult__comb[15:0]);
  assign p2_sel_142754_comb = $signed(p2_or_137814_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__506_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137814_comb[23:9], 1'h0};
  assign p2_sel_142755_comb = $signed(p2_prod__48_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__48_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57966_NarrowedMult_, 1'h0};
  assign p2_sel_142756_comb = $signed(p2_or_137819_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__49_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137819_comb[23:10], 2'h0};
  assign p2_sel_142757_comb = $signed(p2_prod__50_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__50_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57970_NarrowedMult_, 1'h0};
  assign p2_sel_142758_comb = $signed(p2_or_137824_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__51_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137824_comb[23:10], 2'h0};
  assign p2_sel_142759_comb = $signed(p2_or_137827_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__52_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137827_comb[23:10], 2'h0};
  assign p2_sel_142760_comb = $signed(p2_prod__53_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__53_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57976_NarrowedMult_, 1'h0};
  assign p2_sel_142761_comb = $signed(p2_or_137832_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__54_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137832_comb[23:10], 2'h0};
  assign p2_sel_142762_comb = $signed(p2_prod__55_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__55_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57980_NarrowedMult_, 1'h0};
  assign p2_sel_142763_comb = $signed(p2_prod__91_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__91_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57982_NarrowedMult_, 1'h0};
  assign p2_sel_142764_comb = $signed(p2_or_137839_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__98_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137839_comb[23:10], 2'h0};
  assign p2_sel_142765_comb = $signed(p2_prod__105_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__105_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57986_NarrowedMult_, 1'h0};
  assign p2_sel_142766_comb = $signed(p2_or_137844_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__111_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137844_comb[23:10], 2'h0};
  assign p2_sel_142767_comb = $signed(p2_or_137847_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__116_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137847_comb[23:10], 2'h0};
  assign p2_sel_142768_comb = $signed(p2_prod__120_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__120_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57992_NarrowedMult_, 1'h0};
  assign p2_sel_142769_comb = $signed(p2_or_137852_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__123_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137852_comb[23:10], 2'h0};
  assign p2_sel_142770_comb = $signed(p2_prod__125_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__125_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57996_NarrowedMult_, 1'h0};
  assign p2_sel_142771_comb = $signed(p2_prod__219_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__219_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58014_NarrowedMult_, 1'h0};
  assign p2_sel_142772_comb = $signed(p2_or_137859_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__226_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137859_comb[23:10], 2'h0};
  assign p2_sel_142773_comb = $signed(p2_prod__233_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__233_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58018_NarrowedMult_, 1'h0};
  assign p2_sel_142774_comb = $signed(p2_or_137864_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__239_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137864_comb[23:10], 2'h0};
  assign p2_sel_142775_comb = $signed(p2_or_137867_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__244_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137867_comb[23:10], 2'h0};
  assign p2_sel_142776_comb = $signed(p2_prod__248_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__248_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58024_NarrowedMult_, 1'h0};
  assign p2_sel_142777_comb = $signed(p2_or_137872_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__251_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137872_comb[23:10], 2'h0};
  assign p2_sel_142778_comb = $signed(p2_prod__253_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__253_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58028_NarrowedMult_, 1'h0};
  assign p2_sel_142779_comb = $signed(p2_prod__283_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__283_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58030_NarrowedMult_, 1'h0};
  assign p2_sel_142780_comb = $signed(p2_or_137879_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__290_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137879_comb[23:10], 2'h0};
  assign p2_sel_142781_comb = $signed(p2_prod__297_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__297_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58034_NarrowedMult_, 1'h0};
  assign p2_sel_142782_comb = $signed(p2_or_137884_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__303_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137884_comb[23:10], 2'h0};
  assign p2_sel_142783_comb = $signed(p2_or_137887_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__308_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137887_comb[23:10], 2'h0};
  assign p2_sel_142784_comb = $signed(p2_prod__312_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__312_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58040_NarrowedMult_, 1'h0};
  assign p2_sel_142785_comb = $signed(p2_or_137892_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__315_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137892_comb[23:10], 2'h0};
  assign p2_sel_142786_comb = $signed(p2_prod__317_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__317_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58044_NarrowedMult_, 1'h0};
  assign p2_sel_142787_comb = $signed(p2_prod__411_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__411_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58062_NarrowedMult_, 1'h0};
  assign p2_sel_142788_comb = $signed(p2_or_137899_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__418_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137899_comb[23:10], 2'h0};
  assign p2_sel_142789_comb = $signed(p2_prod__425_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__425_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58066_NarrowedMult_, 1'h0};
  assign p2_sel_142790_comb = $signed(p2_or_137904_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__431_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137904_comb[23:10], 2'h0};
  assign p2_sel_142791_comb = $signed(p2_or_137907_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__436_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137907_comb[23:10], 2'h0};
  assign p2_sel_142792_comb = $signed(p2_prod__440_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__440_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58072_NarrowedMult_, 1'h0};
  assign p2_sel_142793_comb = $signed(p2_or_137912_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__443_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137912_comb[23:10], 2'h0};
  assign p2_sel_142794_comb = $signed(p2_prod__445_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__445_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58076_NarrowedMult_, 1'h0};
  assign p2_sel_142795_comb = $signed(p2_prod__475_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__475_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58078_NarrowedMult_, 1'h0};
  assign p2_sel_142796_comb = $signed(p2_or_137919_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__482_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137919_comb[23:10], 2'h0};
  assign p2_sel_142797_comb = $signed(p2_prod__489_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__489_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58082_NarrowedMult_, 1'h0};
  assign p2_sel_142798_comb = $signed(p2_or_137924_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__495_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137924_comb[23:10], 2'h0};
  assign p2_sel_142799_comb = $signed(p2_or_137927_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__500_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137927_comb[23:10], 2'h0};
  assign p2_sel_142800_comb = $signed(p2_prod__504_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__504_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58088_NarrowedMult_, 1'h0};
  assign p2_sel_142801_comb = $signed(p2_or_137932_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__507_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p2_or_137932_comb[23:10], 2'h0};
  assign p2_sel_142802_comb = $signed(p2_prod__509_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__509_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58092_NarrowedMult_, 1'h0};
  assign p2_sel_142803_comb = $signed(p2_or_139011_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139011_comb[23:9], 1'h0};
  assign p2_sel_142804_comb = $signed(p2_or_137939_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__57_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137939_comb[23:9], 1'h0};
  assign p2_sel_142805_comb = $signed(p2_smul_58098_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58098_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58098_NarrowedMult__comb[15:0]);
  assign p2_sel_142806_comb = $signed(p2_smul_58100_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58100_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58100_NarrowedMult__comb[15:0]);
  assign p2_sel_142807_comb = $signed(p2_smul_58102_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58102_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58102_NarrowedMult__comb[15:0]);
  assign p2_sel_142808_comb = $signed(p2_smul_58104_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58104_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58104_NarrowedMult__comb[15:0]);
  assign p2_sel_142809_comb = $signed(p2_or_137946_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__62_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137946_comb[23:9], 1'h0};
  assign p2_sel_142810_comb = $signed(p2_or_139026_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139026_comb[23:9], 1'h0};
  assign p2_sel_142811_comb = $signed(p2_or_139027_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139027_comb[23:9], 1'h0};
  assign p2_sel_142812_comb = $signed(p2_or_137953_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__106_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137953_comb[23:9], 1'h0};
  assign p2_sel_142813_comb = $signed(p2_smul_58114_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58114_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58114_NarrowedMult__comb[15:0]);
  assign p2_sel_142814_comb = $signed(p2_smul_58116_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58116_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58116_NarrowedMult__comb[15:0]);
  assign p2_sel_142815_comb = $signed(p2_smul_58118_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58118_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58118_NarrowedMult__comb[15:0]);
  assign p2_sel_142816_comb = $signed(p2_smul_58120_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58120_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58120_NarrowedMult__comb[15:0]);
  assign p2_sel_142817_comb = $signed(p2_or_137960_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__126_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137960_comb[23:9], 1'h0};
  assign p2_sel_142818_comb = $signed(p2_or_139042_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139042_comb[23:9], 1'h0};
  assign p2_sel_142835_comb = $signed(p2_or_139075_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139075_comb[23:9], 1'h0};
  assign p2_sel_142836_comb = $signed(p2_or_137995_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__426_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_137995_comb[23:9], 1'h0};
  assign p2_sel_142837_comb = $signed(p2_smul_58194_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58194_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58194_NarrowedMult__comb[15:0]);
  assign p2_sel_142838_comb = $signed(p2_smul_58196_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58196_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58196_NarrowedMult__comb[15:0]);
  assign p2_sel_142839_comb = $signed(p2_smul_58198_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58198_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58198_NarrowedMult__comb[15:0]);
  assign p2_sel_142840_comb = $signed(p2_smul_58200_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58200_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58200_NarrowedMult__comb[15:0]);
  assign p2_sel_142841_comb = $signed(p2_or_138002_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__446_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_138002_comb[23:9], 1'h0};
  assign p2_sel_142842_comb = $signed(p2_or_139090_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139090_comb[23:9], 1'h0};
  assign p2_sel_142843_comb = $signed(p2_or_139091_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139091_comb[23:9], 1'h0};
  assign p2_sel_142844_comb = $signed(p2_or_138009_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__490_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_138009_comb[23:9], 1'h0};
  assign p2_sel_142845_comb = $signed(p2_smul_58210_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58210_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58210_NarrowedMult__comb[15:0]);
  assign p2_sel_142846_comb = $signed(p2_smul_58212_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58212_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58212_NarrowedMult__comb[15:0]);
  assign p2_sel_142847_comb = $signed(p2_smul_58214_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58214_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58214_NarrowedMult__comb[15:0]);
  assign p2_sel_142848_comb = $signed(p2_smul_58216_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p2_smul_58216_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p2_smul_58216_NarrowedMult__comb[15:0]);
  assign p2_sel_142849_comb = $signed(p2_or_138016_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p2_prod__510_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p2_or_138016_comb[23:9], 1'h0};
  assign p2_sel_142850_comb = $signed(p2_or_139106_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p2_or_139106_comb[23:9], 1'h0};
  assign p2_sum__989_comb = {{15{p2_add_142371_comb[16]}}, p2_add_142371_comb};
  assign p2_sum__990_comb = {{15{p2_add_142372_comb[16]}}, p2_add_142372_comb};
  assign p2_sum__991_comb = {{15{p2_add_142373_comb[16]}}, p2_add_142373_comb};
  assign p2_sum__992_comb = {{15{p2_add_142374_comb[16]}}, p2_add_142374_comb};
  assign p2_sum__884_comb = {{15{p2_add_142375_comb[16]}}, p2_add_142375_comb};
  assign p2_sum__885_comb = {{15{p2_add_142376_comb[16]}}, p2_add_142376_comb};
  assign p2_sum__886_comb = {{15{p2_add_142377_comb[16]}}, p2_add_142377_comb};
  assign p2_sum__887_comb = {{15{p2_add_142378_comb[16]}}, p2_add_142378_comb};
  assign p2_sum__1017_comb = {{15{p2_add_142491_comb[16]}}, p2_add_142491_comb};
  assign p2_sum__1018_comb = {{15{p2_add_142492_comb[16]}}, p2_add_142492_comb};
  assign p2_sum__1019_comb = {{15{p2_add_142493_comb[16]}}, p2_add_142493_comb};
  assign p2_sum__1020_comb = {{15{p2_add_142494_comb[16]}}, p2_add_142494_comb};
  assign p2_sum__1010_comb = {{15{p2_add_142495_comb[16]}}, p2_add_142495_comb};
  assign p2_sum__1011_comb = {{15{p2_add_142496_comb[16]}}, p2_add_142496_comb};
  assign p2_sum__1012_comb = {{15{p2_add_142497_comb[16]}}, p2_add_142497_comb};
  assign p2_sum__1013_comb = {{15{p2_add_142498_comb[16]}}, p2_add_142498_comb};
  assign p2_sum__961_comb = {{15{p2_add_142499_comb[16]}}, p2_add_142499_comb};
  assign p2_sum__962_comb = {{15{p2_add_142500_comb[16]}}, p2_add_142500_comb};
  assign p2_sum__963_comb = {{15{p2_add_142501_comb[16]}}, p2_add_142501_comb};
  assign p2_sum__964_comb = {{15{p2_add_142502_comb[16]}}, p2_add_142502_comb};
  assign p2_sum__926_comb = {{15{p2_add_142503_comb[16]}}, p2_add_142503_comb};
  assign p2_sum__927_comb = {{15{p2_add_142504_comb[16]}}, p2_add_142504_comb};
  assign p2_sum__928_comb = {{15{p2_add_142505_comb[16]}}, p2_add_142505_comb};
  assign p2_sum__929_comb = {{15{p2_add_142506_comb[16]}}, p2_add_142506_comb};
  assign p2_sum__835_comb = {{15{p2_add_142507_comb[16]}}, p2_add_142507_comb};
  assign p2_sum__836_comb = {{15{p2_add_142508_comb[16]}}, p2_add_142508_comb};
  assign p2_sum__837_comb = {{15{p2_add_142509_comb[16]}}, p2_add_142509_comb};
  assign p2_sum__838_comb = {{15{p2_add_142510_comb[16]}}, p2_add_142510_comb};
  assign p2_sum__779_comb = {{15{p2_add_142511_comb[16]}}, p2_add_142511_comb};
  assign p2_sum__780_comb = {{15{p2_add_142512_comb[16]}}, p2_add_142512_comb};
  assign p2_sum__781_comb = {{15{p2_add_142513_comb[16]}}, p2_add_142513_comb};
  assign p2_sum__782_comb = {{15{p2_add_142514_comb[16]}}, p2_add_142514_comb};
  assign p2_add_143359_comb = {{1{p2_sel_142427_comb[15]}}, p2_sel_142427_comb} + {{1{p2_sel_142428_comb[15]}}, p2_sel_142428_comb};
  assign p2_add_143360_comb = {{1{p2_sel_142429_comb[15]}}, p2_sel_142429_comb} + {{1{p2_sel_142430_comb[15]}}, p2_sel_142430_comb};
  assign p2_add_143361_comb = {{1{p2_sel_142431_comb[15]}}, p2_sel_142431_comb} + {{1{p2_sel_142432_comb[15]}}, p2_sel_142432_comb};
  assign p2_add_143362_comb = {{1{p2_sel_142433_comb[15]}}, p2_sel_142433_comb} + {{1{p2_sel_142434_comb[15]}}, p2_sel_142434_comb};
  assign p2_add_143363_comb = {{1{p2_sel_142435_comb[15]}}, p2_sel_142435_comb} + {{1{p2_sel_142436_comb[15]}}, p2_sel_142436_comb};
  assign p2_add_143364_comb = {{1{p2_sel_142437_comb[15]}}, p2_sel_142437_comb} + {{1{p2_sel_142438_comb[15]}}, p2_sel_142438_comb};
  assign p2_add_143365_comb = {{1{p2_sel_142439_comb[15]}}, p2_sel_142439_comb} + {{1{p2_sel_142440_comb[15]}}, p2_sel_142440_comb};
  assign p2_add_143366_comb = {{1{p2_sel_142441_comb[15]}}, p2_sel_142441_comb} + {{1{p2_sel_142442_comb[15]}}, p2_sel_142442_comb};
  assign p2_add_143475_comb = {{1{p2_sel_142659_comb[15]}}, p2_sel_142659_comb} + {{1{p2_sel_142660_comb[15]}}, p2_sel_142660_comb};
  assign p2_add_143476_comb = {{1{p2_sel_142661_comb[15]}}, p2_sel_142661_comb} + {{1{p2_sel_142662_comb[15]}}, p2_sel_142662_comb};
  assign p2_add_143477_comb = {{1{p2_sel_142663_comb[15]}}, p2_sel_142663_comb} + {{1{p2_sel_142664_comb[15]}}, p2_sel_142664_comb};
  assign p2_add_143478_comb = {{1{p2_sel_142665_comb[15]}}, p2_sel_142665_comb} + {{1{p2_sel_142666_comb[15]}}, p2_sel_142666_comb};
  assign p2_add_143479_comb = {{1{p2_sel_142667_comb[15]}}, p2_sel_142667_comb} + {{1{p2_sel_142668_comb[15]}}, p2_sel_142668_comb};
  assign p2_add_143480_comb = {{1{p2_sel_142669_comb[15]}}, p2_sel_142669_comb} + {{1{p2_sel_142670_comb[15]}}, p2_sel_142670_comb};
  assign p2_add_143481_comb = {{1{p2_sel_142671_comb[15]}}, p2_sel_142671_comb} + {{1{p2_sel_142672_comb[15]}}, p2_sel_142672_comb};
  assign p2_add_143482_comb = {{1{p2_sel_142673_comb[15]}}, p2_sel_142673_comb} + {{1{p2_sel_142674_comb[15]}}, p2_sel_142674_comb};
  assign p2_add_143483_comb = {{1{p2_sel_142675_comb[15]}}, p2_sel_142675_comb} + {{1{p2_sel_142676_comb[15]}}, p2_sel_142676_comb};
  assign p2_add_143484_comb = {{1{p2_sel_142677_comb[15]}}, p2_sel_142677_comb} + {{1{p2_sel_142678_comb[15]}}, p2_sel_142678_comb};
  assign p2_add_143485_comb = {{1{p2_sel_142679_comb[15]}}, p2_sel_142679_comb} + {{1{p2_sel_142680_comb[15]}}, p2_sel_142680_comb};
  assign p2_add_143486_comb = {{1{p2_sel_142681_comb[15]}}, p2_sel_142681_comb} + {{1{p2_sel_142682_comb[15]}}, p2_sel_142682_comb};
  assign p2_add_143487_comb = {{1{p2_sel_142683_comb[15]}}, p2_sel_142683_comb} + {{1{p2_sel_142684_comb[15]}}, p2_sel_142684_comb};
  assign p2_add_143488_comb = {{1{p2_sel_142685_comb[15]}}, p2_sel_142685_comb} + {{1{p2_sel_142686_comb[15]}}, p2_sel_142686_comb};
  assign p2_add_143489_comb = {{1{p2_sel_142687_comb[15]}}, p2_sel_142687_comb} + {{1{p2_sel_142688_comb[15]}}, p2_sel_142688_comb};
  assign p2_add_143490_comb = {{1{p2_sel_142689_comb[15]}}, p2_sel_142689_comb} + {{1{p2_sel_142690_comb[15]}}, p2_sel_142690_comb};
  assign p2_add_143491_comb = {{1{p2_sel_142691_comb[15]}}, p2_sel_142691_comb} + {{1{p2_sel_142692_comb[15]}}, p2_sel_142692_comb};
  assign p2_add_143492_comb = {{1{p2_sel_142693_comb[15]}}, p2_sel_142693_comb} + {{1{p2_sel_142694_comb[15]}}, p2_sel_142694_comb};
  assign p2_add_143493_comb = {{1{p2_sel_142695_comb[15]}}, p2_sel_142695_comb} + {{1{p2_sel_142696_comb[15]}}, p2_sel_142696_comb};
  assign p2_add_143494_comb = {{1{p2_sel_142697_comb[15]}}, p2_sel_142697_comb} + {{1{p2_sel_142698_comb[15]}}, p2_sel_142698_comb};
  assign p2_add_143495_comb = {{1{p2_sel_142699_comb[15]}}, p2_sel_142699_comb} + {{1{p2_sel_142700_comb[15]}}, p2_sel_142700_comb};
  assign p2_add_143496_comb = {{1{p2_sel_142701_comb[15]}}, p2_sel_142701_comb} + {{1{p2_sel_142702_comb[15]}}, p2_sel_142702_comb};
  assign p2_add_143497_comb = {{1{p2_sel_142703_comb[15]}}, p2_sel_142703_comb} + {{1{p2_sel_142704_comb[15]}}, p2_sel_142704_comb};
  assign p2_add_143498_comb = {{1{p2_sel_142705_comb[15]}}, p2_sel_142705_comb} + {{1{p2_sel_142706_comb[15]}}, p2_sel_142706_comb};
  assign p2_sum__993_comb = p2_sum__989_comb + p2_sum__990_comb;
  assign p2_sum__994_comb = p2_sum__991_comb + p2_sum__992_comb;
  assign p2_sum__888_comb = p2_sum__884_comb + p2_sum__885_comb;
  assign p2_sum__889_comb = p2_sum__886_comb + p2_sum__887_comb;
  assign p2_sum__1021_comb = p2_sum__1017_comb + p2_sum__1018_comb;
  assign p2_sum__1022_comb = p2_sum__1019_comb + p2_sum__1020_comb;
  assign p2_sum__1014_comb = p2_sum__1010_comb + p2_sum__1011_comb;
  assign p2_sum__1015_comb = p2_sum__1012_comb + p2_sum__1013_comb;
  assign p2_sum__965_comb = p2_sum__961_comb + p2_sum__962_comb;
  assign p2_sum__966_comb = p2_sum__963_comb + p2_sum__964_comb;
  assign p2_sum__930_comb = p2_sum__926_comb + p2_sum__927_comb;
  assign p2_sum__931_comb = p2_sum__928_comb + p2_sum__929_comb;
  assign p2_sum__839_comb = p2_sum__835_comb + p2_sum__836_comb;
  assign p2_sum__840_comb = p2_sum__837_comb + p2_sum__838_comb;
  assign p2_sum__783_comb = p2_sum__779_comb + p2_sum__780_comb;
  assign p2_sum__784_comb = p2_sum__781_comb + p2_sum__782_comb;
  assign p2_add_143411_comb = {{1{p2_sel_142531_comb[15]}}, p2_sel_142531_comb} + {{1{p2_sel_142532_comb[15]}}, p2_sel_142532_comb};
  assign p2_add_143412_comb = {{1{p2_sel_142533_comb[15]}}, p2_sel_142533_comb} + {{1{p2_sel_142534_comb[15]}}, p2_sel_142534_comb};
  assign p2_add_143413_comb = {{1{p2_sel_142535_comb[15]}}, p2_sel_142535_comb} + {{1{p2_sel_142536_comb[15]}}, p2_sel_142536_comb};
  assign p2_add_143414_comb = {{1{p2_sel_142537_comb[15]}}, p2_sel_142537_comb} + {{1{p2_sel_142538_comb[15]}}, p2_sel_142538_comb};
  assign p2_add_143415_comb = {{1{p2_sel_142539_comb[15]}}, p2_sel_142539_comb} + {{1{p2_sel_142540_comb[15]}}, p2_sel_142540_comb};
  assign p2_add_143416_comb = {{1{p2_sel_142541_comb[15]}}, p2_sel_142541_comb} + {{1{p2_sel_142542_comb[15]}}, p2_sel_142542_comb};
  assign p2_add_143417_comb = {{1{p2_sel_142543_comb[15]}}, p2_sel_142543_comb} + {{1{p2_sel_142544_comb[15]}}, p2_sel_142544_comb};
  assign p2_add_143418_comb = {{1{p2_sel_142545_comb[15]}}, p2_sel_142545_comb} + {{1{p2_sel_142546_comb[15]}}, p2_sel_142546_comb};
  assign p2_add_143459_comb = {{1{p2_sel_142627_comb[15]}}, p2_sel_142627_comb} + {{1{p2_sel_142628_comb[15]}}, p2_sel_142628_comb};
  assign p2_add_143460_comb = {{1{p2_sel_142629_comb[15]}}, p2_sel_142629_comb} + {{1{p2_sel_142630_comb[15]}}, p2_sel_142630_comb};
  assign p2_add_143461_comb = {{1{p2_sel_142631_comb[15]}}, p2_sel_142631_comb} + {{1{p2_sel_142632_comb[15]}}, p2_sel_142632_comb};
  assign p2_add_143462_comb = {{1{p2_sel_142633_comb[15]}}, p2_sel_142633_comb} + {{1{p2_sel_142634_comb[15]}}, p2_sel_142634_comb};
  assign p2_add_143463_comb = {{1{p2_sel_142635_comb[15]}}, p2_sel_142635_comb} + {{1{p2_sel_142636_comb[15]}}, p2_sel_142636_comb};
  assign p2_add_143464_comb = {{1{p2_sel_142637_comb[15]}}, p2_sel_142637_comb} + {{1{p2_sel_142638_comb[15]}}, p2_sel_142638_comb};
  assign p2_add_143465_comb = {{1{p2_sel_142639_comb[15]}}, p2_sel_142639_comb} + {{1{p2_sel_142640_comb[15]}}, p2_sel_142640_comb};
  assign p2_add_143466_comb = {{1{p2_sel_142641_comb[15]}}, p2_sel_142641_comb} + {{1{p2_sel_142642_comb[15]}}, p2_sel_142642_comb};
  assign p2_add_143507_comb = {{1{p2_sel_142723_comb[15]}}, p2_sel_142723_comb} + {{1{p2_sel_142724_comb[15]}}, p2_sel_142724_comb};
  assign p2_add_143508_comb = {{1{p2_sel_142725_comb[15]}}, p2_sel_142725_comb} + {{1{p2_sel_142726_comb[15]}}, p2_sel_142726_comb};
  assign p2_add_143509_comb = {{1{p2_sel_142727_comb[15]}}, p2_sel_142727_comb} + {{1{p2_sel_142728_comb[15]}}, p2_sel_142728_comb};
  assign p2_add_143510_comb = {{1{p2_sel_142729_comb[15]}}, p2_sel_142729_comb} + {{1{p2_sel_142730_comb[15]}}, p2_sel_142730_comb};
  assign p2_add_143511_comb = {{1{p2_sel_142731_comb[15]}}, p2_sel_142731_comb} + {{1{p2_sel_142732_comb[15]}}, p2_sel_142732_comb};
  assign p2_add_143512_comb = {{1{p2_sel_142733_comb[15]}}, p2_sel_142733_comb} + {{1{p2_sel_142734_comb[15]}}, p2_sel_142734_comb};
  assign p2_add_143513_comb = {{1{p2_sel_142735_comb[15]}}, p2_sel_142735_comb} + {{1{p2_sel_142736_comb[15]}}, p2_sel_142736_comb};
  assign p2_add_143514_comb = {{1{p2_sel_142737_comb[15]}}, p2_sel_142737_comb} + {{1{p2_sel_142738_comb[15]}}, p2_sel_142738_comb};
  assign p2_add_143555_comb = {{1{p2_sel_142819_comb[15]}}, p2_sel_142819_comb} + {{1{p2_sel_142820_comb[15]}}, p2_sel_142820_comb};
  assign p2_add_143556_comb = {{1{p2_sel_142821_comb[15]}}, p2_sel_142821_comb} + {{1{p2_sel_142822_comb[15]}}, p2_sel_142822_comb};
  assign p2_add_143557_comb = {{1{p2_sel_142823_comb[15]}}, p2_sel_142823_comb} + {{1{p2_sel_142824_comb[15]}}, p2_sel_142824_comb};
  assign p2_add_143558_comb = {{1{p2_sel_142825_comb[15]}}, p2_sel_142825_comb} + {{1{p2_sel_142826_comb[15]}}, p2_sel_142826_comb};
  assign p2_add_143559_comb = {{1{p2_sel_142827_comb[15]}}, p2_sel_142827_comb} + {{1{p2_sel_142828_comb[15]}}, p2_sel_142828_comb};
  assign p2_add_143560_comb = {{1{p2_sel_142829_comb[15]}}, p2_sel_142829_comb} + {{1{p2_sel_142830_comb[15]}}, p2_sel_142830_comb};
  assign p2_add_143561_comb = {{1{p2_sel_142831_comb[15]}}, p2_sel_142831_comb} + {{1{p2_sel_142832_comb[15]}}, p2_sel_142832_comb};
  assign p2_add_143562_comb = {{1{p2_sel_142833_comb[15]}}, p2_sel_142833_comb} + {{1{p2_sel_142834_comb[15]}}, p2_sel_142834_comb};
  assign p2_sum__1736_comb = {{8{p2_add_143359_comb[16]}}, p2_add_143359_comb};
  assign p2_sum__1737_comb = {{8{p2_add_143360_comb[16]}}, p2_add_143360_comb};
  assign p2_sum__1738_comb = {{8{p2_add_143361_comb[16]}}, p2_add_143361_comb};
  assign p2_sum__1739_comb = {{8{p2_add_143362_comb[16]}}, p2_add_143362_comb};
  assign p2_sum__1652_comb = {{8{p2_add_143363_comb[16]}}, p2_add_143363_comb};
  assign p2_sum__1653_comb = {{8{p2_add_143364_comb[16]}}, p2_add_143364_comb};
  assign p2_sum__1654_comb = {{8{p2_add_143365_comb[16]}}, p2_add_143365_comb};
  assign p2_sum__1655_comb = {{8{p2_add_143366_comb[16]}}, p2_add_143366_comb};
  assign p2_sum__1780_comb = {{8{p2_add_143475_comb[16]}}, p2_add_143475_comb};
  assign p2_sum__1781_comb = {{8{p2_add_143476_comb[16]}}, p2_add_143476_comb};
  assign p2_sum__1782_comb = {{8{p2_add_143477_comb[16]}}, p2_add_143477_comb};
  assign p2_sum__1783_comb = {{8{p2_add_143478_comb[16]}}, p2_add_143478_comb};
  assign p2_sum__1760_comb = {{8{p2_add_143479_comb[16]}}, p2_add_143479_comb};
  assign p2_sum__1761_comb = {{8{p2_add_143480_comb[16]}}, p2_add_143480_comb};
  assign p2_sum__1762_comb = {{8{p2_add_143481_comb[16]}}, p2_add_143481_comb};
  assign p2_sum__1763_comb = {{8{p2_add_143482_comb[16]}}, p2_add_143482_comb};
  assign p2_sum__1708_comb = {{8{p2_add_143483_comb[16]}}, p2_add_143483_comb};
  assign p2_sum__1709_comb = {{8{p2_add_143484_comb[16]}}, p2_add_143484_comb};
  assign p2_sum__1710_comb = {{8{p2_add_143485_comb[16]}}, p2_add_143485_comb};
  assign p2_sum__1711_comb = {{8{p2_add_143486_comb[16]}}, p2_add_143486_comb};
  assign p2_sum__1680_comb = {{8{p2_add_143487_comb[16]}}, p2_add_143487_comb};
  assign p2_sum__1681_comb = {{8{p2_add_143488_comb[16]}}, p2_add_143488_comb};
  assign p2_sum__1682_comb = {{8{p2_add_143489_comb[16]}}, p2_add_143489_comb};
  assign p2_sum__1683_comb = {{8{p2_add_143490_comb[16]}}, p2_add_143490_comb};
  assign p2_sum__1628_comb = {{8{p2_add_143491_comb[16]}}, p2_add_143491_comb};
  assign p2_sum__1629_comb = {{8{p2_add_143492_comb[16]}}, p2_add_143492_comb};
  assign p2_sum__1630_comb = {{8{p2_add_143493_comb[16]}}, p2_add_143493_comb};
  assign p2_sum__1631_comb = {{8{p2_add_143494_comb[16]}}, p2_add_143494_comb};
  assign p2_sum__1608_comb = {{8{p2_add_143495_comb[16]}}, p2_add_143495_comb};
  assign p2_sum__1609_comb = {{8{p2_add_143496_comb[16]}}, p2_add_143496_comb};
  assign p2_sum__1610_comb = {{8{p2_add_143497_comb[16]}}, p2_add_143497_comb};
  assign p2_sum__1611_comb = {{8{p2_add_143498_comb[16]}}, p2_add_143498_comb};
  assign p2_add_143335_comb = {{1{p2_sel_142379_comb[15]}}, p2_sel_142379_comb} + {{1{p2_sel_142380_comb[15]}}, p2_sel_142380_comb};
  assign p2_add_143336_comb = {{1{p2_sel_142381_comb[15]}}, p2_sel_142381_comb} + {{1{p2_sel_142382_comb[15]}}, p2_sel_142382_comb};
  assign p2_add_143337_comb = {{1{p2_sel_142383_comb[15]}}, p2_sel_142383_comb} + {{1{p2_sel_142384_comb[15]}}, p2_sel_142384_comb};
  assign p2_add_143338_comb = {{1{p2_sel_142385_comb[15]}}, p2_sel_142385_comb} + {{1{p2_sel_142386_comb[15]}}, p2_sel_142386_comb};
  assign p2_add_143339_comb = {{1{p2_sel_142387_comb[15]}}, p2_sel_142387_comb} + {{1{p2_sel_142388_comb[15]}}, p2_sel_142388_comb};
  assign p2_add_143340_comb = {{1{p2_sel_142389_comb[15]}}, p2_sel_142389_comb} + {{1{p2_sel_142390_comb[15]}}, p2_sel_142390_comb};
  assign p2_add_143341_comb = {{1{p2_sel_142391_comb[15]}}, p2_sel_142391_comb} + {{1{p2_sel_142392_comb[15]}}, p2_sel_142392_comb};
  assign p2_add_143342_comb = {{1{p2_sel_142393_comb[15]}}, p2_sel_142393_comb} + {{1{p2_sel_142394_comb[15]}}, p2_sel_142394_comb};
  assign p2_add_143343_comb = {{1{p2_sel_142395_comb[15]}}, p2_sel_142395_comb} + {{1{p2_sel_142396_comb[15]}}, p2_sel_142396_comb};
  assign p2_add_143344_comb = {{1{p2_sel_142397_comb[15]}}, p2_sel_142397_comb} + {{1{p2_sel_142398_comb[15]}}, p2_sel_142398_comb};
  assign p2_add_143345_comb = {{1{p2_sel_142399_comb[15]}}, p2_sel_142399_comb} + {{1{p2_sel_142400_comb[15]}}, p2_sel_142400_comb};
  assign p2_add_143346_comb = {{1{p2_sel_142401_comb[15]}}, p2_sel_142401_comb} + {{1{p2_sel_142402_comb[15]}}, p2_sel_142402_comb};
  assign p2_add_143347_comb = {{1{p2_sel_142403_comb[15]}}, p2_sel_142403_comb} + {{1{p2_sel_142404_comb[15]}}, p2_sel_142404_comb};
  assign p2_add_143348_comb = {{1{p2_sel_142405_comb[15]}}, p2_sel_142405_comb} + {{1{p2_sel_142406_comb[15]}}, p2_sel_142406_comb};
  assign p2_add_143349_comb = {{1{p2_sel_142407_comb[15]}}, p2_sel_142407_comb} + {{1{p2_sel_142408_comb[15]}}, p2_sel_142408_comb};
  assign p2_add_143350_comb = {{1{p2_sel_142409_comb[15]}}, p2_sel_142409_comb} + {{1{p2_sel_142410_comb[15]}}, p2_sel_142410_comb};
  assign p2_add_143351_comb = {{1{p2_sel_142411_comb[15]}}, p2_sel_142411_comb} + {{1{p2_sel_142412_comb[15]}}, p2_sel_142412_comb};
  assign p2_add_143352_comb = {{1{p2_sel_142413_comb[15]}}, p2_sel_142413_comb} + {{1{p2_sel_142414_comb[15]}}, p2_sel_142414_comb};
  assign p2_add_143353_comb = {{1{p2_sel_142415_comb[15]}}, p2_sel_142415_comb} + {{1{p2_sel_142416_comb[15]}}, p2_sel_142416_comb};
  assign p2_add_143354_comb = {{1{p2_sel_142417_comb[15]}}, p2_sel_142417_comb} + {{1{p2_sel_142418_comb[15]}}, p2_sel_142418_comb};
  assign p2_add_143355_comb = {{1{p2_sel_142419_comb[15]}}, p2_sel_142419_comb} + {{1{p2_sel_142420_comb[15]}}, p2_sel_142420_comb};
  assign p2_add_143356_comb = {{1{p2_sel_142421_comb[15]}}, p2_sel_142421_comb} + {{1{p2_sel_142422_comb[15]}}, p2_sel_142422_comb};
  assign p2_add_143357_comb = {{1{p2_sel_142423_comb[15]}}, p2_sel_142423_comb} + {{1{p2_sel_142424_comb[15]}}, p2_sel_142424_comb};
  assign p2_add_143358_comb = {{1{p2_sel_142425_comb[15]}}, p2_sel_142425_comb} + {{1{p2_sel_142426_comb[15]}}, p2_sel_142426_comb};
  assign p2_add_143367_comb = {{1{p2_sel_142443_comb[15]}}, p2_sel_142443_comb} + {{1{p2_sel_142444_comb[15]}}, p2_sel_142444_comb};
  assign p2_add_143368_comb = {{1{p2_sel_142445_comb[15]}}, p2_sel_142445_comb} + {{1{p2_sel_142446_comb[15]}}, p2_sel_142446_comb};
  assign p2_add_143369_comb = {{1{p2_sel_142447_comb[15]}}, p2_sel_142447_comb} + {{1{p2_sel_142448_comb[15]}}, p2_sel_142448_comb};
  assign p2_add_143370_comb = {{1{p2_sel_142449_comb[15]}}, p2_sel_142449_comb} + {{1{p2_sel_142450_comb[15]}}, p2_sel_142450_comb};
  assign p2_add_143371_comb = {{1{p2_sel_142451_comb[15]}}, p2_sel_142451_comb} + {{1{p2_sel_142452_comb[15]}}, p2_sel_142452_comb};
  assign p2_add_143372_comb = {{1{p2_sel_142453_comb[15]}}, p2_sel_142453_comb} + {{1{p2_sel_142454_comb[15]}}, p2_sel_142454_comb};
  assign p2_add_143373_comb = {{1{p2_sel_142455_comb[15]}}, p2_sel_142455_comb} + {{1{p2_sel_142456_comb[15]}}, p2_sel_142456_comb};
  assign p2_add_143374_comb = {{1{p2_sel_142457_comb[15]}}, p2_sel_142457_comb} + {{1{p2_sel_142458_comb[15]}}, p2_sel_142458_comb};
  assign p2_add_143375_comb = {{1{p2_sel_142459_comb[15]}}, p2_sel_142459_comb} + {{1{p2_sel_142460_comb[15]}}, p2_sel_142460_comb};
  assign p2_add_143376_comb = {{1{p2_sel_142461_comb[15]}}, p2_sel_142461_comb} + {{1{p2_sel_142462_comb[15]}}, p2_sel_142462_comb};
  assign p2_add_143377_comb = {{1{p2_sel_142463_comb[15]}}, p2_sel_142463_comb} + {{1{p2_sel_142464_comb[15]}}, p2_sel_142464_comb};
  assign p2_add_143378_comb = {{1{p2_sel_142465_comb[15]}}, p2_sel_142465_comb} + {{1{p2_sel_142466_comb[15]}}, p2_sel_142466_comb};
  assign p2_add_143379_comb = {{1{p2_sel_142467_comb[15]}}, p2_sel_142467_comb} + {{1{p2_sel_142468_comb[15]}}, p2_sel_142468_comb};
  assign p2_add_143380_comb = {{1{p2_sel_142469_comb[15]}}, p2_sel_142469_comb} + {{1{p2_sel_142470_comb[15]}}, p2_sel_142470_comb};
  assign p2_add_143381_comb = {{1{p2_sel_142471_comb[15]}}, p2_sel_142471_comb} + {{1{p2_sel_142472_comb[15]}}, p2_sel_142472_comb};
  assign p2_add_143382_comb = {{1{p2_sel_142473_comb[15]}}, p2_sel_142473_comb} + {{1{p2_sel_142474_comb[15]}}, p2_sel_142474_comb};
  assign p2_add_143383_comb = {{1{p2_sel_142475_comb[15]}}, p2_sel_142475_comb} + {{1{p2_sel_142476_comb[15]}}, p2_sel_142476_comb};
  assign p2_add_143384_comb = {{1{p2_sel_142477_comb[15]}}, p2_sel_142477_comb} + {{1{p2_sel_142478_comb[15]}}, p2_sel_142478_comb};
  assign p2_add_143385_comb = {{1{p2_sel_142479_comb[15]}}, p2_sel_142479_comb} + {{1{p2_sel_142480_comb[15]}}, p2_sel_142480_comb};
  assign p2_add_143386_comb = {{1{p2_sel_142481_comb[15]}}, p2_sel_142481_comb} + {{1{p2_sel_142482_comb[15]}}, p2_sel_142482_comb};
  assign p2_add_143387_comb = {{1{p2_sel_142483_comb[15]}}, p2_sel_142483_comb} + {{1{p2_sel_142484_comb[15]}}, p2_sel_142484_comb};
  assign p2_add_143388_comb = {{1{p2_sel_142485_comb[15]}}, p2_sel_142485_comb} + {{1{p2_sel_142486_comb[15]}}, p2_sel_142486_comb};
  assign p2_add_143389_comb = {{1{p2_sel_142487_comb[15]}}, p2_sel_142487_comb} + {{1{p2_sel_142488_comb[15]}}, p2_sel_142488_comb};
  assign p2_add_143390_comb = {{1{p2_sel_142489_comb[15]}}, p2_sel_142489_comb} + {{1{p2_sel_142490_comb[15]}}, p2_sel_142490_comb};
  assign p2_add_143403_comb = {{1{p2_sel_142515_comb[15]}}, p2_sel_142515_comb} + {{1{p2_sel_142516_comb[15]}}, p2_sel_142516_comb};
  assign p2_add_143404_comb = {{1{p2_sel_142517_comb[15]}}, p2_sel_142517_comb} + {{1{p2_sel_142518_comb[15]}}, p2_sel_142518_comb};
  assign p2_add_143405_comb = {{1{p2_sel_142519_comb[15]}}, p2_sel_142519_comb} + {{1{p2_sel_142520_comb[15]}}, p2_sel_142520_comb};
  assign p2_add_143406_comb = {{1{p2_sel_142521_comb[15]}}, p2_sel_142521_comb} + {{1{p2_sel_142522_comb[15]}}, p2_sel_142522_comb};
  assign p2_add_143407_comb = {{1{p2_sel_142523_comb[15]}}, p2_sel_142523_comb} + {{1{p2_sel_142524_comb[15]}}, p2_sel_142524_comb};
  assign p2_add_143408_comb = {{1{p2_sel_142525_comb[15]}}, p2_sel_142525_comb} + {{1{p2_sel_142526_comb[15]}}, p2_sel_142526_comb};
  assign p2_add_143409_comb = {{1{p2_sel_142527_comb[15]}}, p2_sel_142527_comb} + {{1{p2_sel_142528_comb[15]}}, p2_sel_142528_comb};
  assign p2_add_143410_comb = {{1{p2_sel_142529_comb[15]}}, p2_sel_142529_comb} + {{1{p2_sel_142530_comb[15]}}, p2_sel_142530_comb};
  assign p2_add_143419_comb = {{1{p2_sel_142547_comb[15]}}, p2_sel_142547_comb} + {{1{p2_sel_142548_comb[15]}}, p2_sel_142548_comb};
  assign p2_add_143420_comb = {{1{p2_sel_142549_comb[15]}}, p2_sel_142549_comb} + {{1{p2_sel_142550_comb[15]}}, p2_sel_142550_comb};
  assign p2_add_143421_comb = {{1{p2_sel_142551_comb[15]}}, p2_sel_142551_comb} + {{1{p2_sel_142552_comb[15]}}, p2_sel_142552_comb};
  assign p2_add_143422_comb = {{1{p2_sel_142553_comb[15]}}, p2_sel_142553_comb} + {{1{p2_sel_142554_comb[15]}}, p2_sel_142554_comb};
  assign p2_add_143423_comb = {{1{p2_sel_142555_comb[15]}}, p2_sel_142555_comb} + {{1{p2_sel_142556_comb[15]}}, p2_sel_142556_comb};
  assign p2_add_143424_comb = {{1{p2_sel_142557_comb[15]}}, p2_sel_142557_comb} + {{1{p2_sel_142558_comb[15]}}, p2_sel_142558_comb};
  assign p2_add_143425_comb = {{1{p2_sel_142559_comb[15]}}, p2_sel_142559_comb} + {{1{p2_sel_142560_comb[15]}}, p2_sel_142560_comb};
  assign p2_add_143426_comb = {{1{p2_sel_142561_comb[15]}}, p2_sel_142561_comb} + {{1{p2_sel_142562_comb[15]}}, p2_sel_142562_comb};
  assign p2_add_143427_comb = {{1{p2_sel_142563_comb[15]}}, p2_sel_142563_comb} + {{1{p2_sel_142564_comb[15]}}, p2_sel_142564_comb};
  assign p2_add_143428_comb = {{1{p2_sel_142565_comb[15]}}, p2_sel_142565_comb} + {{1{p2_sel_142566_comb[15]}}, p2_sel_142566_comb};
  assign p2_add_143429_comb = {{1{p2_sel_142567_comb[15]}}, p2_sel_142567_comb} + {{1{p2_sel_142568_comb[15]}}, p2_sel_142568_comb};
  assign p2_add_143430_comb = {{1{p2_sel_142569_comb[15]}}, p2_sel_142569_comb} + {{1{p2_sel_142570_comb[15]}}, p2_sel_142570_comb};
  assign p2_add_143431_comb = {{1{p2_sel_142571_comb[15]}}, p2_sel_142571_comb} + {{1{p2_sel_142572_comb[15]}}, p2_sel_142572_comb};
  assign p2_add_143432_comb = {{1{p2_sel_142573_comb[15]}}, p2_sel_142573_comb} + {{1{p2_sel_142574_comb[15]}}, p2_sel_142574_comb};
  assign p2_add_143433_comb = {{1{p2_sel_142575_comb[15]}}, p2_sel_142575_comb} + {{1{p2_sel_142576_comb[15]}}, p2_sel_142576_comb};
  assign p2_add_143434_comb = {{1{p2_sel_142577_comb[15]}}, p2_sel_142577_comb} + {{1{p2_sel_142578_comb[15]}}, p2_sel_142578_comb};
  assign p2_add_143435_comb = {{1{p2_sel_142579_comb[15]}}, p2_sel_142579_comb} + {{1{p2_sel_142580_comb[15]}}, p2_sel_142580_comb};
  assign p2_add_143436_comb = {{1{p2_sel_142581_comb[15]}}, p2_sel_142581_comb} + {{1{p2_sel_142582_comb[15]}}, p2_sel_142582_comb};
  assign p2_add_143437_comb = {{1{p2_sel_142583_comb[15]}}, p2_sel_142583_comb} + {{1{p2_sel_142584_comb[15]}}, p2_sel_142584_comb};
  assign p2_add_143438_comb = {{1{p2_sel_142585_comb[15]}}, p2_sel_142585_comb} + {{1{p2_sel_142586_comb[15]}}, p2_sel_142586_comb};
  assign p2_add_143439_comb = {{1{p2_sel_142587_comb[15]}}, p2_sel_142587_comb} + {{1{p2_sel_142588_comb[15]}}, p2_sel_142588_comb};
  assign p2_add_143440_comb = {{1{p2_sel_142589_comb[15]}}, p2_sel_142589_comb} + {{1{p2_sel_142590_comb[15]}}, p2_sel_142590_comb};
  assign p2_add_143441_comb = {{1{p2_sel_142591_comb[15]}}, p2_sel_142591_comb} + {{1{p2_sel_142592_comb[15]}}, p2_sel_142592_comb};
  assign p2_add_143442_comb = {{1{p2_sel_142593_comb[15]}}, p2_sel_142593_comb} + {{1{p2_sel_142594_comb[15]}}, p2_sel_142594_comb};
  assign p2_add_143443_comb = {{1{p2_sel_142595_comb[15]}}, p2_sel_142595_comb} + {{1{p2_sel_142596_comb[15]}}, p2_sel_142596_comb};
  assign p2_add_143444_comb = {{1{p2_sel_142597_comb[15]}}, p2_sel_142597_comb} + {{1{p2_sel_142598_comb[15]}}, p2_sel_142598_comb};
  assign p2_add_143445_comb = {{1{p2_sel_142599_comb[15]}}, p2_sel_142599_comb} + {{1{p2_sel_142600_comb[15]}}, p2_sel_142600_comb};
  assign p2_add_143446_comb = {{1{p2_sel_142601_comb[15]}}, p2_sel_142601_comb} + {{1{p2_sel_142602_comb[15]}}, p2_sel_142602_comb};
  assign p2_add_143447_comb = {{1{p2_sel_142603_comb[15]}}, p2_sel_142603_comb} + {{1{p2_sel_142604_comb[15]}}, p2_sel_142604_comb};
  assign p2_add_143448_comb = {{1{p2_sel_142605_comb[15]}}, p2_sel_142605_comb} + {{1{p2_sel_142606_comb[15]}}, p2_sel_142606_comb};
  assign p2_add_143449_comb = {{1{p2_sel_142607_comb[15]}}, p2_sel_142607_comb} + {{1{p2_sel_142608_comb[15]}}, p2_sel_142608_comb};
  assign p2_add_143450_comb = {{1{p2_sel_142609_comb[15]}}, p2_sel_142609_comb} + {{1{p2_sel_142610_comb[15]}}, p2_sel_142610_comb};
  assign p2_add_143451_comb = {{1{p2_sel_142611_comb[15]}}, p2_sel_142611_comb} + {{1{p2_sel_142612_comb[15]}}, p2_sel_142612_comb};
  assign p2_add_143452_comb = {{1{p2_sel_142613_comb[15]}}, p2_sel_142613_comb} + {{1{p2_sel_142614_comb[15]}}, p2_sel_142614_comb};
  assign p2_add_143453_comb = {{1{p2_sel_142615_comb[15]}}, p2_sel_142615_comb} + {{1{p2_sel_142616_comb[15]}}, p2_sel_142616_comb};
  assign p2_add_143454_comb = {{1{p2_sel_142617_comb[15]}}, p2_sel_142617_comb} + {{1{p2_sel_142618_comb[15]}}, p2_sel_142618_comb};
  assign p2_add_143455_comb = {{1{p2_sel_142619_comb[15]}}, p2_sel_142619_comb} + {{1{p2_sel_142620_comb[15]}}, p2_sel_142620_comb};
  assign p2_add_143456_comb = {{1{p2_sel_142621_comb[15]}}, p2_sel_142621_comb} + {{1{p2_sel_142622_comb[15]}}, p2_sel_142622_comb};
  assign p2_add_143457_comb = {{1{p2_sel_142623_comb[15]}}, p2_sel_142623_comb} + {{1{p2_sel_142624_comb[15]}}, p2_sel_142624_comb};
  assign p2_add_143458_comb = {{1{p2_sel_142625_comb[15]}}, p2_sel_142625_comb} + {{1{p2_sel_142626_comb[15]}}, p2_sel_142626_comb};
  assign p2_add_143467_comb = {{1{p2_sel_142643_comb[15]}}, p2_sel_142643_comb} + {{1{p2_sel_142644_comb[15]}}, p2_sel_142644_comb};
  assign p2_add_143468_comb = {{1{p2_sel_142645_comb[15]}}, p2_sel_142645_comb} + {{1{p2_sel_142646_comb[15]}}, p2_sel_142646_comb};
  assign p2_add_143469_comb = {{1{p2_sel_142647_comb[15]}}, p2_sel_142647_comb} + {{1{p2_sel_142648_comb[15]}}, p2_sel_142648_comb};
  assign p2_add_143470_comb = {{1{p2_sel_142649_comb[15]}}, p2_sel_142649_comb} + {{1{p2_sel_142650_comb[15]}}, p2_sel_142650_comb};
  assign p2_add_143471_comb = {{1{p2_sel_142651_comb[15]}}, p2_sel_142651_comb} + {{1{p2_sel_142652_comb[15]}}, p2_sel_142652_comb};
  assign p2_add_143472_comb = {{1{p2_sel_142653_comb[15]}}, p2_sel_142653_comb} + {{1{p2_sel_142654_comb[15]}}, p2_sel_142654_comb};
  assign p2_add_143473_comb = {{1{p2_sel_142655_comb[15]}}, p2_sel_142655_comb} + {{1{p2_sel_142656_comb[15]}}, p2_sel_142656_comb};
  assign p2_add_143474_comb = {{1{p2_sel_142657_comb[15]}}, p2_sel_142657_comb} + {{1{p2_sel_142658_comb[15]}}, p2_sel_142658_comb};
  assign p2_add_143499_comb = {{1{p2_sel_142707_comb[15]}}, p2_sel_142707_comb} + {{1{p2_sel_142708_comb[15]}}, p2_sel_142708_comb};
  assign p2_add_143500_comb = {{1{p2_sel_142709_comb[15]}}, p2_sel_142709_comb} + {{1{p2_sel_142710_comb[15]}}, p2_sel_142710_comb};
  assign p2_add_143501_comb = {{1{p2_sel_142711_comb[15]}}, p2_sel_142711_comb} + {{1{p2_sel_142712_comb[15]}}, p2_sel_142712_comb};
  assign p2_add_143502_comb = {{1{p2_sel_142713_comb[15]}}, p2_sel_142713_comb} + {{1{p2_sel_142714_comb[15]}}, p2_sel_142714_comb};
  assign p2_add_143503_comb = {{1{p2_sel_142715_comb[15]}}, p2_sel_142715_comb} + {{1{p2_sel_142716_comb[15]}}, p2_sel_142716_comb};
  assign p2_add_143504_comb = {{1{p2_sel_142717_comb[15]}}, p2_sel_142717_comb} + {{1{p2_sel_142718_comb[15]}}, p2_sel_142718_comb};
  assign p2_add_143505_comb = {{1{p2_sel_142719_comb[15]}}, p2_sel_142719_comb} + {{1{p2_sel_142720_comb[15]}}, p2_sel_142720_comb};
  assign p2_add_143506_comb = {{1{p2_sel_142721_comb[15]}}, p2_sel_142721_comb} + {{1{p2_sel_142722_comb[15]}}, p2_sel_142722_comb};
  assign p2_add_143515_comb = {{1{p2_sel_142739_comb[15]}}, p2_sel_142739_comb} + {{1{p2_sel_142740_comb[15]}}, p2_sel_142740_comb};
  assign p2_add_143516_comb = {{1{p2_sel_142741_comb[15]}}, p2_sel_142741_comb} + {{1{p2_sel_142742_comb[15]}}, p2_sel_142742_comb};
  assign p2_add_143517_comb = {{1{p2_sel_142743_comb[15]}}, p2_sel_142743_comb} + {{1{p2_sel_142744_comb[15]}}, p2_sel_142744_comb};
  assign p2_add_143518_comb = {{1{p2_sel_142745_comb[15]}}, p2_sel_142745_comb} + {{1{p2_sel_142746_comb[15]}}, p2_sel_142746_comb};
  assign p2_add_143519_comb = {{1{p2_sel_142747_comb[15]}}, p2_sel_142747_comb} + {{1{p2_sel_142748_comb[15]}}, p2_sel_142748_comb};
  assign p2_add_143520_comb = {{1{p2_sel_142749_comb[15]}}, p2_sel_142749_comb} + {{1{p2_sel_142750_comb[15]}}, p2_sel_142750_comb};
  assign p2_add_143521_comb = {{1{p2_sel_142751_comb[15]}}, p2_sel_142751_comb} + {{1{p2_sel_142752_comb[15]}}, p2_sel_142752_comb};
  assign p2_add_143522_comb = {{1{p2_sel_142753_comb[15]}}, p2_sel_142753_comb} + {{1{p2_sel_142754_comb[15]}}, p2_sel_142754_comb};
  assign p2_add_143523_comb = {{1{p2_sel_142755_comb[15]}}, p2_sel_142755_comb} + {{1{p2_sel_142756_comb[15]}}, p2_sel_142756_comb};
  assign p2_add_143524_comb = {{1{p2_sel_142757_comb[15]}}, p2_sel_142757_comb} + {{1{p2_sel_142758_comb[15]}}, p2_sel_142758_comb};
  assign p2_add_143525_comb = {{1{p2_sel_142759_comb[15]}}, p2_sel_142759_comb} + {{1{p2_sel_142760_comb[15]}}, p2_sel_142760_comb};
  assign p2_add_143526_comb = {{1{p2_sel_142761_comb[15]}}, p2_sel_142761_comb} + {{1{p2_sel_142762_comb[15]}}, p2_sel_142762_comb};
  assign p2_add_143527_comb = {{1{p2_sel_142763_comb[15]}}, p2_sel_142763_comb} + {{1{p2_sel_142764_comb[15]}}, p2_sel_142764_comb};
  assign p2_add_143528_comb = {{1{p2_sel_142765_comb[15]}}, p2_sel_142765_comb} + {{1{p2_sel_142766_comb[15]}}, p2_sel_142766_comb};
  assign p2_add_143529_comb = {{1{p2_sel_142767_comb[15]}}, p2_sel_142767_comb} + {{1{p2_sel_142768_comb[15]}}, p2_sel_142768_comb};
  assign p2_add_143530_comb = {{1{p2_sel_142769_comb[15]}}, p2_sel_142769_comb} + {{1{p2_sel_142770_comb[15]}}, p2_sel_142770_comb};
  assign p2_add_143531_comb = {{1{p2_sel_142771_comb[15]}}, p2_sel_142771_comb} + {{1{p2_sel_142772_comb[15]}}, p2_sel_142772_comb};
  assign p2_add_143532_comb = {{1{p2_sel_142773_comb[15]}}, p2_sel_142773_comb} + {{1{p2_sel_142774_comb[15]}}, p2_sel_142774_comb};
  assign p2_add_143533_comb = {{1{p2_sel_142775_comb[15]}}, p2_sel_142775_comb} + {{1{p2_sel_142776_comb[15]}}, p2_sel_142776_comb};
  assign p2_add_143534_comb = {{1{p2_sel_142777_comb[15]}}, p2_sel_142777_comb} + {{1{p2_sel_142778_comb[15]}}, p2_sel_142778_comb};
  assign p2_add_143535_comb = {{1{p2_sel_142779_comb[15]}}, p2_sel_142779_comb} + {{1{p2_sel_142780_comb[15]}}, p2_sel_142780_comb};
  assign p2_add_143536_comb = {{1{p2_sel_142781_comb[15]}}, p2_sel_142781_comb} + {{1{p2_sel_142782_comb[15]}}, p2_sel_142782_comb};
  assign p2_add_143537_comb = {{1{p2_sel_142783_comb[15]}}, p2_sel_142783_comb} + {{1{p2_sel_142784_comb[15]}}, p2_sel_142784_comb};
  assign p2_add_143538_comb = {{1{p2_sel_142785_comb[15]}}, p2_sel_142785_comb} + {{1{p2_sel_142786_comb[15]}}, p2_sel_142786_comb};
  assign p2_add_143539_comb = {{1{p2_sel_142787_comb[15]}}, p2_sel_142787_comb} + {{1{p2_sel_142788_comb[15]}}, p2_sel_142788_comb};
  assign p2_add_143540_comb = {{1{p2_sel_142789_comb[15]}}, p2_sel_142789_comb} + {{1{p2_sel_142790_comb[15]}}, p2_sel_142790_comb};
  assign p2_add_143541_comb = {{1{p2_sel_142791_comb[15]}}, p2_sel_142791_comb} + {{1{p2_sel_142792_comb[15]}}, p2_sel_142792_comb};
  assign p2_add_143542_comb = {{1{p2_sel_142793_comb[15]}}, p2_sel_142793_comb} + {{1{p2_sel_142794_comb[15]}}, p2_sel_142794_comb};
  assign p2_add_143543_comb = {{1{p2_sel_142795_comb[15]}}, p2_sel_142795_comb} + {{1{p2_sel_142796_comb[15]}}, p2_sel_142796_comb};
  assign p2_add_143544_comb = {{1{p2_sel_142797_comb[15]}}, p2_sel_142797_comb} + {{1{p2_sel_142798_comb[15]}}, p2_sel_142798_comb};
  assign p2_add_143545_comb = {{1{p2_sel_142799_comb[15]}}, p2_sel_142799_comb} + {{1{p2_sel_142800_comb[15]}}, p2_sel_142800_comb};
  assign p2_add_143546_comb = {{1{p2_sel_142801_comb[15]}}, p2_sel_142801_comb} + {{1{p2_sel_142802_comb[15]}}, p2_sel_142802_comb};
  assign p2_add_143547_comb = {{1{p2_sel_142803_comb[15]}}, p2_sel_142803_comb} + {{1{p2_sel_142804_comb[15]}}, p2_sel_142804_comb};
  assign p2_add_143548_comb = {{1{p2_sel_142805_comb[15]}}, p2_sel_142805_comb} + {{1{p2_sel_142806_comb[15]}}, p2_sel_142806_comb};
  assign p2_add_143549_comb = {{1{p2_sel_142807_comb[15]}}, p2_sel_142807_comb} + {{1{p2_sel_142808_comb[15]}}, p2_sel_142808_comb};
  assign p2_add_143550_comb = {{1{p2_sel_142809_comb[15]}}, p2_sel_142809_comb} + {{1{p2_sel_142810_comb[15]}}, p2_sel_142810_comb};
  assign p2_add_143551_comb = {{1{p2_sel_142811_comb[15]}}, p2_sel_142811_comb} + {{1{p2_sel_142812_comb[15]}}, p2_sel_142812_comb};
  assign p2_add_143552_comb = {{1{p2_sel_142813_comb[15]}}, p2_sel_142813_comb} + {{1{p2_sel_142814_comb[15]}}, p2_sel_142814_comb};
  assign p2_add_143553_comb = {{1{p2_sel_142815_comb[15]}}, p2_sel_142815_comb} + {{1{p2_sel_142816_comb[15]}}, p2_sel_142816_comb};
  assign p2_add_143554_comb = {{1{p2_sel_142817_comb[15]}}, p2_sel_142817_comb} + {{1{p2_sel_142818_comb[15]}}, p2_sel_142818_comb};
  assign p2_add_143563_comb = {{1{p2_sel_142835_comb[15]}}, p2_sel_142835_comb} + {{1{p2_sel_142836_comb[15]}}, p2_sel_142836_comb};
  assign p2_add_143564_comb = {{1{p2_sel_142837_comb[15]}}, p2_sel_142837_comb} + {{1{p2_sel_142838_comb[15]}}, p2_sel_142838_comb};
  assign p2_add_143565_comb = {{1{p2_sel_142839_comb[15]}}, p2_sel_142839_comb} + {{1{p2_sel_142840_comb[15]}}, p2_sel_142840_comb};
  assign p2_add_143566_comb = {{1{p2_sel_142841_comb[15]}}, p2_sel_142841_comb} + {{1{p2_sel_142842_comb[15]}}, p2_sel_142842_comb};
  assign p2_add_143567_comb = {{1{p2_sel_142843_comb[15]}}, p2_sel_142843_comb} + {{1{p2_sel_142844_comb[15]}}, p2_sel_142844_comb};
  assign p2_add_143568_comb = {{1{p2_sel_142845_comb[15]}}, p2_sel_142845_comb} + {{1{p2_sel_142846_comb[15]}}, p2_sel_142846_comb};
  assign p2_add_143569_comb = {{1{p2_sel_142847_comb[15]}}, p2_sel_142847_comb} + {{1{p2_sel_142848_comb[15]}}, p2_sel_142848_comb};
  assign p2_add_143570_comb = {{1{p2_sel_142849_comb[15]}}, p2_sel_142849_comb} + {{1{p2_sel_142850_comb[15]}}, p2_sel_142850_comb};
  assign p2_sum__995_comb = p2_sum__993_comb + p2_sum__994_comb;
  assign p2_sum__890_comb = p2_sum__888_comb + p2_sum__889_comb;
  assign p2_sum__1023_comb = p2_sum__1021_comb + p2_sum__1022_comb;
  assign p2_sum__1016_comb = p2_sum__1014_comb + p2_sum__1015_comb;
  assign p2_sum__967_comb = p2_sum__965_comb + p2_sum__966_comb;
  assign p2_sum__932_comb = p2_sum__930_comb + p2_sum__931_comb;
  assign p2_sum__841_comb = p2_sum__839_comb + p2_sum__840_comb;
  assign p2_sum__785_comb = p2_sum__783_comb + p2_sum__784_comb;
  assign p2_sum__1768_comb = {{8{p2_add_143411_comb[16]}}, p2_add_143411_comb};
  assign p2_sum__1769_comb = {{8{p2_add_143412_comb[16]}}, p2_add_143412_comb};
  assign p2_sum__1770_comb = {{8{p2_add_143413_comb[16]}}, p2_add_143413_comb};
  assign p2_sum__1771_comb = {{8{p2_add_143414_comb[16]}}, p2_add_143414_comb};
  assign p2_sum__1748_comb = {{8{p2_add_143415_comb[16]}}, p2_add_143415_comb};
  assign p2_sum__1749_comb = {{8{p2_add_143416_comb[16]}}, p2_add_143416_comb};
  assign p2_sum__1750_comb = {{8{p2_add_143417_comb[16]}}, p2_add_143417_comb};
  assign p2_sum__1751_comb = {{8{p2_add_143418_comb[16]}}, p2_add_143418_comb};
  assign p2_sum__1732_comb = {{8{p2_add_143459_comb[16]}}, p2_add_143459_comb};
  assign p2_sum__1733_comb = {{8{p2_add_143460_comb[16]}}, p2_add_143460_comb};
  assign p2_sum__1734_comb = {{8{p2_add_143461_comb[16]}}, p2_add_143461_comb};
  assign p2_sum__1735_comb = {{8{p2_add_143462_comb[16]}}, p2_add_143462_comb};
  assign p2_sum__1704_comb = {{8{p2_add_143463_comb[16]}}, p2_add_143463_comb};
  assign p2_sum__1705_comb = {{8{p2_add_143464_comb[16]}}, p2_add_143464_comb};
  assign p2_sum__1706_comb = {{8{p2_add_143465_comb[16]}}, p2_add_143465_comb};
  assign p2_sum__1707_comb = {{8{p2_add_143466_comb[16]}}, p2_add_143466_comb};
  assign p2_sum__1684_comb = {{8{p2_add_143507_comb[16]}}, p2_add_143507_comb};
  assign p2_sum__1685_comb = {{8{p2_add_143508_comb[16]}}, p2_add_143508_comb};
  assign p2_sum__1686_comb = {{8{p2_add_143509_comb[16]}}, p2_add_143509_comb};
  assign p2_sum__1687_comb = {{8{p2_add_143510_comb[16]}}, p2_add_143510_comb};
  assign p2_sum__1656_comb = {{8{p2_add_143511_comb[16]}}, p2_add_143511_comb};
  assign p2_sum__1657_comb = {{8{p2_add_143512_comb[16]}}, p2_add_143512_comb};
  assign p2_sum__1658_comb = {{8{p2_add_143513_comb[16]}}, p2_add_143513_comb};
  assign p2_sum__1659_comb = {{8{p2_add_143514_comb[16]}}, p2_add_143514_comb};
  assign p2_sum__1640_comb = {{8{p2_add_143555_comb[16]}}, p2_add_143555_comb};
  assign p2_sum__1641_comb = {{8{p2_add_143556_comb[16]}}, p2_add_143556_comb};
  assign p2_sum__1642_comb = {{8{p2_add_143557_comb[16]}}, p2_add_143557_comb};
  assign p2_sum__1643_comb = {{8{p2_add_143558_comb[16]}}, p2_add_143558_comb};
  assign p2_sum__1620_comb = {{8{p2_add_143559_comb[16]}}, p2_add_143559_comb};
  assign p2_sum__1621_comb = {{8{p2_add_143560_comb[16]}}, p2_add_143560_comb};
  assign p2_sum__1622_comb = {{8{p2_add_143561_comb[16]}}, p2_add_143561_comb};
  assign p2_sum__1623_comb = {{8{p2_add_143562_comb[16]}}, p2_add_143562_comb};
  assign p2_sum__1324_comb = p2_sum__1736_comb + p2_sum__1737_comb;
  assign p2_sum__1325_comb = p2_sum__1738_comb + p2_sum__1739_comb;
  assign p2_sum__1282_comb = p2_sum__1652_comb + p2_sum__1653_comb;
  assign p2_sum__1283_comb = p2_sum__1654_comb + p2_sum__1655_comb;
  assign p2_sum__1346_comb = p2_sum__1780_comb + p2_sum__1781_comb;
  assign p2_sum__1347_comb = p2_sum__1782_comb + p2_sum__1783_comb;
  assign p2_sum__1336_comb = p2_sum__1760_comb + p2_sum__1761_comb;
  assign p2_sum__1337_comb = p2_sum__1762_comb + p2_sum__1763_comb;
  assign p2_sum__1310_comb = p2_sum__1708_comb + p2_sum__1709_comb;
  assign p2_sum__1311_comb = p2_sum__1710_comb + p2_sum__1711_comb;
  assign p2_sum__1296_comb = p2_sum__1680_comb + p2_sum__1681_comb;
  assign p2_sum__1297_comb = p2_sum__1682_comb + p2_sum__1683_comb;
  assign p2_sum__1270_comb = p2_sum__1628_comb + p2_sum__1629_comb;
  assign p2_sum__1271_comb = p2_sum__1630_comb + p2_sum__1631_comb;
  assign p2_sum__1260_comb = p2_sum__1608_comb + p2_sum__1609_comb;
  assign p2_sum__1261_comb = p2_sum__1610_comb + p2_sum__1611_comb;

  // Registers for pipe stage 2:
  reg [16:0] p2_add_143335;
  reg [16:0] p2_add_143336;
  reg [16:0] p2_add_143337;
  reg [16:0] p2_add_143338;
  reg [16:0] p2_add_143339;
  reg [16:0] p2_add_143340;
  reg [16:0] p2_add_143341;
  reg [16:0] p2_add_143342;
  reg [16:0] p2_add_143343;
  reg [16:0] p2_add_143344;
  reg [16:0] p2_add_143345;
  reg [16:0] p2_add_143346;
  reg [16:0] p2_add_143347;
  reg [16:0] p2_add_143348;
  reg [16:0] p2_add_143349;
  reg [16:0] p2_add_143350;
  reg [16:0] p2_add_143351;
  reg [16:0] p2_add_143352;
  reg [16:0] p2_add_143353;
  reg [16:0] p2_add_143354;
  reg [16:0] p2_add_143355;
  reg [16:0] p2_add_143356;
  reg [16:0] p2_add_143357;
  reg [16:0] p2_add_143358;
  reg [16:0] p2_add_143367;
  reg [16:0] p2_add_143368;
  reg [16:0] p2_add_143369;
  reg [16:0] p2_add_143370;
  reg [16:0] p2_add_143371;
  reg [16:0] p2_add_143372;
  reg [16:0] p2_add_143373;
  reg [16:0] p2_add_143374;
  reg [16:0] p2_add_143375;
  reg [16:0] p2_add_143376;
  reg [16:0] p2_add_143377;
  reg [16:0] p2_add_143378;
  reg [16:0] p2_add_143379;
  reg [16:0] p2_add_143380;
  reg [16:0] p2_add_143381;
  reg [16:0] p2_add_143382;
  reg [16:0] p2_add_143383;
  reg [16:0] p2_add_143384;
  reg [16:0] p2_add_143385;
  reg [16:0] p2_add_143386;
  reg [16:0] p2_add_143387;
  reg [16:0] p2_add_143388;
  reg [16:0] p2_add_143389;
  reg [16:0] p2_add_143390;
  reg [16:0] p2_add_143403;
  reg [16:0] p2_add_143404;
  reg [16:0] p2_add_143405;
  reg [16:0] p2_add_143406;
  reg [16:0] p2_add_143407;
  reg [16:0] p2_add_143408;
  reg [16:0] p2_add_143409;
  reg [16:0] p2_add_143410;
  reg [16:0] p2_add_143419;
  reg [16:0] p2_add_143420;
  reg [16:0] p2_add_143421;
  reg [16:0] p2_add_143422;
  reg [16:0] p2_add_143423;
  reg [16:0] p2_add_143424;
  reg [16:0] p2_add_143425;
  reg [16:0] p2_add_143426;
  reg [16:0] p2_add_143427;
  reg [16:0] p2_add_143428;
  reg [16:0] p2_add_143429;
  reg [16:0] p2_add_143430;
  reg [16:0] p2_add_143431;
  reg [16:0] p2_add_143432;
  reg [16:0] p2_add_143433;
  reg [16:0] p2_add_143434;
  reg [16:0] p2_add_143435;
  reg [16:0] p2_add_143436;
  reg [16:0] p2_add_143437;
  reg [16:0] p2_add_143438;
  reg [16:0] p2_add_143439;
  reg [16:0] p2_add_143440;
  reg [16:0] p2_add_143441;
  reg [16:0] p2_add_143442;
  reg [16:0] p2_add_143443;
  reg [16:0] p2_add_143444;
  reg [16:0] p2_add_143445;
  reg [16:0] p2_add_143446;
  reg [16:0] p2_add_143447;
  reg [16:0] p2_add_143448;
  reg [16:0] p2_add_143449;
  reg [16:0] p2_add_143450;
  reg [16:0] p2_add_143451;
  reg [16:0] p2_add_143452;
  reg [16:0] p2_add_143453;
  reg [16:0] p2_add_143454;
  reg [16:0] p2_add_143455;
  reg [16:0] p2_add_143456;
  reg [16:0] p2_add_143457;
  reg [16:0] p2_add_143458;
  reg [16:0] p2_add_143467;
  reg [16:0] p2_add_143468;
  reg [16:0] p2_add_143469;
  reg [16:0] p2_add_143470;
  reg [16:0] p2_add_143471;
  reg [16:0] p2_add_143472;
  reg [16:0] p2_add_143473;
  reg [16:0] p2_add_143474;
  reg [16:0] p2_add_143499;
  reg [16:0] p2_add_143500;
  reg [16:0] p2_add_143501;
  reg [16:0] p2_add_143502;
  reg [16:0] p2_add_143503;
  reg [16:0] p2_add_143504;
  reg [16:0] p2_add_143505;
  reg [16:0] p2_add_143506;
  reg [16:0] p2_add_143515;
  reg [16:0] p2_add_143516;
  reg [16:0] p2_add_143517;
  reg [16:0] p2_add_143518;
  reg [16:0] p2_add_143519;
  reg [16:0] p2_add_143520;
  reg [16:0] p2_add_143521;
  reg [16:0] p2_add_143522;
  reg [16:0] p2_add_143523;
  reg [16:0] p2_add_143524;
  reg [16:0] p2_add_143525;
  reg [16:0] p2_add_143526;
  reg [16:0] p2_add_143527;
  reg [16:0] p2_add_143528;
  reg [16:0] p2_add_143529;
  reg [16:0] p2_add_143530;
  reg [16:0] p2_add_143531;
  reg [16:0] p2_add_143532;
  reg [16:0] p2_add_143533;
  reg [16:0] p2_add_143534;
  reg [16:0] p2_add_143535;
  reg [16:0] p2_add_143536;
  reg [16:0] p2_add_143537;
  reg [16:0] p2_add_143538;
  reg [16:0] p2_add_143539;
  reg [16:0] p2_add_143540;
  reg [16:0] p2_add_143541;
  reg [16:0] p2_add_143542;
  reg [16:0] p2_add_143543;
  reg [16:0] p2_add_143544;
  reg [16:0] p2_add_143545;
  reg [16:0] p2_add_143546;
  reg [16:0] p2_add_143547;
  reg [16:0] p2_add_143548;
  reg [16:0] p2_add_143549;
  reg [16:0] p2_add_143550;
  reg [16:0] p2_add_143551;
  reg [16:0] p2_add_143552;
  reg [16:0] p2_add_143553;
  reg [16:0] p2_add_143554;
  reg [16:0] p2_add_143563;
  reg [16:0] p2_add_143564;
  reg [16:0] p2_add_143565;
  reg [16:0] p2_add_143566;
  reg [16:0] p2_add_143567;
  reg [16:0] p2_add_143568;
  reg [16:0] p2_add_143569;
  reg [16:0] p2_add_143570;
  reg [31:0] p2_sum__995;
  reg [31:0] p2_sum__890;
  reg [31:0] p2_sum__1023;
  reg [31:0] p2_sum__1016;
  reg [31:0] p2_sum__967;
  reg [31:0] p2_sum__932;
  reg [31:0] p2_sum__841;
  reg [31:0] p2_sum__785;
  reg [24:0] p2_sum__1768;
  reg [24:0] p2_sum__1769;
  reg [24:0] p2_sum__1770;
  reg [24:0] p2_sum__1771;
  reg [24:0] p2_sum__1748;
  reg [24:0] p2_sum__1749;
  reg [24:0] p2_sum__1750;
  reg [24:0] p2_sum__1751;
  reg [24:0] p2_sum__1732;
  reg [24:0] p2_sum__1733;
  reg [24:0] p2_sum__1734;
  reg [24:0] p2_sum__1735;
  reg [24:0] p2_sum__1704;
  reg [24:0] p2_sum__1705;
  reg [24:0] p2_sum__1706;
  reg [24:0] p2_sum__1707;
  reg [24:0] p2_sum__1684;
  reg [24:0] p2_sum__1685;
  reg [24:0] p2_sum__1686;
  reg [24:0] p2_sum__1687;
  reg [24:0] p2_sum__1656;
  reg [24:0] p2_sum__1657;
  reg [24:0] p2_sum__1658;
  reg [24:0] p2_sum__1659;
  reg [24:0] p2_sum__1640;
  reg [24:0] p2_sum__1641;
  reg [24:0] p2_sum__1642;
  reg [24:0] p2_sum__1643;
  reg [24:0] p2_sum__1620;
  reg [24:0] p2_sum__1621;
  reg [24:0] p2_sum__1622;
  reg [24:0] p2_sum__1623;
  reg [24:0] p2_sum__1324;
  reg [24:0] p2_sum__1325;
  reg [24:0] p2_sum__1282;
  reg [24:0] p2_sum__1283;
  reg [24:0] p2_sum__1346;
  reg [24:0] p2_sum__1347;
  reg [24:0] p2_sum__1336;
  reg [24:0] p2_sum__1337;
  reg [24:0] p2_sum__1310;
  reg [24:0] p2_sum__1311;
  reg [24:0] p2_sum__1296;
  reg [24:0] p2_sum__1297;
  reg [24:0] p2_sum__1270;
  reg [24:0] p2_sum__1271;
  reg [24:0] p2_sum__1260;
  reg [24:0] p2_sum__1261;
  always @ (posedge clk) begin
    p2_add_143335 <= p2_add_143335_comb;
    p2_add_143336 <= p2_add_143336_comb;
    p2_add_143337 <= p2_add_143337_comb;
    p2_add_143338 <= p2_add_143338_comb;
    p2_add_143339 <= p2_add_143339_comb;
    p2_add_143340 <= p2_add_143340_comb;
    p2_add_143341 <= p2_add_143341_comb;
    p2_add_143342 <= p2_add_143342_comb;
    p2_add_143343 <= p2_add_143343_comb;
    p2_add_143344 <= p2_add_143344_comb;
    p2_add_143345 <= p2_add_143345_comb;
    p2_add_143346 <= p2_add_143346_comb;
    p2_add_143347 <= p2_add_143347_comb;
    p2_add_143348 <= p2_add_143348_comb;
    p2_add_143349 <= p2_add_143349_comb;
    p2_add_143350 <= p2_add_143350_comb;
    p2_add_143351 <= p2_add_143351_comb;
    p2_add_143352 <= p2_add_143352_comb;
    p2_add_143353 <= p2_add_143353_comb;
    p2_add_143354 <= p2_add_143354_comb;
    p2_add_143355 <= p2_add_143355_comb;
    p2_add_143356 <= p2_add_143356_comb;
    p2_add_143357 <= p2_add_143357_comb;
    p2_add_143358 <= p2_add_143358_comb;
    p2_add_143367 <= p2_add_143367_comb;
    p2_add_143368 <= p2_add_143368_comb;
    p2_add_143369 <= p2_add_143369_comb;
    p2_add_143370 <= p2_add_143370_comb;
    p2_add_143371 <= p2_add_143371_comb;
    p2_add_143372 <= p2_add_143372_comb;
    p2_add_143373 <= p2_add_143373_comb;
    p2_add_143374 <= p2_add_143374_comb;
    p2_add_143375 <= p2_add_143375_comb;
    p2_add_143376 <= p2_add_143376_comb;
    p2_add_143377 <= p2_add_143377_comb;
    p2_add_143378 <= p2_add_143378_comb;
    p2_add_143379 <= p2_add_143379_comb;
    p2_add_143380 <= p2_add_143380_comb;
    p2_add_143381 <= p2_add_143381_comb;
    p2_add_143382 <= p2_add_143382_comb;
    p2_add_143383 <= p2_add_143383_comb;
    p2_add_143384 <= p2_add_143384_comb;
    p2_add_143385 <= p2_add_143385_comb;
    p2_add_143386 <= p2_add_143386_comb;
    p2_add_143387 <= p2_add_143387_comb;
    p2_add_143388 <= p2_add_143388_comb;
    p2_add_143389 <= p2_add_143389_comb;
    p2_add_143390 <= p2_add_143390_comb;
    p2_add_143403 <= p2_add_143403_comb;
    p2_add_143404 <= p2_add_143404_comb;
    p2_add_143405 <= p2_add_143405_comb;
    p2_add_143406 <= p2_add_143406_comb;
    p2_add_143407 <= p2_add_143407_comb;
    p2_add_143408 <= p2_add_143408_comb;
    p2_add_143409 <= p2_add_143409_comb;
    p2_add_143410 <= p2_add_143410_comb;
    p2_add_143419 <= p2_add_143419_comb;
    p2_add_143420 <= p2_add_143420_comb;
    p2_add_143421 <= p2_add_143421_comb;
    p2_add_143422 <= p2_add_143422_comb;
    p2_add_143423 <= p2_add_143423_comb;
    p2_add_143424 <= p2_add_143424_comb;
    p2_add_143425 <= p2_add_143425_comb;
    p2_add_143426 <= p2_add_143426_comb;
    p2_add_143427 <= p2_add_143427_comb;
    p2_add_143428 <= p2_add_143428_comb;
    p2_add_143429 <= p2_add_143429_comb;
    p2_add_143430 <= p2_add_143430_comb;
    p2_add_143431 <= p2_add_143431_comb;
    p2_add_143432 <= p2_add_143432_comb;
    p2_add_143433 <= p2_add_143433_comb;
    p2_add_143434 <= p2_add_143434_comb;
    p2_add_143435 <= p2_add_143435_comb;
    p2_add_143436 <= p2_add_143436_comb;
    p2_add_143437 <= p2_add_143437_comb;
    p2_add_143438 <= p2_add_143438_comb;
    p2_add_143439 <= p2_add_143439_comb;
    p2_add_143440 <= p2_add_143440_comb;
    p2_add_143441 <= p2_add_143441_comb;
    p2_add_143442 <= p2_add_143442_comb;
    p2_add_143443 <= p2_add_143443_comb;
    p2_add_143444 <= p2_add_143444_comb;
    p2_add_143445 <= p2_add_143445_comb;
    p2_add_143446 <= p2_add_143446_comb;
    p2_add_143447 <= p2_add_143447_comb;
    p2_add_143448 <= p2_add_143448_comb;
    p2_add_143449 <= p2_add_143449_comb;
    p2_add_143450 <= p2_add_143450_comb;
    p2_add_143451 <= p2_add_143451_comb;
    p2_add_143452 <= p2_add_143452_comb;
    p2_add_143453 <= p2_add_143453_comb;
    p2_add_143454 <= p2_add_143454_comb;
    p2_add_143455 <= p2_add_143455_comb;
    p2_add_143456 <= p2_add_143456_comb;
    p2_add_143457 <= p2_add_143457_comb;
    p2_add_143458 <= p2_add_143458_comb;
    p2_add_143467 <= p2_add_143467_comb;
    p2_add_143468 <= p2_add_143468_comb;
    p2_add_143469 <= p2_add_143469_comb;
    p2_add_143470 <= p2_add_143470_comb;
    p2_add_143471 <= p2_add_143471_comb;
    p2_add_143472 <= p2_add_143472_comb;
    p2_add_143473 <= p2_add_143473_comb;
    p2_add_143474 <= p2_add_143474_comb;
    p2_add_143499 <= p2_add_143499_comb;
    p2_add_143500 <= p2_add_143500_comb;
    p2_add_143501 <= p2_add_143501_comb;
    p2_add_143502 <= p2_add_143502_comb;
    p2_add_143503 <= p2_add_143503_comb;
    p2_add_143504 <= p2_add_143504_comb;
    p2_add_143505 <= p2_add_143505_comb;
    p2_add_143506 <= p2_add_143506_comb;
    p2_add_143515 <= p2_add_143515_comb;
    p2_add_143516 <= p2_add_143516_comb;
    p2_add_143517 <= p2_add_143517_comb;
    p2_add_143518 <= p2_add_143518_comb;
    p2_add_143519 <= p2_add_143519_comb;
    p2_add_143520 <= p2_add_143520_comb;
    p2_add_143521 <= p2_add_143521_comb;
    p2_add_143522 <= p2_add_143522_comb;
    p2_add_143523 <= p2_add_143523_comb;
    p2_add_143524 <= p2_add_143524_comb;
    p2_add_143525 <= p2_add_143525_comb;
    p2_add_143526 <= p2_add_143526_comb;
    p2_add_143527 <= p2_add_143527_comb;
    p2_add_143528 <= p2_add_143528_comb;
    p2_add_143529 <= p2_add_143529_comb;
    p2_add_143530 <= p2_add_143530_comb;
    p2_add_143531 <= p2_add_143531_comb;
    p2_add_143532 <= p2_add_143532_comb;
    p2_add_143533 <= p2_add_143533_comb;
    p2_add_143534 <= p2_add_143534_comb;
    p2_add_143535 <= p2_add_143535_comb;
    p2_add_143536 <= p2_add_143536_comb;
    p2_add_143537 <= p2_add_143537_comb;
    p2_add_143538 <= p2_add_143538_comb;
    p2_add_143539 <= p2_add_143539_comb;
    p2_add_143540 <= p2_add_143540_comb;
    p2_add_143541 <= p2_add_143541_comb;
    p2_add_143542 <= p2_add_143542_comb;
    p2_add_143543 <= p2_add_143543_comb;
    p2_add_143544 <= p2_add_143544_comb;
    p2_add_143545 <= p2_add_143545_comb;
    p2_add_143546 <= p2_add_143546_comb;
    p2_add_143547 <= p2_add_143547_comb;
    p2_add_143548 <= p2_add_143548_comb;
    p2_add_143549 <= p2_add_143549_comb;
    p2_add_143550 <= p2_add_143550_comb;
    p2_add_143551 <= p2_add_143551_comb;
    p2_add_143552 <= p2_add_143552_comb;
    p2_add_143553 <= p2_add_143553_comb;
    p2_add_143554 <= p2_add_143554_comb;
    p2_add_143563 <= p2_add_143563_comb;
    p2_add_143564 <= p2_add_143564_comb;
    p2_add_143565 <= p2_add_143565_comb;
    p2_add_143566 <= p2_add_143566_comb;
    p2_add_143567 <= p2_add_143567_comb;
    p2_add_143568 <= p2_add_143568_comb;
    p2_add_143569 <= p2_add_143569_comb;
    p2_add_143570 <= p2_add_143570_comb;
    p2_sum__995 <= p2_sum__995_comb;
    p2_sum__890 <= p2_sum__890_comb;
    p2_sum__1023 <= p2_sum__1023_comb;
    p2_sum__1016 <= p2_sum__1016_comb;
    p2_sum__967 <= p2_sum__967_comb;
    p2_sum__932 <= p2_sum__932_comb;
    p2_sum__841 <= p2_sum__841_comb;
    p2_sum__785 <= p2_sum__785_comb;
    p2_sum__1768 <= p2_sum__1768_comb;
    p2_sum__1769 <= p2_sum__1769_comb;
    p2_sum__1770 <= p2_sum__1770_comb;
    p2_sum__1771 <= p2_sum__1771_comb;
    p2_sum__1748 <= p2_sum__1748_comb;
    p2_sum__1749 <= p2_sum__1749_comb;
    p2_sum__1750 <= p2_sum__1750_comb;
    p2_sum__1751 <= p2_sum__1751_comb;
    p2_sum__1732 <= p2_sum__1732_comb;
    p2_sum__1733 <= p2_sum__1733_comb;
    p2_sum__1734 <= p2_sum__1734_comb;
    p2_sum__1735 <= p2_sum__1735_comb;
    p2_sum__1704 <= p2_sum__1704_comb;
    p2_sum__1705 <= p2_sum__1705_comb;
    p2_sum__1706 <= p2_sum__1706_comb;
    p2_sum__1707 <= p2_sum__1707_comb;
    p2_sum__1684 <= p2_sum__1684_comb;
    p2_sum__1685 <= p2_sum__1685_comb;
    p2_sum__1686 <= p2_sum__1686_comb;
    p2_sum__1687 <= p2_sum__1687_comb;
    p2_sum__1656 <= p2_sum__1656_comb;
    p2_sum__1657 <= p2_sum__1657_comb;
    p2_sum__1658 <= p2_sum__1658_comb;
    p2_sum__1659 <= p2_sum__1659_comb;
    p2_sum__1640 <= p2_sum__1640_comb;
    p2_sum__1641 <= p2_sum__1641_comb;
    p2_sum__1642 <= p2_sum__1642_comb;
    p2_sum__1643 <= p2_sum__1643_comb;
    p2_sum__1620 <= p2_sum__1620_comb;
    p2_sum__1621 <= p2_sum__1621_comb;
    p2_sum__1622 <= p2_sum__1622_comb;
    p2_sum__1623 <= p2_sum__1623_comb;
    p2_sum__1324 <= p2_sum__1324_comb;
    p2_sum__1325 <= p2_sum__1325_comb;
    p2_sum__1282 <= p2_sum__1282_comb;
    p2_sum__1283 <= p2_sum__1283_comb;
    p2_sum__1346 <= p2_sum__1346_comb;
    p2_sum__1347 <= p2_sum__1347_comb;
    p2_sum__1336 <= p2_sum__1336_comb;
    p2_sum__1337 <= p2_sum__1337_comb;
    p2_sum__1310 <= p2_sum__1310_comb;
    p2_sum__1311 <= p2_sum__1311_comb;
    p2_sum__1296 <= p2_sum__1296_comb;
    p2_sum__1297 <= p2_sum__1297_comb;
    p2_sum__1270 <= p2_sum__1270_comb;
    p2_sum__1271 <= p2_sum__1271_comb;
    p2_sum__1260 <= p2_sum__1260_comb;
    p2_sum__1261 <= p2_sum__1261_comb;
  end

  // ===== Pipe stage 3:
  wire [24:0] p3_sum__1784_comb;
  wire [24:0] p3_sum__1785_comb;
  wire [24:0] p3_sum__1786_comb;
  wire [24:0] p3_sum__1787_comb;
  wire [24:0] p3_sum__1724_comb;
  wire [24:0] p3_sum__1725_comb;
  wire [24:0] p3_sum__1726_comb;
  wire [24:0] p3_sum__1727_comb;
  wire [24:0] p3_sum__1772_comb;
  wire [24:0] p3_sum__1773_comb;
  wire [24:0] p3_sum__1774_comb;
  wire [24:0] p3_sum__1775_comb;
  wire [24:0] p3_sum__1700_comb;
  wire [24:0] p3_sum__1701_comb;
  wire [24:0] p3_sum__1702_comb;
  wire [24:0] p3_sum__1703_comb;
  wire [24:0] p3_sum__1756_comb;
  wire [24:0] p3_sum__1757_comb;
  wire [24:0] p3_sum__1758_comb;
  wire [24:0] p3_sum__1759_comb;
  wire [24:0] p3_sum__1676_comb;
  wire [24:0] p3_sum__1677_comb;
  wire [24:0] p3_sum__1678_comb;
  wire [24:0] p3_sum__1679_comb;
  wire [24:0] p3_sum__1712_comb;
  wire [24:0] p3_sum__1713_comb;
  wire [24:0] p3_sum__1714_comb;
  wire [24:0] p3_sum__1715_comb;
  wire [24:0] p3_sum__1632_comb;
  wire [24:0] p3_sum__1633_comb;
  wire [24:0] p3_sum__1634_comb;
  wire [24:0] p3_sum__1635_comb;
  wire [24:0] p3_sum__1688_comb;
  wire [24:0] p3_sum__1689_comb;
  wire [24:0] p3_sum__1690_comb;
  wire [24:0] p3_sum__1691_comb;
  wire [24:0] p3_sum__1616_comb;
  wire [24:0] p3_sum__1617_comb;
  wire [24:0] p3_sum__1618_comb;
  wire [24:0] p3_sum__1619_comb;
  wire [24:0] p3_sum__1664_comb;
  wire [24:0] p3_sum__1665_comb;
  wire [24:0] p3_sum__1666_comb;
  wire [24:0] p3_sum__1667_comb;
  wire [24:0] p3_sum__1604_comb;
  wire [24:0] p3_sum__1605_comb;
  wire [24:0] p3_sum__1606_comb;
  wire [24:0] p3_sum__1607_comb;
  wire [24:0] p3_sum__1804_comb;
  wire [24:0] p3_sum__1805_comb;
  wire [24:0] p3_sum__1806_comb;
  wire [24:0] p3_sum__1807_comb;
  wire [24:0] p3_sum__1796_comb;
  wire [24:0] p3_sum__1797_comb;
  wire [24:0] p3_sum__1798_comb;
  wire [24:0] p3_sum__1799_comb;
  wire [24:0] p3_sum__1696_comb;
  wire [24:0] p3_sum__1697_comb;
  wire [24:0] p3_sum__1698_comb;
  wire [24:0] p3_sum__1699_comb;
  wire [24:0] p3_sum__1668_comb;
  wire [24:0] p3_sum__1669_comb;
  wire [24:0] p3_sum__1670_comb;
  wire [24:0] p3_sum__1671_comb;
  wire [24:0] p3_sum__1800_comb;
  wire [24:0] p3_sum__1801_comb;
  wire [24:0] p3_sum__1802_comb;
  wire [24:0] p3_sum__1803_comb;
  wire [24:0] p3_sum__1788_comb;
  wire [24:0] p3_sum__1789_comb;
  wire [24:0] p3_sum__1790_comb;
  wire [24:0] p3_sum__1791_comb;
  wire [24:0] p3_sum__1752_comb;
  wire [24:0] p3_sum__1753_comb;
  wire [24:0] p3_sum__1754_comb;
  wire [24:0] p3_sum__1755_comb;
  wire [24:0] p3_sum__1728_comb;
  wire [24:0] p3_sum__1729_comb;
  wire [24:0] p3_sum__1730_comb;
  wire [24:0] p3_sum__1731_comb;
  wire [24:0] p3_sum__1672_comb;
  wire [24:0] p3_sum__1673_comb;
  wire [24:0] p3_sum__1674_comb;
  wire [24:0] p3_sum__1675_comb;
  wire [24:0] p3_sum__1644_comb;
  wire [24:0] p3_sum__1645_comb;
  wire [24:0] p3_sum__1646_comb;
  wire [24:0] p3_sum__1647_comb;
  wire [24:0] p3_sum__1792_comb;
  wire [24:0] p3_sum__1793_comb;
  wire [24:0] p3_sum__1794_comb;
  wire [24:0] p3_sum__1795_comb;
  wire [24:0] p3_sum__1776_comb;
  wire [24:0] p3_sum__1777_comb;
  wire [24:0] p3_sum__1778_comb;
  wire [24:0] p3_sum__1779_comb;
  wire [24:0] p3_sum__1648_comb;
  wire [24:0] p3_sum__1649_comb;
  wire [24:0] p3_sum__1650_comb;
  wire [24:0] p3_sum__1651_comb;
  wire [24:0] p3_sum__1624_comb;
  wire [24:0] p3_sum__1625_comb;
  wire [24:0] p3_sum__1626_comb;
  wire [24:0] p3_sum__1627_comb;
  wire [24:0] p3_sum__1764_comb;
  wire [24:0] p3_sum__1765_comb;
  wire [24:0] p3_sum__1766_comb;
  wire [24:0] p3_sum__1767_comb;
  wire [24:0] p3_sum__1740_comb;
  wire [24:0] p3_sum__1741_comb;
  wire [24:0] p3_sum__1742_comb;
  wire [24:0] p3_sum__1743_comb;
  wire [24:0] p3_sum__1612_comb;
  wire [24:0] p3_sum__1613_comb;
  wire [24:0] p3_sum__1614_comb;
  wire [24:0] p3_sum__1615_comb;
  wire [24:0] p3_sum__1596_comb;
  wire [24:0] p3_sum__1597_comb;
  wire [24:0] p3_sum__1598_comb;
  wire [24:0] p3_sum__1599_comb;
  wire [24:0] p3_sum__1744_comb;
  wire [24:0] p3_sum__1745_comb;
  wire [24:0] p3_sum__1746_comb;
  wire [24:0] p3_sum__1747_comb;
  wire [24:0] p3_sum__1716_comb;
  wire [24:0] p3_sum__1717_comb;
  wire [24:0] p3_sum__1718_comb;
  wire [24:0] p3_sum__1719_comb;
  wire [24:0] p3_sum__1660_comb;
  wire [24:0] p3_sum__1661_comb;
  wire [24:0] p3_sum__1662_comb;
  wire [24:0] p3_sum__1663_comb;
  wire [24:0] p3_sum__1636_comb;
  wire [24:0] p3_sum__1637_comb;
  wire [24:0] p3_sum__1638_comb;
  wire [24:0] p3_sum__1639_comb;
  wire [24:0] p3_sum__1600_comb;
  wire [24:0] p3_sum__1601_comb;
  wire [24:0] p3_sum__1602_comb;
  wire [24:0] p3_sum__1603_comb;
  wire [24:0] p3_sum__1588_comb;
  wire [24:0] p3_sum__1589_comb;
  wire [24:0] p3_sum__1590_comb;
  wire [24:0] p3_sum__1591_comb;
  wire [24:0] p3_sum__1720_comb;
  wire [24:0] p3_sum__1721_comb;
  wire [24:0] p3_sum__1722_comb;
  wire [24:0] p3_sum__1723_comb;
  wire [24:0] p3_sum__1692_comb;
  wire [24:0] p3_sum__1693_comb;
  wire [24:0] p3_sum__1694_comb;
  wire [24:0] p3_sum__1695_comb;
  wire [24:0] p3_sum__1592_comb;
  wire [24:0] p3_sum__1593_comb;
  wire [24:0] p3_sum__1594_comb;
  wire [24:0] p3_sum__1595_comb;
  wire [24:0] p3_sum__1584_comb;
  wire [24:0] p3_sum__1585_comb;
  wire [24:0] p3_sum__1586_comb;
  wire [24:0] p3_sum__1587_comb;
  wire [31:0] p3_umul_144259_comb;
  wire [31:0] p3_umul_144260_comb;
  wire [31:0] p3_umul_144285_comb;
  wire [31:0] p3_umul_144286_comb;
  wire [31:0] p3_umul_144287_comb;
  wire [31:0] p3_umul_144288_comb;
  wire [31:0] p3_umul_144289_comb;
  wire [31:0] p3_umul_144290_comb;
  wire [24:0] p3_sum__1340_comb;
  wire [24:0] p3_sum__1341_comb;
  wire [24:0] p3_sum__1330_comb;
  wire [24:0] p3_sum__1331_comb;
  wire [24:0] p3_sum__1322_comb;
  wire [24:0] p3_sum__1323_comb;
  wire [24:0] p3_sum__1308_comb;
  wire [24:0] p3_sum__1309_comb;
  wire [24:0] p3_sum__1298_comb;
  wire [24:0] p3_sum__1299_comb;
  wire [24:0] p3_sum__1284_comb;
  wire [24:0] p3_sum__1285_comb;
  wire [24:0] p3_sum__1276_comb;
  wire [24:0] p3_sum__1277_comb;
  wire [24:0] p3_sum__1266_comb;
  wire [24:0] p3_sum__1267_comb;
  wire [24:0] p3_sum__1118_comb;
  wire [24:0] p3_sum__1097_comb;
  wire [24:0] p3_sum__1129_comb;
  wire [24:0] p3_sum__1124_comb;
  wire [24:0] p3_sum__1111_comb;
  wire [24:0] p3_sum__1104_comb;
  wire [24:0] p3_sum__1091_comb;
  wire [24:0] p3_sum__1086_comb;
  wire [24:0] p3_sum__1348_comb;
  wire [24:0] p3_sum__1349_comb;
  wire [24:0] p3_sum__1318_comb;
  wire [24:0] p3_sum__1319_comb;
  wire [24:0] p3_sum__1342_comb;
  wire [24:0] p3_sum__1343_comb;
  wire [24:0] p3_sum__1306_comb;
  wire [24:0] p3_sum__1307_comb;
  wire [24:0] p3_sum__1334_comb;
  wire [24:0] p3_sum__1335_comb;
  wire [24:0] p3_sum__1294_comb;
  wire [24:0] p3_sum__1295_comb;
  wire [24:0] p3_sum__1312_comb;
  wire [24:0] p3_sum__1313_comb;
  wire [24:0] p3_sum__1272_comb;
  wire [24:0] p3_sum__1273_comb;
  wire [24:0] p3_sum__1300_comb;
  wire [24:0] p3_sum__1301_comb;
  wire [24:0] p3_sum__1264_comb;
  wire [24:0] p3_sum__1265_comb;
  wire [24:0] p3_sum__1288_comb;
  wire [24:0] p3_sum__1289_comb;
  wire [24:0] p3_sum__1258_comb;
  wire [24:0] p3_sum__1259_comb;
  wire [24:0] p3_sum__1358_comb;
  wire [24:0] p3_sum__1359_comb;
  wire [24:0] p3_sum__1354_comb;
  wire [24:0] p3_sum__1355_comb;
  wire [24:0] p3_sum__1304_comb;
  wire [24:0] p3_sum__1305_comb;
  wire [24:0] p3_sum__1290_comb;
  wire [24:0] p3_sum__1291_comb;
  wire [24:0] p3_sum__1356_comb;
  wire [24:0] p3_sum__1357_comb;
  wire [24:0] p3_sum__1350_comb;
  wire [24:0] p3_sum__1351_comb;
  wire [24:0] p3_sum__1332_comb;
  wire [24:0] p3_sum__1333_comb;
  wire [24:0] p3_sum__1320_comb;
  wire [24:0] p3_sum__1321_comb;
  wire [24:0] p3_sum__1292_comb;
  wire [24:0] p3_sum__1293_comb;
  wire [24:0] p3_sum__1278_comb;
  wire [24:0] p3_sum__1279_comb;
  wire [24:0] p3_sum__1352_comb;
  wire [24:0] p3_sum__1353_comb;
  wire [24:0] p3_sum__1344_comb;
  wire [24:0] p3_sum__1345_comb;
  wire [24:0] p3_sum__1280_comb;
  wire [24:0] p3_sum__1281_comb;
  wire [24:0] p3_sum__1268_comb;
  wire [24:0] p3_sum__1269_comb;
  wire [24:0] p3_sum__1338_comb;
  wire [24:0] p3_sum__1339_comb;
  wire [24:0] p3_sum__1326_comb;
  wire [24:0] p3_sum__1327_comb;
  wire [24:0] p3_sum__1262_comb;
  wire [24:0] p3_sum__1263_comb;
  wire [24:0] p3_sum__1254_comb;
  wire [24:0] p3_sum__1255_comb;
  wire [24:0] p3_sum__1328_comb;
  wire [24:0] p3_sum__1329_comb;
  wire [24:0] p3_sum__1314_comb;
  wire [24:0] p3_sum__1315_comb;
  wire [24:0] p3_sum__1286_comb;
  wire [24:0] p3_sum__1287_comb;
  wire [24:0] p3_sum__1274_comb;
  wire [24:0] p3_sum__1275_comb;
  wire [24:0] p3_sum__1256_comb;
  wire [24:0] p3_sum__1257_comb;
  wire [24:0] p3_sum__1250_comb;
  wire [24:0] p3_sum__1251_comb;
  wire [24:0] p3_sum__1316_comb;
  wire [24:0] p3_sum__1317_comb;
  wire [24:0] p3_sum__1302_comb;
  wire [24:0] p3_sum__1303_comb;
  wire [24:0] p3_sum__1252_comb;
  wire [24:0] p3_sum__1253_comb;
  wire [24:0] p3_sum__1248_comb;
  wire [24:0] p3_sum__1249_comb;
  wire [24:0] p3_sum__1126_comb;
  wire [24:0] p3_sum__1121_comb;
  wire [24:0] p3_sum__1117_comb;
  wire [24:0] p3_sum__1110_comb;
  wire [24:0] p3_sum__1105_comb;
  wire [24:0] p3_sum__1098_comb;
  wire [24:0] p3_sum__1094_comb;
  wire [24:0] p3_sum__1089_comb;
  wire [24:0] p3_add_144499_comb;
  wire [24:0] p3_add_144500_comb;
  wire [24:0] p3_add_144531_comb;
  wire [24:0] p3_add_144532_comb;
  wire [24:0] p3_add_144533_comb;
  wire [24:0] p3_add_144534_comb;
  wire [24:0] p3_add_144535_comb;
  wire [24:0] p3_add_144536_comb;
  wire [24:0] p3_sum__1130_comb;
  wire [24:0] p3_sum__1115_comb;
  wire [24:0] p3_sum__1127_comb;
  wire [24:0] p3_sum__1109_comb;
  wire [24:0] p3_sum__1123_comb;
  wire [24:0] p3_sum__1103_comb;
  wire [24:0] p3_sum__1112_comb;
  wire [24:0] p3_sum__1092_comb;
  wire [24:0] p3_sum__1106_comb;
  wire [24:0] p3_sum__1088_comb;
  wire [24:0] p3_sum__1100_comb;
  wire [24:0] p3_sum__1085_comb;
  wire [24:0] p3_sum__1135_comb;
  wire [24:0] p3_sum__1133_comb;
  wire [24:0] p3_sum__1108_comb;
  wire [24:0] p3_sum__1101_comb;
  wire [24:0] p3_sum__1134_comb;
  wire [24:0] p3_sum__1131_comb;
  wire [24:0] p3_sum__1122_comb;
  wire [24:0] p3_sum__1116_comb;
  wire [24:0] p3_sum__1102_comb;
  wire [24:0] p3_sum__1095_comb;
  wire [24:0] p3_sum__1132_comb;
  wire [24:0] p3_sum__1128_comb;
  wire [24:0] p3_sum__1096_comb;
  wire [24:0] p3_sum__1090_comb;
  wire [24:0] p3_sum__1125_comb;
  wire [24:0] p3_sum__1119_comb;
  wire [24:0] p3_sum__1087_comb;
  wire [24:0] p3_sum__1083_comb;
  wire [24:0] p3_sum__1120_comb;
  wire [24:0] p3_sum__1113_comb;
  wire [24:0] p3_sum__1099_comb;
  wire [24:0] p3_sum__1093_comb;
  wire [24:0] p3_sum__1084_comb;
  wire [24:0] p3_sum__1081_comb;
  wire [24:0] p3_sum__1114_comb;
  wire [24:0] p3_sum__1107_comb;
  wire [24:0] p3_sum__1082_comb;
  wire [24:0] p3_sum__1080_comb;
  wire [24:0] p3_add_144491_comb;
  wire [24:0] p3_add_144492_comb;
  wire [24:0] p3_add_144507_comb;
  wire [24:0] p3_add_144508_comb;
  wire [24:0] p3_add_144509_comb;
  wire [24:0] p3_add_144510_comb;
  wire [24:0] p3_add_144511_comb;
  wire [24:0] p3_add_144512_comb;
  wire [24:0] p3_add_144515_comb;
  wire [24:0] p3_add_144516_comb;
  wire [24:0] p3_add_144527_comb;
  wire [24:0] p3_add_144528_comb;
  wire [24:0] p3_add_144539_comb;
  wire [24:0] p3_add_144540_comb;
  wire [24:0] p3_add_144551_comb;
  wire [24:0] p3_add_144552_comb;
  wire [24:0] p3_add_144493_comb;
  wire [24:0] p3_add_144494_comb;
  wire [24:0] p3_add_144495_comb;
  wire [24:0] p3_add_144496_comb;
  wire [24:0] p3_add_144497_comb;
  wire [24:0] p3_add_144498_comb;
  wire [24:0] p3_add_144501_comb;
  wire [24:0] p3_add_144502_comb;
  wire [24:0] p3_add_144503_comb;
  wire [24:0] p3_add_144504_comb;
  wire [24:0] p3_add_144505_comb;
  wire [24:0] p3_add_144506_comb;
  wire [24:0] p3_add_144513_comb;
  wire [24:0] p3_add_144514_comb;
  wire [24:0] p3_add_144517_comb;
  wire [24:0] p3_add_144518_comb;
  wire [24:0] p3_add_144519_comb;
  wire [24:0] p3_add_144520_comb;
  wire [24:0] p3_add_144521_comb;
  wire [24:0] p3_add_144522_comb;
  wire [24:0] p3_add_144523_comb;
  wire [24:0] p3_add_144524_comb;
  wire [24:0] p3_add_144525_comb;
  wire [24:0] p3_add_144526_comb;
  wire [24:0] p3_add_144529_comb;
  wire [24:0] p3_add_144530_comb;
  wire [24:0] p3_add_144537_comb;
  wire [24:0] p3_add_144538_comb;
  wire [24:0] p3_add_144541_comb;
  wire [24:0] p3_add_144542_comb;
  wire [24:0] p3_add_144543_comb;
  wire [24:0] p3_add_144544_comb;
  wire [24:0] p3_add_144545_comb;
  wire [24:0] p3_add_144546_comb;
  wire [24:0] p3_add_144547_comb;
  wire [24:0] p3_add_144548_comb;
  wire [24:0] p3_add_144549_comb;
  wire [24:0] p3_add_144550_comb;
  wire [24:0] p3_add_144553_comb;
  wire [24:0] p3_add_144554_comb;
  wire [8:0] p3_clipped__272_comb;
  wire [8:0] p3_clipped__275_comb;
  wire [8:0] p3_clipped__304_comb;
  wire [8:0] p3_clipped__305_comb;
  wire [8:0] p3_clipped__273_comb;
  wire [8:0] p3_clipped__274_comb;
  wire [8:0] p3_clipped__306_comb;
  wire [8:0] p3_clipped__307_comb;
  wire [8:0] p3_clipped__256_comb;
  wire [8:0] p3_clipped__259_comb;
  wire [8:0] p3_clipped__288_comb;
  wire [8:0] p3_clipped__289_comb;
  wire [8:0] p3_clipped__257_comb;
  wire [8:0] p3_clipped__258_comb;
  wire [8:0] p3_clipped__290_comb;
  wire [8:0] p3_clipped__291_comb;
  wire [8:0] p3_clipped__261_comb;
  wire [8:0] p3_clipped__262_comb;
  wire [8:0] p3_clipped__269_comb;
  wire [8:0] p3_clipped__270_comb;
  wire [8:0] p3_clipped__277_comb;
  wire [8:0] p3_clipped__278_comb;
  wire [8:0] p3_clipped__285_comb;
  wire [8:0] p3_clipped__286_comb;
  wire [8:0] p3_clipped__260_comb;
  wire [8:0] p3_clipped__263_comb;
  wire [8:0] p3_clipped__264_comb;
  wire [8:0] p3_clipped__267_comb;
  wire [8:0] p3_clipped__268_comb;
  wire [8:0] p3_clipped__271_comb;
  wire [8:0] p3_clipped__276_comb;
  wire [8:0] p3_clipped__279_comb;
  wire [8:0] p3_clipped__280_comb;
  wire [8:0] p3_clipped__283_comb;
  wire [8:0] p3_clipped__284_comb;
  wire [8:0] p3_clipped__287_comb;
  wire [8:0] p3_clipped__292_comb;
  wire [8:0] p3_clipped__293_comb;
  wire [8:0] p3_clipped__294_comb;
  wire [8:0] p3_clipped__295_comb;
  wire [8:0] p3_clipped__296_comb;
  wire [8:0] p3_clipped__297_comb;
  wire [8:0] p3_clipped__265_comb;
  wire [8:0] p3_clipped__266_comb;
  wire [8:0] p3_clipped__298_comb;
  wire [8:0] p3_clipped__299_comb;
  wire [8:0] p3_clipped__300_comb;
  wire [8:0] p3_clipped__301_comb;
  wire [8:0] p3_clipped__302_comb;
  wire [8:0] p3_clipped__303_comb;
  wire [8:0] p3_clipped__308_comb;
  wire [8:0] p3_clipped__309_comb;
  wire [8:0] p3_clipped__310_comb;
  wire [8:0] p3_clipped__311_comb;
  wire [8:0] p3_clipped__312_comb;
  wire [8:0] p3_clipped__313_comb;
  wire [8:0] p3_clipped__281_comb;
  wire [8:0] p3_clipped__282_comb;
  wire [8:0] p3_clipped__314_comb;
  wire [8:0] p3_clipped__315_comb;
  wire [8:0] p3_clipped__316_comb;
  wire [8:0] p3_clipped__317_comb;
  wire [8:0] p3_clipped__318_comb;
  wire [8:0] p3_clipped__319_comb;
  wire [9:0] p3_sign_ext_145195_comb;
  wire [9:0] p3_sign_ext_145196_comb;
  wire [9:0] p3_sign_ext_145201_comb;
  wire [9:0] p3_sign_ext_145202_comb;
  wire [9:0] p3_sign_ext_145203_comb;
  wire [9:0] p3_sign_ext_145204_comb;
  wire [9:0] p3_sign_ext_145205_comb;
  wire [9:0] p3_sign_ext_145206_comb;
  wire [9:0] p3_sign_ext_145207_comb;
  wire [9:0] p3_sign_ext_145208_comb;
  wire [9:0] p3_sign_ext_145209_comb;
  wire [9:0] p3_sign_ext_145210_comb;
  wire [9:0] p3_sign_ext_145223_comb;
  wire [9:0] p3_sign_ext_145224_comb;
  wire [9:0] p3_sign_ext_145225_comb;
  wire [9:0] p3_sign_ext_145226_comb;
  wire [9:0] p3_add_145227_comb;
  wire [9:0] p3_add_145228_comb;
  wire [9:0] p3_add_145229_comb;
  wire [9:0] p3_add_145230_comb;
  wire [9:0] p3_add_145231_comb;
  wire [9:0] p3_add_145232_comb;
  wire [9:0] p3_add_145233_comb;
  wire [9:0] p3_add_145234_comb;
  assign p3_sum__1784_comb = {{8{p2_add_143335[16]}}, p2_add_143335};
  assign p3_sum__1785_comb = {{8{p2_add_143336[16]}}, p2_add_143336};
  assign p3_sum__1786_comb = {{8{p2_add_143337[16]}}, p2_add_143337};
  assign p3_sum__1787_comb = {{8{p2_add_143338[16]}}, p2_add_143338};
  assign p3_sum__1724_comb = {{8{p2_add_143339[16]}}, p2_add_143339};
  assign p3_sum__1725_comb = {{8{p2_add_143340[16]}}, p2_add_143340};
  assign p3_sum__1726_comb = {{8{p2_add_143341[16]}}, p2_add_143341};
  assign p3_sum__1727_comb = {{8{p2_add_143342[16]}}, p2_add_143342};
  assign p3_sum__1772_comb = {{8{p2_add_143343[16]}}, p2_add_143343};
  assign p3_sum__1773_comb = {{8{p2_add_143344[16]}}, p2_add_143344};
  assign p3_sum__1774_comb = {{8{p2_add_143345[16]}}, p2_add_143345};
  assign p3_sum__1775_comb = {{8{p2_add_143346[16]}}, p2_add_143346};
  assign p3_sum__1700_comb = {{8{p2_add_143347[16]}}, p2_add_143347};
  assign p3_sum__1701_comb = {{8{p2_add_143348[16]}}, p2_add_143348};
  assign p3_sum__1702_comb = {{8{p2_add_143349[16]}}, p2_add_143349};
  assign p3_sum__1703_comb = {{8{p2_add_143350[16]}}, p2_add_143350};
  assign p3_sum__1756_comb = {{8{p2_add_143351[16]}}, p2_add_143351};
  assign p3_sum__1757_comb = {{8{p2_add_143352[16]}}, p2_add_143352};
  assign p3_sum__1758_comb = {{8{p2_add_143353[16]}}, p2_add_143353};
  assign p3_sum__1759_comb = {{8{p2_add_143354[16]}}, p2_add_143354};
  assign p3_sum__1676_comb = {{8{p2_add_143355[16]}}, p2_add_143355};
  assign p3_sum__1677_comb = {{8{p2_add_143356[16]}}, p2_add_143356};
  assign p3_sum__1678_comb = {{8{p2_add_143357[16]}}, p2_add_143357};
  assign p3_sum__1679_comb = {{8{p2_add_143358[16]}}, p2_add_143358};
  assign p3_sum__1712_comb = {{8{p2_add_143367[16]}}, p2_add_143367};
  assign p3_sum__1713_comb = {{8{p2_add_143368[16]}}, p2_add_143368};
  assign p3_sum__1714_comb = {{8{p2_add_143369[16]}}, p2_add_143369};
  assign p3_sum__1715_comb = {{8{p2_add_143370[16]}}, p2_add_143370};
  assign p3_sum__1632_comb = {{8{p2_add_143371[16]}}, p2_add_143371};
  assign p3_sum__1633_comb = {{8{p2_add_143372[16]}}, p2_add_143372};
  assign p3_sum__1634_comb = {{8{p2_add_143373[16]}}, p2_add_143373};
  assign p3_sum__1635_comb = {{8{p2_add_143374[16]}}, p2_add_143374};
  assign p3_sum__1688_comb = {{8{p2_add_143375[16]}}, p2_add_143375};
  assign p3_sum__1689_comb = {{8{p2_add_143376[16]}}, p2_add_143376};
  assign p3_sum__1690_comb = {{8{p2_add_143377[16]}}, p2_add_143377};
  assign p3_sum__1691_comb = {{8{p2_add_143378[16]}}, p2_add_143378};
  assign p3_sum__1616_comb = {{8{p2_add_143379[16]}}, p2_add_143379};
  assign p3_sum__1617_comb = {{8{p2_add_143380[16]}}, p2_add_143380};
  assign p3_sum__1618_comb = {{8{p2_add_143381[16]}}, p2_add_143381};
  assign p3_sum__1619_comb = {{8{p2_add_143382[16]}}, p2_add_143382};
  assign p3_sum__1664_comb = {{8{p2_add_143383[16]}}, p2_add_143383};
  assign p3_sum__1665_comb = {{8{p2_add_143384[16]}}, p2_add_143384};
  assign p3_sum__1666_comb = {{8{p2_add_143385[16]}}, p2_add_143385};
  assign p3_sum__1667_comb = {{8{p2_add_143386[16]}}, p2_add_143386};
  assign p3_sum__1604_comb = {{8{p2_add_143387[16]}}, p2_add_143387};
  assign p3_sum__1605_comb = {{8{p2_add_143388[16]}}, p2_add_143388};
  assign p3_sum__1606_comb = {{8{p2_add_143389[16]}}, p2_add_143389};
  assign p3_sum__1607_comb = {{8{p2_add_143390[16]}}, p2_add_143390};
  assign p3_sum__1804_comb = {{8{p2_add_143403[16]}}, p2_add_143403};
  assign p3_sum__1805_comb = {{8{p2_add_143404[16]}}, p2_add_143404};
  assign p3_sum__1806_comb = {{8{p2_add_143405[16]}}, p2_add_143405};
  assign p3_sum__1807_comb = {{8{p2_add_143406[16]}}, p2_add_143406};
  assign p3_sum__1796_comb = {{8{p2_add_143407[16]}}, p2_add_143407};
  assign p3_sum__1797_comb = {{8{p2_add_143408[16]}}, p2_add_143408};
  assign p3_sum__1798_comb = {{8{p2_add_143409[16]}}, p2_add_143409};
  assign p3_sum__1799_comb = {{8{p2_add_143410[16]}}, p2_add_143410};
  assign p3_sum__1696_comb = {{8{p2_add_143419[16]}}, p2_add_143419};
  assign p3_sum__1697_comb = {{8{p2_add_143420[16]}}, p2_add_143420};
  assign p3_sum__1698_comb = {{8{p2_add_143421[16]}}, p2_add_143421};
  assign p3_sum__1699_comb = {{8{p2_add_143422[16]}}, p2_add_143422};
  assign p3_sum__1668_comb = {{8{p2_add_143423[16]}}, p2_add_143423};
  assign p3_sum__1669_comb = {{8{p2_add_143424[16]}}, p2_add_143424};
  assign p3_sum__1670_comb = {{8{p2_add_143425[16]}}, p2_add_143425};
  assign p3_sum__1671_comb = {{8{p2_add_143426[16]}}, p2_add_143426};
  assign p3_sum__1800_comb = {{8{p2_add_143427[16]}}, p2_add_143427};
  assign p3_sum__1801_comb = {{8{p2_add_143428[16]}}, p2_add_143428};
  assign p3_sum__1802_comb = {{8{p2_add_143429[16]}}, p2_add_143429};
  assign p3_sum__1803_comb = {{8{p2_add_143430[16]}}, p2_add_143430};
  assign p3_sum__1788_comb = {{8{p2_add_143431[16]}}, p2_add_143431};
  assign p3_sum__1789_comb = {{8{p2_add_143432[16]}}, p2_add_143432};
  assign p3_sum__1790_comb = {{8{p2_add_143433[16]}}, p2_add_143433};
  assign p3_sum__1791_comb = {{8{p2_add_143434[16]}}, p2_add_143434};
  assign p3_sum__1752_comb = {{8{p2_add_143435[16]}}, p2_add_143435};
  assign p3_sum__1753_comb = {{8{p2_add_143436[16]}}, p2_add_143436};
  assign p3_sum__1754_comb = {{8{p2_add_143437[16]}}, p2_add_143437};
  assign p3_sum__1755_comb = {{8{p2_add_143438[16]}}, p2_add_143438};
  assign p3_sum__1728_comb = {{8{p2_add_143439[16]}}, p2_add_143439};
  assign p3_sum__1729_comb = {{8{p2_add_143440[16]}}, p2_add_143440};
  assign p3_sum__1730_comb = {{8{p2_add_143441[16]}}, p2_add_143441};
  assign p3_sum__1731_comb = {{8{p2_add_143442[16]}}, p2_add_143442};
  assign p3_sum__1672_comb = {{8{p2_add_143443[16]}}, p2_add_143443};
  assign p3_sum__1673_comb = {{8{p2_add_143444[16]}}, p2_add_143444};
  assign p3_sum__1674_comb = {{8{p2_add_143445[16]}}, p2_add_143445};
  assign p3_sum__1675_comb = {{8{p2_add_143446[16]}}, p2_add_143446};
  assign p3_sum__1644_comb = {{8{p2_add_143447[16]}}, p2_add_143447};
  assign p3_sum__1645_comb = {{8{p2_add_143448[16]}}, p2_add_143448};
  assign p3_sum__1646_comb = {{8{p2_add_143449[16]}}, p2_add_143449};
  assign p3_sum__1647_comb = {{8{p2_add_143450[16]}}, p2_add_143450};
  assign p3_sum__1792_comb = {{8{p2_add_143451[16]}}, p2_add_143451};
  assign p3_sum__1793_comb = {{8{p2_add_143452[16]}}, p2_add_143452};
  assign p3_sum__1794_comb = {{8{p2_add_143453[16]}}, p2_add_143453};
  assign p3_sum__1795_comb = {{8{p2_add_143454[16]}}, p2_add_143454};
  assign p3_sum__1776_comb = {{8{p2_add_143455[16]}}, p2_add_143455};
  assign p3_sum__1777_comb = {{8{p2_add_143456[16]}}, p2_add_143456};
  assign p3_sum__1778_comb = {{8{p2_add_143457[16]}}, p2_add_143457};
  assign p3_sum__1779_comb = {{8{p2_add_143458[16]}}, p2_add_143458};
  assign p3_sum__1648_comb = {{8{p2_add_143467[16]}}, p2_add_143467};
  assign p3_sum__1649_comb = {{8{p2_add_143468[16]}}, p2_add_143468};
  assign p3_sum__1650_comb = {{8{p2_add_143469[16]}}, p2_add_143469};
  assign p3_sum__1651_comb = {{8{p2_add_143470[16]}}, p2_add_143470};
  assign p3_sum__1624_comb = {{8{p2_add_143471[16]}}, p2_add_143471};
  assign p3_sum__1625_comb = {{8{p2_add_143472[16]}}, p2_add_143472};
  assign p3_sum__1626_comb = {{8{p2_add_143473[16]}}, p2_add_143473};
  assign p3_sum__1627_comb = {{8{p2_add_143474[16]}}, p2_add_143474};
  assign p3_sum__1764_comb = {{8{p2_add_143499[16]}}, p2_add_143499};
  assign p3_sum__1765_comb = {{8{p2_add_143500[16]}}, p2_add_143500};
  assign p3_sum__1766_comb = {{8{p2_add_143501[16]}}, p2_add_143501};
  assign p3_sum__1767_comb = {{8{p2_add_143502[16]}}, p2_add_143502};
  assign p3_sum__1740_comb = {{8{p2_add_143503[16]}}, p2_add_143503};
  assign p3_sum__1741_comb = {{8{p2_add_143504[16]}}, p2_add_143504};
  assign p3_sum__1742_comb = {{8{p2_add_143505[16]}}, p2_add_143505};
  assign p3_sum__1743_comb = {{8{p2_add_143506[16]}}, p2_add_143506};
  assign p3_sum__1612_comb = {{8{p2_add_143515[16]}}, p2_add_143515};
  assign p3_sum__1613_comb = {{8{p2_add_143516[16]}}, p2_add_143516};
  assign p3_sum__1614_comb = {{8{p2_add_143517[16]}}, p2_add_143517};
  assign p3_sum__1615_comb = {{8{p2_add_143518[16]}}, p2_add_143518};
  assign p3_sum__1596_comb = {{8{p2_add_143519[16]}}, p2_add_143519};
  assign p3_sum__1597_comb = {{8{p2_add_143520[16]}}, p2_add_143520};
  assign p3_sum__1598_comb = {{8{p2_add_143521[16]}}, p2_add_143521};
  assign p3_sum__1599_comb = {{8{p2_add_143522[16]}}, p2_add_143522};
  assign p3_sum__1744_comb = {{8{p2_add_143523[16]}}, p2_add_143523};
  assign p3_sum__1745_comb = {{8{p2_add_143524[16]}}, p2_add_143524};
  assign p3_sum__1746_comb = {{8{p2_add_143525[16]}}, p2_add_143525};
  assign p3_sum__1747_comb = {{8{p2_add_143526[16]}}, p2_add_143526};
  assign p3_sum__1716_comb = {{8{p2_add_143527[16]}}, p2_add_143527};
  assign p3_sum__1717_comb = {{8{p2_add_143528[16]}}, p2_add_143528};
  assign p3_sum__1718_comb = {{8{p2_add_143529[16]}}, p2_add_143529};
  assign p3_sum__1719_comb = {{8{p2_add_143530[16]}}, p2_add_143530};
  assign p3_sum__1660_comb = {{8{p2_add_143531[16]}}, p2_add_143531};
  assign p3_sum__1661_comb = {{8{p2_add_143532[16]}}, p2_add_143532};
  assign p3_sum__1662_comb = {{8{p2_add_143533[16]}}, p2_add_143533};
  assign p3_sum__1663_comb = {{8{p2_add_143534[16]}}, p2_add_143534};
  assign p3_sum__1636_comb = {{8{p2_add_143535[16]}}, p2_add_143535};
  assign p3_sum__1637_comb = {{8{p2_add_143536[16]}}, p2_add_143536};
  assign p3_sum__1638_comb = {{8{p2_add_143537[16]}}, p2_add_143537};
  assign p3_sum__1639_comb = {{8{p2_add_143538[16]}}, p2_add_143538};
  assign p3_sum__1600_comb = {{8{p2_add_143539[16]}}, p2_add_143539};
  assign p3_sum__1601_comb = {{8{p2_add_143540[16]}}, p2_add_143540};
  assign p3_sum__1602_comb = {{8{p2_add_143541[16]}}, p2_add_143541};
  assign p3_sum__1603_comb = {{8{p2_add_143542[16]}}, p2_add_143542};
  assign p3_sum__1588_comb = {{8{p2_add_143543[16]}}, p2_add_143543};
  assign p3_sum__1589_comb = {{8{p2_add_143544[16]}}, p2_add_143544};
  assign p3_sum__1590_comb = {{8{p2_add_143545[16]}}, p2_add_143545};
  assign p3_sum__1591_comb = {{8{p2_add_143546[16]}}, p2_add_143546};
  assign p3_sum__1720_comb = {{8{p2_add_143547[16]}}, p2_add_143547};
  assign p3_sum__1721_comb = {{8{p2_add_143548[16]}}, p2_add_143548};
  assign p3_sum__1722_comb = {{8{p2_add_143549[16]}}, p2_add_143549};
  assign p3_sum__1723_comb = {{8{p2_add_143550[16]}}, p2_add_143550};
  assign p3_sum__1692_comb = {{8{p2_add_143551[16]}}, p2_add_143551};
  assign p3_sum__1693_comb = {{8{p2_add_143552[16]}}, p2_add_143552};
  assign p3_sum__1694_comb = {{8{p2_add_143553[16]}}, p2_add_143553};
  assign p3_sum__1695_comb = {{8{p2_add_143554[16]}}, p2_add_143554};
  assign p3_sum__1592_comb = {{8{p2_add_143563[16]}}, p2_add_143563};
  assign p3_sum__1593_comb = {{8{p2_add_143564[16]}}, p2_add_143564};
  assign p3_sum__1594_comb = {{8{p2_add_143565[16]}}, p2_add_143565};
  assign p3_sum__1595_comb = {{8{p2_add_143566[16]}}, p2_add_143566};
  assign p3_sum__1584_comb = {{8{p2_add_143567[16]}}, p2_add_143567};
  assign p3_sum__1585_comb = {{8{p2_add_143568[16]}}, p2_add_143568};
  assign p3_sum__1586_comb = {{8{p2_add_143569[16]}}, p2_add_143569};
  assign p3_sum__1587_comb = {{8{p2_add_143570[16]}}, p2_add_143570};
  assign p3_umul_144259_comb = umul32b_32b_x_7b(p2_sum__995, 7'h5b);
  assign p3_umul_144260_comb = umul32b_32b_x_7b(p2_sum__890, 7'h5b);
  assign p3_umul_144285_comb = umul32b_32b_x_7b(p2_sum__1023, 7'h5b);
  assign p3_umul_144286_comb = umul32b_32b_x_7b(p2_sum__1016, 7'h5b);
  assign p3_umul_144287_comb = umul32b_32b_x_7b(p2_sum__967, 7'h5b);
  assign p3_umul_144288_comb = umul32b_32b_x_7b(p2_sum__932, 7'h5b);
  assign p3_umul_144289_comb = umul32b_32b_x_7b(p2_sum__841, 7'h5b);
  assign p3_umul_144290_comb = umul32b_32b_x_7b(p2_sum__785, 7'h5b);
  assign p3_sum__1340_comb = p2_sum__1768 + p2_sum__1769;
  assign p3_sum__1341_comb = p2_sum__1770 + p2_sum__1771;
  assign p3_sum__1330_comb = p2_sum__1748 + p2_sum__1749;
  assign p3_sum__1331_comb = p2_sum__1750 + p2_sum__1751;
  assign p3_sum__1322_comb = p2_sum__1732 + p2_sum__1733;
  assign p3_sum__1323_comb = p2_sum__1734 + p2_sum__1735;
  assign p3_sum__1308_comb = p2_sum__1704 + p2_sum__1705;
  assign p3_sum__1309_comb = p2_sum__1706 + p2_sum__1707;
  assign p3_sum__1298_comb = p2_sum__1684 + p2_sum__1685;
  assign p3_sum__1299_comb = p2_sum__1686 + p2_sum__1687;
  assign p3_sum__1284_comb = p2_sum__1656 + p2_sum__1657;
  assign p3_sum__1285_comb = p2_sum__1658 + p2_sum__1659;
  assign p3_sum__1276_comb = p2_sum__1640 + p2_sum__1641;
  assign p3_sum__1277_comb = p2_sum__1642 + p2_sum__1643;
  assign p3_sum__1266_comb = p2_sum__1620 + p2_sum__1621;
  assign p3_sum__1267_comb = p2_sum__1622 + p2_sum__1623;
  assign p3_sum__1118_comb = p2_sum__1324 + p2_sum__1325;
  assign p3_sum__1097_comb = p2_sum__1282 + p2_sum__1283;
  assign p3_sum__1129_comb = p2_sum__1346 + p2_sum__1347;
  assign p3_sum__1124_comb = p2_sum__1336 + p2_sum__1337;
  assign p3_sum__1111_comb = p2_sum__1310 + p2_sum__1311;
  assign p3_sum__1104_comb = p2_sum__1296 + p2_sum__1297;
  assign p3_sum__1091_comb = p2_sum__1270 + p2_sum__1271;
  assign p3_sum__1086_comb = p2_sum__1260 + p2_sum__1261;
  assign p3_sum__1348_comb = p3_sum__1784_comb + p3_sum__1785_comb;
  assign p3_sum__1349_comb = p3_sum__1786_comb + p3_sum__1787_comb;
  assign p3_sum__1318_comb = p3_sum__1724_comb + p3_sum__1725_comb;
  assign p3_sum__1319_comb = p3_sum__1726_comb + p3_sum__1727_comb;
  assign p3_sum__1342_comb = p3_sum__1772_comb + p3_sum__1773_comb;
  assign p3_sum__1343_comb = p3_sum__1774_comb + p3_sum__1775_comb;
  assign p3_sum__1306_comb = p3_sum__1700_comb + p3_sum__1701_comb;
  assign p3_sum__1307_comb = p3_sum__1702_comb + p3_sum__1703_comb;
  assign p3_sum__1334_comb = p3_sum__1756_comb + p3_sum__1757_comb;
  assign p3_sum__1335_comb = p3_sum__1758_comb + p3_sum__1759_comb;
  assign p3_sum__1294_comb = p3_sum__1676_comb + p3_sum__1677_comb;
  assign p3_sum__1295_comb = p3_sum__1678_comb + p3_sum__1679_comb;
  assign p3_sum__1312_comb = p3_sum__1712_comb + p3_sum__1713_comb;
  assign p3_sum__1313_comb = p3_sum__1714_comb + p3_sum__1715_comb;
  assign p3_sum__1272_comb = p3_sum__1632_comb + p3_sum__1633_comb;
  assign p3_sum__1273_comb = p3_sum__1634_comb + p3_sum__1635_comb;
  assign p3_sum__1300_comb = p3_sum__1688_comb + p3_sum__1689_comb;
  assign p3_sum__1301_comb = p3_sum__1690_comb + p3_sum__1691_comb;
  assign p3_sum__1264_comb = p3_sum__1616_comb + p3_sum__1617_comb;
  assign p3_sum__1265_comb = p3_sum__1618_comb + p3_sum__1619_comb;
  assign p3_sum__1288_comb = p3_sum__1664_comb + p3_sum__1665_comb;
  assign p3_sum__1289_comb = p3_sum__1666_comb + p3_sum__1667_comb;
  assign p3_sum__1258_comb = p3_sum__1604_comb + p3_sum__1605_comb;
  assign p3_sum__1259_comb = p3_sum__1606_comb + p3_sum__1607_comb;
  assign p3_sum__1358_comb = p3_sum__1804_comb + p3_sum__1805_comb;
  assign p3_sum__1359_comb = p3_sum__1806_comb + p3_sum__1807_comb;
  assign p3_sum__1354_comb = p3_sum__1796_comb + p3_sum__1797_comb;
  assign p3_sum__1355_comb = p3_sum__1798_comb + p3_sum__1799_comb;
  assign p3_sum__1304_comb = p3_sum__1696_comb + p3_sum__1697_comb;
  assign p3_sum__1305_comb = p3_sum__1698_comb + p3_sum__1699_comb;
  assign p3_sum__1290_comb = p3_sum__1668_comb + p3_sum__1669_comb;
  assign p3_sum__1291_comb = p3_sum__1670_comb + p3_sum__1671_comb;
  assign p3_sum__1356_comb = p3_sum__1800_comb + p3_sum__1801_comb;
  assign p3_sum__1357_comb = p3_sum__1802_comb + p3_sum__1803_comb;
  assign p3_sum__1350_comb = p3_sum__1788_comb + p3_sum__1789_comb;
  assign p3_sum__1351_comb = p3_sum__1790_comb + p3_sum__1791_comb;
  assign p3_sum__1332_comb = p3_sum__1752_comb + p3_sum__1753_comb;
  assign p3_sum__1333_comb = p3_sum__1754_comb + p3_sum__1755_comb;
  assign p3_sum__1320_comb = p3_sum__1728_comb + p3_sum__1729_comb;
  assign p3_sum__1321_comb = p3_sum__1730_comb + p3_sum__1731_comb;
  assign p3_sum__1292_comb = p3_sum__1672_comb + p3_sum__1673_comb;
  assign p3_sum__1293_comb = p3_sum__1674_comb + p3_sum__1675_comb;
  assign p3_sum__1278_comb = p3_sum__1644_comb + p3_sum__1645_comb;
  assign p3_sum__1279_comb = p3_sum__1646_comb + p3_sum__1647_comb;
  assign p3_sum__1352_comb = p3_sum__1792_comb + p3_sum__1793_comb;
  assign p3_sum__1353_comb = p3_sum__1794_comb + p3_sum__1795_comb;
  assign p3_sum__1344_comb = p3_sum__1776_comb + p3_sum__1777_comb;
  assign p3_sum__1345_comb = p3_sum__1778_comb + p3_sum__1779_comb;
  assign p3_sum__1280_comb = p3_sum__1648_comb + p3_sum__1649_comb;
  assign p3_sum__1281_comb = p3_sum__1650_comb + p3_sum__1651_comb;
  assign p3_sum__1268_comb = p3_sum__1624_comb + p3_sum__1625_comb;
  assign p3_sum__1269_comb = p3_sum__1626_comb + p3_sum__1627_comb;
  assign p3_sum__1338_comb = p3_sum__1764_comb + p3_sum__1765_comb;
  assign p3_sum__1339_comb = p3_sum__1766_comb + p3_sum__1767_comb;
  assign p3_sum__1326_comb = p3_sum__1740_comb + p3_sum__1741_comb;
  assign p3_sum__1327_comb = p3_sum__1742_comb + p3_sum__1743_comb;
  assign p3_sum__1262_comb = p3_sum__1612_comb + p3_sum__1613_comb;
  assign p3_sum__1263_comb = p3_sum__1614_comb + p3_sum__1615_comb;
  assign p3_sum__1254_comb = p3_sum__1596_comb + p3_sum__1597_comb;
  assign p3_sum__1255_comb = p3_sum__1598_comb + p3_sum__1599_comb;
  assign p3_sum__1328_comb = p3_sum__1744_comb + p3_sum__1745_comb;
  assign p3_sum__1329_comb = p3_sum__1746_comb + p3_sum__1747_comb;
  assign p3_sum__1314_comb = p3_sum__1716_comb + p3_sum__1717_comb;
  assign p3_sum__1315_comb = p3_sum__1718_comb + p3_sum__1719_comb;
  assign p3_sum__1286_comb = p3_sum__1660_comb + p3_sum__1661_comb;
  assign p3_sum__1287_comb = p3_sum__1662_comb + p3_sum__1663_comb;
  assign p3_sum__1274_comb = p3_sum__1636_comb + p3_sum__1637_comb;
  assign p3_sum__1275_comb = p3_sum__1638_comb + p3_sum__1639_comb;
  assign p3_sum__1256_comb = p3_sum__1600_comb + p3_sum__1601_comb;
  assign p3_sum__1257_comb = p3_sum__1602_comb + p3_sum__1603_comb;
  assign p3_sum__1250_comb = p3_sum__1588_comb + p3_sum__1589_comb;
  assign p3_sum__1251_comb = p3_sum__1590_comb + p3_sum__1591_comb;
  assign p3_sum__1316_comb = p3_sum__1720_comb + p3_sum__1721_comb;
  assign p3_sum__1317_comb = p3_sum__1722_comb + p3_sum__1723_comb;
  assign p3_sum__1302_comb = p3_sum__1692_comb + p3_sum__1693_comb;
  assign p3_sum__1303_comb = p3_sum__1694_comb + p3_sum__1695_comb;
  assign p3_sum__1252_comb = p3_sum__1592_comb + p3_sum__1593_comb;
  assign p3_sum__1253_comb = p3_sum__1594_comb + p3_sum__1595_comb;
  assign p3_sum__1248_comb = p3_sum__1584_comb + p3_sum__1585_comb;
  assign p3_sum__1249_comb = p3_sum__1586_comb + p3_sum__1587_comb;
  assign p3_sum__1126_comb = p3_sum__1340_comb + p3_sum__1341_comb;
  assign p3_sum__1121_comb = p3_sum__1330_comb + p3_sum__1331_comb;
  assign p3_sum__1117_comb = p3_sum__1322_comb + p3_sum__1323_comb;
  assign p3_sum__1110_comb = p3_sum__1308_comb + p3_sum__1309_comb;
  assign p3_sum__1105_comb = p3_sum__1298_comb + p3_sum__1299_comb;
  assign p3_sum__1098_comb = p3_sum__1284_comb + p3_sum__1285_comb;
  assign p3_sum__1094_comb = p3_sum__1276_comb + p3_sum__1277_comb;
  assign p3_sum__1089_comb = p3_sum__1266_comb + p3_sum__1267_comb;
  assign p3_add_144499_comb = p3_sum__1118_comb + 25'h000_0001;
  assign p3_add_144500_comb = p3_sum__1097_comb + 25'h000_0001;
  assign p3_add_144531_comb = p3_sum__1129_comb + 25'h000_0001;
  assign p3_add_144532_comb = p3_sum__1124_comb + 25'h000_0001;
  assign p3_add_144533_comb = p3_sum__1111_comb + 25'h000_0001;
  assign p3_add_144534_comb = p3_sum__1104_comb + 25'h000_0001;
  assign p3_add_144535_comb = p3_sum__1091_comb + 25'h000_0001;
  assign p3_add_144536_comb = p3_sum__1086_comb + 25'h000_0001;
  assign p3_sum__1130_comb = p3_sum__1348_comb + p3_sum__1349_comb;
  assign p3_sum__1115_comb = p3_sum__1318_comb + p3_sum__1319_comb;
  assign p3_sum__1127_comb = p3_sum__1342_comb + p3_sum__1343_comb;
  assign p3_sum__1109_comb = p3_sum__1306_comb + p3_sum__1307_comb;
  assign p3_sum__1123_comb = p3_sum__1334_comb + p3_sum__1335_comb;
  assign p3_sum__1103_comb = p3_sum__1294_comb + p3_sum__1295_comb;
  assign p3_sum__1112_comb = p3_sum__1312_comb + p3_sum__1313_comb;
  assign p3_sum__1092_comb = p3_sum__1272_comb + p3_sum__1273_comb;
  assign p3_sum__1106_comb = p3_sum__1300_comb + p3_sum__1301_comb;
  assign p3_sum__1088_comb = p3_sum__1264_comb + p3_sum__1265_comb;
  assign p3_sum__1100_comb = p3_sum__1288_comb + p3_sum__1289_comb;
  assign p3_sum__1085_comb = p3_sum__1258_comb + p3_sum__1259_comb;
  assign p3_sum__1135_comb = p3_sum__1358_comb + p3_sum__1359_comb;
  assign p3_sum__1133_comb = p3_sum__1354_comb + p3_sum__1355_comb;
  assign p3_sum__1108_comb = p3_sum__1304_comb + p3_sum__1305_comb;
  assign p3_sum__1101_comb = p3_sum__1290_comb + p3_sum__1291_comb;
  assign p3_sum__1134_comb = p3_sum__1356_comb + p3_sum__1357_comb;
  assign p3_sum__1131_comb = p3_sum__1350_comb + p3_sum__1351_comb;
  assign p3_sum__1122_comb = p3_sum__1332_comb + p3_sum__1333_comb;
  assign p3_sum__1116_comb = p3_sum__1320_comb + p3_sum__1321_comb;
  assign p3_sum__1102_comb = p3_sum__1292_comb + p3_sum__1293_comb;
  assign p3_sum__1095_comb = p3_sum__1278_comb + p3_sum__1279_comb;
  assign p3_sum__1132_comb = p3_sum__1352_comb + p3_sum__1353_comb;
  assign p3_sum__1128_comb = p3_sum__1344_comb + p3_sum__1345_comb;
  assign p3_sum__1096_comb = p3_sum__1280_comb + p3_sum__1281_comb;
  assign p3_sum__1090_comb = p3_sum__1268_comb + p3_sum__1269_comb;
  assign p3_sum__1125_comb = p3_sum__1338_comb + p3_sum__1339_comb;
  assign p3_sum__1119_comb = p3_sum__1326_comb + p3_sum__1327_comb;
  assign p3_sum__1087_comb = p3_sum__1262_comb + p3_sum__1263_comb;
  assign p3_sum__1083_comb = p3_sum__1254_comb + p3_sum__1255_comb;
  assign p3_sum__1120_comb = p3_sum__1328_comb + p3_sum__1329_comb;
  assign p3_sum__1113_comb = p3_sum__1314_comb + p3_sum__1315_comb;
  assign p3_sum__1099_comb = p3_sum__1286_comb + p3_sum__1287_comb;
  assign p3_sum__1093_comb = p3_sum__1274_comb + p3_sum__1275_comb;
  assign p3_sum__1084_comb = p3_sum__1256_comb + p3_sum__1257_comb;
  assign p3_sum__1081_comb = p3_sum__1250_comb + p3_sum__1251_comb;
  assign p3_sum__1114_comb = p3_sum__1316_comb + p3_sum__1317_comb;
  assign p3_sum__1107_comb = p3_sum__1302_comb + p3_sum__1303_comb;
  assign p3_sum__1082_comb = p3_sum__1252_comb + p3_sum__1253_comb;
  assign p3_sum__1080_comb = p3_sum__1248_comb + p3_sum__1249_comb;
  assign p3_add_144491_comb = p3_umul_144259_comb[31:7] + 25'h000_0001;
  assign p3_add_144492_comb = p3_umul_144260_comb[31:7] + 25'h000_0001;
  assign p3_add_144507_comb = p3_umul_144285_comb[31:7] + 25'h000_0001;
  assign p3_add_144508_comb = p3_umul_144286_comb[31:7] + 25'h000_0001;
  assign p3_add_144509_comb = p3_umul_144287_comb[31:7] + 25'h000_0001;
  assign p3_add_144510_comb = p3_umul_144288_comb[31:7] + 25'h000_0001;
  assign p3_add_144511_comb = p3_umul_144289_comb[31:7] + 25'h000_0001;
  assign p3_add_144512_comb = p3_umul_144290_comb[31:7] + 25'h000_0001;
  assign p3_add_144515_comb = p3_sum__1126_comb + 25'h000_0001;
  assign p3_add_144516_comb = p3_sum__1121_comb + 25'h000_0001;
  assign p3_add_144527_comb = p3_sum__1117_comb + 25'h000_0001;
  assign p3_add_144528_comb = p3_sum__1110_comb + 25'h000_0001;
  assign p3_add_144539_comb = p3_sum__1105_comb + 25'h000_0001;
  assign p3_add_144540_comb = p3_sum__1098_comb + 25'h000_0001;
  assign p3_add_144551_comb = p3_sum__1094_comb + 25'h000_0001;
  assign p3_add_144552_comb = p3_sum__1089_comb + 25'h000_0001;
  assign p3_add_144493_comb = p3_sum__1130_comb + 25'h000_0001;
  assign p3_add_144494_comb = p3_sum__1115_comb + 25'h000_0001;
  assign p3_add_144495_comb = p3_sum__1127_comb + 25'h000_0001;
  assign p3_add_144496_comb = p3_sum__1109_comb + 25'h000_0001;
  assign p3_add_144497_comb = p3_sum__1123_comb + 25'h000_0001;
  assign p3_add_144498_comb = p3_sum__1103_comb + 25'h000_0001;
  assign p3_add_144501_comb = p3_sum__1112_comb + 25'h000_0001;
  assign p3_add_144502_comb = p3_sum__1092_comb + 25'h000_0001;
  assign p3_add_144503_comb = p3_sum__1106_comb + 25'h000_0001;
  assign p3_add_144504_comb = p3_sum__1088_comb + 25'h000_0001;
  assign p3_add_144505_comb = p3_sum__1100_comb + 25'h000_0001;
  assign p3_add_144506_comb = p3_sum__1085_comb + 25'h000_0001;
  assign p3_add_144513_comb = p3_sum__1135_comb + 25'h000_0001;
  assign p3_add_144514_comb = p3_sum__1133_comb + 25'h000_0001;
  assign p3_add_144517_comb = p3_sum__1108_comb + 25'h000_0001;
  assign p3_add_144518_comb = p3_sum__1101_comb + 25'h000_0001;
  assign p3_add_144519_comb = p3_sum__1134_comb + 25'h000_0001;
  assign p3_add_144520_comb = p3_sum__1131_comb + 25'h000_0001;
  assign p3_add_144521_comb = p3_sum__1122_comb + 25'h000_0001;
  assign p3_add_144522_comb = p3_sum__1116_comb + 25'h000_0001;
  assign p3_add_144523_comb = p3_sum__1102_comb + 25'h000_0001;
  assign p3_add_144524_comb = p3_sum__1095_comb + 25'h000_0001;
  assign p3_add_144525_comb = p3_sum__1132_comb + 25'h000_0001;
  assign p3_add_144526_comb = p3_sum__1128_comb + 25'h000_0001;
  assign p3_add_144529_comb = p3_sum__1096_comb + 25'h000_0001;
  assign p3_add_144530_comb = p3_sum__1090_comb + 25'h000_0001;
  assign p3_add_144537_comb = p3_sum__1125_comb + 25'h000_0001;
  assign p3_add_144538_comb = p3_sum__1119_comb + 25'h000_0001;
  assign p3_add_144541_comb = p3_sum__1087_comb + 25'h000_0001;
  assign p3_add_144542_comb = p3_sum__1083_comb + 25'h000_0001;
  assign p3_add_144543_comb = p3_sum__1120_comb + 25'h000_0001;
  assign p3_add_144544_comb = p3_sum__1113_comb + 25'h000_0001;
  assign p3_add_144545_comb = p3_sum__1099_comb + 25'h000_0001;
  assign p3_add_144546_comb = p3_sum__1093_comb + 25'h000_0001;
  assign p3_add_144547_comb = p3_sum__1084_comb + 25'h000_0001;
  assign p3_add_144548_comb = p3_sum__1081_comb + 25'h000_0001;
  assign p3_add_144549_comb = p3_sum__1114_comb + 25'h000_0001;
  assign p3_add_144550_comb = p3_sum__1107_comb + 25'h000_0001;
  assign p3_add_144553_comb = p3_sum__1082_comb + 25'h000_0001;
  assign p3_add_144554_comb = p3_sum__1080_comb + 25'h000_0001;
  assign p3_clipped__272_comb = $signed(p3_add_144499_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144499_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144499_comb[16:8]);
  assign p3_clipped__275_comb = $signed(p3_add_144500_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144500_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144500_comb[16:8]);
  assign p3_clipped__304_comb = $signed(p3_add_144531_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144531_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144531_comb[16:8]);
  assign p3_clipped__305_comb = $signed(p3_add_144532_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144532_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144532_comb[16:8]);
  assign p3_clipped__273_comb = $signed(p3_add_144533_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144533_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144533_comb[16:8]);
  assign p3_clipped__274_comb = $signed(p3_add_144534_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144534_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144534_comb[16:8]);
  assign p3_clipped__306_comb = $signed(p3_add_144535_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144535_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144535_comb[16:8]);
  assign p3_clipped__307_comb = $signed(p3_add_144536_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144536_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144536_comb[16:8]);
  assign p3_clipped__256_comb = $signed(p3_add_144491_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144491_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144491_comb[16:8]);
  assign p3_clipped__259_comb = $signed(p3_add_144492_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144492_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144492_comb[16:8]);
  assign p3_clipped__288_comb = $signed(p3_add_144507_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144507_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144507_comb[16:8]);
  assign p3_clipped__289_comb = $signed(p3_add_144508_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144508_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144508_comb[16:8]);
  assign p3_clipped__257_comb = $signed(p3_add_144509_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144509_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144509_comb[16:8]);
  assign p3_clipped__258_comb = $signed(p3_add_144510_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144510_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144510_comb[16:8]);
  assign p3_clipped__290_comb = $signed(p3_add_144511_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144511_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144511_comb[16:8]);
  assign p3_clipped__291_comb = $signed(p3_add_144512_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144512_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144512_comb[16:8]);
  assign p3_clipped__261_comb = $signed(p3_add_144515_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144515_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144515_comb[16:8]);
  assign p3_clipped__262_comb = $signed(p3_add_144516_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144516_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144516_comb[16:8]);
  assign p3_clipped__269_comb = $signed(p3_add_144527_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144527_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144527_comb[16:8]);
  assign p3_clipped__270_comb = $signed(p3_add_144528_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144528_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144528_comb[16:8]);
  assign p3_clipped__277_comb = $signed(p3_add_144539_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144539_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144539_comb[16:8]);
  assign p3_clipped__278_comb = $signed(p3_add_144540_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144540_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144540_comb[16:8]);
  assign p3_clipped__285_comb = $signed(p3_add_144551_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144551_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144551_comb[16:8]);
  assign p3_clipped__286_comb = $signed(p3_add_144552_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144552_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144552_comb[16:8]);
  assign p3_clipped__260_comb = $signed(p3_add_144493_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144493_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144493_comb[16:8]);
  assign p3_clipped__263_comb = $signed(p3_add_144494_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144494_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144494_comb[16:8]);
  assign p3_clipped__264_comb = $signed(p3_add_144495_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144495_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144495_comb[16:8]);
  assign p3_clipped__267_comb = $signed(p3_add_144496_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144496_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144496_comb[16:8]);
  assign p3_clipped__268_comb = $signed(p3_add_144497_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144497_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144497_comb[16:8]);
  assign p3_clipped__271_comb = $signed(p3_add_144498_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144498_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144498_comb[16:8]);
  assign p3_clipped__276_comb = $signed(p3_add_144501_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144501_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144501_comb[16:8]);
  assign p3_clipped__279_comb = $signed(p3_add_144502_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144502_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144502_comb[16:8]);
  assign p3_clipped__280_comb = $signed(p3_add_144503_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144503_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144503_comb[16:8]);
  assign p3_clipped__283_comb = $signed(p3_add_144504_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144504_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144504_comb[16:8]);
  assign p3_clipped__284_comb = $signed(p3_add_144505_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144505_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144505_comb[16:8]);
  assign p3_clipped__287_comb = $signed(p3_add_144506_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144506_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144506_comb[16:8]);
  assign p3_clipped__292_comb = $signed(p3_add_144513_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144513_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144513_comb[16:8]);
  assign p3_clipped__293_comb = $signed(p3_add_144514_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144514_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144514_comb[16:8]);
  assign p3_clipped__294_comb = $signed(p3_add_144517_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144517_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144517_comb[16:8]);
  assign p3_clipped__295_comb = $signed(p3_add_144518_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144518_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144518_comb[16:8]);
  assign p3_clipped__296_comb = $signed(p3_add_144519_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144519_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144519_comb[16:8]);
  assign p3_clipped__297_comb = $signed(p3_add_144520_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144520_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144520_comb[16:8]);
  assign p3_clipped__265_comb = $signed(p3_add_144521_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144521_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144521_comb[16:8]);
  assign p3_clipped__266_comb = $signed(p3_add_144522_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144522_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144522_comb[16:8]);
  assign p3_clipped__298_comb = $signed(p3_add_144523_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144523_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144523_comb[16:8]);
  assign p3_clipped__299_comb = $signed(p3_add_144524_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144524_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144524_comb[16:8]);
  assign p3_clipped__300_comb = $signed(p3_add_144525_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144525_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144525_comb[16:8]);
  assign p3_clipped__301_comb = $signed(p3_add_144526_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144526_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144526_comb[16:8]);
  assign p3_clipped__302_comb = $signed(p3_add_144529_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144529_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144529_comb[16:8]);
  assign p3_clipped__303_comb = $signed(p3_add_144530_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144530_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144530_comb[16:8]);
  assign p3_clipped__308_comb = $signed(p3_add_144537_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144537_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144537_comb[16:8]);
  assign p3_clipped__309_comb = $signed(p3_add_144538_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144538_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144538_comb[16:8]);
  assign p3_clipped__310_comb = $signed(p3_add_144541_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144541_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144541_comb[16:8]);
  assign p3_clipped__311_comb = $signed(p3_add_144542_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144542_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144542_comb[16:8]);
  assign p3_clipped__312_comb = $signed(p3_add_144543_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144543_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144543_comb[16:8]);
  assign p3_clipped__313_comb = $signed(p3_add_144544_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144544_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144544_comb[16:8]);
  assign p3_clipped__281_comb = $signed(p3_add_144545_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144545_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144545_comb[16:8]);
  assign p3_clipped__282_comb = $signed(p3_add_144546_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144546_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144546_comb[16:8]);
  assign p3_clipped__314_comb = $signed(p3_add_144547_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144547_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144547_comb[16:8]);
  assign p3_clipped__315_comb = $signed(p3_add_144548_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144548_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144548_comb[16:8]);
  assign p3_clipped__316_comb = $signed(p3_add_144549_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144549_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144549_comb[16:8]);
  assign p3_clipped__317_comb = $signed(p3_add_144550_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144550_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144550_comb[16:8]);
  assign p3_clipped__318_comb = $signed(p3_add_144553_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144553_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144553_comb[16:8]);
  assign p3_clipped__319_comb = $signed(p3_add_144554_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p3_add_144554_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p3_add_144554_comb[16:8]);
  assign p3_sign_ext_145195_comb = {{1{p3_clipped__256_comb[8]}}, p3_clipped__256_comb};
  assign p3_sign_ext_145196_comb = {{1{p3_clipped__259_comb[8]}}, p3_clipped__259_comb};
  assign p3_sign_ext_145201_comb = {{1{p3_clipped__288_comb[8]}}, p3_clipped__288_comb};
  assign p3_sign_ext_145202_comb = {{1{p3_clipped__289_comb[8]}}, p3_clipped__289_comb};
  assign p3_sign_ext_145203_comb = {{1{p3_clipped__257_comb[8]}}, p3_clipped__257_comb};
  assign p3_sign_ext_145204_comb = {{1{p3_clipped__258_comb[8]}}, p3_clipped__258_comb};
  assign p3_sign_ext_145205_comb = {{1{p3_clipped__290_comb[8]}}, p3_clipped__290_comb};
  assign p3_sign_ext_145206_comb = {{1{p3_clipped__291_comb[8]}}, p3_clipped__291_comb};
  assign p3_sign_ext_145207_comb = {{1{p3_clipped__261_comb[8]}}, p3_clipped__261_comb};
  assign p3_sign_ext_145208_comb = {{1{p3_clipped__262_comb[8]}}, p3_clipped__262_comb};
  assign p3_sign_ext_145209_comb = {{1{p3_clipped__269_comb[8]}}, p3_clipped__269_comb};
  assign p3_sign_ext_145210_comb = {{1{p3_clipped__270_comb[8]}}, p3_clipped__270_comb};
  assign p3_sign_ext_145223_comb = {{1{p3_clipped__277_comb[8]}}, p3_clipped__277_comb};
  assign p3_sign_ext_145224_comb = {{1{p3_clipped__278_comb[8]}}, p3_clipped__278_comb};
  assign p3_sign_ext_145225_comb = {{1{p3_clipped__285_comb[8]}}, p3_clipped__285_comb};
  assign p3_sign_ext_145226_comb = {{1{p3_clipped__286_comb[8]}}, p3_clipped__286_comb};
  assign p3_add_145227_comb = {{1{p3_clipped__272_comb[8]}}, p3_clipped__272_comb} + 10'h001;
  assign p3_add_145228_comb = {{1{p3_clipped__275_comb[8]}}, p3_clipped__275_comb} + 10'h001;
  assign p3_add_145229_comb = {{1{p3_clipped__304_comb[8]}}, p3_clipped__304_comb} + 10'h001;
  assign p3_add_145230_comb = {{1{p3_clipped__305_comb[8]}}, p3_clipped__305_comb} + 10'h001;
  assign p3_add_145231_comb = {{1{p3_clipped__273_comb[8]}}, p3_clipped__273_comb} + 10'h001;
  assign p3_add_145232_comb = {{1{p3_clipped__274_comb[8]}}, p3_clipped__274_comb} + 10'h001;
  assign p3_add_145233_comb = {{1{p3_clipped__306_comb[8]}}, p3_clipped__306_comb} + 10'h001;
  assign p3_add_145234_comb = {{1{p3_clipped__307_comb[8]}}, p3_clipped__307_comb} + 10'h001;

  // Registers for pipe stage 3:
  reg [8:0] p3_clipped__260;
  reg [8:0] p3_clipped__263;
  reg [8:0] p3_clipped__264;
  reg [8:0] p3_clipped__267;
  reg [8:0] p3_clipped__268;
  reg [8:0] p3_clipped__271;
  reg [8:0] p3_clipped__276;
  reg [8:0] p3_clipped__279;
  reg [8:0] p3_clipped__280;
  reg [8:0] p3_clipped__283;
  reg [8:0] p3_clipped__284;
  reg [8:0] p3_clipped__287;
  reg [8:0] p3_clipped__292;
  reg [8:0] p3_clipped__293;
  reg [8:0] p3_clipped__294;
  reg [8:0] p3_clipped__295;
  reg [8:0] p3_clipped__296;
  reg [8:0] p3_clipped__297;
  reg [8:0] p3_clipped__265;
  reg [8:0] p3_clipped__266;
  reg [8:0] p3_clipped__298;
  reg [8:0] p3_clipped__299;
  reg [8:0] p3_clipped__300;
  reg [8:0] p3_clipped__301;
  reg [8:0] p3_clipped__302;
  reg [8:0] p3_clipped__303;
  reg [8:0] p3_clipped__308;
  reg [8:0] p3_clipped__309;
  reg [8:0] p3_clipped__310;
  reg [8:0] p3_clipped__311;
  reg [8:0] p3_clipped__312;
  reg [8:0] p3_clipped__313;
  reg [8:0] p3_clipped__281;
  reg [8:0] p3_clipped__282;
  reg [8:0] p3_clipped__314;
  reg [8:0] p3_clipped__315;
  reg [8:0] p3_clipped__316;
  reg [8:0] p3_clipped__317;
  reg [8:0] p3_clipped__318;
  reg [8:0] p3_clipped__319;
  reg [9:0] p3_sign_ext_145195;
  reg [9:0] p3_sign_ext_145196;
  reg [9:0] p3_sign_ext_145201;
  reg [9:0] p3_sign_ext_145202;
  reg [9:0] p3_sign_ext_145203;
  reg [9:0] p3_sign_ext_145204;
  reg [9:0] p3_sign_ext_145205;
  reg [9:0] p3_sign_ext_145206;
  reg [9:0] p3_sign_ext_145207;
  reg [9:0] p3_sign_ext_145208;
  reg [9:0] p3_sign_ext_145209;
  reg [9:0] p3_sign_ext_145210;
  reg [9:0] p3_sign_ext_145223;
  reg [9:0] p3_sign_ext_145224;
  reg [9:0] p3_sign_ext_145225;
  reg [9:0] p3_sign_ext_145226;
  reg [9:0] p3_add_145227;
  reg [9:0] p3_add_145228;
  reg [9:0] p3_add_145229;
  reg [9:0] p3_add_145230;
  reg [9:0] p3_add_145231;
  reg [9:0] p3_add_145232;
  reg [9:0] p3_add_145233;
  reg [9:0] p3_add_145234;
  always @ (posedge clk) begin
    p3_clipped__260 <= p3_clipped__260_comb;
    p3_clipped__263 <= p3_clipped__263_comb;
    p3_clipped__264 <= p3_clipped__264_comb;
    p3_clipped__267 <= p3_clipped__267_comb;
    p3_clipped__268 <= p3_clipped__268_comb;
    p3_clipped__271 <= p3_clipped__271_comb;
    p3_clipped__276 <= p3_clipped__276_comb;
    p3_clipped__279 <= p3_clipped__279_comb;
    p3_clipped__280 <= p3_clipped__280_comb;
    p3_clipped__283 <= p3_clipped__283_comb;
    p3_clipped__284 <= p3_clipped__284_comb;
    p3_clipped__287 <= p3_clipped__287_comb;
    p3_clipped__292 <= p3_clipped__292_comb;
    p3_clipped__293 <= p3_clipped__293_comb;
    p3_clipped__294 <= p3_clipped__294_comb;
    p3_clipped__295 <= p3_clipped__295_comb;
    p3_clipped__296 <= p3_clipped__296_comb;
    p3_clipped__297 <= p3_clipped__297_comb;
    p3_clipped__265 <= p3_clipped__265_comb;
    p3_clipped__266 <= p3_clipped__266_comb;
    p3_clipped__298 <= p3_clipped__298_comb;
    p3_clipped__299 <= p3_clipped__299_comb;
    p3_clipped__300 <= p3_clipped__300_comb;
    p3_clipped__301 <= p3_clipped__301_comb;
    p3_clipped__302 <= p3_clipped__302_comb;
    p3_clipped__303 <= p3_clipped__303_comb;
    p3_clipped__308 <= p3_clipped__308_comb;
    p3_clipped__309 <= p3_clipped__309_comb;
    p3_clipped__310 <= p3_clipped__310_comb;
    p3_clipped__311 <= p3_clipped__311_comb;
    p3_clipped__312 <= p3_clipped__312_comb;
    p3_clipped__313 <= p3_clipped__313_comb;
    p3_clipped__281 <= p3_clipped__281_comb;
    p3_clipped__282 <= p3_clipped__282_comb;
    p3_clipped__314 <= p3_clipped__314_comb;
    p3_clipped__315 <= p3_clipped__315_comb;
    p3_clipped__316 <= p3_clipped__316_comb;
    p3_clipped__317 <= p3_clipped__317_comb;
    p3_clipped__318 <= p3_clipped__318_comb;
    p3_clipped__319 <= p3_clipped__319_comb;
    p3_sign_ext_145195 <= p3_sign_ext_145195_comb;
    p3_sign_ext_145196 <= p3_sign_ext_145196_comb;
    p3_sign_ext_145201 <= p3_sign_ext_145201_comb;
    p3_sign_ext_145202 <= p3_sign_ext_145202_comb;
    p3_sign_ext_145203 <= p3_sign_ext_145203_comb;
    p3_sign_ext_145204 <= p3_sign_ext_145204_comb;
    p3_sign_ext_145205 <= p3_sign_ext_145205_comb;
    p3_sign_ext_145206 <= p3_sign_ext_145206_comb;
    p3_sign_ext_145207 <= p3_sign_ext_145207_comb;
    p3_sign_ext_145208 <= p3_sign_ext_145208_comb;
    p3_sign_ext_145209 <= p3_sign_ext_145209_comb;
    p3_sign_ext_145210 <= p3_sign_ext_145210_comb;
    p3_sign_ext_145223 <= p3_sign_ext_145223_comb;
    p3_sign_ext_145224 <= p3_sign_ext_145224_comb;
    p3_sign_ext_145225 <= p3_sign_ext_145225_comb;
    p3_sign_ext_145226 <= p3_sign_ext_145226_comb;
    p3_add_145227 <= p3_add_145227_comb;
    p3_add_145228 <= p3_add_145228_comb;
    p3_add_145229 <= p3_add_145229_comb;
    p3_add_145230 <= p3_add_145230_comb;
    p3_add_145231 <= p3_add_145231_comb;
    p3_add_145232 <= p3_add_145232_comb;
    p3_add_145233 <= p3_add_145233_comb;
    p3_add_145234 <= p3_add_145234_comb;
  end

  // ===== Pipe stage 4:
  wire [9:0] p4_add_145459_comb;
  wire [9:0] p4_add_145460_comb;
  wire [9:0] p4_add_145473_comb;
  wire [9:0] p4_add_145474_comb;
  wire [9:0] p4_add_145475_comb;
  wire [9:0] p4_add_145476_comb;
  wire [9:0] p4_add_145477_comb;
  wire [9:0] p4_add_145478_comb;
  wire [9:0] p4_add_145481_comb;
  wire [9:0] p4_add_145482_comb;
  wire [9:0] p4_add_145493_comb;
  wire [9:0] p4_add_145494_comb;
  wire [9:0] p4_add_145499_comb;
  wire [9:0] p4_add_145500_comb;
  wire [9:0] p4_add_145511_comb;
  wire [9:0] p4_add_145512_comb;
  wire [1:0] p4_bit_slice_145523_comb;
  wire [1:0] p4_bit_slice_145524_comb;
  wire [1:0] p4_bit_slice_145555_comb;
  wire [1:0] p4_bit_slice_145556_comb;
  wire [1:0] p4_bit_slice_145557_comb;
  wire [1:0] p4_bit_slice_145558_comb;
  wire [1:0] p4_bit_slice_145559_comb;
  wire [1:0] p4_bit_slice_145560_comb;
  wire [9:0] p4_add_145461_comb;
  wire [9:0] p4_add_145462_comb;
  wire [9:0] p4_add_145463_comb;
  wire [9:0] p4_add_145464_comb;
  wire [9:0] p4_add_145465_comb;
  wire [9:0] p4_add_145466_comb;
  wire [9:0] p4_add_145467_comb;
  wire [9:0] p4_add_145468_comb;
  wire [9:0] p4_add_145469_comb;
  wire [9:0] p4_add_145470_comb;
  wire [9:0] p4_add_145471_comb;
  wire [9:0] p4_add_145472_comb;
  wire [9:0] p4_add_145479_comb;
  wire [9:0] p4_add_145480_comb;
  wire [9:0] p4_add_145483_comb;
  wire [9:0] p4_add_145484_comb;
  wire [9:0] p4_add_145485_comb;
  wire [9:0] p4_add_145486_comb;
  wire [9:0] p4_add_145487_comb;
  wire [9:0] p4_add_145488_comb;
  wire [9:0] p4_add_145489_comb;
  wire [9:0] p4_add_145490_comb;
  wire [9:0] p4_add_145491_comb;
  wire [9:0] p4_add_145492_comb;
  wire [9:0] p4_add_145495_comb;
  wire [9:0] p4_add_145496_comb;
  wire [9:0] p4_add_145497_comb;
  wire [9:0] p4_add_145498_comb;
  wire [9:0] p4_add_145501_comb;
  wire [9:0] p4_add_145502_comb;
  wire [9:0] p4_add_145503_comb;
  wire [9:0] p4_add_145504_comb;
  wire [9:0] p4_add_145505_comb;
  wire [9:0] p4_add_145506_comb;
  wire [9:0] p4_add_145507_comb;
  wire [9:0] p4_add_145508_comb;
  wire [9:0] p4_add_145509_comb;
  wire [9:0] p4_add_145510_comb;
  wire [9:0] p4_add_145513_comb;
  wire [9:0] p4_add_145514_comb;
  wire [1:0] p4_bit_slice_145515_comb;
  wire [1:0] p4_bit_slice_145516_comb;
  wire [1:0] p4_bit_slice_145531_comb;
  wire [1:0] p4_bit_slice_145532_comb;
  wire [1:0] p4_bit_slice_145533_comb;
  wire [1:0] p4_bit_slice_145534_comb;
  wire [1:0] p4_bit_slice_145535_comb;
  wire [1:0] p4_bit_slice_145536_comb;
  wire [1:0] p4_bit_slice_145539_comb;
  wire [1:0] p4_bit_slice_145540_comb;
  wire [1:0] p4_bit_slice_145551_comb;
  wire [1:0] p4_bit_slice_145552_comb;
  wire [1:0] p4_bit_slice_145563_comb;
  wire [1:0] p4_bit_slice_145564_comb;
  wire [1:0] p4_bit_slice_145575_comb;
  wire [1:0] p4_bit_slice_145576_comb;
  wire [1:0] p4_bit_slice_145517_comb;
  wire [1:0] p4_bit_slice_145518_comb;
  wire [1:0] p4_bit_slice_145519_comb;
  wire [1:0] p4_bit_slice_145520_comb;
  wire [1:0] p4_bit_slice_145521_comb;
  wire [1:0] p4_bit_slice_145522_comb;
  wire [1:0] p4_bit_slice_145525_comb;
  wire [1:0] p4_bit_slice_145526_comb;
  wire [1:0] p4_bit_slice_145527_comb;
  wire [1:0] p4_bit_slice_145528_comb;
  wire [1:0] p4_bit_slice_145529_comb;
  wire [1:0] p4_bit_slice_145530_comb;
  wire [1:0] p4_bit_slice_145537_comb;
  wire [1:0] p4_bit_slice_145538_comb;
  wire [1:0] p4_bit_slice_145541_comb;
  wire [1:0] p4_bit_slice_145542_comb;
  wire [1:0] p4_bit_slice_145543_comb;
  wire [1:0] p4_bit_slice_145544_comb;
  wire [1:0] p4_bit_slice_145545_comb;
  wire [1:0] p4_bit_slice_145546_comb;
  wire [1:0] p4_bit_slice_145547_comb;
  wire [1:0] p4_bit_slice_145548_comb;
  wire [1:0] p4_bit_slice_145549_comb;
  wire [1:0] p4_bit_slice_145550_comb;
  wire [1:0] p4_bit_slice_145553_comb;
  wire [1:0] p4_bit_slice_145554_comb;
  wire [1:0] p4_bit_slice_145561_comb;
  wire [1:0] p4_bit_slice_145562_comb;
  wire [1:0] p4_bit_slice_145565_comb;
  wire [1:0] p4_bit_slice_145566_comb;
  wire [1:0] p4_bit_slice_145567_comb;
  wire [1:0] p4_bit_slice_145568_comb;
  wire [1:0] p4_bit_slice_145569_comb;
  wire [1:0] p4_bit_slice_145570_comb;
  wire [1:0] p4_bit_slice_145571_comb;
  wire [1:0] p4_bit_slice_145572_comb;
  wire [1:0] p4_bit_slice_145573_comb;
  wire [1:0] p4_bit_slice_145574_comb;
  wire [1:0] p4_bit_slice_145577_comb;
  wire [1:0] p4_bit_slice_145578_comb;
  wire [2:0] p4_add_145715_comb;
  wire [2:0] p4_add_145716_comb;
  wire [2:0] p4_add_145747_comb;
  wire [2:0] p4_add_145748_comb;
  wire [2:0] p4_add_145749_comb;
  wire [2:0] p4_add_145750_comb;
  wire [2:0] p4_add_145751_comb;
  wire [2:0] p4_add_145752_comb;
  wire [2:0] p4_add_145707_comb;
  wire [2:0] p4_add_145708_comb;
  wire [2:0] p4_add_145723_comb;
  wire [2:0] p4_add_145724_comb;
  wire [2:0] p4_add_145725_comb;
  wire [2:0] p4_add_145726_comb;
  wire [2:0] p4_add_145727_comb;
  wire [2:0] p4_add_145728_comb;
  wire [2:0] p4_add_145731_comb;
  wire [2:0] p4_add_145732_comb;
  wire [2:0] p4_add_145743_comb;
  wire [2:0] p4_add_145744_comb;
  wire [2:0] p4_add_145755_comb;
  wire [2:0] p4_add_145756_comb;
  wire [2:0] p4_add_145767_comb;
  wire [2:0] p4_add_145768_comb;
  wire [2:0] p4_add_145709_comb;
  wire [2:0] p4_add_145710_comb;
  wire [2:0] p4_add_145711_comb;
  wire [2:0] p4_add_145712_comb;
  wire [2:0] p4_add_145713_comb;
  wire [2:0] p4_add_145714_comb;
  wire [2:0] p4_add_145717_comb;
  wire [2:0] p4_add_145718_comb;
  wire [2:0] p4_add_145719_comb;
  wire [2:0] p4_add_145720_comb;
  wire [2:0] p4_add_145721_comb;
  wire [2:0] p4_add_145722_comb;
  wire [2:0] p4_add_145729_comb;
  wire [2:0] p4_add_145730_comb;
  wire [2:0] p4_add_145733_comb;
  wire [2:0] p4_add_145734_comb;
  wire [2:0] p4_add_145735_comb;
  wire [2:0] p4_add_145736_comb;
  wire [2:0] p4_add_145737_comb;
  wire [2:0] p4_add_145738_comb;
  wire [2:0] p4_add_145739_comb;
  wire [2:0] p4_add_145740_comb;
  wire [2:0] p4_add_145741_comb;
  wire [2:0] p4_add_145742_comb;
  wire [2:0] p4_add_145745_comb;
  wire [2:0] p4_add_145746_comb;
  wire [2:0] p4_add_145753_comb;
  wire [2:0] p4_add_145754_comb;
  wire [2:0] p4_add_145757_comb;
  wire [2:0] p4_add_145758_comb;
  wire [2:0] p4_add_145759_comb;
  wire [2:0] p4_add_145760_comb;
  wire [2:0] p4_add_145761_comb;
  wire [2:0] p4_add_145762_comb;
  wire [2:0] p4_add_145763_comb;
  wire [2:0] p4_add_145764_comb;
  wire [2:0] p4_add_145765_comb;
  wire [2:0] p4_add_145766_comb;
  wire [2:0] p4_add_145769_comb;
  wire [2:0] p4_add_145770_comb;
  wire [7:0] p4_clipped__44_comb;
  wire [7:0] p4_clipped__92_comb;
  wire [7:0] p4_clipped__12_comb;
  wire [7:0] p4_clipped__28_comb;
  wire [7:0] p4_clipped__60_comb;
  wire [7:0] p4_clipped__76_comb;
  wire [7:0] p4_clipped__108_comb;
  wire [7:0] p4_clipped__124_comb;
  wire [7:0] p4_clipped__40_comb;
  wire [7:0] p4_clipped__88_comb;
  wire [7:0] p4_clipped__8_comb;
  wire [7:0] p4_clipped__24_comb;
  wire [7:0] p4_clipped__56_comb;
  wire [7:0] p4_clipped__72_comb;
  wire [7:0] p4_clipped__104_comb;
  wire [7:0] p4_clipped__120_comb;
  wire [7:0] p4_clipped__57_comb;
  wire [7:0] p4_clipped__73_comb;
  wire [7:0] p4_clipped__59_comb;
  wire [7:0] p4_clipped__75_comb;
  wire [7:0] p4_clipped__61_comb;
  wire [7:0] p4_clipped__77_comb;
  wire [7:0] p4_clipped__63_comb;
  wire [7:0] p4_clipped__79_comb;
  wire [7:0] p4_clipped__41_comb;
  wire [7:0] p4_clipped__89_comb;
  wire [7:0] p4_clipped__42_comb;
  wire [7:0] p4_clipped__90_comb;
  wire [7:0] p4_clipped__43_comb;
  wire [7:0] p4_clipped__91_comb;
  wire [7:0] p4_clipped__45_comb;
  wire [7:0] p4_clipped__93_comb;
  wire [7:0] p4_clipped__46_comb;
  wire [7:0] p4_clipped__94_comb;
  wire [7:0] p4_clipped__47_comb;
  wire [7:0] p4_clipped__95_comb;
  wire [7:0] p4_clipped__9_comb;
  wire [7:0] p4_clipped__25_comb;
  wire [7:0] p4_clipped__105_comb;
  wire [7:0] p4_clipped__121_comb;
  wire [7:0] p4_clipped__10_comb;
  wire [7:0] p4_clipped__26_comb;
  wire [7:0] p4_clipped__58_comb;
  wire [7:0] p4_clipped__74_comb;
  wire [7:0] p4_clipped__106_comb;
  wire [7:0] p4_clipped__122_comb;
  wire [7:0] p4_clipped__11_comb;
  wire [7:0] p4_clipped__27_comb;
  wire [7:0] p4_clipped__107_comb;
  wire [7:0] p4_clipped__123_comb;
  wire [7:0] p4_clipped__13_comb;
  wire [7:0] p4_clipped__29_comb;
  wire [7:0] p4_clipped__109_comb;
  wire [7:0] p4_clipped__125_comb;
  wire [7:0] p4_clipped__14_comb;
  wire [7:0] p4_clipped__30_comb;
  wire [7:0] p4_clipped__62_comb;
  wire [7:0] p4_clipped__78_comb;
  wire [7:0] p4_clipped__110_comb;
  wire [7:0] p4_clipped__126_comb;
  wire [7:0] p4_clipped__15_comb;
  wire [7:0] p4_clipped__31_comb;
  wire [7:0] p4_clipped__111_comb;
  wire [7:0] p4_clipped__127_comb;
  wire p4_bit_slice_146155_comb;
  wire p4_bit_slice_146156_comb;
  wire p4_bit_slice_146159_comb;
  wire p4_bit_slice_146160_comb;
  wire p4_bit_slice_146161_comb;
  wire p4_bit_slice_146162_comb;
  wire p4_bit_slice_146163_comb;
  wire p4_bit_slice_146164_comb;
  wire p4_bit_slice_146165_comb;
  wire p4_bit_slice_146166_comb;
  wire p4_bit_slice_146167_comb;
  wire p4_bit_slice_146168_comb;
  wire p4_bit_slice_146175_comb;
  wire p4_bit_slice_146176_comb;
  wire p4_bit_slice_146177_comb;
  wire p4_bit_slice_146178_comb;
  wire [6:0] p4_bit_slice_146179_comb;
  wire [6:0] p4_bit_slice_146180_comb;
  wire p4_not_146181_comb;
  wire [6:0] p4_bit_slice_146182_comb;
  wire p4_not_146183_comb;
  wire [6:0] p4_bit_slice_146184_comb;
  wire [6:0] p4_bit_slice_146185_comb;
  wire [6:0] p4_bit_slice_146186_comb;
  wire [6:0] p4_bit_slice_146187_comb;
  wire [6:0] p4_bit_slice_146188_comb;
  wire [6:0] p4_bit_slice_146189_comb;
  wire [6:0] p4_bit_slice_146190_comb;
  wire [6:0] p4_bit_slice_146191_comb;
  wire [6:0] p4_bit_slice_146192_comb;
  wire [6:0] p4_bit_slice_146193_comb;
  wire [6:0] p4_bit_slice_146194_comb;
  wire p4_not_146195_comb;
  wire [6:0] p4_bit_slice_146196_comb;
  wire p4_not_146197_comb;
  wire [6:0] p4_bit_slice_146198_comb;
  wire p4_not_146199_comb;
  wire [6:0] p4_bit_slice_146200_comb;
  wire p4_not_146201_comb;
  wire [6:0] p4_bit_slice_146202_comb;
  wire p4_not_146203_comb;
  wire [6:0] p4_bit_slice_146204_comb;
  wire p4_not_146205_comb;
  wire [6:0] p4_bit_slice_146206_comb;
  wire [6:0] p4_bit_slice_146207_comb;
  wire [6:0] p4_bit_slice_146208_comb;
  wire [6:0] p4_bit_slice_146209_comb;
  wire [6:0] p4_bit_slice_146210_comb;
  assign p4_add_145459_comb = p3_sign_ext_145195 + 10'h001;
  assign p4_add_145460_comb = p3_sign_ext_145196 + 10'h001;
  assign p4_add_145473_comb = p3_sign_ext_145201 + 10'h001;
  assign p4_add_145474_comb = p3_sign_ext_145202 + 10'h001;
  assign p4_add_145475_comb = p3_sign_ext_145203 + 10'h001;
  assign p4_add_145476_comb = p3_sign_ext_145204 + 10'h001;
  assign p4_add_145477_comb = p3_sign_ext_145205 + 10'h001;
  assign p4_add_145478_comb = p3_sign_ext_145206 + 10'h001;
  assign p4_add_145481_comb = p3_sign_ext_145207 + 10'h001;
  assign p4_add_145482_comb = p3_sign_ext_145208 + 10'h001;
  assign p4_add_145493_comb = p3_sign_ext_145209 + 10'h001;
  assign p4_add_145494_comb = p3_sign_ext_145210 + 10'h001;
  assign p4_add_145499_comb = p3_sign_ext_145223 + 10'h001;
  assign p4_add_145500_comb = p3_sign_ext_145224 + 10'h001;
  assign p4_add_145511_comb = p3_sign_ext_145225 + 10'h001;
  assign p4_add_145512_comb = p3_sign_ext_145226 + 10'h001;
  assign p4_bit_slice_145523_comb = p3_add_145227[9:8];
  assign p4_bit_slice_145524_comb = p3_add_145228[9:8];
  assign p4_bit_slice_145555_comb = p3_add_145229[9:8];
  assign p4_bit_slice_145556_comb = p3_add_145230[9:8];
  assign p4_bit_slice_145557_comb = p3_add_145231[9:8];
  assign p4_bit_slice_145558_comb = p3_add_145232[9:8];
  assign p4_bit_slice_145559_comb = p3_add_145233[9:8];
  assign p4_bit_slice_145560_comb = p3_add_145234[9:8];
  assign p4_add_145461_comb = {{1{p3_clipped__260[8]}}, p3_clipped__260} + 10'h001;
  assign p4_add_145462_comb = {{1{p3_clipped__263[8]}}, p3_clipped__263} + 10'h001;
  assign p4_add_145463_comb = {{1{p3_clipped__264[8]}}, p3_clipped__264} + 10'h001;
  assign p4_add_145464_comb = {{1{p3_clipped__267[8]}}, p3_clipped__267} + 10'h001;
  assign p4_add_145465_comb = {{1{p3_clipped__268[8]}}, p3_clipped__268} + 10'h001;
  assign p4_add_145466_comb = {{1{p3_clipped__271[8]}}, p3_clipped__271} + 10'h001;
  assign p4_add_145467_comb = {{1{p3_clipped__276[8]}}, p3_clipped__276} + 10'h001;
  assign p4_add_145468_comb = {{1{p3_clipped__279[8]}}, p3_clipped__279} + 10'h001;
  assign p4_add_145469_comb = {{1{p3_clipped__280[8]}}, p3_clipped__280} + 10'h001;
  assign p4_add_145470_comb = {{1{p3_clipped__283[8]}}, p3_clipped__283} + 10'h001;
  assign p4_add_145471_comb = {{1{p3_clipped__284[8]}}, p3_clipped__284} + 10'h001;
  assign p4_add_145472_comb = {{1{p3_clipped__287[8]}}, p3_clipped__287} + 10'h001;
  assign p4_add_145479_comb = {{1{p3_clipped__292[8]}}, p3_clipped__292} + 10'h001;
  assign p4_add_145480_comb = {{1{p3_clipped__293[8]}}, p3_clipped__293} + 10'h001;
  assign p4_add_145483_comb = {{1{p3_clipped__294[8]}}, p3_clipped__294} + 10'h001;
  assign p4_add_145484_comb = {{1{p3_clipped__295[8]}}, p3_clipped__295} + 10'h001;
  assign p4_add_145485_comb = {{1{p3_clipped__296[8]}}, p3_clipped__296} + 10'h001;
  assign p4_add_145486_comb = {{1{p3_clipped__297[8]}}, p3_clipped__297} + 10'h001;
  assign p4_add_145487_comb = {{1{p3_clipped__265[8]}}, p3_clipped__265} + 10'h001;
  assign p4_add_145488_comb = {{1{p3_clipped__266[8]}}, p3_clipped__266} + 10'h001;
  assign p4_add_145489_comb = {{1{p3_clipped__298[8]}}, p3_clipped__298} + 10'h001;
  assign p4_add_145490_comb = {{1{p3_clipped__299[8]}}, p3_clipped__299} + 10'h001;
  assign p4_add_145491_comb = {{1{p3_clipped__300[8]}}, p3_clipped__300} + 10'h001;
  assign p4_add_145492_comb = {{1{p3_clipped__301[8]}}, p3_clipped__301} + 10'h001;
  assign p4_add_145495_comb = {{1{p3_clipped__302[8]}}, p3_clipped__302} + 10'h001;
  assign p4_add_145496_comb = {{1{p3_clipped__303[8]}}, p3_clipped__303} + 10'h001;
  assign p4_add_145497_comb = {{1{p3_clipped__308[8]}}, p3_clipped__308} + 10'h001;
  assign p4_add_145498_comb = {{1{p3_clipped__309[8]}}, p3_clipped__309} + 10'h001;
  assign p4_add_145501_comb = {{1{p3_clipped__310[8]}}, p3_clipped__310} + 10'h001;
  assign p4_add_145502_comb = {{1{p3_clipped__311[8]}}, p3_clipped__311} + 10'h001;
  assign p4_add_145503_comb = {{1{p3_clipped__312[8]}}, p3_clipped__312} + 10'h001;
  assign p4_add_145504_comb = {{1{p3_clipped__313[8]}}, p3_clipped__313} + 10'h001;
  assign p4_add_145505_comb = {{1{p3_clipped__281[8]}}, p3_clipped__281} + 10'h001;
  assign p4_add_145506_comb = {{1{p3_clipped__282[8]}}, p3_clipped__282} + 10'h001;
  assign p4_add_145507_comb = {{1{p3_clipped__314[8]}}, p3_clipped__314} + 10'h001;
  assign p4_add_145508_comb = {{1{p3_clipped__315[8]}}, p3_clipped__315} + 10'h001;
  assign p4_add_145509_comb = {{1{p3_clipped__316[8]}}, p3_clipped__316} + 10'h001;
  assign p4_add_145510_comb = {{1{p3_clipped__317[8]}}, p3_clipped__317} + 10'h001;
  assign p4_add_145513_comb = {{1{p3_clipped__318[8]}}, p3_clipped__318} + 10'h001;
  assign p4_add_145514_comb = {{1{p3_clipped__319[8]}}, p3_clipped__319} + 10'h001;
  assign p4_bit_slice_145515_comb = p4_add_145459_comb[9:8];
  assign p4_bit_slice_145516_comb = p4_add_145460_comb[9:8];
  assign p4_bit_slice_145531_comb = p4_add_145473_comb[9:8];
  assign p4_bit_slice_145532_comb = p4_add_145474_comb[9:8];
  assign p4_bit_slice_145533_comb = p4_add_145475_comb[9:8];
  assign p4_bit_slice_145534_comb = p4_add_145476_comb[9:8];
  assign p4_bit_slice_145535_comb = p4_add_145477_comb[9:8];
  assign p4_bit_slice_145536_comb = p4_add_145478_comb[9:8];
  assign p4_bit_slice_145539_comb = p4_add_145481_comb[9:8];
  assign p4_bit_slice_145540_comb = p4_add_145482_comb[9:8];
  assign p4_bit_slice_145551_comb = p4_add_145493_comb[9:8];
  assign p4_bit_slice_145552_comb = p4_add_145494_comb[9:8];
  assign p4_bit_slice_145563_comb = p4_add_145499_comb[9:8];
  assign p4_bit_slice_145564_comb = p4_add_145500_comb[9:8];
  assign p4_bit_slice_145575_comb = p4_add_145511_comb[9:8];
  assign p4_bit_slice_145576_comb = p4_add_145512_comb[9:8];
  assign p4_bit_slice_145517_comb = p4_add_145461_comb[9:8];
  assign p4_bit_slice_145518_comb = p4_add_145462_comb[9:8];
  assign p4_bit_slice_145519_comb = p4_add_145463_comb[9:8];
  assign p4_bit_slice_145520_comb = p4_add_145464_comb[9:8];
  assign p4_bit_slice_145521_comb = p4_add_145465_comb[9:8];
  assign p4_bit_slice_145522_comb = p4_add_145466_comb[9:8];
  assign p4_bit_slice_145525_comb = p4_add_145467_comb[9:8];
  assign p4_bit_slice_145526_comb = p4_add_145468_comb[9:8];
  assign p4_bit_slice_145527_comb = p4_add_145469_comb[9:8];
  assign p4_bit_slice_145528_comb = p4_add_145470_comb[9:8];
  assign p4_bit_slice_145529_comb = p4_add_145471_comb[9:8];
  assign p4_bit_slice_145530_comb = p4_add_145472_comb[9:8];
  assign p4_bit_slice_145537_comb = p4_add_145479_comb[9:8];
  assign p4_bit_slice_145538_comb = p4_add_145480_comb[9:8];
  assign p4_bit_slice_145541_comb = p4_add_145483_comb[9:8];
  assign p4_bit_slice_145542_comb = p4_add_145484_comb[9:8];
  assign p4_bit_slice_145543_comb = p4_add_145485_comb[9:8];
  assign p4_bit_slice_145544_comb = p4_add_145486_comb[9:8];
  assign p4_bit_slice_145545_comb = p4_add_145487_comb[9:8];
  assign p4_bit_slice_145546_comb = p4_add_145488_comb[9:8];
  assign p4_bit_slice_145547_comb = p4_add_145489_comb[9:8];
  assign p4_bit_slice_145548_comb = p4_add_145490_comb[9:8];
  assign p4_bit_slice_145549_comb = p4_add_145491_comb[9:8];
  assign p4_bit_slice_145550_comb = p4_add_145492_comb[9:8];
  assign p4_bit_slice_145553_comb = p4_add_145495_comb[9:8];
  assign p4_bit_slice_145554_comb = p4_add_145496_comb[9:8];
  assign p4_bit_slice_145561_comb = p4_add_145497_comb[9:8];
  assign p4_bit_slice_145562_comb = p4_add_145498_comb[9:8];
  assign p4_bit_slice_145565_comb = p4_add_145501_comb[9:8];
  assign p4_bit_slice_145566_comb = p4_add_145502_comb[9:8];
  assign p4_bit_slice_145567_comb = p4_add_145503_comb[9:8];
  assign p4_bit_slice_145568_comb = p4_add_145504_comb[9:8];
  assign p4_bit_slice_145569_comb = p4_add_145505_comb[9:8];
  assign p4_bit_slice_145570_comb = p4_add_145506_comb[9:8];
  assign p4_bit_slice_145571_comb = p4_add_145507_comb[9:8];
  assign p4_bit_slice_145572_comb = p4_add_145508_comb[9:8];
  assign p4_bit_slice_145573_comb = p4_add_145509_comb[9:8];
  assign p4_bit_slice_145574_comb = p4_add_145510_comb[9:8];
  assign p4_bit_slice_145577_comb = p4_add_145513_comb[9:8];
  assign p4_bit_slice_145578_comb = p4_add_145514_comb[9:8];
  assign p4_add_145715_comb = {{1{p4_bit_slice_145523_comb[1]}}, p4_bit_slice_145523_comb} + 3'h1;
  assign p4_add_145716_comb = {{1{p4_bit_slice_145524_comb[1]}}, p4_bit_slice_145524_comb} + 3'h1;
  assign p4_add_145747_comb = {{1{p4_bit_slice_145555_comb[1]}}, p4_bit_slice_145555_comb} + 3'h1;
  assign p4_add_145748_comb = {{1{p4_bit_slice_145556_comb[1]}}, p4_bit_slice_145556_comb} + 3'h1;
  assign p4_add_145749_comb = {{1{p4_bit_slice_145557_comb[1]}}, p4_bit_slice_145557_comb} + 3'h1;
  assign p4_add_145750_comb = {{1{p4_bit_slice_145558_comb[1]}}, p4_bit_slice_145558_comb} + 3'h1;
  assign p4_add_145751_comb = {{1{p4_bit_slice_145559_comb[1]}}, p4_bit_slice_145559_comb} + 3'h1;
  assign p4_add_145752_comb = {{1{p4_bit_slice_145560_comb[1]}}, p4_bit_slice_145560_comb} + 3'h1;
  assign p4_add_145707_comb = {{1{p4_bit_slice_145515_comb[1]}}, p4_bit_slice_145515_comb} + 3'h1;
  assign p4_add_145708_comb = {{1{p4_bit_slice_145516_comb[1]}}, p4_bit_slice_145516_comb} + 3'h1;
  assign p4_add_145723_comb = {{1{p4_bit_slice_145531_comb[1]}}, p4_bit_slice_145531_comb} + 3'h1;
  assign p4_add_145724_comb = {{1{p4_bit_slice_145532_comb[1]}}, p4_bit_slice_145532_comb} + 3'h1;
  assign p4_add_145725_comb = {{1{p4_bit_slice_145533_comb[1]}}, p4_bit_slice_145533_comb} + 3'h1;
  assign p4_add_145726_comb = {{1{p4_bit_slice_145534_comb[1]}}, p4_bit_slice_145534_comb} + 3'h1;
  assign p4_add_145727_comb = {{1{p4_bit_slice_145535_comb[1]}}, p4_bit_slice_145535_comb} + 3'h1;
  assign p4_add_145728_comb = {{1{p4_bit_slice_145536_comb[1]}}, p4_bit_slice_145536_comb} + 3'h1;
  assign p4_add_145731_comb = {{1{p4_bit_slice_145539_comb[1]}}, p4_bit_slice_145539_comb} + 3'h1;
  assign p4_add_145732_comb = {{1{p4_bit_slice_145540_comb[1]}}, p4_bit_slice_145540_comb} + 3'h1;
  assign p4_add_145743_comb = {{1{p4_bit_slice_145551_comb[1]}}, p4_bit_slice_145551_comb} + 3'h1;
  assign p4_add_145744_comb = {{1{p4_bit_slice_145552_comb[1]}}, p4_bit_slice_145552_comb} + 3'h1;
  assign p4_add_145755_comb = {{1{p4_bit_slice_145563_comb[1]}}, p4_bit_slice_145563_comb} + 3'h1;
  assign p4_add_145756_comb = {{1{p4_bit_slice_145564_comb[1]}}, p4_bit_slice_145564_comb} + 3'h1;
  assign p4_add_145767_comb = {{1{p4_bit_slice_145575_comb[1]}}, p4_bit_slice_145575_comb} + 3'h1;
  assign p4_add_145768_comb = {{1{p4_bit_slice_145576_comb[1]}}, p4_bit_slice_145576_comb} + 3'h1;
  assign p4_add_145709_comb = {{1{p4_bit_slice_145517_comb[1]}}, p4_bit_slice_145517_comb} + 3'h1;
  assign p4_add_145710_comb = {{1{p4_bit_slice_145518_comb[1]}}, p4_bit_slice_145518_comb} + 3'h1;
  assign p4_add_145711_comb = {{1{p4_bit_slice_145519_comb[1]}}, p4_bit_slice_145519_comb} + 3'h1;
  assign p4_add_145712_comb = {{1{p4_bit_slice_145520_comb[1]}}, p4_bit_slice_145520_comb} + 3'h1;
  assign p4_add_145713_comb = {{1{p4_bit_slice_145521_comb[1]}}, p4_bit_slice_145521_comb} + 3'h1;
  assign p4_add_145714_comb = {{1{p4_bit_slice_145522_comb[1]}}, p4_bit_slice_145522_comb} + 3'h1;
  assign p4_add_145717_comb = {{1{p4_bit_slice_145525_comb[1]}}, p4_bit_slice_145525_comb} + 3'h1;
  assign p4_add_145718_comb = {{1{p4_bit_slice_145526_comb[1]}}, p4_bit_slice_145526_comb} + 3'h1;
  assign p4_add_145719_comb = {{1{p4_bit_slice_145527_comb[1]}}, p4_bit_slice_145527_comb} + 3'h1;
  assign p4_add_145720_comb = {{1{p4_bit_slice_145528_comb[1]}}, p4_bit_slice_145528_comb} + 3'h1;
  assign p4_add_145721_comb = {{1{p4_bit_slice_145529_comb[1]}}, p4_bit_slice_145529_comb} + 3'h1;
  assign p4_add_145722_comb = {{1{p4_bit_slice_145530_comb[1]}}, p4_bit_slice_145530_comb} + 3'h1;
  assign p4_add_145729_comb = {{1{p4_bit_slice_145537_comb[1]}}, p4_bit_slice_145537_comb} + 3'h1;
  assign p4_add_145730_comb = {{1{p4_bit_slice_145538_comb[1]}}, p4_bit_slice_145538_comb} + 3'h1;
  assign p4_add_145733_comb = {{1{p4_bit_slice_145541_comb[1]}}, p4_bit_slice_145541_comb} + 3'h1;
  assign p4_add_145734_comb = {{1{p4_bit_slice_145542_comb[1]}}, p4_bit_slice_145542_comb} + 3'h1;
  assign p4_add_145735_comb = {{1{p4_bit_slice_145543_comb[1]}}, p4_bit_slice_145543_comb} + 3'h1;
  assign p4_add_145736_comb = {{1{p4_bit_slice_145544_comb[1]}}, p4_bit_slice_145544_comb} + 3'h1;
  assign p4_add_145737_comb = {{1{p4_bit_slice_145545_comb[1]}}, p4_bit_slice_145545_comb} + 3'h1;
  assign p4_add_145738_comb = {{1{p4_bit_slice_145546_comb[1]}}, p4_bit_slice_145546_comb} + 3'h1;
  assign p4_add_145739_comb = {{1{p4_bit_slice_145547_comb[1]}}, p4_bit_slice_145547_comb} + 3'h1;
  assign p4_add_145740_comb = {{1{p4_bit_slice_145548_comb[1]}}, p4_bit_slice_145548_comb} + 3'h1;
  assign p4_add_145741_comb = {{1{p4_bit_slice_145549_comb[1]}}, p4_bit_slice_145549_comb} + 3'h1;
  assign p4_add_145742_comb = {{1{p4_bit_slice_145550_comb[1]}}, p4_bit_slice_145550_comb} + 3'h1;
  assign p4_add_145745_comb = {{1{p4_bit_slice_145553_comb[1]}}, p4_bit_slice_145553_comb} + 3'h1;
  assign p4_add_145746_comb = {{1{p4_bit_slice_145554_comb[1]}}, p4_bit_slice_145554_comb} + 3'h1;
  assign p4_add_145753_comb = {{1{p4_bit_slice_145561_comb[1]}}, p4_bit_slice_145561_comb} + 3'h1;
  assign p4_add_145754_comb = {{1{p4_bit_slice_145562_comb[1]}}, p4_bit_slice_145562_comb} + 3'h1;
  assign p4_add_145757_comb = {{1{p4_bit_slice_145565_comb[1]}}, p4_bit_slice_145565_comb} + 3'h1;
  assign p4_add_145758_comb = {{1{p4_bit_slice_145566_comb[1]}}, p4_bit_slice_145566_comb} + 3'h1;
  assign p4_add_145759_comb = {{1{p4_bit_slice_145567_comb[1]}}, p4_bit_slice_145567_comb} + 3'h1;
  assign p4_add_145760_comb = {{1{p4_bit_slice_145568_comb[1]}}, p4_bit_slice_145568_comb} + 3'h1;
  assign p4_add_145761_comb = {{1{p4_bit_slice_145569_comb[1]}}, p4_bit_slice_145569_comb} + 3'h1;
  assign p4_add_145762_comb = {{1{p4_bit_slice_145570_comb[1]}}, p4_bit_slice_145570_comb} + 3'h1;
  assign p4_add_145763_comb = {{1{p4_bit_slice_145571_comb[1]}}, p4_bit_slice_145571_comb} + 3'h1;
  assign p4_add_145764_comb = {{1{p4_bit_slice_145572_comb[1]}}, p4_bit_slice_145572_comb} + 3'h1;
  assign p4_add_145765_comb = {{1{p4_bit_slice_145573_comb[1]}}, p4_bit_slice_145573_comb} + 3'h1;
  assign p4_add_145766_comb = {{1{p4_bit_slice_145574_comb[1]}}, p4_bit_slice_145574_comb} + 3'h1;
  assign p4_add_145769_comb = {{1{p4_bit_slice_145577_comb[1]}}, p4_bit_slice_145577_comb} + 3'h1;
  assign p4_add_145770_comb = {{1{p4_bit_slice_145578_comb[1]}}, p4_bit_slice_145578_comb} + 3'h1;
  assign p4_clipped__44_comb = p4_add_145715_comb[1] ? 8'hff : {p4_add_145715_comb[0], p3_add_145227[7:1]};
  assign p4_clipped__92_comb = p4_add_145716_comb[1] ? 8'hff : {p4_add_145716_comb[0], p3_add_145228[7:1]};
  assign p4_clipped__12_comb = p4_add_145747_comb[1] ? 8'hff : {p4_add_145747_comb[0], p3_add_145229[7:1]};
  assign p4_clipped__28_comb = p4_add_145748_comb[1] ? 8'hff : {p4_add_145748_comb[0], p3_add_145230[7:1]};
  assign p4_clipped__60_comb = p4_add_145749_comb[1] ? 8'hff : {p4_add_145749_comb[0], p3_add_145231[7:1]};
  assign p4_clipped__76_comb = p4_add_145750_comb[1] ? 8'hff : {p4_add_145750_comb[0], p3_add_145232[7:1]};
  assign p4_clipped__108_comb = p4_add_145751_comb[1] ? 8'hff : {p4_add_145751_comb[0], p3_add_145233[7:1]};
  assign p4_clipped__124_comb = p4_add_145752_comb[1] ? 8'hff : {p4_add_145752_comb[0], p3_add_145234[7:1]};
  assign p4_clipped__40_comb = p4_add_145707_comb[1] ? 8'hff : {p4_add_145707_comb[0], p4_add_145459_comb[7:1]};
  assign p4_clipped__88_comb = p4_add_145708_comb[1] ? 8'hff : {p4_add_145708_comb[0], p4_add_145460_comb[7:1]};
  assign p4_clipped__8_comb = p4_add_145723_comb[1] ? 8'hff : {p4_add_145723_comb[0], p4_add_145473_comb[7:1]};
  assign p4_clipped__24_comb = p4_add_145724_comb[1] ? 8'hff : {p4_add_145724_comb[0], p4_add_145474_comb[7:1]};
  assign p4_clipped__56_comb = p4_add_145725_comb[1] ? 8'hff : {p4_add_145725_comb[0], p4_add_145475_comb[7:1]};
  assign p4_clipped__72_comb = p4_add_145726_comb[1] ? 8'hff : {p4_add_145726_comb[0], p4_add_145476_comb[7:1]};
  assign p4_clipped__104_comb = p4_add_145727_comb[1] ? 8'hff : {p4_add_145727_comb[0], p4_add_145477_comb[7:1]};
  assign p4_clipped__120_comb = p4_add_145728_comb[1] ? 8'hff : {p4_add_145728_comb[0], p4_add_145478_comb[7:1]};
  assign p4_clipped__57_comb = p4_add_145731_comb[1] ? 8'hff : {p4_add_145731_comb[0], p4_add_145481_comb[7:1]};
  assign p4_clipped__73_comb = p4_add_145732_comb[1] ? 8'hff : {p4_add_145732_comb[0], p4_add_145482_comb[7:1]};
  assign p4_clipped__59_comb = p4_add_145743_comb[1] ? 8'hff : {p4_add_145743_comb[0], p4_add_145493_comb[7:1]};
  assign p4_clipped__75_comb = p4_add_145744_comb[1] ? 8'hff : {p4_add_145744_comb[0], p4_add_145494_comb[7:1]};
  assign p4_clipped__61_comb = p4_add_145755_comb[1] ? 8'hff : {p4_add_145755_comb[0], p4_add_145499_comb[7:1]};
  assign p4_clipped__77_comb = p4_add_145756_comb[1] ? 8'hff : {p4_add_145756_comb[0], p4_add_145500_comb[7:1]};
  assign p4_clipped__63_comb = p4_add_145767_comb[1] ? 8'hff : {p4_add_145767_comb[0], p4_add_145511_comb[7:1]};
  assign p4_clipped__79_comb = p4_add_145768_comb[1] ? 8'hff : {p4_add_145768_comb[0], p4_add_145512_comb[7:1]};
  assign p4_clipped__41_comb = p4_add_145709_comb[1] ? 8'hff : {p4_add_145709_comb[0], p4_add_145461_comb[7:1]};
  assign p4_clipped__89_comb = p4_add_145710_comb[1] ? 8'hff : {p4_add_145710_comb[0], p4_add_145462_comb[7:1]};
  assign p4_clipped__42_comb = p4_add_145711_comb[1] ? 8'hff : {p4_add_145711_comb[0], p4_add_145463_comb[7:1]};
  assign p4_clipped__90_comb = p4_add_145712_comb[1] ? 8'hff : {p4_add_145712_comb[0], p4_add_145464_comb[7:1]};
  assign p4_clipped__43_comb = p4_add_145713_comb[1] ? 8'hff : {p4_add_145713_comb[0], p4_add_145465_comb[7:1]};
  assign p4_clipped__91_comb = p4_add_145714_comb[1] ? 8'hff : {p4_add_145714_comb[0], p4_add_145466_comb[7:1]};
  assign p4_clipped__45_comb = p4_add_145717_comb[1] ? 8'hff : {p4_add_145717_comb[0], p4_add_145467_comb[7:1]};
  assign p4_clipped__93_comb = p4_add_145718_comb[1] ? 8'hff : {p4_add_145718_comb[0], p4_add_145468_comb[7:1]};
  assign p4_clipped__46_comb = p4_add_145719_comb[1] ? 8'hff : {p4_add_145719_comb[0], p4_add_145469_comb[7:1]};
  assign p4_clipped__94_comb = p4_add_145720_comb[1] ? 8'hff : {p4_add_145720_comb[0], p4_add_145470_comb[7:1]};
  assign p4_clipped__47_comb = p4_add_145721_comb[1] ? 8'hff : {p4_add_145721_comb[0], p4_add_145471_comb[7:1]};
  assign p4_clipped__95_comb = p4_add_145722_comb[1] ? 8'hff : {p4_add_145722_comb[0], p4_add_145472_comb[7:1]};
  assign p4_clipped__9_comb = p4_add_145729_comb[1] ? 8'hff : {p4_add_145729_comb[0], p4_add_145479_comb[7:1]};
  assign p4_clipped__25_comb = p4_add_145730_comb[1] ? 8'hff : {p4_add_145730_comb[0], p4_add_145480_comb[7:1]};
  assign p4_clipped__105_comb = p4_add_145733_comb[1] ? 8'hff : {p4_add_145733_comb[0], p4_add_145483_comb[7:1]};
  assign p4_clipped__121_comb = p4_add_145734_comb[1] ? 8'hff : {p4_add_145734_comb[0], p4_add_145484_comb[7:1]};
  assign p4_clipped__10_comb = p4_add_145735_comb[1] ? 8'hff : {p4_add_145735_comb[0], p4_add_145485_comb[7:1]};
  assign p4_clipped__26_comb = p4_add_145736_comb[1] ? 8'hff : {p4_add_145736_comb[0], p4_add_145486_comb[7:1]};
  assign p4_clipped__58_comb = p4_add_145737_comb[1] ? 8'hff : {p4_add_145737_comb[0], p4_add_145487_comb[7:1]};
  assign p4_clipped__74_comb = p4_add_145738_comb[1] ? 8'hff : {p4_add_145738_comb[0], p4_add_145488_comb[7:1]};
  assign p4_clipped__106_comb = p4_add_145739_comb[1] ? 8'hff : {p4_add_145739_comb[0], p4_add_145489_comb[7:1]};
  assign p4_clipped__122_comb = p4_add_145740_comb[1] ? 8'hff : {p4_add_145740_comb[0], p4_add_145490_comb[7:1]};
  assign p4_clipped__11_comb = p4_add_145741_comb[1] ? 8'hff : {p4_add_145741_comb[0], p4_add_145491_comb[7:1]};
  assign p4_clipped__27_comb = p4_add_145742_comb[1] ? 8'hff : {p4_add_145742_comb[0], p4_add_145492_comb[7:1]};
  assign p4_clipped__107_comb = p4_add_145745_comb[1] ? 8'hff : {p4_add_145745_comb[0], p4_add_145495_comb[7:1]};
  assign p4_clipped__123_comb = p4_add_145746_comb[1] ? 8'hff : {p4_add_145746_comb[0], p4_add_145496_comb[7:1]};
  assign p4_clipped__13_comb = p4_add_145753_comb[1] ? 8'hff : {p4_add_145753_comb[0], p4_add_145497_comb[7:1]};
  assign p4_clipped__29_comb = p4_add_145754_comb[1] ? 8'hff : {p4_add_145754_comb[0], p4_add_145498_comb[7:1]};
  assign p4_clipped__109_comb = p4_add_145757_comb[1] ? 8'hff : {p4_add_145757_comb[0], p4_add_145501_comb[7:1]};
  assign p4_clipped__125_comb = p4_add_145758_comb[1] ? 8'hff : {p4_add_145758_comb[0], p4_add_145502_comb[7:1]};
  assign p4_clipped__14_comb = p4_add_145759_comb[1] ? 8'hff : {p4_add_145759_comb[0], p4_add_145503_comb[7:1]};
  assign p4_clipped__30_comb = p4_add_145760_comb[1] ? 8'hff : {p4_add_145760_comb[0], p4_add_145504_comb[7:1]};
  assign p4_clipped__62_comb = p4_add_145761_comb[1] ? 8'hff : {p4_add_145761_comb[0], p4_add_145505_comb[7:1]};
  assign p4_clipped__78_comb = p4_add_145762_comb[1] ? 8'hff : {p4_add_145762_comb[0], p4_add_145506_comb[7:1]};
  assign p4_clipped__110_comb = p4_add_145763_comb[1] ? 8'hff : {p4_add_145763_comb[0], p4_add_145507_comb[7:1]};
  assign p4_clipped__126_comb = p4_add_145764_comb[1] ? 8'hff : {p4_add_145764_comb[0], p4_add_145508_comb[7:1]};
  assign p4_clipped__15_comb = p4_add_145765_comb[1] ? 8'hff : {p4_add_145765_comb[0], p4_add_145509_comb[7:1]};
  assign p4_clipped__31_comb = p4_add_145766_comb[1] ? 8'hff : {p4_add_145766_comb[0], p4_add_145510_comb[7:1]};
  assign p4_clipped__111_comb = p4_add_145769_comb[1] ? 8'hff : {p4_add_145769_comb[0], p4_add_145513_comb[7:1]};
  assign p4_clipped__127_comb = p4_add_145770_comb[1] ? 8'hff : {p4_add_145770_comb[0], p4_add_145514_comb[7:1]};
  assign p4_bit_slice_146155_comb = p4_clipped__40_comb[7];
  assign p4_bit_slice_146156_comb = p4_clipped__88_comb[7];
  assign p4_bit_slice_146159_comb = p4_clipped__8_comb[7];
  assign p4_bit_slice_146160_comb = p4_clipped__24_comb[7];
  assign p4_bit_slice_146161_comb = p4_clipped__56_comb[7];
  assign p4_bit_slice_146162_comb = p4_clipped__72_comb[7];
  assign p4_bit_slice_146163_comb = p4_clipped__104_comb[7];
  assign p4_bit_slice_146164_comb = p4_clipped__120_comb[7];
  assign p4_bit_slice_146165_comb = p4_clipped__57_comb[7];
  assign p4_bit_slice_146166_comb = p4_clipped__73_comb[7];
  assign p4_bit_slice_146167_comb = p4_clipped__59_comb[7];
  assign p4_bit_slice_146168_comb = p4_clipped__75_comb[7];
  assign p4_bit_slice_146175_comb = p4_clipped__61_comb[7];
  assign p4_bit_slice_146176_comb = p4_clipped__77_comb[7];
  assign p4_bit_slice_146177_comb = p4_clipped__63_comb[7];
  assign p4_bit_slice_146178_comb = p4_clipped__79_comb[7];
  assign p4_bit_slice_146179_comb = p4_clipped__40_comb[6:0];
  assign p4_bit_slice_146180_comb = p4_clipped__88_comb[6:0];
  assign p4_not_146181_comb = ~p4_clipped__44_comb[7];
  assign p4_bit_slice_146182_comb = p4_clipped__44_comb[6:0];
  assign p4_not_146183_comb = ~p4_clipped__92_comb[7];
  assign p4_bit_slice_146184_comb = p4_clipped__92_comb[6:0];
  assign p4_bit_slice_146185_comb = p4_clipped__8_comb[6:0];
  assign p4_bit_slice_146186_comb = p4_clipped__24_comb[6:0];
  assign p4_bit_slice_146187_comb = p4_clipped__56_comb[6:0];
  assign p4_bit_slice_146188_comb = p4_clipped__72_comb[6:0];
  assign p4_bit_slice_146189_comb = p4_clipped__104_comb[6:0];
  assign p4_bit_slice_146190_comb = p4_clipped__120_comb[6:0];
  assign p4_bit_slice_146191_comb = p4_clipped__57_comb[6:0];
  assign p4_bit_slice_146192_comb = p4_clipped__73_comb[6:0];
  assign p4_bit_slice_146193_comb = p4_clipped__59_comb[6:0];
  assign p4_bit_slice_146194_comb = p4_clipped__75_comb[6:0];
  assign p4_not_146195_comb = ~p4_clipped__12_comb[7];
  assign p4_bit_slice_146196_comb = p4_clipped__12_comb[6:0];
  assign p4_not_146197_comb = ~p4_clipped__28_comb[7];
  assign p4_bit_slice_146198_comb = p4_clipped__28_comb[6:0];
  assign p4_not_146199_comb = ~p4_clipped__60_comb[7];
  assign p4_bit_slice_146200_comb = p4_clipped__60_comb[6:0];
  assign p4_not_146201_comb = ~p4_clipped__76_comb[7];
  assign p4_bit_slice_146202_comb = p4_clipped__76_comb[6:0];
  assign p4_not_146203_comb = ~p4_clipped__108_comb[7];
  assign p4_bit_slice_146204_comb = p4_clipped__108_comb[6:0];
  assign p4_not_146205_comb = ~p4_clipped__124_comb[7];
  assign p4_bit_slice_146206_comb = p4_clipped__124_comb[6:0];
  assign p4_bit_slice_146207_comb = p4_clipped__61_comb[6:0];
  assign p4_bit_slice_146208_comb = p4_clipped__77_comb[6:0];
  assign p4_bit_slice_146209_comb = p4_clipped__63_comb[6:0];
  assign p4_bit_slice_146210_comb = p4_clipped__79_comb[6:0];

  // Registers for pipe stage 4:
  reg [7:0] p4_clipped__41;
  reg [7:0] p4_clipped__89;
  reg [7:0] p4_clipped__42;
  reg [7:0] p4_clipped__90;
  reg [7:0] p4_clipped__43;
  reg [7:0] p4_clipped__91;
  reg [7:0] p4_clipped__45;
  reg [7:0] p4_clipped__93;
  reg [7:0] p4_clipped__46;
  reg [7:0] p4_clipped__94;
  reg [7:0] p4_clipped__47;
  reg [7:0] p4_clipped__95;
  reg [7:0] p4_clipped__9;
  reg [7:0] p4_clipped__25;
  reg [7:0] p4_clipped__105;
  reg [7:0] p4_clipped__121;
  reg [7:0] p4_clipped__10;
  reg [7:0] p4_clipped__26;
  reg [7:0] p4_clipped__58;
  reg [7:0] p4_clipped__74;
  reg [7:0] p4_clipped__106;
  reg [7:0] p4_clipped__122;
  reg [7:0] p4_clipped__11;
  reg [7:0] p4_clipped__27;
  reg [7:0] p4_clipped__107;
  reg [7:0] p4_clipped__123;
  reg [7:0] p4_clipped__13;
  reg [7:0] p4_clipped__29;
  reg [7:0] p4_clipped__109;
  reg [7:0] p4_clipped__125;
  reg [7:0] p4_clipped__14;
  reg [7:0] p4_clipped__30;
  reg [7:0] p4_clipped__62;
  reg [7:0] p4_clipped__78;
  reg [7:0] p4_clipped__110;
  reg [7:0] p4_clipped__126;
  reg [7:0] p4_clipped__15;
  reg [7:0] p4_clipped__31;
  reg [7:0] p4_clipped__111;
  reg [7:0] p4_clipped__127;
  reg p4_bit_slice_146155;
  reg p4_bit_slice_146156;
  reg p4_bit_slice_146159;
  reg p4_bit_slice_146160;
  reg p4_bit_slice_146161;
  reg p4_bit_slice_146162;
  reg p4_bit_slice_146163;
  reg p4_bit_slice_146164;
  reg p4_bit_slice_146165;
  reg p4_bit_slice_146166;
  reg p4_bit_slice_146167;
  reg p4_bit_slice_146168;
  reg p4_bit_slice_146175;
  reg p4_bit_slice_146176;
  reg p4_bit_slice_146177;
  reg p4_bit_slice_146178;
  reg [6:0] p4_bit_slice_146179;
  reg [6:0] p4_bit_slice_146180;
  reg p4_not_146181;
  reg [6:0] p4_bit_slice_146182;
  reg p4_not_146183;
  reg [6:0] p4_bit_slice_146184;
  reg [6:0] p4_bit_slice_146185;
  reg [6:0] p4_bit_slice_146186;
  reg [6:0] p4_bit_slice_146187;
  reg [6:0] p4_bit_slice_146188;
  reg [6:0] p4_bit_slice_146189;
  reg [6:0] p4_bit_slice_146190;
  reg [6:0] p4_bit_slice_146191;
  reg [6:0] p4_bit_slice_146192;
  reg [6:0] p4_bit_slice_146193;
  reg [6:0] p4_bit_slice_146194;
  reg p4_not_146195;
  reg [6:0] p4_bit_slice_146196;
  reg p4_not_146197;
  reg [6:0] p4_bit_slice_146198;
  reg p4_not_146199;
  reg [6:0] p4_bit_slice_146200;
  reg p4_not_146201;
  reg [6:0] p4_bit_slice_146202;
  reg p4_not_146203;
  reg [6:0] p4_bit_slice_146204;
  reg p4_not_146205;
  reg [6:0] p4_bit_slice_146206;
  reg [6:0] p4_bit_slice_146207;
  reg [6:0] p4_bit_slice_146208;
  reg [6:0] p4_bit_slice_146209;
  reg [6:0] p4_bit_slice_146210;
  always @ (posedge clk) begin
    p4_clipped__41 <= p4_clipped__41_comb;
    p4_clipped__89 <= p4_clipped__89_comb;
    p4_clipped__42 <= p4_clipped__42_comb;
    p4_clipped__90 <= p4_clipped__90_comb;
    p4_clipped__43 <= p4_clipped__43_comb;
    p4_clipped__91 <= p4_clipped__91_comb;
    p4_clipped__45 <= p4_clipped__45_comb;
    p4_clipped__93 <= p4_clipped__93_comb;
    p4_clipped__46 <= p4_clipped__46_comb;
    p4_clipped__94 <= p4_clipped__94_comb;
    p4_clipped__47 <= p4_clipped__47_comb;
    p4_clipped__95 <= p4_clipped__95_comb;
    p4_clipped__9 <= p4_clipped__9_comb;
    p4_clipped__25 <= p4_clipped__25_comb;
    p4_clipped__105 <= p4_clipped__105_comb;
    p4_clipped__121 <= p4_clipped__121_comb;
    p4_clipped__10 <= p4_clipped__10_comb;
    p4_clipped__26 <= p4_clipped__26_comb;
    p4_clipped__58 <= p4_clipped__58_comb;
    p4_clipped__74 <= p4_clipped__74_comb;
    p4_clipped__106 <= p4_clipped__106_comb;
    p4_clipped__122 <= p4_clipped__122_comb;
    p4_clipped__11 <= p4_clipped__11_comb;
    p4_clipped__27 <= p4_clipped__27_comb;
    p4_clipped__107 <= p4_clipped__107_comb;
    p4_clipped__123 <= p4_clipped__123_comb;
    p4_clipped__13 <= p4_clipped__13_comb;
    p4_clipped__29 <= p4_clipped__29_comb;
    p4_clipped__109 <= p4_clipped__109_comb;
    p4_clipped__125 <= p4_clipped__125_comb;
    p4_clipped__14 <= p4_clipped__14_comb;
    p4_clipped__30 <= p4_clipped__30_comb;
    p4_clipped__62 <= p4_clipped__62_comb;
    p4_clipped__78 <= p4_clipped__78_comb;
    p4_clipped__110 <= p4_clipped__110_comb;
    p4_clipped__126 <= p4_clipped__126_comb;
    p4_clipped__15 <= p4_clipped__15_comb;
    p4_clipped__31 <= p4_clipped__31_comb;
    p4_clipped__111 <= p4_clipped__111_comb;
    p4_clipped__127 <= p4_clipped__127_comb;
    p4_bit_slice_146155 <= p4_bit_slice_146155_comb;
    p4_bit_slice_146156 <= p4_bit_slice_146156_comb;
    p4_bit_slice_146159 <= p4_bit_slice_146159_comb;
    p4_bit_slice_146160 <= p4_bit_slice_146160_comb;
    p4_bit_slice_146161 <= p4_bit_slice_146161_comb;
    p4_bit_slice_146162 <= p4_bit_slice_146162_comb;
    p4_bit_slice_146163 <= p4_bit_slice_146163_comb;
    p4_bit_slice_146164 <= p4_bit_slice_146164_comb;
    p4_bit_slice_146165 <= p4_bit_slice_146165_comb;
    p4_bit_slice_146166 <= p4_bit_slice_146166_comb;
    p4_bit_slice_146167 <= p4_bit_slice_146167_comb;
    p4_bit_slice_146168 <= p4_bit_slice_146168_comb;
    p4_bit_slice_146175 <= p4_bit_slice_146175_comb;
    p4_bit_slice_146176 <= p4_bit_slice_146176_comb;
    p4_bit_slice_146177 <= p4_bit_slice_146177_comb;
    p4_bit_slice_146178 <= p4_bit_slice_146178_comb;
    p4_bit_slice_146179 <= p4_bit_slice_146179_comb;
    p4_bit_slice_146180 <= p4_bit_slice_146180_comb;
    p4_not_146181 <= p4_not_146181_comb;
    p4_bit_slice_146182 <= p4_bit_slice_146182_comb;
    p4_not_146183 <= p4_not_146183_comb;
    p4_bit_slice_146184 <= p4_bit_slice_146184_comb;
    p4_bit_slice_146185 <= p4_bit_slice_146185_comb;
    p4_bit_slice_146186 <= p4_bit_slice_146186_comb;
    p4_bit_slice_146187 <= p4_bit_slice_146187_comb;
    p4_bit_slice_146188 <= p4_bit_slice_146188_comb;
    p4_bit_slice_146189 <= p4_bit_slice_146189_comb;
    p4_bit_slice_146190 <= p4_bit_slice_146190_comb;
    p4_bit_slice_146191 <= p4_bit_slice_146191_comb;
    p4_bit_slice_146192 <= p4_bit_slice_146192_comb;
    p4_bit_slice_146193 <= p4_bit_slice_146193_comb;
    p4_bit_slice_146194 <= p4_bit_slice_146194_comb;
    p4_not_146195 <= p4_not_146195_comb;
    p4_bit_slice_146196 <= p4_bit_slice_146196_comb;
    p4_not_146197 <= p4_not_146197_comb;
    p4_bit_slice_146198 <= p4_bit_slice_146198_comb;
    p4_not_146199 <= p4_not_146199_comb;
    p4_bit_slice_146200 <= p4_bit_slice_146200_comb;
    p4_not_146201 <= p4_not_146201_comb;
    p4_bit_slice_146202 <= p4_bit_slice_146202_comb;
    p4_not_146203 <= p4_not_146203_comb;
    p4_bit_slice_146204 <= p4_bit_slice_146204_comb;
    p4_not_146205 <= p4_not_146205_comb;
    p4_bit_slice_146206 <= p4_bit_slice_146206_comb;
    p4_bit_slice_146207 <= p4_bit_slice_146207_comb;
    p4_bit_slice_146208 <= p4_bit_slice_146208_comb;
    p4_bit_slice_146209 <= p4_bit_slice_146209_comb;
    p4_bit_slice_146210 <= p4_bit_slice_146210_comb;
  end

  // ===== Pipe stage 5:
  wire [7:0] p5_shifted__99_squeezed_comb;
  wire [7:0] p5_shifted__100_squeezed_comb;
  wire [7:0] p5_shifted__97_squeezed_comb;
  wire [7:0] p5_shifted__102_squeezed_comb;
  wire [7:0] p5_shifted__98_squeezed_comb;
  wire [7:0] p5_shifted__101_squeezed_comb;
  wire [7:0] p5_shifted__96_squeezed_comb;
  wire [7:0] p5_shifted__103_squeezed_comb;
  wire [7:0] p5_shifted__66_squeezed_comb;
  wire [7:0] p5_shifted__69_squeezed_comb;
  wire [7:0] p5_shifted__64_squeezed_comb;
  wire [7:0] p5_shifted__65_squeezed_comb;
  wire [7:0] p5_shifted__67_squeezed_comb;
  wire [7:0] p5_shifted__68_squeezed_comb;
  wire [7:0] p5_shifted__70_squeezed_comb;
  wire [7:0] p5_shifted__71_squeezed_comb;
  wire [7:0] p5_shifted__75_squeezed_comb;
  wire [7:0] p5_shifted__76_squeezed_comb;
  wire [7:0] p5_shifted__91_squeezed_comb;
  wire [7:0] p5_shifted__92_squeezed_comb;
  wire [7:0] p5_shifted__107_squeezed_comb;
  wire [7:0] p5_shifted__108_squeezed_comb;
  wire [7:0] p5_shifted__123_squeezed_comb;
  wire [7:0] p5_shifted__124_squeezed_comb;
  wire [13:0] p5_smul_58292_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___209_comb;
  wire [13:0] p5_smul_58294_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___210_comb;
  wire [13:0] p5_smul_58544_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___272_comb;
  wire [13:0] p5_smul_58554_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___275_comb;
  wire [13:0] p5_smul_58802_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___305_comb;
  wire [13:0] p5_smul_58808_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___306_comb;
  wire [13:0] p5_smul_59054_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___368_comb;
  wire [13:0] p5_smul_59068_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___371_comb;
  wire [7:0] p5_shifted__74_squeezed_comb;
  wire [7:0] p5_shifted__77_squeezed_comb;
  wire [7:0] p5_shifted__82_squeezed_comb;
  wire [7:0] p5_shifted__85_squeezed_comb;
  wire [7:0] p5_shifted__90_squeezed_comb;
  wire [7:0] p5_shifted__93_squeezed_comb;
  wire [7:0] p5_shifted__106_squeezed_comb;
  wire [7:0] p5_shifted__109_squeezed_comb;
  wire [7:0] p5_shifted__114_squeezed_comb;
  wire [7:0] p5_shifted__117_squeezed_comb;
  wire [7:0] p5_shifted__122_squeezed_comb;
  wire [7:0] p5_shifted__125_squeezed_comb;
  wire [7:0] p5_shifted__72_squeezed_comb;
  wire [7:0] p5_shifted__73_squeezed_comb;
  wire [7:0] p5_shifted__78_squeezed_comb;
  wire [7:0] p5_shifted__79_squeezed_comb;
  wire [7:0] p5_shifted__80_squeezed_comb;
  wire [7:0] p5_shifted__81_squeezed_comb;
  wire [7:0] p5_shifted__83_squeezed_comb;
  wire [7:0] p5_shifted__84_squeezed_comb;
  wire [7:0] p5_shifted__86_squeezed_comb;
  wire [7:0] p5_shifted__87_squeezed_comb;
  wire [7:0] p5_shifted__88_squeezed_comb;
  wire [7:0] p5_shifted__89_squeezed_comb;
  wire [7:0] p5_shifted__94_squeezed_comb;
  wire [7:0] p5_shifted__95_squeezed_comb;
  wire [7:0] p5_shifted__104_squeezed_comb;
  wire [7:0] p5_shifted__105_squeezed_comb;
  wire [7:0] p5_shifted__110_squeezed_comb;
  wire [7:0] p5_shifted__111_squeezed_comb;
  wire [7:0] p5_shifted__112_squeezed_comb;
  wire [7:0] p5_shifted__113_squeezed_comb;
  wire [7:0] p5_shifted__115_squeezed_comb;
  wire [7:0] p5_shifted__116_squeezed_comb;
  wire [7:0] p5_shifted__118_squeezed_comb;
  wire [7:0] p5_shifted__119_squeezed_comb;
  wire [7:0] p5_shifted__120_squeezed_comb;
  wire [7:0] p5_shifted__121_squeezed_comb;
  wire [7:0] p5_shifted__126_squeezed_comb;
  wire [7:0] p5_shifted__127_squeezed_comb;
  wire [15:0] p5_smul_58226_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___192_comb;
  wire [15:0] p5_smul_58232_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___195_comb;
  wire [15:0] p5_smul_58290_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___208_comb;
  wire [15:0] p5_smul_58296_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___211_comb;
  wire [14:0] p5_smul_58350_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___64_comb;
  wire [14:0] p5_smul_58352_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___224_comb;
  wire [14:0] p5_smul_58354_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___225_comb;
  wire [14:0] p5_smul_58356_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___65_comb;
  wire [14:0] p5_smul_58358_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___66_comb;
  wire [14:0] p5_smul_58360_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___226_comb;
  wire [14:0] p5_smul_58362_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___227_comb;
  wire [14:0] p5_smul_58364_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___67_comb;
  wire [14:0] p5_smul_58372_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___69_comb;
  wire [14:0] p5_smul_58374_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___70_comb;
  wire [14:0] p5_smul_58404_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___77_comb;
  wire [14:0] p5_smul_58406_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___78_comb;
  wire [14:0] p5_smul_58414_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___80_comb;
  wire [14:0] p5_smul_58416_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___240_comb;
  wire [14:0] p5_smul_58418_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___241_comb;
  wire [14:0] p5_smul_58420_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___81_comb;
  wire [14:0] p5_smul_58422_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___82_comb;
  wire [14:0] p5_smul_58424_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___242_comb;
  wire [14:0] p5_smul_58426_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___243_comb;
  wire [14:0] p5_smul_58428_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___83_comb;
  wire [14:0] p5_smul_58436_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___85_comb;
  wire [14:0] p5_smul_58438_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___86_comb;
  wire [14:0] p5_smul_58468_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___93_comb;
  wire [14:0] p5_smul_58470_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___94_comb;
  wire [15:0] p5_smul_58484_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___257_comb;
  wire [15:0] p5_smul_58486_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___258_comb;
  wire [15:0] p5_smul_58500_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___261_comb;
  wire [15:0] p5_smul_58502_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___262_comb;
  wire [15:0] p5_smul_58532_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___269_comb;
  wire [15:0] p5_smul_58534_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___270_comb;
  wire [15:0] p5_smul_58548_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___273_comb;
  wire [15:0] p5_smul_58550_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___274_comb;
  wire [15:0] p5_smul_58564_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___277_comb;
  wire [15:0] p5_smul_58566_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___278_comb;
  wire [15:0] p5_smul_58596_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___285_comb;
  wire [15:0] p5_smul_58598_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___286_comb;
  wire [15:0] p5_smul_58734_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___288_comb;
  wire [15:0] p5_smul_58748_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___291_comb;
  wire [15:0] p5_smul_58798_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___304_comb;
  wire [15:0] p5_smul_58812_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___307_comb;
  wire [14:0] p5_smul_58862_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___320_comb;
  wire [14:0] p5_smul_58864_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___96_comb;
  wire [14:0] p5_smul_58866_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___321_comb;
  wire [14:0] p5_smul_58868_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___97_comb;
  wire [14:0] p5_smul_58870_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___98_comb;
  wire [14:0] p5_smul_58872_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___322_comb;
  wire [14:0] p5_smul_58874_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___99_comb;
  wire [14:0] p5_smul_58876_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___323_comb;
  wire [14:0] p5_smul_58884_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___101_comb;
  wire [14:0] p5_smul_58886_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___102_comb;
  wire [14:0] p5_smul_58916_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___109_comb;
  wire [14:0] p5_smul_58918_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___110_comb;
  wire [14:0] p5_smul_58926_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___336_comb;
  wire [14:0] p5_smul_58928_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___112_comb;
  wire [14:0] p5_smul_58930_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___337_comb;
  wire [14:0] p5_smul_58932_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___113_comb;
  wire [14:0] p5_smul_58934_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___114_comb;
  wire [14:0] p5_smul_58936_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___338_comb;
  wire [14:0] p5_smul_58938_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___115_comb;
  wire [14:0] p5_smul_58940_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___339_comb;
  wire [14:0] p5_smul_58948_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___117_comb;
  wire [14:0] p5_smul_58950_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___118_comb;
  wire [14:0] p5_smul_58980_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___125_comb;
  wire [14:0] p5_smul_58982_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___126_comb;
  wire [15:0] p5_smul_58992_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___353_comb;
  wire [15:0] p5_smul_59002_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___354_comb;
  wire [15:0] p5_smul_59056_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___369_comb;
  wire [15:0] p5_smul_59066_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___370_comb;
  wire [13:0] p5_smul_58228_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___193_comb;
  wire [13:0] p5_smul_58230_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___194_comb;
  wire [13:0] p5_smul_58244_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___197_comb;
  wire [13:0] p5_smul_58246_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___198_comb;
  wire [13:0] p5_smul_58276_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___205_comb;
  wire [13:0] p5_smul_58278_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___206_comb;
  wire [13:0] p5_smul_58308_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___213_comb;
  wire [13:0] p5_smul_58310_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___214_comb;
  wire [13:0] p5_smul_58340_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___221_comb;
  wire [13:0] p5_smul_58342_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___222_comb;
  wire [13:0] p5_smul_58480_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___256_comb;
  wire [13:0] p5_smul_58490_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___259_comb;
  wire [13:0] p5_smul_58738_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___289_comb;
  wire [13:0] p5_smul_58744_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___290_comb;
  wire [13:0] p5_smul_58990_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___352_comb;
  wire [13:0] p5_smul_59004_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___355_comb;
  wire [7:0] p5_smul_57326_TrailingBits___192_comb;
  wire [7:0] p5_smul_57326_TrailingBits___193_comb;
  wire [7:0] p5_smul_57326_TrailingBits___194_comb;
  wire [7:0] p5_smul_57326_TrailingBits___195_comb;
  wire [7:0] p5_smul_57326_TrailingBits___196_comb;
  wire [7:0] p5_smul_57326_TrailingBits___197_comb;
  wire [7:0] p5_smul_57326_TrailingBits___198_comb;
  wire [7:0] p5_smul_57326_TrailingBits___199_comb;
  wire [7:0] p5_smul_57326_TrailingBits___224_comb;
  wire [7:0] p5_smul_57326_TrailingBits___225_comb;
  wire [7:0] p5_smul_57326_TrailingBits___226_comb;
  wire [7:0] p5_smul_57326_TrailingBits___227_comb;
  wire [7:0] p5_smul_57326_TrailingBits___228_comb;
  wire [7:0] p5_smul_57326_TrailingBits___229_comb;
  wire [7:0] p5_smul_57326_TrailingBits___230_comb;
  wire [7:0] p5_smul_57326_TrailingBits___231_comb;
  wire [22:0] p5_concat_147829_comb;
  wire [22:0] p5_concat_147830_comb;
  wire [22:0] p5_concat_147971_comb;
  wire [22:0] p5_concat_147976_comb;
  wire [22:0] p5_concat_148021_comb;
  wire [22:0] p5_concat_148022_comb;
  wire [22:0] p5_concat_148163_comb;
  wire [22:0] p5_concat_148168_comb;
  wire [15:0] p5_smul_58242_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___196_comb;
  wire [15:0] p5_smul_58248_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___199_comb;
  wire [15:0] p5_smul_58258_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___200_comb;
  wire [15:0] p5_smul_58264_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___203_comb;
  wire [15:0] p5_smul_58274_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___204_comb;
  wire [15:0] p5_smul_58280_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___207_comb;
  wire [15:0] p5_smul_58306_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___212_comb;
  wire [15:0] p5_smul_58312_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___215_comb;
  wire [15:0] p5_smul_58322_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___216_comb;
  wire [15:0] p5_smul_58328_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___219_comb;
  wire [15:0] p5_smul_58338_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___220_comb;
  wire [15:0] p5_smul_58344_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___223_comb;
  wire [14:0] p5_smul_58366_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___68_comb;
  wire [14:0] p5_smul_58368_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___228_comb;
  wire [14:0] p5_smul_58370_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___229_comb;
  wire [14:0] p5_smul_58376_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___230_comb;
  wire [14:0] p5_smul_58378_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___231_comb;
  wire [14:0] p5_smul_58380_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___71_comb;
  wire [14:0] p5_smul_58382_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___72_comb;
  wire [14:0] p5_smul_58384_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___232_comb;
  wire [14:0] p5_smul_58386_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___233_comb;
  wire [14:0] p5_smul_58388_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___73_comb;
  wire [14:0] p5_smul_58390_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___74_comb;
  wire [14:0] p5_smul_58392_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___234_comb;
  wire [14:0] p5_smul_58394_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___235_comb;
  wire [14:0] p5_smul_58396_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___75_comb;
  wire [14:0] p5_smul_58398_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___76_comb;
  wire [14:0] p5_smul_58400_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___236_comb;
  wire [14:0] p5_smul_58402_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___237_comb;
  wire [14:0] p5_smul_58408_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___238_comb;
  wire [14:0] p5_smul_58410_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___239_comb;
  wire [14:0] p5_smul_58412_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___79_comb;
  wire [14:0] p5_smul_58430_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___84_comb;
  wire [14:0] p5_smul_58432_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___244_comb;
  wire [14:0] p5_smul_58434_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___245_comb;
  wire [14:0] p5_smul_58440_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___246_comb;
  wire [14:0] p5_smul_58442_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___247_comb;
  wire [14:0] p5_smul_58444_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___87_comb;
  wire [14:0] p5_smul_58446_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___88_comb;
  wire [14:0] p5_smul_58448_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___248_comb;
  wire [14:0] p5_smul_58450_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___249_comb;
  wire [14:0] p5_smul_58452_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___89_comb;
  wire [14:0] p5_smul_58454_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___90_comb;
  wire [14:0] p5_smul_58456_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___250_comb;
  wire [14:0] p5_smul_58458_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___251_comb;
  wire [14:0] p5_smul_58460_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___91_comb;
  wire [14:0] p5_smul_58462_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___92_comb;
  wire [14:0] p5_smul_58464_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___252_comb;
  wire [14:0] p5_smul_58466_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___253_comb;
  wire [14:0] p5_smul_58472_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___254_comb;
  wire [14:0] p5_smul_58474_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___255_comb;
  wire [14:0] p5_smul_58476_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___95_comb;
  wire [15:0] p5_smul_58516_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___265_comb;
  wire [15:0] p5_smul_58518_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___266_comb;
  wire [15:0] p5_smul_58580_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___281_comb;
  wire [15:0] p5_smul_58582_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___282_comb;
  wire [15:0] p5_smul_58750_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___292_comb;
  wire [15:0] p5_smul_58764_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___295_comb;
  wire [15:0] p5_smul_58766_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___296_comb;
  wire [15:0] p5_smul_58780_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___299_comb;
  wire [15:0] p5_smul_58782_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___300_comb;
  wire [15:0] p5_smul_58796_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___303_comb;
  wire [15:0] p5_smul_58814_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___308_comb;
  wire [15:0] p5_smul_58828_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___311_comb;
  wire [15:0] p5_smul_58830_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___312_comb;
  wire [15:0] p5_smul_58844_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___315_comb;
  wire [15:0] p5_smul_58846_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___316_comb;
  wire [15:0] p5_smul_58860_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___319_comb;
  wire [14:0] p5_smul_58878_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___324_comb;
  wire [14:0] p5_smul_58880_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___100_comb;
  wire [14:0] p5_smul_58882_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___325_comb;
  wire [14:0] p5_smul_58888_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___326_comb;
  wire [14:0] p5_smul_58890_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___103_comb;
  wire [14:0] p5_smul_58892_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___327_comb;
  wire [14:0] p5_smul_58894_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___328_comb;
  wire [14:0] p5_smul_58896_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___104_comb;
  wire [14:0] p5_smul_58898_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___329_comb;
  wire [14:0] p5_smul_58900_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___105_comb;
  wire [14:0] p5_smul_58902_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___106_comb;
  wire [14:0] p5_smul_58904_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___330_comb;
  wire [14:0] p5_smul_58906_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___107_comb;
  wire [14:0] p5_smul_58908_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___331_comb;
  wire [14:0] p5_smul_58910_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___332_comb;
  wire [14:0] p5_smul_58912_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___108_comb;
  wire [14:0] p5_smul_58914_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___333_comb;
  wire [14:0] p5_smul_58920_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___334_comb;
  wire [14:0] p5_smul_58922_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___111_comb;
  wire [14:0] p5_smul_58924_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___335_comb;
  wire [14:0] p5_smul_58942_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___340_comb;
  wire [14:0] p5_smul_58944_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___116_comb;
  wire [14:0] p5_smul_58946_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___341_comb;
  wire [14:0] p5_smul_58952_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___342_comb;
  wire [14:0] p5_smul_58954_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___119_comb;
  wire [14:0] p5_smul_58956_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___343_comb;
  wire [14:0] p5_smul_58958_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___344_comb;
  wire [14:0] p5_smul_58960_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___120_comb;
  wire [14:0] p5_smul_58962_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___345_comb;
  wire [14:0] p5_smul_58964_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___121_comb;
  wire [14:0] p5_smul_58966_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___122_comb;
  wire [14:0] p5_smul_58968_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___346_comb;
  wire [14:0] p5_smul_58970_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___123_comb;
  wire [14:0] p5_smul_58972_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___347_comb;
  wire [14:0] p5_smul_58974_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___348_comb;
  wire [14:0] p5_smul_58976_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___124_comb;
  wire [14:0] p5_smul_58978_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___349_comb;
  wire [14:0] p5_smul_58984_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___350_comb;
  wire [14:0] p5_smul_58986_NarrowedMult__comb;
  wire [9:0] p5_smul_57454_TrailingBits___127_comb;
  wire [14:0] p5_smul_58988_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___351_comb;
  wire [15:0] p5_smul_59008_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___357_comb;
  wire [15:0] p5_smul_59018_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___358_comb;
  wire [15:0] p5_smul_59024_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___361_comb;
  wire [15:0] p5_smul_59034_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___362_comb;
  wire [15:0] p5_smul_59040_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___365_comb;
  wire [15:0] p5_smul_59050_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___366_comb;
  wire [15:0] p5_smul_59072_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___373_comb;
  wire [15:0] p5_smul_59082_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___374_comb;
  wire [15:0] p5_smul_59088_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___377_comb;
  wire [15:0] p5_smul_59098_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___378_comb;
  wire [15:0] p5_smul_59104_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___381_comb;
  wire [15:0] p5_smul_59114_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___382_comb;
  wire [24:0] p5_concat_147291_comb;
  wire [24:0] p5_concat_147296_comb;
  wire [24:0] p5_concat_147315_comb;
  wire [24:0] p5_concat_147320_comb;
  wire [24:0] p5_concat_147339_comb;
  wire [23:0] p5_concat_147340_comb;
  wire [23:0] p5_concat_147341_comb;
  wire [24:0] p5_concat_147342_comb;
  wire [24:0] p5_concat_147343_comb;
  wire [23:0] p5_concat_147344_comb;
  wire [23:0] p5_concat_147345_comb;
  wire [24:0] p5_concat_147346_comb;
  wire [24:0] p5_concat_147350_comb;
  wire [24:0] p5_concat_147351_comb;
  wire [24:0] p5_concat_147366_comb;
  wire [24:0] p5_concat_147367_comb;
  wire [24:0] p5_concat_147371_comb;
  wire [23:0] p5_concat_147372_comb;
  wire [23:0] p5_concat_147373_comb;
  wire [24:0] p5_concat_147374_comb;
  wire [24:0] p5_concat_147375_comb;
  wire [23:0] p5_concat_147376_comb;
  wire [23:0] p5_concat_147377_comb;
  wire [24:0] p5_concat_147378_comb;
  wire [24:0] p5_concat_147382_comb;
  wire [24:0] p5_concat_147383_comb;
  wire [24:0] p5_concat_147398_comb;
  wire [24:0] p5_concat_147399_comb;
  wire [24:0] p5_concat_147405_comb;
  wire [24:0] p5_concat_147406_comb;
  wire [24:0] p5_concat_147411_comb;
  wire [24:0] p5_concat_147412_comb;
  wire [24:0] p5_concat_147423_comb;
  wire [24:0] p5_concat_147424_comb;
  wire [24:0] p5_concat_147429_comb;
  wire [24:0] p5_concat_147430_comb;
  wire [24:0] p5_concat_147435_comb;
  wire [24:0] p5_concat_147436_comb;
  wire [24:0] p5_concat_147447_comb;
  wire [24:0] p5_concat_147448_comb;
  wire [24:0] p5_concat_147451_comb;
  wire [24:0] p5_concat_147456_comb;
  wire [24:0] p5_concat_147475_comb;
  wire [24:0] p5_concat_147480_comb;
  wire [23:0] p5_concat_147499_comb;
  wire [24:0] p5_concat_147500_comb;
  wire [23:0] p5_concat_147501_comb;
  wire [24:0] p5_concat_147502_comb;
  wire [24:0] p5_concat_147503_comb;
  wire [23:0] p5_concat_147504_comb;
  wire [24:0] p5_concat_147505_comb;
  wire [23:0] p5_concat_147506_comb;
  wire [24:0] p5_concat_147510_comb;
  wire [24:0] p5_concat_147511_comb;
  wire [24:0] p5_concat_147526_comb;
  wire [24:0] p5_concat_147527_comb;
  wire [23:0] p5_concat_147531_comb;
  wire [24:0] p5_concat_147532_comb;
  wire [23:0] p5_concat_147533_comb;
  wire [24:0] p5_concat_147534_comb;
  wire [24:0] p5_concat_147535_comb;
  wire [23:0] p5_concat_147536_comb;
  wire [24:0] p5_concat_147537_comb;
  wire [23:0] p5_concat_147538_comb;
  wire [24:0] p5_concat_147542_comb;
  wire [24:0] p5_concat_147543_comb;
  wire [24:0] p5_concat_147558_comb;
  wire [24:0] p5_concat_147559_comb;
  wire [24:0] p5_concat_147565_comb;
  wire [24:0] p5_concat_147566_comb;
  wire [24:0] p5_concat_147589_comb;
  wire [24:0] p5_concat_147590_comb;
  wire [22:0] p5_concat_147805_comb;
  wire [22:0] p5_concat_147806_comb;
  wire [22:0] p5_concat_147811_comb;
  wire [22:0] p5_concat_147812_comb;
  wire [22:0] p5_concat_147823_comb;
  wire [22:0] p5_concat_147824_comb;
  wire [22:0] p5_concat_147835_comb;
  wire [22:0] p5_concat_147836_comb;
  wire [22:0] p5_concat_147847_comb;
  wire [22:0] p5_concat_147848_comb;
  wire [22:0] p5_concat_147947_comb;
  wire [22:0] p5_concat_147952_comb;
  wire [22:0] p5_concat_147997_comb;
  wire [22:0] p5_concat_147998_comb;
  wire [22:0] p5_concat_148139_comb;
  wire [22:0] p5_concat_148144_comb;
  wire [15:0] p5_shifted__64_comb;
  wire [7:0] p5_smul_57326_TrailingBits___64_comb;
  wire [15:0] p5_shifted__65_comb;
  wire [7:0] p5_smul_57326_TrailingBits___65_comb;
  wire [15:0] p5_shifted__66_comb;
  wire [7:0] p5_smul_57326_TrailingBits___66_comb;
  wire [15:0] p5_shifted__67_comb;
  wire [7:0] p5_smul_57326_TrailingBits___67_comb;
  wire [15:0] p5_shifted__68_comb;
  wire [7:0] p5_smul_57326_TrailingBits___68_comb;
  wire [15:0] p5_shifted__69_comb;
  wire [7:0] p5_smul_57326_TrailingBits___69_comb;
  wire [15:0] p5_shifted__70_comb;
  wire [7:0] p5_smul_57326_TrailingBits___70_comb;
  wire [15:0] p5_shifted__71_comb;
  wire [7:0] p5_smul_57326_TrailingBits___71_comb;
  wire [15:0] p5_shifted__96_comb;
  wire [7:0] p5_smul_57326_TrailingBits___96_comb;
  wire [15:0] p5_shifted__97_comb;
  wire [7:0] p5_smul_57326_TrailingBits___97_comb;
  wire [15:0] p5_shifted__98_comb;
  wire [7:0] p5_smul_57326_TrailingBits___98_comb;
  wire [15:0] p5_shifted__99_comb;
  wire [7:0] p5_smul_57326_TrailingBits___99_comb;
  wire [15:0] p5_shifted__100_comb;
  wire [7:0] p5_smul_57326_TrailingBits___100_comb;
  wire [15:0] p5_shifted__101_comb;
  wire [7:0] p5_smul_57326_TrailingBits___101_comb;
  wire [15:0] p5_shifted__102_comb;
  wire [7:0] p5_smul_57326_TrailingBits___102_comb;
  wire [15:0] p5_shifted__103_comb;
  wire [7:0] p5_smul_57326_TrailingBits___103_comb;
  wire [31:0] p5_prod__779_comb;
  wire [31:0] p5_prod__784_comb;
  wire [31:0] p5_prod__781_comb;
  wire [31:0] p5_prod__812_comb;
  wire [31:0] p5_prod__801_comb;
  wire [31:0] p5_prod__819_comb;
  wire [31:0] p5_prod__803_comb;
  wire [31:0] p5_prod__831_comb;
  wire [24:0] p5_concat_147297_comb;
  wire [24:0] p5_concat_147302_comb;
  wire [24:0] p5_concat_147303_comb;
  wire [13:0] p5_smul_58260_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___201_comb;
  wire [13:0] p5_smul_58262_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___202_comb;
  wire [24:0] p5_concat_147308_comb;
  wire [24:0] p5_concat_147309_comb;
  wire [24:0] p5_concat_147314_comb;
  wire [24:0] p5_concat_147321_comb;
  wire [24:0] p5_concat_147326_comb;
  wire [24:0] p5_concat_147327_comb;
  wire [13:0] p5_smul_58324_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___217_comb;
  wire [13:0] p5_smul_58326_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___218_comb;
  wire [24:0] p5_concat_147332_comb;
  wire [24:0] p5_concat_147333_comb;
  wire [24:0] p5_concat_147338_comb;
  wire [24:0] p5_concat_147347_comb;
  wire [23:0] p5_concat_147348_comb;
  wire [23:0] p5_concat_147349_comb;
  wire [23:0] p5_concat_147352_comb;
  wire [23:0] p5_concat_147353_comb;
  wire [24:0] p5_concat_147354_comb;
  wire [24:0] p5_concat_147355_comb;
  wire [23:0] p5_concat_147356_comb;
  wire [23:0] p5_concat_147357_comb;
  wire [24:0] p5_concat_147358_comb;
  wire [24:0] p5_concat_147359_comb;
  wire [23:0] p5_concat_147360_comb;
  wire [23:0] p5_concat_147361_comb;
  wire [24:0] p5_concat_147362_comb;
  wire [24:0] p5_concat_147363_comb;
  wire [23:0] p5_concat_147364_comb;
  wire [23:0] p5_concat_147365_comb;
  wire [23:0] p5_concat_147368_comb;
  wire [23:0] p5_concat_147369_comb;
  wire [24:0] p5_concat_147370_comb;
  wire [24:0] p5_concat_147379_comb;
  wire [23:0] p5_concat_147380_comb;
  wire [23:0] p5_concat_147381_comb;
  wire [23:0] p5_concat_147384_comb;
  wire [23:0] p5_concat_147385_comb;
  wire [24:0] p5_concat_147386_comb;
  wire [24:0] p5_concat_147387_comb;
  wire [23:0] p5_concat_147388_comb;
  wire [23:0] p5_concat_147389_comb;
  wire [24:0] p5_concat_147390_comb;
  wire [24:0] p5_concat_147391_comb;
  wire [23:0] p5_concat_147392_comb;
  wire [23:0] p5_concat_147393_comb;
  wire [24:0] p5_concat_147394_comb;
  wire [24:0] p5_concat_147395_comb;
  wire [23:0] p5_concat_147396_comb;
  wire [23:0] p5_concat_147397_comb;
  wire [23:0] p5_concat_147400_comb;
  wire [23:0] p5_concat_147401_comb;
  wire [24:0] p5_concat_147402_comb;
  wire [13:0] p5_smul_58496_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___260_comb;
  wire [13:0] p5_smul_58506_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___263_comb;
  wire [13:0] p5_smul_58512_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___264_comb;
  wire [24:0] p5_concat_147417_comb;
  wire [24:0] p5_concat_147418_comb;
  wire [13:0] p5_smul_58522_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___267_comb;
  wire [13:0] p5_smul_58528_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___268_comb;
  wire [13:0] p5_smul_58538_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___271_comb;
  wire [13:0] p5_smul_58560_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___276_comb;
  wire [13:0] p5_smul_58570_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___279_comb;
  wire [13:0] p5_smul_58576_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___280_comb;
  wire [24:0] p5_concat_147441_comb;
  wire [24:0] p5_concat_147442_comb;
  wire [13:0] p5_smul_58586_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___283_comb;
  wire [13:0] p5_smul_58592_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___284_comb;
  wire [13:0] p5_smul_58602_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___287_comb;
  wire [24:0] p5_concat_147457_comb;
  wire [13:0] p5_smul_58754_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___293_comb;
  wire [13:0] p5_smul_58760_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___294_comb;
  wire [24:0] p5_concat_147462_comb;
  wire [24:0] p5_concat_147463_comb;
  wire [13:0] p5_smul_58770_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___297_comb;
  wire [13:0] p5_smul_58776_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___298_comb;
  wire [24:0] p5_concat_147468_comb;
  wire [24:0] p5_concat_147469_comb;
  wire [13:0] p5_smul_58786_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___301_comb;
  wire [13:0] p5_smul_58792_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___302_comb;
  wire [24:0] p5_concat_147474_comb;
  wire [24:0] p5_concat_147481_comb;
  wire [13:0] p5_smul_58818_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___309_comb;
  wire [13:0] p5_smul_58824_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___310_comb;
  wire [24:0] p5_concat_147486_comb;
  wire [24:0] p5_concat_147487_comb;
  wire [13:0] p5_smul_58834_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___313_comb;
  wire [13:0] p5_smul_58840_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___314_comb;
  wire [24:0] p5_concat_147492_comb;
  wire [24:0] p5_concat_147493_comb;
  wire [13:0] p5_smul_58850_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___317_comb;
  wire [13:0] p5_smul_58856_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___318_comb;
  wire [24:0] p5_concat_147498_comb;
  wire [23:0] p5_concat_147507_comb;
  wire [24:0] p5_concat_147508_comb;
  wire [23:0] p5_concat_147509_comb;
  wire [23:0] p5_concat_147512_comb;
  wire [24:0] p5_concat_147513_comb;
  wire [23:0] p5_concat_147514_comb;
  wire [23:0] p5_concat_147515_comb;
  wire [24:0] p5_concat_147516_comb;
  wire [23:0] p5_concat_147517_comb;
  wire [24:0] p5_concat_147518_comb;
  wire [24:0] p5_concat_147519_comb;
  wire [23:0] p5_concat_147520_comb;
  wire [24:0] p5_concat_147521_comb;
  wire [23:0] p5_concat_147522_comb;
  wire [23:0] p5_concat_147523_comb;
  wire [24:0] p5_concat_147524_comb;
  wire [23:0] p5_concat_147525_comb;
  wire [23:0] p5_concat_147528_comb;
  wire [24:0] p5_concat_147529_comb;
  wire [23:0] p5_concat_147530_comb;
  wire [23:0] p5_concat_147539_comb;
  wire [24:0] p5_concat_147540_comb;
  wire [23:0] p5_concat_147541_comb;
  wire [23:0] p5_concat_147544_comb;
  wire [24:0] p5_concat_147545_comb;
  wire [23:0] p5_concat_147546_comb;
  wire [23:0] p5_concat_147547_comb;
  wire [24:0] p5_concat_147548_comb;
  wire [23:0] p5_concat_147549_comb;
  wire [24:0] p5_concat_147550_comb;
  wire [24:0] p5_concat_147551_comb;
  wire [23:0] p5_concat_147552_comb;
  wire [24:0] p5_concat_147553_comb;
  wire [23:0] p5_concat_147554_comb;
  wire [23:0] p5_concat_147555_comb;
  wire [24:0] p5_concat_147556_comb;
  wire [23:0] p5_concat_147557_comb;
  wire [23:0] p5_concat_147560_comb;
  wire [24:0] p5_concat_147561_comb;
  wire [23:0] p5_concat_147562_comb;
  wire [13:0] p5_smul_59006_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___356_comb;
  wire [24:0] p5_concat_147571_comb;
  wire [24:0] p5_concat_147572_comb;
  wire [13:0] p5_smul_59020_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___359_comb;
  wire [13:0] p5_smul_59022_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___360_comb;
  wire [24:0] p5_concat_147577_comb;
  wire [24:0] p5_concat_147578_comb;
  wire [13:0] p5_smul_59036_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___363_comb;
  wire [13:0] p5_smul_59038_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___364_comb;
  wire [24:0] p5_concat_147583_comb;
  wire [24:0] p5_concat_147584_comb;
  wire [13:0] p5_smul_59052_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___367_comb;
  wire [13:0] p5_smul_59070_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___372_comb;
  wire [24:0] p5_concat_147595_comb;
  wire [24:0] p5_concat_147596_comb;
  wire [13:0] p5_smul_59084_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___375_comb;
  wire [13:0] p5_smul_59086_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___376_comb;
  wire [24:0] p5_concat_147601_comb;
  wire [24:0] p5_concat_147602_comb;
  wire [13:0] p5_smul_59100_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___379_comb;
  wire [13:0] p5_smul_59102_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___380_comb;
  wire [24:0] p5_concat_147607_comb;
  wire [24:0] p5_concat_147608_comb;
  wire [13:0] p5_smul_59116_NarrowedMult__comb;
  wire [8:0] p5_smul_57330_TrailingBits___383_comb;
  wire [31:0] p5_prod__519_comb;
  wire [31:0] p5_prod__534_comb;
  wire [31:0] p5_prod__775_comb;
  wire [31:0] p5_prod__790_comb;
  wire [31:0] p5_prod__517_comb;
  wire [31:0] p5_prod__520_comb;
  wire [31:0] p5_prod__524_comb;
  wire [31:0] p5_prod__529_comb;
  wire [31:0] p5_prod__535_comb;
  wire [31:0] p5_prod__542_comb;
  wire [31:0] p5_prod__549_comb;
  wire [31:0] p5_prod__555_comb;
  wire [31:0] p5_prod__593_comb;
  wire [31:0] p5_prod__599_comb;
  wire [31:0] p5_prod__721_comb;
  wire [31:0] p5_prod__727_comb;
  wire [31:0] p5_prod__773_comb;
  wire [31:0] p5_prod__776_comb;
  wire [31:0] p5_prod__780_comb;
  wire [31:0] p5_prod__785_comb;
  wire [31:0] p5_prod__791_comb;
  wire [31:0] p5_prod__798_comb;
  wire [31:0] p5_prod__805_comb;
  wire [31:0] p5_prod__811_comb;
  wire [31:0] p5_prod__849_comb;
  wire [31:0] p5_prod__855_comb;
  wire [31:0] p5_prod__977_comb;
  wire [31:0] p5_prod__983_comb;
  wire [31:0] p5_prod__536_comb;
  wire [31:0] p5_prod__543_comb;
  wire [31:0] p5_prod__600_comb;
  wire [31:0] p5_prod__607_comb;
  wire [31:0] p5_prod__728_comb;
  wire [31:0] p5_prod__735_comb;
  wire [31:0] p5_prod__792_comb;
  wire [31:0] p5_prod__799_comb;
  wire [31:0] p5_prod__856_comb;
  wire [31:0] p5_prod__863_comb;
  wire [31:0] p5_prod__984_comb;
  wire [31:0] p5_prod__991_comb;
  wire [31:0] p5_prod__532_comb;
  wire [31:0] p5_prod__570_comb;
  wire [31:0] p5_prod__788_comb;
  wire [31:0] p5_prod__826_comb;
  wire [31:0] p5_prod__539_comb;
  wire [31:0] p5_prod__546_comb;
  wire [31:0] p5_prod__553_comb;
  wire [31:0] p5_prod__559_comb;
  wire [31:0] p5_prod__564_comb;
  wire [31:0] p5_prod__568_comb;
  wire [31:0] p5_prod__571_comb;
  wire [31:0] p5_prod__573_comb;
  wire [31:0] p5_prod__623_comb;
  wire [31:0] p5_prod__628_comb;
  wire [31:0] p5_prod__751_comb;
  wire [31:0] p5_prod__756_comb;
  wire [31:0] p5_prod__795_comb;
  wire [31:0] p5_prod__802_comb;
  wire [31:0] p5_prod__809_comb;
  wire [31:0] p5_prod__815_comb;
  wire [31:0] p5_prod__820_comb;
  wire [31:0] p5_prod__824_comb;
  wire [31:0] p5_prod__827_comb;
  wire [31:0] p5_prod__829_comb;
  wire [31:0] p5_prod__879_comb;
  wire [31:0] p5_prod__884_comb;
  wire [31:0] p5_prod__1007_comb;
  wire [31:0] p5_prod__1012_comb;
  wire [31:0] p5_prod__554_comb;
  wire [31:0] p5_prod__574_comb;
  wire [31:0] p5_prod__810_comb;
  wire [31:0] p5_prod__830_comb;
  wire [31:0] p5_prod__523_comb;
  wire [31:0] p5_prod__528_comb;
  wire [31:0] p5_prod__587_comb;
  wire [31:0] p5_prod__592_comb;
  wire [31:0] p5_prod__715_comb;
  wire [31:0] p5_prod__720_comb;
  wire [31:0] p5_prod__843_comb;
  wire [31:0] p5_prod__848_comb;
  wire [31:0] p5_prod__971_comb;
  wire [31:0] p5_prod__976_comb;
  wire [31:0] p5_prod__525_comb;
  wire [31:0] p5_prod__556_comb;
  wire [31:0] p5_prod__545_comb;
  wire [31:0] p5_prod__563_comb;
  wire [31:0] p5_prod__547_comb;
  wire [31:0] p5_prod__575_comb;
  wire [31:0] p5_or_149154_comb;
  wire [31:0] p5_or_149155_comb;
  wire [31:0] p5_or_149319_comb;
  wire [31:0] p5_or_149326_comb;
  wire [31:0] p5_or_149370_comb;
  wire [31:0] p5_or_149371_comb;
  wire [31:0] p5_or_149527_comb;
  wire [31:0] p5_or_149534_comb;
  wire [7:0] p5_smul_57326_TrailingBits___200_comb;
  wire [7:0] p5_smul_57326_TrailingBits___201_comb;
  wire [7:0] p5_smul_57326_TrailingBits___202_comb;
  wire [7:0] p5_smul_57326_TrailingBits___203_comb;
  wire [7:0] p5_smul_57326_TrailingBits___204_comb;
  wire [7:0] p5_smul_57326_TrailingBits___205_comb;
  wire [7:0] p5_smul_57326_TrailingBits___206_comb;
  wire [7:0] p5_smul_57326_TrailingBits___207_comb;
  wire [7:0] p5_smul_57326_TrailingBits___208_comb;
  wire [7:0] p5_smul_57326_TrailingBits___209_comb;
  wire [7:0] p5_smul_57326_TrailingBits___210_comb;
  wire [7:0] p5_smul_57326_TrailingBits___211_comb;
  wire [7:0] p5_smul_57326_TrailingBits___212_comb;
  wire [7:0] p5_smul_57326_TrailingBits___213_comb;
  wire [7:0] p5_smul_57326_TrailingBits___214_comb;
  wire [7:0] p5_smul_57326_TrailingBits___215_comb;
  wire [7:0] p5_smul_57326_TrailingBits___216_comb;
  wire [7:0] p5_smul_57326_TrailingBits___217_comb;
  wire [7:0] p5_smul_57326_TrailingBits___218_comb;
  wire [7:0] p5_smul_57326_TrailingBits___219_comb;
  wire [7:0] p5_smul_57326_TrailingBits___220_comb;
  wire [7:0] p5_smul_57326_TrailingBits___221_comb;
  wire [7:0] p5_smul_57326_TrailingBits___222_comb;
  wire [7:0] p5_smul_57326_TrailingBits___223_comb;
  wire [7:0] p5_smul_57326_TrailingBits___232_comb;
  wire [7:0] p5_smul_57326_TrailingBits___233_comb;
  wire [7:0] p5_smul_57326_TrailingBits___234_comb;
  wire [7:0] p5_smul_57326_TrailingBits___235_comb;
  wire [7:0] p5_smul_57326_TrailingBits___236_comb;
  wire [7:0] p5_smul_57326_TrailingBits___237_comb;
  wire [7:0] p5_smul_57326_TrailingBits___238_comb;
  wire [7:0] p5_smul_57326_TrailingBits___239_comb;
  wire [7:0] p5_smul_57326_TrailingBits___240_comb;
  wire [7:0] p5_smul_57326_TrailingBits___241_comb;
  wire [7:0] p5_smul_57326_TrailingBits___242_comb;
  wire [7:0] p5_smul_57326_TrailingBits___243_comb;
  wire [7:0] p5_smul_57326_TrailingBits___244_comb;
  wire [7:0] p5_smul_57326_TrailingBits___245_comb;
  wire [7:0] p5_smul_57326_TrailingBits___246_comb;
  wire [7:0] p5_smul_57326_TrailingBits___247_comb;
  wire [7:0] p5_smul_57326_TrailingBits___248_comb;
  wire [7:0] p5_smul_57326_TrailingBits___249_comb;
  wire [7:0] p5_smul_57326_TrailingBits___250_comb;
  wire [7:0] p5_smul_57326_TrailingBits___251_comb;
  wire [7:0] p5_smul_57326_TrailingBits___252_comb;
  wire [7:0] p5_smul_57326_TrailingBits___253_comb;
  wire [7:0] p5_smul_57326_TrailingBits___254_comb;
  wire [7:0] p5_smul_57326_TrailingBits___255_comb;
  wire [31:0] p5_prod__583_comb;
  wire [31:0] p5_prod__598_comb;
  wire [31:0] p5_prod__647_comb;
  wire [22:0] p5_concat_147817_comb;
  wire [22:0] p5_concat_147818_comb;
  wire [31:0] p5_prod__662_comb;
  wire [31:0] p5_prod__711_comb;
  wire [31:0] p5_prod__726_comb;
  wire [31:0] p5_prod__839_comb;
  wire [31:0] p5_prod__854_comb;
  wire [31:0] p5_prod__903_comb;
  wire [22:0] p5_concat_147841_comb;
  wire [22:0] p5_concat_147842_comb;
  wire [31:0] p5_prod__918_comb;
  wire [31:0] p5_prod__967_comb;
  wire [31:0] p5_prod__982_comb;
  wire [31:0] p5_prod__581_comb;
  wire [31:0] p5_prod__584_comb;
  wire [31:0] p5_prod__588_comb;
  wire [31:0] p5_prod__606_comb;
  wire [31:0] p5_prod__613_comb;
  wire [31:0] p5_prod__619_comb;
  wire [31:0] p5_prod__645_comb;
  wire [31:0] p5_prod__648_comb;
  wire [31:0] p5_prod__652_comb;
  wire [31:0] p5_prod__657_comb;
  wire [31:0] p5_prod__663_comb;
  wire [31:0] p5_prod__670_comb;
  wire [31:0] p5_prod__677_comb;
  wire [31:0] p5_prod__683_comb;
  wire [31:0] p5_prod__709_comb;
  wire [31:0] p5_prod__712_comb;
  wire [31:0] p5_prod__716_comb;
  wire [31:0] p5_prod__734_comb;
  wire [31:0] p5_prod__741_comb;
  wire [31:0] p5_prod__747_comb;
  wire [31:0] p5_prod__837_comb;
  wire [31:0] p5_prod__840_comb;
  wire [31:0] p5_prod__844_comb;
  wire [31:0] p5_prod__862_comb;
  wire [31:0] p5_prod__869_comb;
  wire [31:0] p5_prod__875_comb;
  wire [31:0] p5_prod__901_comb;
  wire [31:0] p5_prod__904_comb;
  wire [31:0] p5_prod__908_comb;
  wire [31:0] p5_prod__913_comb;
  wire [31:0] p5_prod__919_comb;
  wire [31:0] p5_prod__926_comb;
  wire [31:0] p5_prod__933_comb;
  wire [31:0] p5_prod__939_comb;
  wire [31:0] p5_prod__965_comb;
  wire [31:0] p5_prod__968_comb;
  wire [31:0] p5_prod__972_comb;
  wire [31:0] p5_prod__990_comb;
  wire [31:0] p5_prod__997_comb;
  wire [31:0] p5_prod__1003_comb;
  wire [22:0] p5_concat_147953_comb;
  wire [22:0] p5_concat_147958_comb;
  wire [22:0] p5_concat_147959_comb;
  wire [31:0] p5_prod__664_comb;
  wire [31:0] p5_prod__671_comb;
  wire [22:0] p5_concat_147964_comb;
  wire [22:0] p5_concat_147965_comb;
  wire [22:0] p5_concat_147970_comb;
  wire [22:0] p5_concat_147977_comb;
  wire [22:0] p5_concat_147982_comb;
  wire [22:0] p5_concat_147983_comb;
  wire [31:0] p5_prod__920_comb;
  wire [31:0] p5_prod__927_comb;
  wire [22:0] p5_concat_147988_comb;
  wire [22:0] p5_concat_147989_comb;
  wire [22:0] p5_concat_147994_comb;
  wire [31:0] p5_prod__596_comb;
  wire [22:0] p5_concat_148003_comb;
  wire [22:0] p5_concat_148004_comb;
  wire [31:0] p5_prod__634_comb;
  wire [31:0] p5_prod__660_comb;
  wire [22:0] p5_concat_148009_comb;
  wire [22:0] p5_concat_148010_comb;
  wire [31:0] p5_prod__698_comb;
  wire [31:0] p5_prod__724_comb;
  wire [22:0] p5_concat_148015_comb;
  wire [22:0] p5_concat_148016_comb;
  wire [31:0] p5_prod__762_comb;
  wire [31:0] p5_prod__852_comb;
  wire [22:0] p5_concat_148027_comb;
  wire [22:0] p5_concat_148028_comb;
  wire [31:0] p5_prod__890_comb;
  wire [31:0] p5_prod__916_comb;
  wire [22:0] p5_concat_148033_comb;
  wire [22:0] p5_concat_148034_comb;
  wire [31:0] p5_prod__954_comb;
  wire [31:0] p5_prod__980_comb;
  wire [22:0] p5_concat_148039_comb;
  wire [22:0] p5_concat_148040_comb;
  wire [31:0] p5_prod__1018_comb;
  wire [31:0] p5_prod__603_comb;
  wire [31:0] p5_prod__610_comb;
  wire [31:0] p5_prod__617_comb;
  wire [31:0] p5_prod__632_comb;
  wire [31:0] p5_prod__635_comb;
  wire [31:0] p5_prod__637_comb;
  wire [31:0] p5_prod__667_comb;
  wire [31:0] p5_prod__674_comb;
  wire [31:0] p5_prod__681_comb;
  wire [31:0] p5_prod__687_comb;
  wire [31:0] p5_prod__692_comb;
  wire [31:0] p5_prod__696_comb;
  wire [31:0] p5_prod__699_comb;
  wire [31:0] p5_prod__701_comb;
  wire [31:0] p5_prod__731_comb;
  wire [31:0] p5_prod__738_comb;
  wire [31:0] p5_prod__745_comb;
  wire [31:0] p5_prod__760_comb;
  wire [31:0] p5_prod__763_comb;
  wire [31:0] p5_prod__765_comb;
  wire [31:0] p5_prod__859_comb;
  wire [31:0] p5_prod__866_comb;
  wire [31:0] p5_prod__873_comb;
  wire [31:0] p5_prod__888_comb;
  wire [31:0] p5_prod__891_comb;
  wire [31:0] p5_prod__893_comb;
  wire [31:0] p5_prod__923_comb;
  wire [31:0] p5_prod__930_comb;
  wire [31:0] p5_prod__937_comb;
  wire [31:0] p5_prod__943_comb;
  wire [31:0] p5_prod__948_comb;
  wire [31:0] p5_prod__952_comb;
  wire [31:0] p5_prod__955_comb;
  wire [31:0] p5_prod__957_comb;
  wire [31:0] p5_prod__987_comb;
  wire [31:0] p5_prod__994_comb;
  wire [31:0] p5_prod__1001_comb;
  wire [31:0] p5_prod__1016_comb;
  wire [31:0] p5_prod__1019_comb;
  wire [31:0] p5_prod__1021_comb;
  wire [22:0] p5_concat_148145_comb;
  wire [31:0] p5_prod__618_comb;
  wire [31:0] p5_prod__638_comb;
  wire [22:0] p5_concat_148150_comb;
  wire [22:0] p5_concat_148151_comb;
  wire [31:0] p5_prod__682_comb;
  wire [31:0] p5_prod__702_comb;
  wire [22:0] p5_concat_148156_comb;
  wire [22:0] p5_concat_148157_comb;
  wire [31:0] p5_prod__746_comb;
  wire [31:0] p5_prod__766_comb;
  wire [22:0] p5_concat_148162_comb;
  wire [22:0] p5_concat_148169_comb;
  wire [31:0] p5_prod__874_comb;
  wire [31:0] p5_prod__894_comb;
  wire [22:0] p5_concat_148174_comb;
  wire [22:0] p5_concat_148175_comb;
  wire [31:0] p5_prod__938_comb;
  wire [31:0] p5_prod__958_comb;
  wire [22:0] p5_concat_148180_comb;
  wire [22:0] p5_concat_148181_comb;
  wire [31:0] p5_prod__1002_comb;
  wire [31:0] p5_prod__1022_comb;
  wire [22:0] p5_concat_148186_comb;
  wire [31:0] p5_or_148397_comb;
  wire [31:0] p5_or_148404_comb;
  wire [31:0] p5_or_148437_comb;
  wire [31:0] p5_or_148444_comb;
  wire [31:0] p5_or_148477_comb;
  wire [31:0] p5_or_148484_comb;
  wire [31:0] p5_or_148487_comb;
  wire [31:0] p5_or_148494_comb;
  wire [31:0] p5_or_148504_comb;
  wire [31:0] p5_or_148507_comb;
  wire [31:0] p5_or_148544_comb;
  wire [31:0] p5_or_148547_comb;
  wire [31:0] p5_or_148557_comb;
  wire [31:0] p5_or_148564_comb;
  wire [31:0] p5_or_148567_comb;
  wire [31:0] p5_or_148574_comb;
  wire [31:0] p5_or_148584_comb;
  wire [31:0] p5_or_148587_comb;
  wire [31:0] p5_or_148624_comb;
  wire [31:0] p5_or_148627_comb;
  wire [31:0] p5_or_148639_comb;
  wire [31:0] p5_or_148642_comb;
  wire [31:0] p5_or_148649_comb;
  wire [31:0] p5_or_148652_comb;
  wire [31:0] p5_or_148669_comb;
  wire [31:0] p5_or_148672_comb;
  wire [31:0] p5_or_148679_comb;
  wire [31:0] p5_or_148682_comb;
  wire [31:0] p5_or_148689_comb;
  wire [31:0] p5_or_148692_comb;
  wire [31:0] p5_or_148709_comb;
  wire [31:0] p5_or_148712_comb;
  wire [31:0] p5_or_148717_comb;
  wire [31:0] p5_or_148724_comb;
  wire [31:0] p5_or_148757_comb;
  wire [31:0] p5_or_148764_comb;
  wire [31:0] p5_or_148799_comb;
  wire [31:0] p5_or_148804_comb;
  wire [31:0] p5_or_148807_comb;
  wire [31:0] p5_or_148812_comb;
  wire [31:0] p5_or_148824_comb;
  wire [31:0] p5_or_148827_comb;
  wire [31:0] p5_or_148864_comb;
  wire [31:0] p5_or_148867_comb;
  wire [31:0] p5_or_148879_comb;
  wire [31:0] p5_or_148884_comb;
  wire [31:0] p5_or_148887_comb;
  wire [31:0] p5_or_148892_comb;
  wire [31:0] p5_or_148904_comb;
  wire [31:0] p5_or_148907_comb;
  wire [31:0] p5_or_148944_comb;
  wire [31:0] p5_or_148947_comb;
  wire [31:0] p5_or_148959_comb;
  wire [31:0] p5_or_148962_comb;
  wire [31:0] p5_or_148999_comb;
  wire [31:0] p5_or_149002_comb;
  wire [31:0] p5_or_149134_comb;
  wire [31:0] p5_or_149135_comb;
  wire [31:0] p5_or_149140_comb;
  wire [31:0] p5_or_149141_comb;
  wire [31:0] p5_or_149148_comb;
  wire [31:0] p5_or_149149_comb;
  wire [31:0] p5_or_149160_comb;
  wire [31:0] p5_or_149161_comb;
  wire [31:0] p5_or_149168_comb;
  wire [31:0] p5_or_149169_comb;
  wire [31:0] p5_or_149291_comb;
  wire [31:0] p5_or_149298_comb;
  wire [31:0] p5_or_149350_comb;
  wire [31:0] p5_or_149351_comb;
  wire [31:0] p5_or_149507_comb;
  wire [31:0] p5_or_149514_comb;
  wire [15:0] p5_sel_149547_comb;
  wire [15:0] p5_sel_149548_comb;
  wire [15:0] p5_sel_149549_comb;
  wire [15:0] p5_sel_149550_comb;
  wire [15:0] p5_sel_149551_comb;
  wire [15:0] p5_sel_149552_comb;
  wire [15:0] p5_sel_149553_comb;
  wire [15:0] p5_sel_149554_comb;
  wire [15:0] p5_sel_149555_comb;
  wire [15:0] p5_sel_149556_comb;
  wire [15:0] p5_sel_149557_comb;
  wire [15:0] p5_sel_149558_comb;
  wire [15:0] p5_sel_149559_comb;
  wire [15:0] p5_sel_149560_comb;
  wire [15:0] p5_sel_149561_comb;
  wire [15:0] p5_sel_149562_comb;
  wire [15:0] p5_shifted__72_comb;
  wire [15:0] p5_shifted__73_comb;
  wire [15:0] p5_shifted__74_comb;
  wire [15:0] p5_shifted__75_comb;
  wire [15:0] p5_shifted__76_comb;
  wire [15:0] p5_shifted__77_comb;
  wire [15:0] p5_shifted__78_comb;
  wire [15:0] p5_shifted__79_comb;
  wire [15:0] p5_shifted__80_comb;
  wire [15:0] p5_shifted__81_comb;
  wire [15:0] p5_shifted__82_comb;
  wire [15:0] p5_shifted__83_comb;
  wire [15:0] p5_shifted__84_comb;
  wire [15:0] p5_shifted__85_comb;
  wire [15:0] p5_shifted__86_comb;
  wire [15:0] p5_shifted__87_comb;
  wire [15:0] p5_shifted__88_comb;
  wire [15:0] p5_shifted__89_comb;
  wire [15:0] p5_shifted__90_comb;
  wire [15:0] p5_shifted__91_comb;
  wire [15:0] p5_shifted__92_comb;
  wire [15:0] p5_shifted__93_comb;
  wire [15:0] p5_shifted__94_comb;
  wire [15:0] p5_shifted__95_comb;
  wire [15:0] p5_shifted__104_comb;
  wire [15:0] p5_shifted__105_comb;
  wire [15:0] p5_shifted__106_comb;
  wire [15:0] p5_shifted__107_comb;
  wire [15:0] p5_shifted__108_comb;
  wire [15:0] p5_shifted__109_comb;
  wire [15:0] p5_shifted__110_comb;
  wire [15:0] p5_shifted__111_comb;
  wire [15:0] p5_shifted__112_comb;
  wire [15:0] p5_shifted__113_comb;
  wire [15:0] p5_shifted__114_comb;
  wire [15:0] p5_shifted__115_comb;
  wire [15:0] p5_shifted__116_comb;
  wire [15:0] p5_shifted__117_comb;
  wire [15:0] p5_shifted__118_comb;
  wire [15:0] p5_shifted__119_comb;
  wire [15:0] p5_shifted__120_comb;
  wire [15:0] p5_shifted__121_comb;
  wire [15:0] p5_shifted__122_comb;
  wire [15:0] p5_shifted__123_comb;
  wire [15:0] p5_shifted__124_comb;
  wire [15:0] p5_shifted__125_comb;
  wire [15:0] p5_shifted__126_comb;
  wire [15:0] p5_shifted__127_comb;
  wire [31:0] p5_prod__651_comb;
  wire [31:0] p5_prod__656_comb;
  wire [31:0] p5_prod__907_comb;
  wire [31:0] p5_prod__912_comb;
  wire [31:0] p5_or_148497_comb;
  wire [31:0] p5_or_148514_comb;
  wire [31:0] p5_or_148517_comb;
  wire [31:0] p5_or_148524_comb;
  wire [31:0] p5_or_148527_comb;
  wire [31:0] p5_or_148534_comb;
  wire [31:0] p5_or_148537_comb;
  wire [31:0] p5_or_148554_comb;
  wire [31:0] p5_or_148577_comb;
  wire [31:0] p5_or_148594_comb;
  wire [31:0] p5_or_148597_comb;
  wire [31:0] p5_or_148604_comb;
  wire [31:0] p5_or_148607_comb;
  wire [31:0] p5_or_148614_comb;
  wire [31:0] p5_or_148617_comb;
  wire [31:0] p5_or_148634_comb;
  wire [31:0] p5_prod__589_comb;
  wire [31:0] p5_prod__620_comb;
  wire [31:0] p5_prod__653_comb;
  wire [31:0] p5_prod__684_comb;
  wire [31:0] p5_prod__717_comb;
  wire [31:0] p5_prod__748_comb;
  wire [31:0] p5_prod__845_comb;
  wire [31:0] p5_prod__876_comb;
  wire [31:0] p5_prod__909_comb;
  wire [31:0] p5_prod__940_comb;
  wire [31:0] p5_prod__973_comb;
  wire [31:0] p5_prod__1004_comb;
  wire [31:0] p5_prod__609_comb;
  wire [31:0] p5_prod__627_comb;
  wire [31:0] p5_prod__673_comb;
  wire [31:0] p5_prod__691_comb;
  wire [31:0] p5_prod__737_comb;
  wire [31:0] p5_prod__755_comb;
  wire [31:0] p5_prod__865_comb;
  wire [31:0] p5_prod__883_comb;
  wire [31:0] p5_prod__929_comb;
  wire [31:0] p5_prod__947_comb;
  wire [31:0] p5_prod__993_comb;
  wire [31:0] p5_prod__1011_comb;
  wire [31:0] p5_or_148819_comb;
  wire [31:0] p5_or_148832_comb;
  wire [31:0] p5_or_148839_comb;
  wire [31:0] p5_or_148844_comb;
  wire [31:0] p5_or_148847_comb;
  wire [31:0] p5_or_148852_comb;
  wire [31:0] p5_or_148859_comb;
  wire [31:0] p5_or_148872_comb;
  wire [31:0] p5_or_148899_comb;
  wire [31:0] p5_or_148912_comb;
  wire [31:0] p5_or_148919_comb;
  wire [31:0] p5_or_148924_comb;
  wire [31:0] p5_or_148927_comb;
  wire [31:0] p5_or_148932_comb;
  wire [31:0] p5_or_148939_comb;
  wire [31:0] p5_or_148952_comb;
  wire [31:0] p5_prod__611_comb;
  wire [31:0] p5_prod__639_comb;
  wire [31:0] p5_prod__675_comb;
  wire [31:0] p5_prod__703_comb;
  wire [31:0] p5_prod__739_comb;
  wire [31:0] p5_prod__767_comb;
  wire [31:0] p5_prod__867_comb;
  wire [31:0] p5_prod__895_comb;
  wire [31:0] p5_prod__931_comb;
  wire [31:0] p5_prod__959_comb;
  wire [31:0] p5_prod__995_comb;
  wire [31:0] p5_prod__1023_comb;
  wire [7:0] p5_sel_148221_comb;
  wire [7:0] p5_sel_148224_comb;
  wire [7:0] p5_sel_148227_comb;
  wire [7:0] p5_sel_148230_comb;
  wire [7:0] p5_sel_148233_comb;
  wire [7:0] p5_sel_148236_comb;
  wire [7:0] p5_sel_148239_comb;
  wire [7:0] p5_sel_148242_comb;
  wire [7:0] p5_sel_148245_comb;
  wire [7:0] p5_sel_148248_comb;
  wire [7:0] p5_sel_148251_comb;
  wire [7:0] p5_sel_148254_comb;
  wire [7:0] p5_sel_148257_comb;
  wire [7:0] p5_sel_148260_comb;
  wire [7:0] p5_sel_148263_comb;
  wire [7:0] p5_sel_148266_comb;
  wire [7:0] p5_sel_148269_comb;
  wire [7:0] p5_sel_148272_comb;
  wire [7:0] p5_sel_148275_comb;
  wire [7:0] p5_sel_148278_comb;
  wire [7:0] p5_sel_148281_comb;
  wire [7:0] p5_sel_148284_comb;
  wire [7:0] p5_sel_148287_comb;
  wire [7:0] p5_sel_148290_comb;
  wire [7:0] p5_sel_148325_comb;
  wire [7:0] p5_sel_148328_comb;
  wire [7:0] p5_sel_148331_comb;
  wire [7:0] p5_sel_148334_comb;
  wire [7:0] p5_sel_148337_comb;
  wire [7:0] p5_sel_148340_comb;
  wire [7:0] p5_sel_148343_comb;
  wire [7:0] p5_sel_148346_comb;
  wire [7:0] p5_sel_148349_comb;
  wire [7:0] p5_sel_148352_comb;
  wire [7:0] p5_sel_148355_comb;
  wire [7:0] p5_sel_148358_comb;
  wire [7:0] p5_sel_148361_comb;
  wire [7:0] p5_sel_148364_comb;
  wire [7:0] p5_sel_148367_comb;
  wire [7:0] p5_sel_148370_comb;
  wire [7:0] p5_sel_148373_comb;
  wire [7:0] p5_sel_148376_comb;
  wire [7:0] p5_sel_148379_comb;
  wire [7:0] p5_sel_148382_comb;
  wire [7:0] p5_sel_148385_comb;
  wire [7:0] p5_sel_148388_comb;
  wire [7:0] p5_sel_148391_comb;
  wire [7:0] p5_sel_148394_comb;
  wire [31:0] p5_or_148407_comb;
  wire [31:0] p5_or_148414_comb;
  wire [31:0] p5_or_148417_comb;
  wire [31:0] p5_or_148424_comb;
  wire [31:0] p5_or_148427_comb;
  wire [31:0] p5_or_148434_comb;
  wire [31:0] p5_or_148447_comb;
  wire [31:0] p5_or_148454_comb;
  wire [31:0] p5_or_148457_comb;
  wire [31:0] p5_or_148464_comb;
  wire [31:0] p5_or_148467_comb;
  wire [31:0] p5_or_148474_comb;
  wire [31:0] p5_or_148659_comb;
  wire [31:0] p5_or_148662_comb;
  wire [31:0] p5_or_148699_comb;
  wire [31:0] p5_or_148702_comb;
  wire [31:0] p5_or_148727_comb;
  wire [31:0] p5_or_148734_comb;
  wire [31:0] p5_or_148737_comb;
  wire [31:0] p5_or_148744_comb;
  wire [31:0] p5_or_148747_comb;
  wire [31:0] p5_or_148754_comb;
  wire [31:0] p5_or_148767_comb;
  wire [31:0] p5_or_148774_comb;
  wire [31:0] p5_or_148777_comb;
  wire [31:0] p5_or_148784_comb;
  wire [31:0] p5_or_148787_comb;
  wire [31:0] p5_or_148794_comb;
  wire [31:0] p5_or_148969_comb;
  wire [31:0] p5_or_148972_comb;
  wire [31:0] p5_or_148979_comb;
  wire [31:0] p5_or_148982_comb;
  wire [31:0] p5_or_148989_comb;
  wire [31:0] p5_or_148992_comb;
  wire [31:0] p5_or_149009_comb;
  wire [31:0] p5_or_149012_comb;
  wire [31:0] p5_or_149019_comb;
  wire [31:0] p5_or_149022_comb;
  wire [31:0] p5_or_149029_comb;
  wire [31:0] p5_or_149032_comb;
  wire p5_sgt_149059_comb;
  wire p5_sgt_149060_comb;
  wire p5_sgt_149061_comb;
  wire p5_sgt_149062_comb;
  wire p5_sgt_149063_comb;
  wire p5_sgt_149064_comb;
  wire p5_sgt_149065_comb;
  wire p5_sgt_149066_comb;
  wire p5_sgt_149067_comb;
  wire p5_sgt_149068_comb;
  wire p5_sgt_149069_comb;
  wire p5_sgt_149070_comb;
  wire p5_sgt_149071_comb;
  wire p5_sgt_149072_comb;
  wire p5_sgt_149073_comb;
  wire p5_sgt_149074_comb;
  wire p5_sgt_149075_comb;
  wire p5_sgt_149076_comb;
  wire p5_sgt_149077_comb;
  wire p5_sgt_149078_comb;
  wire p5_sgt_149079_comb;
  wire p5_sgt_149080_comb;
  wire p5_sgt_149081_comb;
  wire p5_sgt_149082_comb;
  wire p5_sgt_149107_comb;
  wire p5_sgt_149108_comb;
  wire p5_sgt_149109_comb;
  wire p5_sgt_149110_comb;
  wire p5_sgt_149111_comb;
  wire p5_sgt_149112_comb;
  wire p5_sgt_149113_comb;
  wire p5_sgt_149114_comb;
  wire p5_sgt_149115_comb;
  wire p5_sgt_149116_comb;
  wire p5_sgt_149117_comb;
  wire p5_sgt_149118_comb;
  wire p5_sgt_149119_comb;
  wire p5_sgt_149120_comb;
  wire p5_sgt_149121_comb;
  wire p5_sgt_149122_comb;
  wire p5_sgt_149123_comb;
  wire p5_sgt_149124_comb;
  wire p5_sgt_149125_comb;
  wire p5_sgt_149126_comb;
  wire p5_sgt_149127_comb;
  wire p5_sgt_149128_comb;
  wire p5_sgt_149129_comb;
  wire p5_sgt_149130_comb;
  wire p5_slt_149139_comb;
  wire p5_slt_149142_comb;
  wire p5_slt_149143_comb;
  wire [31:0] p5_or_149144_comb;
  wire [31:0] p5_or_149145_comb;
  wire p5_slt_149146_comb;
  wire p5_slt_149147_comb;
  wire p5_slt_149150_comb;
  wire p5_slt_149159_comb;
  wire p5_slt_149162_comb;
  wire p5_slt_149163_comb;
  wire [31:0] p5_or_149164_comb;
  wire [31:0] p5_or_149165_comb;
  wire p5_slt_149166_comb;
  wire p5_slt_149167_comb;
  wire p5_slt_149170_comb;
  wire p5_slt_149191_comb;
  wire [13:0] p5_bit_slice_149192_comb;
  wire p5_slt_149193_comb;
  wire p5_slt_149194_comb;
  wire p5_slt_149201_comb;
  wire p5_slt_149202_comb;
  wire p5_slt_149203_comb;
  wire [13:0] p5_bit_slice_149204_comb;
  wire p5_slt_149205_comb;
  wire [13:0] p5_bit_slice_149206_comb;
  wire p5_slt_149207_comb;
  wire p5_slt_149208_comb;
  wire p5_slt_149209_comb;
  wire [13:0] p5_bit_slice_149210_comb;
  wire p5_slt_149211_comb;
  wire [13:0] p5_bit_slice_149212_comb;
  wire p5_slt_149213_comb;
  wire p5_slt_149214_comb;
  wire p5_slt_149215_comb;
  wire [13:0] p5_bit_slice_149216_comb;
  wire p5_slt_149217_comb;
  wire [13:0] p5_bit_slice_149218_comb;
  wire p5_slt_149219_comb;
  wire p5_slt_149220_comb;
  wire p5_slt_149227_comb;
  wire p5_slt_149228_comb;
  wire p5_slt_149229_comb;
  wire [13:0] p5_bit_slice_149230_comb;
  wire p5_slt_149251_comb;
  wire [13:0] p5_bit_slice_149252_comb;
  wire p5_slt_149253_comb;
  wire p5_slt_149254_comb;
  wire p5_slt_149261_comb;
  wire p5_slt_149262_comb;
  wire p5_slt_149263_comb;
  wire [13:0] p5_bit_slice_149264_comb;
  wire p5_slt_149265_comb;
  wire [13:0] p5_bit_slice_149266_comb;
  wire p5_slt_149267_comb;
  wire p5_slt_149268_comb;
  wire p5_slt_149269_comb;
  wire [13:0] p5_bit_slice_149270_comb;
  wire p5_slt_149271_comb;
  wire [13:0] p5_bit_slice_149272_comb;
  wire p5_slt_149273_comb;
  wire p5_slt_149274_comb;
  wire p5_slt_149275_comb;
  wire [13:0] p5_bit_slice_149276_comb;
  wire p5_slt_149277_comb;
  wire [13:0] p5_bit_slice_149278_comb;
  wire p5_slt_149279_comb;
  wire p5_slt_149280_comb;
  wire p5_slt_149287_comb;
  wire p5_slt_149288_comb;
  wire p5_slt_149289_comb;
  wire [13:0] p5_bit_slice_149290_comb;
  wire [31:0] p5_or_149299_comb;
  wire [31:0] p5_or_149306_comb;
  wire [31:0] p5_or_149307_comb;
  wire p5_slt_149308_comb;
  wire p5_slt_149309_comb;
  wire [31:0] p5_or_149310_comb;
  wire [31:0] p5_or_149311_comb;
  wire [31:0] p5_or_149318_comb;
  wire [31:0] p5_or_149327_comb;
  wire [31:0] p5_or_149334_comb;
  wire [31:0] p5_or_149335_comb;
  wire p5_slt_149336_comb;
  wire p5_slt_149337_comb;
  wire [31:0] p5_or_149338_comb;
  wire [31:0] p5_or_149339_comb;
  wire [31:0] p5_or_149346_comb;
  wire p5_slt_149355_comb;
  wire [31:0] p5_or_149356_comb;
  wire [31:0] p5_or_149357_comb;
  wire p5_slt_149358_comb;
  wire p5_slt_149359_comb;
  wire [31:0] p5_or_149360_comb;
  wire [31:0] p5_or_149361_comb;
  wire p5_slt_149362_comb;
  wire p5_slt_149363_comb;
  wire [31:0] p5_or_149364_comb;
  wire [31:0] p5_or_149365_comb;
  wire p5_slt_149366_comb;
  wire p5_slt_149375_comb;
  wire [31:0] p5_or_149376_comb;
  wire [31:0] p5_or_149377_comb;
  wire p5_slt_149378_comb;
  wire p5_slt_149379_comb;
  wire [31:0] p5_or_149380_comb;
  wire [31:0] p5_or_149381_comb;
  wire p5_slt_149382_comb;
  wire p5_slt_149383_comb;
  wire [31:0] p5_or_149384_comb;
  wire [31:0] p5_or_149385_comb;
  wire p5_slt_149386_comb;
  wire p5_slt_149407_comb;
  wire p5_slt_149408_comb;
  wire [13:0] p5_bit_slice_149409_comb;
  wire p5_slt_149410_comb;
  wire p5_slt_149417_comb;
  wire p5_slt_149418_comb;
  wire [13:0] p5_bit_slice_149419_comb;
  wire p5_slt_149420_comb;
  wire p5_slt_149421_comb;
  wire p5_slt_149422_comb;
  wire [13:0] p5_bit_slice_149423_comb;
  wire p5_slt_149424_comb;
  wire p5_slt_149425_comb;
  wire [13:0] p5_bit_slice_149426_comb;
  wire p5_slt_149427_comb;
  wire [13:0] p5_bit_slice_149428_comb;
  wire p5_slt_149429_comb;
  wire p5_slt_149430_comb;
  wire [13:0] p5_bit_slice_149431_comb;
  wire p5_slt_149432_comb;
  wire p5_slt_149433_comb;
  wire p5_slt_149434_comb;
  wire [13:0] p5_bit_slice_149435_comb;
  wire p5_slt_149436_comb;
  wire p5_slt_149443_comb;
  wire p5_slt_149444_comb;
  wire [13:0] p5_bit_slice_149445_comb;
  wire p5_slt_149446_comb;
  wire p5_slt_149467_comb;
  wire p5_slt_149468_comb;
  wire [13:0] p5_bit_slice_149469_comb;
  wire p5_slt_149470_comb;
  wire p5_slt_149477_comb;
  wire p5_slt_149478_comb;
  wire [13:0] p5_bit_slice_149479_comb;
  wire p5_slt_149480_comb;
  wire p5_slt_149481_comb;
  wire p5_slt_149482_comb;
  wire [13:0] p5_bit_slice_149483_comb;
  wire p5_slt_149484_comb;
  wire p5_slt_149485_comb;
  wire [13:0] p5_bit_slice_149486_comb;
  wire p5_slt_149487_comb;
  wire [13:0] p5_bit_slice_149488_comb;
  wire p5_slt_149489_comb;
  wire p5_slt_149490_comb;
  wire [13:0] p5_bit_slice_149491_comb;
  wire p5_slt_149492_comb;
  wire p5_slt_149493_comb;
  wire p5_slt_149494_comb;
  wire [13:0] p5_bit_slice_149495_comb;
  wire p5_slt_149496_comb;
  wire p5_slt_149503_comb;
  wire p5_slt_149504_comb;
  wire [13:0] p5_bit_slice_149505_comb;
  wire p5_slt_149506_comb;
  wire [31:0] p5_or_149515_comb;
  wire p5_slt_149516_comb;
  wire p5_slt_149517_comb;
  wire [31:0] p5_or_149518_comb;
  wire [31:0] p5_or_149519_comb;
  wire p5_slt_149520_comb;
  wire p5_slt_149521_comb;
  wire [31:0] p5_or_149522_comb;
  wire [31:0] p5_or_149523_comb;
  wire p5_slt_149524_comb;
  wire p5_slt_149525_comb;
  wire [31:0] p5_or_149526_comb;
  wire [31:0] p5_or_149535_comb;
  wire p5_slt_149536_comb;
  wire p5_slt_149537_comb;
  wire [31:0] p5_or_149538_comb;
  wire [31:0] p5_or_149539_comb;
  wire p5_slt_149540_comb;
  wire p5_slt_149541_comb;
  wire [31:0] p5_or_149542_comb;
  wire [31:0] p5_or_149543_comb;
  wire p5_slt_149544_comb;
  wire p5_slt_149545_comb;
  wire [31:0] p5_or_149546_comb;
  wire [14:0] p5_sel_149565_comb;
  wire [14:0] p5_bit_slice_149568_comb;
  wire [14:0] p5_bit_slice_149571_comb;
  wire [14:0] p5_sel_149574_comb;
  wire [14:0] p5_bit_slice_149577_comb;
  wire [14:0] p5_bit_slice_149580_comb;
  wire [14:0] p5_bit_slice_149583_comb;
  wire [14:0] p5_bit_slice_149586_comb;
  wire [14:0] p5_sel_149589_comb;
  wire [14:0] p5_sel_149600_comb;
  wire [14:0] p5_bit_slice_149603_comb;
  wire [14:0] p5_bit_slice_149606_comb;
  wire [14:0] p5_bit_slice_149609_comb;
  wire [14:0] p5_bit_slice_149612_comb;
  wire [13:0] p5_sel_149615_comb;
  wire [14:0] p5_sel_149618_comb;
  wire [14:0] p5_sel_149621_comb;
  wire [13:0] p5_sel_149624_comb;
  wire [13:0] p5_sel_149627_comb;
  wire [14:0] p5_sel_149630_comb;
  wire [14:0] p5_sel_149633_comb;
  wire [13:0] p5_sel_149636_comb;
  wire [23:0] p5_bit_slice_149637_comb;
  wire [13:0] p5_sel_149644_comb;
  wire [13:0] p5_sel_149647_comb;
  wire [23:0] p5_bit_slice_149652_comb;
  wire [23:0] p5_bit_slice_149653_comb;
  wire [23:0] p5_bit_slice_149658_comb;
  wire [23:0] p5_bit_slice_149659_comb;
  wire [23:0] p5_bit_slice_149664_comb;
  wire [23:0] p5_bit_slice_149665_comb;
  wire [13:0] p5_sel_149672_comb;
  wire [13:0] p5_sel_149675_comb;
  wire [23:0] p5_bit_slice_149680_comb;
  wire [13:0] p5_sel_149683_comb;
  wire [14:0] p5_sel_149686_comb;
  wire [14:0] p5_sel_149689_comb;
  wire [13:0] p5_sel_149692_comb;
  wire [13:0] p5_sel_149695_comb;
  wire [14:0] p5_sel_149698_comb;
  wire [14:0] p5_sel_149701_comb;
  wire [13:0] p5_sel_149704_comb;
  wire [23:0] p5_bit_slice_149705_comb;
  wire [13:0] p5_sel_149712_comb;
  wire [13:0] p5_sel_149715_comb;
  wire [23:0] p5_bit_slice_149720_comb;
  wire [23:0] p5_bit_slice_149721_comb;
  wire [23:0] p5_bit_slice_149726_comb;
  wire [23:0] p5_bit_slice_149727_comb;
  wire [23:0] p5_bit_slice_149732_comb;
  wire [23:0] p5_bit_slice_149733_comb;
  wire [13:0] p5_sel_149740_comb;
  wire [13:0] p5_sel_149743_comb;
  wire [23:0] p5_bit_slice_149748_comb;
  wire [14:0] p5_bit_slice_149751_comb;
  wire [14:0] p5_sel_149754_comb;
  wire [14:0] p5_sel_149757_comb;
  wire [14:0] p5_bit_slice_149760_comb;
  wire [14:0] p5_sel_149763_comb;
  wire [14:0] p5_sel_149766_comb;
  wire [14:0] p5_sel_149769_comb;
  wire [14:0] p5_sel_149772_comb;
  wire [14:0] p5_sel_149779_comb;
  wire [14:0] p5_sel_149782_comb;
  wire [14:0] p5_sel_149789_comb;
  wire [14:0] p5_sel_149792_comb;
  wire [14:0] p5_sel_149795_comb;
  wire [14:0] p5_sel_149798_comb;
  wire [14:0] p5_sel_149801_comb;
  wire [14:0] p5_bit_slice_149804_comb;
  wire [14:0] p5_bit_slice_149807_comb;
  wire [14:0] p5_sel_149810_comb;
  wire [14:0] p5_sel_149813_comb;
  wire [14:0] p5_sel_149824_comb;
  wire [14:0] p5_sel_149827_comb;
  wire [13:0] p5_sel_149830_comb;
  wire [14:0] p5_sel_149833_comb;
  wire [13:0] p5_sel_149836_comb;
  wire [13:0] p5_sel_149839_comb;
  wire [14:0] p5_sel_149842_comb;
  wire [13:0] p5_sel_149845_comb;
  wire [14:0] p5_sel_149848_comb;
  wire [23:0] p5_bit_slice_149851_comb;
  wire [13:0] p5_sel_149856_comb;
  wire [13:0] p5_sel_149859_comb;
  wire [23:0] p5_bit_slice_149862_comb;
  wire [23:0] p5_bit_slice_149867_comb;
  wire [23:0] p5_bit_slice_149870_comb;
  wire [23:0] p5_bit_slice_149871_comb;
  wire [23:0] p5_bit_slice_149874_comb;
  wire [23:0] p5_bit_slice_149879_comb;
  wire [13:0] p5_sel_149884_comb;
  wire [13:0] p5_sel_149887_comb;
  wire [23:0] p5_bit_slice_149890_comb;
  wire [14:0] p5_sel_149895_comb;
  wire [13:0] p5_sel_149898_comb;
  wire [14:0] p5_sel_149901_comb;
  wire [13:0] p5_sel_149904_comb;
  wire [13:0] p5_sel_149907_comb;
  wire [14:0] p5_sel_149910_comb;
  wire [13:0] p5_sel_149913_comb;
  wire [14:0] p5_sel_149916_comb;
  wire [23:0] p5_bit_slice_149919_comb;
  wire [13:0] p5_sel_149924_comb;
  wire [13:0] p5_sel_149927_comb;
  wire [23:0] p5_bit_slice_149930_comb;
  wire [23:0] p5_bit_slice_149935_comb;
  wire [23:0] p5_bit_slice_149938_comb;
  wire [23:0] p5_bit_slice_149939_comb;
  wire [23:0] p5_bit_slice_149942_comb;
  wire [23:0] p5_bit_slice_149947_comb;
  wire [13:0] p5_sel_149952_comb;
  wire [13:0] p5_sel_149955_comb;
  wire [23:0] p5_bit_slice_149958_comb;
  wire [14:0] p5_bit_slice_149963_comb;
  wire [14:0] p5_sel_149966_comb;
  wire [14:0] p5_sel_149969_comb;
  wire [14:0] p5_bit_slice_149972_comb;
  wire [14:0] p5_sel_149979_comb;
  wire [14:0] p5_sel_149982_comb;
  wire p5_sgt_150003_comb;
  wire p5_sgt_150004_comb;
  wire p5_sgt_150005_comb;
  wire p5_sgt_150006_comb;
  wire p5_sgt_150007_comb;
  wire p5_sgt_150008_comb;
  wire p5_sgt_150009_comb;
  wire p5_sgt_150010_comb;
  wire p5_sgt_150011_comb;
  wire p5_sgt_150018_comb;
  wire p5_sgt_150019_comb;
  wire p5_sgt_150020_comb;
  wire p5_sgt_150021_comb;
  wire p5_sgt_150022_comb;
  wire p5_sgt_150023_comb;
  wire p5_sgt_150024_comb;
  wire p5_sgt_150025_comb;
  wire p5_sgt_150026_comb;
  wire p5_sgt_150027_comb;
  wire p5_sgt_150028_comb;
  wire p5_sgt_150029_comb;
  wire p5_sgt_150030_comb;
  wire p5_sgt_150031_comb;
  wire p5_sgt_150032_comb;
  wire p5_sgt_150033_comb;
  wire p5_sgt_150034_comb;
  wire p5_sgt_150035_comb;
  wire p5_sgt_150036_comb;
  wire p5_sgt_150037_comb;
  wire p5_sgt_150038_comb;
  wire p5_sgt_150039_comb;
  wire p5_sgt_150040_comb;
  wire p5_sgt_150041_comb;
  wire p5_sgt_150042_comb;
  wire p5_sgt_150043_comb;
  wire p5_sgt_150044_comb;
  wire p5_sgt_150045_comb;
  wire p5_sgt_150046_comb;
  wire p5_sgt_150047_comb;
  wire p5_sgt_150048_comb;
  wire p5_sgt_150049_comb;
  wire p5_sgt_150050_comb;
  wire p5_sgt_150051_comb;
  wire p5_sgt_150052_comb;
  wire p5_sgt_150053_comb;
  wire p5_sgt_150054_comb;
  wire p5_sgt_150055_comb;
  wire p5_sgt_150056_comb;
  wire p5_sgt_150057_comb;
  wire p5_sgt_150058_comb;
  wire p5_sgt_150059_comb;
  wire p5_sgt_150060_comb;
  wire p5_sgt_150061_comb;
  wire p5_sgt_150062_comb;
  wire p5_sgt_150063_comb;
  wire p5_sgt_150064_comb;
  wire p5_sgt_150065_comb;
  wire p5_sgt_150066_comb;
  wire p5_sgt_150067_comb;
  wire p5_sgt_150068_comb;
  wire p5_sgt_150069_comb;
  wire p5_sgt_150070_comb;
  wire p5_sgt_150071_comb;
  wire p5_sgt_150072_comb;
  wire p5_sgt_150073_comb;
  wire p5_sgt_150074_comb;
  wire p5_sgt_150075_comb;
  wire p5_sgt_150076_comb;
  wire p5_sgt_150077_comb;
  wire p5_sgt_150078_comb;
  wire p5_sgt_150082_comb;
  wire p5_sgt_150083_comb;
  wire p5_sgt_150087_comb;
  wire p5_sgt_150088_comb;
  wire p5_sgt_150089_comb;
  wire p5_sgt_150090_comb;
  wire p5_sgt_150091_comb;
  wire p5_sgt_150092_comb;
  wire p5_sgt_150093_comb;
  wire p5_sgt_150094_comb;
  wire p5_sgt_150095_comb;
  wire p5_sgt_150102_comb;
  wire p5_sgt_150103_comb;
  wire p5_sgt_150104_comb;
  wire p5_sgt_150105_comb;
  wire p5_sgt_150106_comb;
  wire p5_sgt_150107_comb;
  wire p5_sgt_150108_comb;
  wire p5_sgt_150109_comb;
  wire p5_sgt_150110_comb;
  wire p5_sgt_150111_comb;
  wire p5_sgt_150112_comb;
  wire p5_sgt_150113_comb;
  wire p5_sgt_150114_comb;
  wire p5_sgt_150115_comb;
  wire p5_sgt_150116_comb;
  wire p5_sgt_150117_comb;
  wire p5_sgt_150118_comb;
  wire p5_sgt_150119_comb;
  wire p5_sgt_150120_comb;
  wire p5_sgt_150121_comb;
  wire p5_sgt_150122_comb;
  wire p5_sgt_150123_comb;
  wire p5_sgt_150124_comb;
  wire p5_sgt_150125_comb;
  wire p5_sgt_150126_comb;
  wire p5_sgt_150127_comb;
  wire p5_sgt_150128_comb;
  wire p5_sgt_150129_comb;
  wire p5_sgt_150130_comb;
  wire p5_sgt_150131_comb;
  wire p5_sgt_150132_comb;
  wire p5_sgt_150133_comb;
  wire p5_sgt_150134_comb;
  wire p5_sgt_150135_comb;
  wire p5_sgt_150136_comb;
  wire p5_sgt_150137_comb;
  wire p5_sgt_150138_comb;
  wire p5_sgt_150139_comb;
  wire p5_sgt_150140_comb;
  wire p5_sgt_150141_comb;
  wire p5_sgt_150142_comb;
  wire p5_sgt_150143_comb;
  wire p5_sgt_150144_comb;
  wire p5_sgt_150145_comb;
  wire p5_sgt_150146_comb;
  wire p5_sgt_150147_comb;
  wire p5_sgt_150148_comb;
  wire p5_sgt_150149_comb;
  wire p5_sgt_150150_comb;
  wire p5_sgt_150151_comb;
  wire p5_sgt_150152_comb;
  wire p5_sgt_150153_comb;
  wire p5_sgt_150154_comb;
  wire p5_sgt_150158_comb;
  wire p5_sgt_150159_comb;
  wire [16:0] p5_add_150163_comb;
  wire [16:0] p5_add_150164_comb;
  wire [16:0] p5_add_150165_comb;
  wire [16:0] p5_add_150166_comb;
  wire [16:0] p5_add_150167_comb;
  wire [16:0] p5_add_150168_comb;
  wire [16:0] p5_add_150169_comb;
  wire [16:0] p5_add_150170_comb;
  wire [15:0] p5_sel_150171_comb;
  wire [15:0] p5_sel_150172_comb;
  wire [15:0] p5_sel_150173_comb;
  wire [15:0] p5_sel_150174_comb;
  wire [15:0] p5_sel_150175_comb;
  wire [15:0] p5_sel_150176_comb;
  wire [15:0] p5_sel_150177_comb;
  wire [15:0] p5_sel_150178_comb;
  assign p5_shifted__99_squeezed_comb = {p4_not_146199, p4_bit_slice_146200};
  assign p5_shifted__100_squeezed_comb = {p4_not_146201, p4_bit_slice_146202};
  assign p5_shifted__97_squeezed_comb = {p4_not_146197, p4_bit_slice_146198};
  assign p5_shifted__102_squeezed_comb = {p4_not_146203, p4_bit_slice_146204};
  assign p5_shifted__98_squeezed_comb = {p4_not_146181, p4_bit_slice_146182};
  assign p5_shifted__101_squeezed_comb = {p4_not_146183, p4_bit_slice_146184};
  assign p5_shifted__96_squeezed_comb = {p4_not_146195, p4_bit_slice_146196};
  assign p5_shifted__103_squeezed_comb = {p4_not_146205, p4_bit_slice_146206};
  assign p5_shifted__66_squeezed_comb = {~p4_bit_slice_146155, p4_bit_slice_146179};
  assign p5_shifted__69_squeezed_comb = {~p4_bit_slice_146156, p4_bit_slice_146180};
  assign p5_shifted__64_squeezed_comb = {~p4_bit_slice_146159, p4_bit_slice_146185};
  assign p5_shifted__65_squeezed_comb = {~p4_bit_slice_146160, p4_bit_slice_146186};
  assign p5_shifted__67_squeezed_comb = {~p4_bit_slice_146161, p4_bit_slice_146187};
  assign p5_shifted__68_squeezed_comb = {~p4_bit_slice_146162, p4_bit_slice_146188};
  assign p5_shifted__70_squeezed_comb = {~p4_bit_slice_146163, p4_bit_slice_146189};
  assign p5_shifted__71_squeezed_comb = {~p4_bit_slice_146164, p4_bit_slice_146190};
  assign p5_shifted__75_squeezed_comb = {~p4_bit_slice_146165, p4_bit_slice_146191};
  assign p5_shifted__76_squeezed_comb = {~p4_bit_slice_146166, p4_bit_slice_146192};
  assign p5_shifted__91_squeezed_comb = {~p4_bit_slice_146167, p4_bit_slice_146193};
  assign p5_shifted__92_squeezed_comb = {~p4_bit_slice_146168, p4_bit_slice_146194};
  assign p5_shifted__107_squeezed_comb = {~p4_bit_slice_146175, p4_bit_slice_146207};
  assign p5_shifted__108_squeezed_comb = {~p4_bit_slice_146176, p4_bit_slice_146208};
  assign p5_shifted__123_squeezed_comb = {~p4_bit_slice_146177, p4_bit_slice_146209};
  assign p5_shifted__124_squeezed_comb = {~p4_bit_slice_146178, p4_bit_slice_146210};
  assign p5_smul_58292_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__99_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___209_comb = 9'h000;
  assign p5_smul_58294_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__100_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___210_comb = 9'h000;
  assign p5_smul_58544_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__97_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___272_comb = 9'h000;
  assign p5_smul_58554_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__102_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___275_comb = 9'h000;
  assign p5_smul_58802_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__98_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___305_comb = 9'h000;
  assign p5_smul_58808_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__101_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___306_comb = 9'h000;
  assign p5_smul_59054_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__96_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___368_comb = 9'h000;
  assign p5_smul_59068_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__103_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___371_comb = 9'h000;
  assign p5_shifted__74_squeezed_comb = {~p4_clipped__41[7], p4_clipped__41[6:0]};
  assign p5_shifted__77_squeezed_comb = {~p4_clipped__89[7], p4_clipped__89[6:0]};
  assign p5_shifted__82_squeezed_comb = {~p4_clipped__42[7], p4_clipped__42[6:0]};
  assign p5_shifted__85_squeezed_comb = {~p4_clipped__90[7], p4_clipped__90[6:0]};
  assign p5_shifted__90_squeezed_comb = {~p4_clipped__43[7], p4_clipped__43[6:0]};
  assign p5_shifted__93_squeezed_comb = {~p4_clipped__91[7], p4_clipped__91[6:0]};
  assign p5_shifted__106_squeezed_comb = {~p4_clipped__45[7], p4_clipped__45[6:0]};
  assign p5_shifted__109_squeezed_comb = {~p4_clipped__93[7], p4_clipped__93[6:0]};
  assign p5_shifted__114_squeezed_comb = {~p4_clipped__46[7], p4_clipped__46[6:0]};
  assign p5_shifted__117_squeezed_comb = {~p4_clipped__94[7], p4_clipped__94[6:0]};
  assign p5_shifted__122_squeezed_comb = {~p4_clipped__47[7], p4_clipped__47[6:0]};
  assign p5_shifted__125_squeezed_comb = {~p4_clipped__95[7], p4_clipped__95[6:0]};
  assign p5_shifted__72_squeezed_comb = {~p4_clipped__9[7], p4_clipped__9[6:0]};
  assign p5_shifted__73_squeezed_comb = {~p4_clipped__25[7], p4_clipped__25[6:0]};
  assign p5_shifted__78_squeezed_comb = {~p4_clipped__105[7], p4_clipped__105[6:0]};
  assign p5_shifted__79_squeezed_comb = {~p4_clipped__121[7], p4_clipped__121[6:0]};
  assign p5_shifted__80_squeezed_comb = {~p4_clipped__10[7], p4_clipped__10[6:0]};
  assign p5_shifted__81_squeezed_comb = {~p4_clipped__26[7], p4_clipped__26[6:0]};
  assign p5_shifted__83_squeezed_comb = {~p4_clipped__58[7], p4_clipped__58[6:0]};
  assign p5_shifted__84_squeezed_comb = {~p4_clipped__74[7], p4_clipped__74[6:0]};
  assign p5_shifted__86_squeezed_comb = {~p4_clipped__106[7], p4_clipped__106[6:0]};
  assign p5_shifted__87_squeezed_comb = {~p4_clipped__122[7], p4_clipped__122[6:0]};
  assign p5_shifted__88_squeezed_comb = {~p4_clipped__11[7], p4_clipped__11[6:0]};
  assign p5_shifted__89_squeezed_comb = {~p4_clipped__27[7], p4_clipped__27[6:0]};
  assign p5_shifted__94_squeezed_comb = {~p4_clipped__107[7], p4_clipped__107[6:0]};
  assign p5_shifted__95_squeezed_comb = {~p4_clipped__123[7], p4_clipped__123[6:0]};
  assign p5_shifted__104_squeezed_comb = {~p4_clipped__13[7], p4_clipped__13[6:0]};
  assign p5_shifted__105_squeezed_comb = {~p4_clipped__29[7], p4_clipped__29[6:0]};
  assign p5_shifted__110_squeezed_comb = {~p4_clipped__109[7], p4_clipped__109[6:0]};
  assign p5_shifted__111_squeezed_comb = {~p4_clipped__125[7], p4_clipped__125[6:0]};
  assign p5_shifted__112_squeezed_comb = {~p4_clipped__14[7], p4_clipped__14[6:0]};
  assign p5_shifted__113_squeezed_comb = {~p4_clipped__30[7], p4_clipped__30[6:0]};
  assign p5_shifted__115_squeezed_comb = {~p4_clipped__62[7], p4_clipped__62[6:0]};
  assign p5_shifted__116_squeezed_comb = {~p4_clipped__78[7], p4_clipped__78[6:0]};
  assign p5_shifted__118_squeezed_comb = {~p4_clipped__110[7], p4_clipped__110[6:0]};
  assign p5_shifted__119_squeezed_comb = {~p4_clipped__126[7], p4_clipped__126[6:0]};
  assign p5_shifted__120_squeezed_comb = {~p4_clipped__15[7], p4_clipped__15[6:0]};
  assign p5_shifted__121_squeezed_comb = {~p4_clipped__31[7], p4_clipped__31[6:0]};
  assign p5_shifted__126_squeezed_comb = {~p4_clipped__111[7], p4_clipped__111[6:0]};
  assign p5_shifted__127_squeezed_comb = {~p4_clipped__127[7], p4_clipped__127[6:0]};
  assign p5_smul_58226_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__66_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___192_comb = 9'h000;
  assign p5_smul_58232_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__69_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___195_comb = 9'h000;
  assign p5_smul_58290_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__98_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___208_comb = 9'h000;
  assign p5_smul_58296_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__101_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___211_comb = 9'h000;
  assign p5_smul_58350_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__64_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___64_comb = 10'h000;
  assign p5_smul_58352_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__65_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___224_comb = 9'h000;
  assign p5_smul_58354_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__66_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___225_comb = 9'h000;
  assign p5_smul_58356_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__67_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___65_comb = 10'h000;
  assign p5_smul_58358_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__68_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___66_comb = 10'h000;
  assign p5_smul_58360_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__69_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___226_comb = 9'h000;
  assign p5_smul_58362_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__70_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___227_comb = 9'h000;
  assign p5_smul_58364_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__71_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___67_comb = 10'h000;
  assign p5_smul_58372_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__75_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___69_comb = 10'h000;
  assign p5_smul_58374_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__76_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___70_comb = 10'h000;
  assign p5_smul_58404_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__91_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___77_comb = 10'h000;
  assign p5_smul_58406_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__92_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___78_comb = 10'h000;
  assign p5_smul_58414_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__96_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___80_comb = 10'h000;
  assign p5_smul_58416_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__97_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___240_comb = 9'h000;
  assign p5_smul_58418_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__98_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___241_comb = 9'h000;
  assign p5_smul_58420_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__99_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___81_comb = 10'h000;
  assign p5_smul_58422_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__100_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___82_comb = 10'h000;
  assign p5_smul_58424_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__101_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___242_comb = 9'h000;
  assign p5_smul_58426_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__102_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___243_comb = 9'h000;
  assign p5_smul_58428_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__103_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___83_comb = 10'h000;
  assign p5_smul_58436_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__107_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___85_comb = 10'h000;
  assign p5_smul_58438_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__108_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___86_comb = 10'h000;
  assign p5_smul_58468_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__123_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___93_comb = 10'h000;
  assign p5_smul_58470_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__124_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___94_comb = 10'h000;
  assign p5_smul_58484_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__67_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___257_comb = 9'h000;
  assign p5_smul_58486_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__68_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___258_comb = 9'h000;
  assign p5_smul_58500_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__75_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___261_comb = 9'h000;
  assign p5_smul_58502_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__76_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___262_comb = 9'h000;
  assign p5_smul_58532_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__91_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___269_comb = 9'h000;
  assign p5_smul_58534_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__92_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___270_comb = 9'h000;
  assign p5_smul_58548_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__99_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___273_comb = 9'h000;
  assign p5_smul_58550_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__100_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___274_comb = 9'h000;
  assign p5_smul_58564_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__107_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___277_comb = 9'h000;
  assign p5_smul_58566_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__108_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___278_comb = 9'h000;
  assign p5_smul_58596_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__123_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___285_comb = 9'h000;
  assign p5_smul_58598_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__124_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___286_comb = 9'h000;
  assign p5_smul_58734_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__64_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___288_comb = 9'h000;
  assign p5_smul_58748_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__71_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___291_comb = 9'h000;
  assign p5_smul_58798_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__96_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___304_comb = 9'h000;
  assign p5_smul_58812_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__103_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___307_comb = 9'h000;
  assign p5_smul_58862_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__64_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___320_comb = 9'h000;
  assign p5_smul_58864_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__65_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___96_comb = 10'h000;
  assign p5_smul_58866_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__66_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___321_comb = 9'h000;
  assign p5_smul_58868_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__67_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___97_comb = 10'h000;
  assign p5_smul_58870_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__68_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___98_comb = 10'h000;
  assign p5_smul_58872_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__69_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___322_comb = 9'h000;
  assign p5_smul_58874_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__70_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___99_comb = 10'h000;
  assign p5_smul_58876_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__71_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___323_comb = 9'h000;
  assign p5_smul_58884_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__75_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___101_comb = 10'h000;
  assign p5_smul_58886_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__76_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___102_comb = 10'h000;
  assign p5_smul_58916_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__91_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___109_comb = 10'h000;
  assign p5_smul_58918_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__92_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___110_comb = 10'h000;
  assign p5_smul_58926_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__96_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___336_comb = 9'h000;
  assign p5_smul_58928_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__97_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___112_comb = 10'h000;
  assign p5_smul_58930_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__98_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___337_comb = 9'h000;
  assign p5_smul_58932_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__99_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___113_comb = 10'h000;
  assign p5_smul_58934_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__100_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___114_comb = 10'h000;
  assign p5_smul_58936_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__101_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___338_comb = 9'h000;
  assign p5_smul_58938_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__102_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___115_comb = 10'h000;
  assign p5_smul_58940_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__103_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___339_comb = 9'h000;
  assign p5_smul_58948_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__107_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___117_comb = 10'h000;
  assign p5_smul_58950_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__108_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___118_comb = 10'h000;
  assign p5_smul_58980_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__123_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___125_comb = 10'h000;
  assign p5_smul_58982_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__124_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___126_comb = 10'h000;
  assign p5_smul_58992_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__65_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___353_comb = 9'h000;
  assign p5_smul_59002_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__70_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___354_comb = 9'h000;
  assign p5_smul_59056_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__97_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___369_comb = 9'h000;
  assign p5_smul_59066_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__102_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___370_comb = 9'h000;
  assign p5_smul_58228_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__67_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___193_comb = 9'h000;
  assign p5_smul_58230_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__68_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___194_comb = 9'h000;
  assign p5_smul_58244_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__75_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___197_comb = 9'h000;
  assign p5_smul_58246_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__76_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___198_comb = 9'h000;
  assign p5_smul_58276_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__91_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___205_comb = 9'h000;
  assign p5_smul_58278_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__92_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___206_comb = 9'h000;
  assign p5_smul_58308_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__107_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___213_comb = 9'h000;
  assign p5_smul_58310_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__108_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___214_comb = 9'h000;
  assign p5_smul_58340_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__123_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___221_comb = 9'h000;
  assign p5_smul_58342_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__124_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___222_comb = 9'h000;
  assign p5_smul_58480_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__65_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___256_comb = 9'h000;
  assign p5_smul_58490_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__70_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___259_comb = 9'h000;
  assign p5_smul_58738_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__66_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___289_comb = 9'h000;
  assign p5_smul_58744_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__69_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___290_comb = 9'h000;
  assign p5_smul_58990_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__64_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___352_comb = 9'h000;
  assign p5_smul_59004_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__71_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___355_comb = 9'h000;
  assign p5_smul_57326_TrailingBits___192_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___193_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___194_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___195_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___196_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___197_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___198_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___199_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___224_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___225_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___226_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___227_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___228_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___229_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___230_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___231_comb = 8'h00;
  assign p5_concat_147829_comb = {p5_smul_58292_NarrowedMult__comb, p5_smul_57330_TrailingBits___209_comb};
  assign p5_concat_147830_comb = {p5_smul_58294_NarrowedMult__comb, p5_smul_57330_TrailingBits___210_comb};
  assign p5_concat_147971_comb = {p5_smul_58544_NarrowedMult__comb, p5_smul_57330_TrailingBits___272_comb};
  assign p5_concat_147976_comb = {p5_smul_58554_NarrowedMult__comb, p5_smul_57330_TrailingBits___275_comb};
  assign p5_concat_148021_comb = {p5_smul_58802_NarrowedMult__comb, p5_smul_57330_TrailingBits___305_comb};
  assign p5_concat_148022_comb = {p5_smul_58808_NarrowedMult__comb, p5_smul_57330_TrailingBits___306_comb};
  assign p5_concat_148163_comb = {p5_smul_59054_NarrowedMult__comb, p5_smul_57330_TrailingBits___368_comb};
  assign p5_concat_148168_comb = {p5_smul_59068_NarrowedMult__comb, p5_smul_57330_TrailingBits___371_comb};
  assign p5_smul_58242_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__74_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___196_comb = 9'h000;
  assign p5_smul_58248_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__77_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___199_comb = 9'h000;
  assign p5_smul_58258_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__82_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___200_comb = 9'h000;
  assign p5_smul_58264_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__85_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___203_comb = 9'h000;
  assign p5_smul_58274_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__90_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___204_comb = 9'h000;
  assign p5_smul_58280_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__93_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___207_comb = 9'h000;
  assign p5_smul_58306_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__106_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___212_comb = 9'h000;
  assign p5_smul_58312_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__109_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___215_comb = 9'h000;
  assign p5_smul_58322_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__114_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___216_comb = 9'h000;
  assign p5_smul_58328_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__117_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___219_comb = 9'h000;
  assign p5_smul_58338_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__122_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___220_comb = 9'h000;
  assign p5_smul_58344_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__125_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___223_comb = 9'h000;
  assign p5_smul_58366_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__72_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___68_comb = 10'h000;
  assign p5_smul_58368_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__73_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___228_comb = 9'h000;
  assign p5_smul_58370_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__74_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___229_comb = 9'h000;
  assign p5_smul_58376_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__77_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___230_comb = 9'h000;
  assign p5_smul_58378_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__78_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___231_comb = 9'h000;
  assign p5_smul_58380_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__79_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___71_comb = 10'h000;
  assign p5_smul_58382_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__80_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___72_comb = 10'h000;
  assign p5_smul_58384_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__81_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___232_comb = 9'h000;
  assign p5_smul_58386_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__82_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___233_comb = 9'h000;
  assign p5_smul_58388_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__83_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___73_comb = 10'h000;
  assign p5_smul_58390_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__84_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___74_comb = 10'h000;
  assign p5_smul_58392_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__85_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___234_comb = 9'h000;
  assign p5_smul_58394_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__86_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___235_comb = 9'h000;
  assign p5_smul_58396_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__87_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___75_comb = 10'h000;
  assign p5_smul_58398_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__88_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___76_comb = 10'h000;
  assign p5_smul_58400_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__89_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___236_comb = 9'h000;
  assign p5_smul_58402_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__90_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___237_comb = 9'h000;
  assign p5_smul_58408_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__93_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___238_comb = 9'h000;
  assign p5_smul_58410_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__94_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___239_comb = 9'h000;
  assign p5_smul_58412_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__95_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___79_comb = 10'h000;
  assign p5_smul_58430_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__104_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___84_comb = 10'h000;
  assign p5_smul_58432_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__105_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___244_comb = 9'h000;
  assign p5_smul_58434_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__106_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___245_comb = 9'h000;
  assign p5_smul_58440_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__109_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___246_comb = 9'h000;
  assign p5_smul_58442_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__110_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___247_comb = 9'h000;
  assign p5_smul_58444_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__111_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___87_comb = 10'h000;
  assign p5_smul_58446_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__112_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___88_comb = 10'h000;
  assign p5_smul_58448_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__113_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___248_comb = 9'h000;
  assign p5_smul_58450_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__114_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___249_comb = 9'h000;
  assign p5_smul_58452_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__115_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___89_comb = 10'h000;
  assign p5_smul_58454_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__116_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___90_comb = 10'h000;
  assign p5_smul_58456_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__117_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___250_comb = 9'h000;
  assign p5_smul_58458_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__118_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___251_comb = 9'h000;
  assign p5_smul_58460_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__119_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___91_comb = 10'h000;
  assign p5_smul_58462_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__120_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___92_comb = 10'h000;
  assign p5_smul_58464_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__121_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___252_comb = 9'h000;
  assign p5_smul_58466_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__122_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___253_comb = 9'h000;
  assign p5_smul_58472_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__125_squeezed_comb, 7'h4f);
  assign p5_smul_57330_TrailingBits___254_comb = 9'h000;
  assign p5_smul_58474_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__126_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___255_comb = 9'h000;
  assign p5_smul_58476_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__127_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___95_comb = 10'h000;
  assign p5_smul_58516_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__83_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___265_comb = 9'h000;
  assign p5_smul_58518_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__84_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___266_comb = 9'h000;
  assign p5_smul_58580_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__115_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___281_comb = 9'h000;
  assign p5_smul_58582_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__116_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___282_comb = 9'h000;
  assign p5_smul_58750_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__72_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___292_comb = 9'h000;
  assign p5_smul_58764_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__79_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___295_comb = 9'h000;
  assign p5_smul_58766_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__80_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___296_comb = 9'h000;
  assign p5_smul_58780_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__87_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___299_comb = 9'h000;
  assign p5_smul_58782_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__88_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___300_comb = 9'h000;
  assign p5_smul_58796_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__95_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___303_comb = 9'h000;
  assign p5_smul_58814_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__104_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___308_comb = 9'h000;
  assign p5_smul_58828_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__111_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___311_comb = 9'h000;
  assign p5_smul_58830_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__112_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___312_comb = 9'h000;
  assign p5_smul_58844_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__119_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___315_comb = 9'h000;
  assign p5_smul_58846_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__120_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___316_comb = 9'h000;
  assign p5_smul_58860_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__127_squeezed_comb, 8'h47);
  assign p5_smul_57330_TrailingBits___319_comb = 9'h000;
  assign p5_smul_58878_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__72_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___324_comb = 9'h000;
  assign p5_smul_58880_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__73_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___100_comb = 10'h000;
  assign p5_smul_58882_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__74_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___325_comb = 9'h000;
  assign p5_smul_58888_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__77_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___326_comb = 9'h000;
  assign p5_smul_58890_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__78_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___103_comb = 10'h000;
  assign p5_smul_58892_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__79_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___327_comb = 9'h000;
  assign p5_smul_58894_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__80_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___328_comb = 9'h000;
  assign p5_smul_58896_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__81_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___104_comb = 10'h000;
  assign p5_smul_58898_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__82_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___329_comb = 9'h000;
  assign p5_smul_58900_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__83_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___105_comb = 10'h000;
  assign p5_smul_58902_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__84_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___106_comb = 10'h000;
  assign p5_smul_58904_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__85_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___330_comb = 9'h000;
  assign p5_smul_58906_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__86_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___107_comb = 10'h000;
  assign p5_smul_58908_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__87_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___331_comb = 9'h000;
  assign p5_smul_58910_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__88_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___332_comb = 9'h000;
  assign p5_smul_58912_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__89_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___108_comb = 10'h000;
  assign p5_smul_58914_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__90_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___333_comb = 9'h000;
  assign p5_smul_58920_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__93_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___334_comb = 9'h000;
  assign p5_smul_58922_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__94_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___111_comb = 10'h000;
  assign p5_smul_58924_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__95_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___335_comb = 9'h000;
  assign p5_smul_58942_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__104_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___340_comb = 9'h000;
  assign p5_smul_58944_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__105_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___116_comb = 10'h000;
  assign p5_smul_58946_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__106_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___341_comb = 9'h000;
  assign p5_smul_58952_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__109_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___342_comb = 9'h000;
  assign p5_smul_58954_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__110_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___119_comb = 10'h000;
  assign p5_smul_58956_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__111_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___343_comb = 9'h000;
  assign p5_smul_58958_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__112_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___344_comb = 9'h000;
  assign p5_smul_58960_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__113_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___120_comb = 10'h000;
  assign p5_smul_58962_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__114_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___345_comb = 9'h000;
  assign p5_smul_58964_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__115_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___121_comb = 10'h000;
  assign p5_smul_58966_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__116_squeezed_comb, 7'h3b);
  assign p5_smul_57454_TrailingBits___122_comb = 10'h000;
  assign p5_smul_58968_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__117_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___346_comb = 9'h000;
  assign p5_smul_58970_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__118_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___123_comb = 10'h000;
  assign p5_smul_58972_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__119_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___347_comb = 9'h000;
  assign p5_smul_58974_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__120_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___348_comb = 9'h000;
  assign p5_smul_58976_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__121_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___124_comb = 10'h000;
  assign p5_smul_58978_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__122_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___349_comb = 9'h000;
  assign p5_smul_58984_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__125_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___350_comb = 9'h000;
  assign p5_smul_58986_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__126_squeezed_comb, 7'h45);
  assign p5_smul_57454_TrailingBits___127_comb = 10'h000;
  assign p5_smul_58988_NarrowedMult__comb = smul15b_8b_x_7b(p5_shifted__127_squeezed_comb, 7'h31);
  assign p5_smul_57330_TrailingBits___351_comb = 9'h000;
  assign p5_smul_59008_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__73_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___357_comb = 9'h000;
  assign p5_smul_59018_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__78_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___358_comb = 9'h000;
  assign p5_smul_59024_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__81_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___361_comb = 9'h000;
  assign p5_smul_59034_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__86_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___362_comb = 9'h000;
  assign p5_smul_59040_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__89_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___365_comb = 9'h000;
  assign p5_smul_59050_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__94_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___366_comb = 9'h000;
  assign p5_smul_59072_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__105_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___373_comb = 9'h000;
  assign p5_smul_59082_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__110_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___374_comb = 9'h000;
  assign p5_smul_59088_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__113_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___377_comb = 9'h000;
  assign p5_smul_59098_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__118_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___378_comb = 9'h000;
  assign p5_smul_59104_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__121_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___381_comb = 9'h000;
  assign p5_smul_59114_NarrowedMult__comb = smul16b_8b_x_8b(p5_shifted__126_squeezed_comb, 8'hb9);
  assign p5_smul_57330_TrailingBits___382_comb = 9'h000;
  assign p5_concat_147291_comb = {p5_smul_58226_NarrowedMult__comb, p5_smul_57330_TrailingBits___192_comb};
  assign p5_concat_147296_comb = {p5_smul_58232_NarrowedMult__comb, p5_smul_57330_TrailingBits___195_comb};
  assign p5_concat_147315_comb = {p5_smul_58290_NarrowedMult__comb, p5_smul_57330_TrailingBits___208_comb};
  assign p5_concat_147320_comb = {p5_smul_58296_NarrowedMult__comb, p5_smul_57330_TrailingBits___211_comb};
  assign p5_concat_147339_comb = {p5_smul_58350_NarrowedMult__comb, p5_smul_57454_TrailingBits___64_comb};
  assign p5_concat_147340_comb = {p5_smul_58352_NarrowedMult__comb, p5_smul_57330_TrailingBits___224_comb};
  assign p5_concat_147341_comb = {p5_smul_58354_NarrowedMult__comb, p5_smul_57330_TrailingBits___225_comb};
  assign p5_concat_147342_comb = {p5_smul_58356_NarrowedMult__comb, p5_smul_57454_TrailingBits___65_comb};
  assign p5_concat_147343_comb = {p5_smul_58358_NarrowedMult__comb, p5_smul_57454_TrailingBits___66_comb};
  assign p5_concat_147344_comb = {p5_smul_58360_NarrowedMult__comb, p5_smul_57330_TrailingBits___226_comb};
  assign p5_concat_147345_comb = {p5_smul_58362_NarrowedMult__comb, p5_smul_57330_TrailingBits___227_comb};
  assign p5_concat_147346_comb = {p5_smul_58364_NarrowedMult__comb, p5_smul_57454_TrailingBits___67_comb};
  assign p5_concat_147350_comb = {p5_smul_58372_NarrowedMult__comb, p5_smul_57454_TrailingBits___69_comb};
  assign p5_concat_147351_comb = {p5_smul_58374_NarrowedMult__comb, p5_smul_57454_TrailingBits___70_comb};
  assign p5_concat_147366_comb = {p5_smul_58404_NarrowedMult__comb, p5_smul_57454_TrailingBits___77_comb};
  assign p5_concat_147367_comb = {p5_smul_58406_NarrowedMult__comb, p5_smul_57454_TrailingBits___78_comb};
  assign p5_concat_147371_comb = {p5_smul_58414_NarrowedMult__comb, p5_smul_57454_TrailingBits___80_comb};
  assign p5_concat_147372_comb = {p5_smul_58416_NarrowedMult__comb, p5_smul_57330_TrailingBits___240_comb};
  assign p5_concat_147373_comb = {p5_smul_58418_NarrowedMult__comb, p5_smul_57330_TrailingBits___241_comb};
  assign p5_concat_147374_comb = {p5_smul_58420_NarrowedMult__comb, p5_smul_57454_TrailingBits___81_comb};
  assign p5_concat_147375_comb = {p5_smul_58422_NarrowedMult__comb, p5_smul_57454_TrailingBits___82_comb};
  assign p5_concat_147376_comb = {p5_smul_58424_NarrowedMult__comb, p5_smul_57330_TrailingBits___242_comb};
  assign p5_concat_147377_comb = {p5_smul_58426_NarrowedMult__comb, p5_smul_57330_TrailingBits___243_comb};
  assign p5_concat_147378_comb = {p5_smul_58428_NarrowedMult__comb, p5_smul_57454_TrailingBits___83_comb};
  assign p5_concat_147382_comb = {p5_smul_58436_NarrowedMult__comb, p5_smul_57454_TrailingBits___85_comb};
  assign p5_concat_147383_comb = {p5_smul_58438_NarrowedMult__comb, p5_smul_57454_TrailingBits___86_comb};
  assign p5_concat_147398_comb = {p5_smul_58468_NarrowedMult__comb, p5_smul_57454_TrailingBits___93_comb};
  assign p5_concat_147399_comb = {p5_smul_58470_NarrowedMult__comb, p5_smul_57454_TrailingBits___94_comb};
  assign p5_concat_147405_comb = {p5_smul_58484_NarrowedMult__comb, p5_smul_57330_TrailingBits___257_comb};
  assign p5_concat_147406_comb = {p5_smul_58486_NarrowedMult__comb, p5_smul_57330_TrailingBits___258_comb};
  assign p5_concat_147411_comb = {p5_smul_58500_NarrowedMult__comb, p5_smul_57330_TrailingBits___261_comb};
  assign p5_concat_147412_comb = {p5_smul_58502_NarrowedMult__comb, p5_smul_57330_TrailingBits___262_comb};
  assign p5_concat_147423_comb = {p5_smul_58532_NarrowedMult__comb, p5_smul_57330_TrailingBits___269_comb};
  assign p5_concat_147424_comb = {p5_smul_58534_NarrowedMult__comb, p5_smul_57330_TrailingBits___270_comb};
  assign p5_concat_147429_comb = {p5_smul_58548_NarrowedMult__comb, p5_smul_57330_TrailingBits___273_comb};
  assign p5_concat_147430_comb = {p5_smul_58550_NarrowedMult__comb, p5_smul_57330_TrailingBits___274_comb};
  assign p5_concat_147435_comb = {p5_smul_58564_NarrowedMult__comb, p5_smul_57330_TrailingBits___277_comb};
  assign p5_concat_147436_comb = {p5_smul_58566_NarrowedMult__comb, p5_smul_57330_TrailingBits___278_comb};
  assign p5_concat_147447_comb = {p5_smul_58596_NarrowedMult__comb, p5_smul_57330_TrailingBits___285_comb};
  assign p5_concat_147448_comb = {p5_smul_58598_NarrowedMult__comb, p5_smul_57330_TrailingBits___286_comb};
  assign p5_concat_147451_comb = {p5_smul_58734_NarrowedMult__comb, p5_smul_57330_TrailingBits___288_comb};
  assign p5_concat_147456_comb = {p5_smul_58748_NarrowedMult__comb, p5_smul_57330_TrailingBits___291_comb};
  assign p5_concat_147475_comb = {p5_smul_58798_NarrowedMult__comb, p5_smul_57330_TrailingBits___304_comb};
  assign p5_concat_147480_comb = {p5_smul_58812_NarrowedMult__comb, p5_smul_57330_TrailingBits___307_comb};
  assign p5_concat_147499_comb = {p5_smul_58862_NarrowedMult__comb, p5_smul_57330_TrailingBits___320_comb};
  assign p5_concat_147500_comb = {p5_smul_58864_NarrowedMult__comb, p5_smul_57454_TrailingBits___96_comb};
  assign p5_concat_147501_comb = {p5_smul_58866_NarrowedMult__comb, p5_smul_57330_TrailingBits___321_comb};
  assign p5_concat_147502_comb = {p5_smul_58868_NarrowedMult__comb, p5_smul_57454_TrailingBits___97_comb};
  assign p5_concat_147503_comb = {p5_smul_58870_NarrowedMult__comb, p5_smul_57454_TrailingBits___98_comb};
  assign p5_concat_147504_comb = {p5_smul_58872_NarrowedMult__comb, p5_smul_57330_TrailingBits___322_comb};
  assign p5_concat_147505_comb = {p5_smul_58874_NarrowedMult__comb, p5_smul_57454_TrailingBits___99_comb};
  assign p5_concat_147506_comb = {p5_smul_58876_NarrowedMult__comb, p5_smul_57330_TrailingBits___323_comb};
  assign p5_concat_147510_comb = {p5_smul_58884_NarrowedMult__comb, p5_smul_57454_TrailingBits___101_comb};
  assign p5_concat_147511_comb = {p5_smul_58886_NarrowedMult__comb, p5_smul_57454_TrailingBits___102_comb};
  assign p5_concat_147526_comb = {p5_smul_58916_NarrowedMult__comb, p5_smul_57454_TrailingBits___109_comb};
  assign p5_concat_147527_comb = {p5_smul_58918_NarrowedMult__comb, p5_smul_57454_TrailingBits___110_comb};
  assign p5_concat_147531_comb = {p5_smul_58926_NarrowedMult__comb, p5_smul_57330_TrailingBits___336_comb};
  assign p5_concat_147532_comb = {p5_smul_58928_NarrowedMult__comb, p5_smul_57454_TrailingBits___112_comb};
  assign p5_concat_147533_comb = {p5_smul_58930_NarrowedMult__comb, p5_smul_57330_TrailingBits___337_comb};
  assign p5_concat_147534_comb = {p5_smul_58932_NarrowedMult__comb, p5_smul_57454_TrailingBits___113_comb};
  assign p5_concat_147535_comb = {p5_smul_58934_NarrowedMult__comb, p5_smul_57454_TrailingBits___114_comb};
  assign p5_concat_147536_comb = {p5_smul_58936_NarrowedMult__comb, p5_smul_57330_TrailingBits___338_comb};
  assign p5_concat_147537_comb = {p5_smul_58938_NarrowedMult__comb, p5_smul_57454_TrailingBits___115_comb};
  assign p5_concat_147538_comb = {p5_smul_58940_NarrowedMult__comb, p5_smul_57330_TrailingBits___339_comb};
  assign p5_concat_147542_comb = {p5_smul_58948_NarrowedMult__comb, p5_smul_57454_TrailingBits___117_comb};
  assign p5_concat_147543_comb = {p5_smul_58950_NarrowedMult__comb, p5_smul_57454_TrailingBits___118_comb};
  assign p5_concat_147558_comb = {p5_smul_58980_NarrowedMult__comb, p5_smul_57454_TrailingBits___125_comb};
  assign p5_concat_147559_comb = {p5_smul_58982_NarrowedMult__comb, p5_smul_57454_TrailingBits___126_comb};
  assign p5_concat_147565_comb = {p5_smul_58992_NarrowedMult__comb, p5_smul_57330_TrailingBits___353_comb};
  assign p5_concat_147566_comb = {p5_smul_59002_NarrowedMult__comb, p5_smul_57330_TrailingBits___354_comb};
  assign p5_concat_147589_comb = {p5_smul_59056_NarrowedMult__comb, p5_smul_57330_TrailingBits___369_comb};
  assign p5_concat_147590_comb = {p5_smul_59066_NarrowedMult__comb, p5_smul_57330_TrailingBits___370_comb};
  assign p5_concat_147805_comb = {p5_smul_58228_NarrowedMult__comb, p5_smul_57330_TrailingBits___193_comb};
  assign p5_concat_147806_comb = {p5_smul_58230_NarrowedMult__comb, p5_smul_57330_TrailingBits___194_comb};
  assign p5_concat_147811_comb = {p5_smul_58244_NarrowedMult__comb, p5_smul_57330_TrailingBits___197_comb};
  assign p5_concat_147812_comb = {p5_smul_58246_NarrowedMult__comb, p5_smul_57330_TrailingBits___198_comb};
  assign p5_concat_147823_comb = {p5_smul_58276_NarrowedMult__comb, p5_smul_57330_TrailingBits___205_comb};
  assign p5_concat_147824_comb = {p5_smul_58278_NarrowedMult__comb, p5_smul_57330_TrailingBits___206_comb};
  assign p5_concat_147835_comb = {p5_smul_58308_NarrowedMult__comb, p5_smul_57330_TrailingBits___213_comb};
  assign p5_concat_147836_comb = {p5_smul_58310_NarrowedMult__comb, p5_smul_57330_TrailingBits___214_comb};
  assign p5_concat_147847_comb = {p5_smul_58340_NarrowedMult__comb, p5_smul_57330_TrailingBits___221_comb};
  assign p5_concat_147848_comb = {p5_smul_58342_NarrowedMult__comb, p5_smul_57330_TrailingBits___222_comb};
  assign p5_concat_147947_comb = {p5_smul_58480_NarrowedMult__comb, p5_smul_57330_TrailingBits___256_comb};
  assign p5_concat_147952_comb = {p5_smul_58490_NarrowedMult__comb, p5_smul_57330_TrailingBits___259_comb};
  assign p5_concat_147997_comb = {p5_smul_58738_NarrowedMult__comb, p5_smul_57330_TrailingBits___289_comb};
  assign p5_concat_147998_comb = {p5_smul_58744_NarrowedMult__comb, p5_smul_57330_TrailingBits___290_comb};
  assign p5_concat_148139_comb = {p5_smul_58990_NarrowedMult__comb, p5_smul_57330_TrailingBits___352_comb};
  assign p5_concat_148144_comb = {p5_smul_59004_NarrowedMult__comb, p5_smul_57330_TrailingBits___355_comb};
  assign p5_shifted__64_comb = {~p4_bit_slice_146159, p4_bit_slice_146185, p5_smul_57326_TrailingBits___192_comb};
  assign p5_smul_57326_TrailingBits___64_comb = 8'h00;
  assign p5_shifted__65_comb = {~p4_bit_slice_146160, p4_bit_slice_146186, p5_smul_57326_TrailingBits___193_comb};
  assign p5_smul_57326_TrailingBits___65_comb = 8'h00;
  assign p5_shifted__66_comb = {~p4_bit_slice_146155, p4_bit_slice_146179, p5_smul_57326_TrailingBits___194_comb};
  assign p5_smul_57326_TrailingBits___66_comb = 8'h00;
  assign p5_shifted__67_comb = {~p4_bit_slice_146161, p4_bit_slice_146187, p5_smul_57326_TrailingBits___195_comb};
  assign p5_smul_57326_TrailingBits___67_comb = 8'h00;
  assign p5_shifted__68_comb = {~p4_bit_slice_146162, p4_bit_slice_146188, p5_smul_57326_TrailingBits___196_comb};
  assign p5_smul_57326_TrailingBits___68_comb = 8'h00;
  assign p5_shifted__69_comb = {~p4_bit_slice_146156, p4_bit_slice_146180, p5_smul_57326_TrailingBits___197_comb};
  assign p5_smul_57326_TrailingBits___69_comb = 8'h00;
  assign p5_shifted__70_comb = {~p4_bit_slice_146163, p4_bit_slice_146189, p5_smul_57326_TrailingBits___198_comb};
  assign p5_smul_57326_TrailingBits___70_comb = 8'h00;
  assign p5_shifted__71_comb = {~p4_bit_slice_146164, p4_bit_slice_146190, p5_smul_57326_TrailingBits___199_comb};
  assign p5_smul_57326_TrailingBits___71_comb = 8'h00;
  assign p5_shifted__96_comb = {p4_not_146195, p4_bit_slice_146196, p5_smul_57326_TrailingBits___224_comb};
  assign p5_smul_57326_TrailingBits___96_comb = 8'h00;
  assign p5_shifted__97_comb = {p4_not_146197, p4_bit_slice_146198, p5_smul_57326_TrailingBits___225_comb};
  assign p5_smul_57326_TrailingBits___97_comb = 8'h00;
  assign p5_shifted__98_comb = {p4_not_146181, p4_bit_slice_146182, p5_smul_57326_TrailingBits___226_comb};
  assign p5_smul_57326_TrailingBits___98_comb = 8'h00;
  assign p5_shifted__99_comb = {p4_not_146199, p4_bit_slice_146200, p5_smul_57326_TrailingBits___227_comb};
  assign p5_smul_57326_TrailingBits___99_comb = 8'h00;
  assign p5_shifted__100_comb = {p4_not_146201, p4_bit_slice_146202, p5_smul_57326_TrailingBits___228_comb};
  assign p5_smul_57326_TrailingBits___100_comb = 8'h00;
  assign p5_shifted__101_comb = {p4_not_146183, p4_bit_slice_146184, p5_smul_57326_TrailingBits___229_comb};
  assign p5_smul_57326_TrailingBits___101_comb = 8'h00;
  assign p5_shifted__102_comb = {p4_not_146203, p4_bit_slice_146204, p5_smul_57326_TrailingBits___230_comb};
  assign p5_smul_57326_TrailingBits___102_comb = 8'h00;
  assign p5_shifted__103_comb = {p4_not_146205, p4_bit_slice_146206, p5_smul_57326_TrailingBits___231_comb};
  assign p5_smul_57326_TrailingBits___103_comb = 8'h00;
  assign p5_prod__779_comb = {{9{p5_concat_147829_comb[22]}}, p5_concat_147829_comb};
  assign p5_prod__784_comb = {{9{p5_concat_147830_comb[22]}}, p5_concat_147830_comb};
  assign p5_prod__781_comb = {{9{p5_concat_147971_comb[22]}}, p5_concat_147971_comb};
  assign p5_prod__812_comb = {{9{p5_concat_147976_comb[22]}}, p5_concat_147976_comb};
  assign p5_prod__801_comb = {{9{p5_concat_148021_comb[22]}}, p5_concat_148021_comb};
  assign p5_prod__819_comb = {{9{p5_concat_148022_comb[22]}}, p5_concat_148022_comb};
  assign p5_prod__803_comb = {{9{p5_concat_148163_comb[22]}}, p5_concat_148163_comb};
  assign p5_prod__831_comb = {{9{p5_concat_148168_comb[22]}}, p5_concat_148168_comb};
  assign p5_concat_147297_comb = {p5_smul_58242_NarrowedMult__comb, p5_smul_57330_TrailingBits___196_comb};
  assign p5_concat_147302_comb = {p5_smul_58248_NarrowedMult__comb, p5_smul_57330_TrailingBits___199_comb};
  assign p5_concat_147303_comb = {p5_smul_58258_NarrowedMult__comb, p5_smul_57330_TrailingBits___200_comb};
  assign p5_smul_58260_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__83_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___201_comb = 9'h000;
  assign p5_smul_58262_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__84_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___202_comb = 9'h000;
  assign p5_concat_147308_comb = {p5_smul_58264_NarrowedMult__comb, p5_smul_57330_TrailingBits___203_comb};
  assign p5_concat_147309_comb = {p5_smul_58274_NarrowedMult__comb, p5_smul_57330_TrailingBits___204_comb};
  assign p5_concat_147314_comb = {p5_smul_58280_NarrowedMult__comb, p5_smul_57330_TrailingBits___207_comb};
  assign p5_concat_147321_comb = {p5_smul_58306_NarrowedMult__comb, p5_smul_57330_TrailingBits___212_comb};
  assign p5_concat_147326_comb = {p5_smul_58312_NarrowedMult__comb, p5_smul_57330_TrailingBits___215_comb};
  assign p5_concat_147327_comb = {p5_smul_58322_NarrowedMult__comb, p5_smul_57330_TrailingBits___216_comb};
  assign p5_smul_58324_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__115_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___217_comb = 9'h000;
  assign p5_smul_58326_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__116_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___218_comb = 9'h000;
  assign p5_concat_147332_comb = {p5_smul_58328_NarrowedMult__comb, p5_smul_57330_TrailingBits___219_comb};
  assign p5_concat_147333_comb = {p5_smul_58338_NarrowedMult__comb, p5_smul_57330_TrailingBits___220_comb};
  assign p5_concat_147338_comb = {p5_smul_58344_NarrowedMult__comb, p5_smul_57330_TrailingBits___223_comb};
  assign p5_concat_147347_comb = {p5_smul_58366_NarrowedMult__comb, p5_smul_57454_TrailingBits___68_comb};
  assign p5_concat_147348_comb = {p5_smul_58368_NarrowedMult__comb, p5_smul_57330_TrailingBits___228_comb};
  assign p5_concat_147349_comb = {p5_smul_58370_NarrowedMult__comb, p5_smul_57330_TrailingBits___229_comb};
  assign p5_concat_147352_comb = {p5_smul_58376_NarrowedMult__comb, p5_smul_57330_TrailingBits___230_comb};
  assign p5_concat_147353_comb = {p5_smul_58378_NarrowedMult__comb, p5_smul_57330_TrailingBits___231_comb};
  assign p5_concat_147354_comb = {p5_smul_58380_NarrowedMult__comb, p5_smul_57454_TrailingBits___71_comb};
  assign p5_concat_147355_comb = {p5_smul_58382_NarrowedMult__comb, p5_smul_57454_TrailingBits___72_comb};
  assign p5_concat_147356_comb = {p5_smul_58384_NarrowedMult__comb, p5_smul_57330_TrailingBits___232_comb};
  assign p5_concat_147357_comb = {p5_smul_58386_NarrowedMult__comb, p5_smul_57330_TrailingBits___233_comb};
  assign p5_concat_147358_comb = {p5_smul_58388_NarrowedMult__comb, p5_smul_57454_TrailingBits___73_comb};
  assign p5_concat_147359_comb = {p5_smul_58390_NarrowedMult__comb, p5_smul_57454_TrailingBits___74_comb};
  assign p5_concat_147360_comb = {p5_smul_58392_NarrowedMult__comb, p5_smul_57330_TrailingBits___234_comb};
  assign p5_concat_147361_comb = {p5_smul_58394_NarrowedMult__comb, p5_smul_57330_TrailingBits___235_comb};
  assign p5_concat_147362_comb = {p5_smul_58396_NarrowedMult__comb, p5_smul_57454_TrailingBits___75_comb};
  assign p5_concat_147363_comb = {p5_smul_58398_NarrowedMult__comb, p5_smul_57454_TrailingBits___76_comb};
  assign p5_concat_147364_comb = {p5_smul_58400_NarrowedMult__comb, p5_smul_57330_TrailingBits___236_comb};
  assign p5_concat_147365_comb = {p5_smul_58402_NarrowedMult__comb, p5_smul_57330_TrailingBits___237_comb};
  assign p5_concat_147368_comb = {p5_smul_58408_NarrowedMult__comb, p5_smul_57330_TrailingBits___238_comb};
  assign p5_concat_147369_comb = {p5_smul_58410_NarrowedMult__comb, p5_smul_57330_TrailingBits___239_comb};
  assign p5_concat_147370_comb = {p5_smul_58412_NarrowedMult__comb, p5_smul_57454_TrailingBits___79_comb};
  assign p5_concat_147379_comb = {p5_smul_58430_NarrowedMult__comb, p5_smul_57454_TrailingBits___84_comb};
  assign p5_concat_147380_comb = {p5_smul_58432_NarrowedMult__comb, p5_smul_57330_TrailingBits___244_comb};
  assign p5_concat_147381_comb = {p5_smul_58434_NarrowedMult__comb, p5_smul_57330_TrailingBits___245_comb};
  assign p5_concat_147384_comb = {p5_smul_58440_NarrowedMult__comb, p5_smul_57330_TrailingBits___246_comb};
  assign p5_concat_147385_comb = {p5_smul_58442_NarrowedMult__comb, p5_smul_57330_TrailingBits___247_comb};
  assign p5_concat_147386_comb = {p5_smul_58444_NarrowedMult__comb, p5_smul_57454_TrailingBits___87_comb};
  assign p5_concat_147387_comb = {p5_smul_58446_NarrowedMult__comb, p5_smul_57454_TrailingBits___88_comb};
  assign p5_concat_147388_comb = {p5_smul_58448_NarrowedMult__comb, p5_smul_57330_TrailingBits___248_comb};
  assign p5_concat_147389_comb = {p5_smul_58450_NarrowedMult__comb, p5_smul_57330_TrailingBits___249_comb};
  assign p5_concat_147390_comb = {p5_smul_58452_NarrowedMult__comb, p5_smul_57454_TrailingBits___89_comb};
  assign p5_concat_147391_comb = {p5_smul_58454_NarrowedMult__comb, p5_smul_57454_TrailingBits___90_comb};
  assign p5_concat_147392_comb = {p5_smul_58456_NarrowedMult__comb, p5_smul_57330_TrailingBits___250_comb};
  assign p5_concat_147393_comb = {p5_smul_58458_NarrowedMult__comb, p5_smul_57330_TrailingBits___251_comb};
  assign p5_concat_147394_comb = {p5_smul_58460_NarrowedMult__comb, p5_smul_57454_TrailingBits___91_comb};
  assign p5_concat_147395_comb = {p5_smul_58462_NarrowedMult__comb, p5_smul_57454_TrailingBits___92_comb};
  assign p5_concat_147396_comb = {p5_smul_58464_NarrowedMult__comb, p5_smul_57330_TrailingBits___252_comb};
  assign p5_concat_147397_comb = {p5_smul_58466_NarrowedMult__comb, p5_smul_57330_TrailingBits___253_comb};
  assign p5_concat_147400_comb = {p5_smul_58472_NarrowedMult__comb, p5_smul_57330_TrailingBits___254_comb};
  assign p5_concat_147401_comb = {p5_smul_58474_NarrowedMult__comb, p5_smul_57330_TrailingBits___255_comb};
  assign p5_concat_147402_comb = {p5_smul_58476_NarrowedMult__comb, p5_smul_57454_TrailingBits___95_comb};
  assign p5_smul_58496_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__73_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___260_comb = 9'h000;
  assign p5_smul_58506_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__78_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___263_comb = 9'h000;
  assign p5_smul_58512_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__81_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___264_comb = 9'h000;
  assign p5_concat_147417_comb = {p5_smul_58516_NarrowedMult__comb, p5_smul_57330_TrailingBits___265_comb};
  assign p5_concat_147418_comb = {p5_smul_58518_NarrowedMult__comb, p5_smul_57330_TrailingBits___266_comb};
  assign p5_smul_58522_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__86_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___267_comb = 9'h000;
  assign p5_smul_58528_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__89_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___268_comb = 9'h000;
  assign p5_smul_58538_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__94_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___271_comb = 9'h000;
  assign p5_smul_58560_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__105_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___276_comb = 9'h000;
  assign p5_smul_58570_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__110_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___279_comb = 9'h000;
  assign p5_smul_58576_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__113_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___280_comb = 9'h000;
  assign p5_concat_147441_comb = {p5_smul_58580_NarrowedMult__comb, p5_smul_57330_TrailingBits___281_comb};
  assign p5_concat_147442_comb = {p5_smul_58582_NarrowedMult__comb, p5_smul_57330_TrailingBits___282_comb};
  assign p5_smul_58586_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__118_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___283_comb = 9'h000;
  assign p5_smul_58592_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__121_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___284_comb = 9'h000;
  assign p5_smul_58602_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__126_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___287_comb = 9'h000;
  assign p5_concat_147457_comb = {p5_smul_58750_NarrowedMult__comb, p5_smul_57330_TrailingBits___292_comb};
  assign p5_smul_58754_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__74_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___293_comb = 9'h000;
  assign p5_smul_58760_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__77_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___294_comb = 9'h000;
  assign p5_concat_147462_comb = {p5_smul_58764_NarrowedMult__comb, p5_smul_57330_TrailingBits___295_comb};
  assign p5_concat_147463_comb = {p5_smul_58766_NarrowedMult__comb, p5_smul_57330_TrailingBits___296_comb};
  assign p5_smul_58770_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__82_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___297_comb = 9'h000;
  assign p5_smul_58776_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__85_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___298_comb = 9'h000;
  assign p5_concat_147468_comb = {p5_smul_58780_NarrowedMult__comb, p5_smul_57330_TrailingBits___299_comb};
  assign p5_concat_147469_comb = {p5_smul_58782_NarrowedMult__comb, p5_smul_57330_TrailingBits___300_comb};
  assign p5_smul_58786_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__90_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___301_comb = 9'h000;
  assign p5_smul_58792_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__93_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___302_comb = 9'h000;
  assign p5_concat_147474_comb = {p5_smul_58796_NarrowedMult__comb, p5_smul_57330_TrailingBits___303_comb};
  assign p5_concat_147481_comb = {p5_smul_58814_NarrowedMult__comb, p5_smul_57330_TrailingBits___308_comb};
  assign p5_smul_58818_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__106_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___309_comb = 9'h000;
  assign p5_smul_58824_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__109_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___310_comb = 9'h000;
  assign p5_concat_147486_comb = {p5_smul_58828_NarrowedMult__comb, p5_smul_57330_TrailingBits___311_comb};
  assign p5_concat_147487_comb = {p5_smul_58830_NarrowedMult__comb, p5_smul_57330_TrailingBits___312_comb};
  assign p5_smul_58834_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__114_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___313_comb = 9'h000;
  assign p5_smul_58840_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__117_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___314_comb = 9'h000;
  assign p5_concat_147492_comb = {p5_smul_58844_NarrowedMult__comb, p5_smul_57330_TrailingBits___315_comb};
  assign p5_concat_147493_comb = {p5_smul_58846_NarrowedMult__comb, p5_smul_57330_TrailingBits___316_comb};
  assign p5_smul_58850_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__122_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___317_comb = 9'h000;
  assign p5_smul_58856_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__125_squeezed_comb, 6'h27);
  assign p5_smul_57330_TrailingBits___318_comb = 9'h000;
  assign p5_concat_147498_comb = {p5_smul_58860_NarrowedMult__comb, p5_smul_57330_TrailingBits___319_comb};
  assign p5_concat_147507_comb = {p5_smul_58878_NarrowedMult__comb, p5_smul_57330_TrailingBits___324_comb};
  assign p5_concat_147508_comb = {p5_smul_58880_NarrowedMult__comb, p5_smul_57454_TrailingBits___100_comb};
  assign p5_concat_147509_comb = {p5_smul_58882_NarrowedMult__comb, p5_smul_57330_TrailingBits___325_comb};
  assign p5_concat_147512_comb = {p5_smul_58888_NarrowedMult__comb, p5_smul_57330_TrailingBits___326_comb};
  assign p5_concat_147513_comb = {p5_smul_58890_NarrowedMult__comb, p5_smul_57454_TrailingBits___103_comb};
  assign p5_concat_147514_comb = {p5_smul_58892_NarrowedMult__comb, p5_smul_57330_TrailingBits___327_comb};
  assign p5_concat_147515_comb = {p5_smul_58894_NarrowedMult__comb, p5_smul_57330_TrailingBits___328_comb};
  assign p5_concat_147516_comb = {p5_smul_58896_NarrowedMult__comb, p5_smul_57454_TrailingBits___104_comb};
  assign p5_concat_147517_comb = {p5_smul_58898_NarrowedMult__comb, p5_smul_57330_TrailingBits___329_comb};
  assign p5_concat_147518_comb = {p5_smul_58900_NarrowedMult__comb, p5_smul_57454_TrailingBits___105_comb};
  assign p5_concat_147519_comb = {p5_smul_58902_NarrowedMult__comb, p5_smul_57454_TrailingBits___106_comb};
  assign p5_concat_147520_comb = {p5_smul_58904_NarrowedMult__comb, p5_smul_57330_TrailingBits___330_comb};
  assign p5_concat_147521_comb = {p5_smul_58906_NarrowedMult__comb, p5_smul_57454_TrailingBits___107_comb};
  assign p5_concat_147522_comb = {p5_smul_58908_NarrowedMult__comb, p5_smul_57330_TrailingBits___331_comb};
  assign p5_concat_147523_comb = {p5_smul_58910_NarrowedMult__comb, p5_smul_57330_TrailingBits___332_comb};
  assign p5_concat_147524_comb = {p5_smul_58912_NarrowedMult__comb, p5_smul_57454_TrailingBits___108_comb};
  assign p5_concat_147525_comb = {p5_smul_58914_NarrowedMult__comb, p5_smul_57330_TrailingBits___333_comb};
  assign p5_concat_147528_comb = {p5_smul_58920_NarrowedMult__comb, p5_smul_57330_TrailingBits___334_comb};
  assign p5_concat_147529_comb = {p5_smul_58922_NarrowedMult__comb, p5_smul_57454_TrailingBits___111_comb};
  assign p5_concat_147530_comb = {p5_smul_58924_NarrowedMult__comb, p5_smul_57330_TrailingBits___335_comb};
  assign p5_concat_147539_comb = {p5_smul_58942_NarrowedMult__comb, p5_smul_57330_TrailingBits___340_comb};
  assign p5_concat_147540_comb = {p5_smul_58944_NarrowedMult__comb, p5_smul_57454_TrailingBits___116_comb};
  assign p5_concat_147541_comb = {p5_smul_58946_NarrowedMult__comb, p5_smul_57330_TrailingBits___341_comb};
  assign p5_concat_147544_comb = {p5_smul_58952_NarrowedMult__comb, p5_smul_57330_TrailingBits___342_comb};
  assign p5_concat_147545_comb = {p5_smul_58954_NarrowedMult__comb, p5_smul_57454_TrailingBits___119_comb};
  assign p5_concat_147546_comb = {p5_smul_58956_NarrowedMult__comb, p5_smul_57330_TrailingBits___343_comb};
  assign p5_concat_147547_comb = {p5_smul_58958_NarrowedMult__comb, p5_smul_57330_TrailingBits___344_comb};
  assign p5_concat_147548_comb = {p5_smul_58960_NarrowedMult__comb, p5_smul_57454_TrailingBits___120_comb};
  assign p5_concat_147549_comb = {p5_smul_58962_NarrowedMult__comb, p5_smul_57330_TrailingBits___345_comb};
  assign p5_concat_147550_comb = {p5_smul_58964_NarrowedMult__comb, p5_smul_57454_TrailingBits___121_comb};
  assign p5_concat_147551_comb = {p5_smul_58966_NarrowedMult__comb, p5_smul_57454_TrailingBits___122_comb};
  assign p5_concat_147552_comb = {p5_smul_58968_NarrowedMult__comb, p5_smul_57330_TrailingBits___346_comb};
  assign p5_concat_147553_comb = {p5_smul_58970_NarrowedMult__comb, p5_smul_57454_TrailingBits___123_comb};
  assign p5_concat_147554_comb = {p5_smul_58972_NarrowedMult__comb, p5_smul_57330_TrailingBits___347_comb};
  assign p5_concat_147555_comb = {p5_smul_58974_NarrowedMult__comb, p5_smul_57330_TrailingBits___348_comb};
  assign p5_concat_147556_comb = {p5_smul_58976_NarrowedMult__comb, p5_smul_57454_TrailingBits___124_comb};
  assign p5_concat_147557_comb = {p5_smul_58978_NarrowedMult__comb, p5_smul_57330_TrailingBits___349_comb};
  assign p5_concat_147560_comb = {p5_smul_58984_NarrowedMult__comb, p5_smul_57330_TrailingBits___350_comb};
  assign p5_concat_147561_comb = {p5_smul_58986_NarrowedMult__comb, p5_smul_57454_TrailingBits___127_comb};
  assign p5_concat_147562_comb = {p5_smul_58988_NarrowedMult__comb, p5_smul_57330_TrailingBits___351_comb};
  assign p5_smul_59006_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__72_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___356_comb = 9'h000;
  assign p5_concat_147571_comb = {p5_smul_59008_NarrowedMult__comb, p5_smul_57330_TrailingBits___357_comb};
  assign p5_concat_147572_comb = {p5_smul_59018_NarrowedMult__comb, p5_smul_57330_TrailingBits___358_comb};
  assign p5_smul_59020_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__79_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___359_comb = 9'h000;
  assign p5_smul_59022_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__80_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___360_comb = 9'h000;
  assign p5_concat_147577_comb = {p5_smul_59024_NarrowedMult__comb, p5_smul_57330_TrailingBits___361_comb};
  assign p5_concat_147578_comb = {p5_smul_59034_NarrowedMult__comb, p5_smul_57330_TrailingBits___362_comb};
  assign p5_smul_59036_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__87_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___363_comb = 9'h000;
  assign p5_smul_59038_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__88_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___364_comb = 9'h000;
  assign p5_concat_147583_comb = {p5_smul_59040_NarrowedMult__comb, p5_smul_57330_TrailingBits___365_comb};
  assign p5_concat_147584_comb = {p5_smul_59050_NarrowedMult__comb, p5_smul_57330_TrailingBits___366_comb};
  assign p5_smul_59052_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__95_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___367_comb = 9'h000;
  assign p5_smul_59070_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__104_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___372_comb = 9'h000;
  assign p5_concat_147595_comb = {p5_smul_59072_NarrowedMult__comb, p5_smul_57330_TrailingBits___373_comb};
  assign p5_concat_147596_comb = {p5_smul_59082_NarrowedMult__comb, p5_smul_57330_TrailingBits___374_comb};
  assign p5_smul_59084_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__111_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___375_comb = 9'h000;
  assign p5_smul_59086_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__112_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___376_comb = 9'h000;
  assign p5_concat_147601_comb = {p5_smul_59088_NarrowedMult__comb, p5_smul_57330_TrailingBits___377_comb};
  assign p5_concat_147602_comb = {p5_smul_59098_NarrowedMult__comb, p5_smul_57330_TrailingBits___378_comb};
  assign p5_smul_59100_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__119_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___379_comb = 9'h000;
  assign p5_smul_59102_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__120_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___380_comb = 9'h000;
  assign p5_concat_147607_comb = {p5_smul_59104_NarrowedMult__comb, p5_smul_57330_TrailingBits___381_comb};
  assign p5_concat_147608_comb = {p5_smul_59114_NarrowedMult__comb, p5_smul_57330_TrailingBits___382_comb};
  assign p5_smul_59116_NarrowedMult__comb = smul14b_8b_x_6b(p5_shifted__127_squeezed_comb, 6'h19);
  assign p5_smul_57330_TrailingBits___383_comb = 9'h000;
  assign p5_prod__519_comb = {{7{p5_concat_147291_comb[24]}}, p5_concat_147291_comb};
  assign p5_prod__534_comb = {{7{p5_concat_147296_comb[24]}}, p5_concat_147296_comb};
  assign p5_prod__775_comb = {{7{p5_concat_147315_comb[24]}}, p5_concat_147315_comb};
  assign p5_prod__790_comb = {{7{p5_concat_147320_comb[24]}}, p5_concat_147320_comb};
  assign p5_prod__517_comb = {{7{p5_concat_147339_comb[24]}}, p5_concat_147339_comb};
  assign p5_prod__520_comb = {{8{p5_concat_147340_comb[23]}}, p5_concat_147340_comb};
  assign p5_prod__524_comb = {{8{p5_concat_147341_comb[23]}}, p5_concat_147341_comb};
  assign p5_prod__529_comb = {{7{p5_concat_147342_comb[24]}}, p5_concat_147342_comb};
  assign p5_prod__535_comb = {{7{p5_concat_147343_comb[24]}}, p5_concat_147343_comb};
  assign p5_prod__542_comb = {{8{p5_concat_147344_comb[23]}}, p5_concat_147344_comb};
  assign p5_prod__549_comb = {{8{p5_concat_147345_comb[23]}}, p5_concat_147345_comb};
  assign p5_prod__555_comb = {{7{p5_concat_147346_comb[24]}}, p5_concat_147346_comb};
  assign p5_prod__593_comb = {{7{p5_concat_147350_comb[24]}}, p5_concat_147350_comb};
  assign p5_prod__599_comb = {{7{p5_concat_147351_comb[24]}}, p5_concat_147351_comb};
  assign p5_prod__721_comb = {{7{p5_concat_147366_comb[24]}}, p5_concat_147366_comb};
  assign p5_prod__727_comb = {{7{p5_concat_147367_comb[24]}}, p5_concat_147367_comb};
  assign p5_prod__773_comb = {{7{p5_concat_147371_comb[24]}}, p5_concat_147371_comb};
  assign p5_prod__776_comb = {{8{p5_concat_147372_comb[23]}}, p5_concat_147372_comb};
  assign p5_prod__780_comb = {{8{p5_concat_147373_comb[23]}}, p5_concat_147373_comb};
  assign p5_prod__785_comb = {{7{p5_concat_147374_comb[24]}}, p5_concat_147374_comb};
  assign p5_prod__791_comb = {{7{p5_concat_147375_comb[24]}}, p5_concat_147375_comb};
  assign p5_prod__798_comb = {{8{p5_concat_147376_comb[23]}}, p5_concat_147376_comb};
  assign p5_prod__805_comb = {{8{p5_concat_147377_comb[23]}}, p5_concat_147377_comb};
  assign p5_prod__811_comb = {{7{p5_concat_147378_comb[24]}}, p5_concat_147378_comb};
  assign p5_prod__849_comb = {{7{p5_concat_147382_comb[24]}}, p5_concat_147382_comb};
  assign p5_prod__855_comb = {{7{p5_concat_147383_comb[24]}}, p5_concat_147383_comb};
  assign p5_prod__977_comb = {{7{p5_concat_147398_comb[24]}}, p5_concat_147398_comb};
  assign p5_prod__983_comb = {{7{p5_concat_147399_comb[24]}}, p5_concat_147399_comb};
  assign p5_prod__536_comb = {{7{p5_concat_147405_comb[24]}}, p5_concat_147405_comb};
  assign p5_prod__543_comb = {{7{p5_concat_147406_comb[24]}}, p5_concat_147406_comb};
  assign p5_prod__600_comb = {{7{p5_concat_147411_comb[24]}}, p5_concat_147411_comb};
  assign p5_prod__607_comb = {{7{p5_concat_147412_comb[24]}}, p5_concat_147412_comb};
  assign p5_prod__728_comb = {{7{p5_concat_147423_comb[24]}}, p5_concat_147423_comb};
  assign p5_prod__735_comb = {{7{p5_concat_147424_comb[24]}}, p5_concat_147424_comb};
  assign p5_prod__792_comb = {{7{p5_concat_147429_comb[24]}}, p5_concat_147429_comb};
  assign p5_prod__799_comb = {{7{p5_concat_147430_comb[24]}}, p5_concat_147430_comb};
  assign p5_prod__856_comb = {{7{p5_concat_147435_comb[24]}}, p5_concat_147435_comb};
  assign p5_prod__863_comb = {{7{p5_concat_147436_comb[24]}}, p5_concat_147436_comb};
  assign p5_prod__984_comb = {{7{p5_concat_147447_comb[24]}}, p5_concat_147447_comb};
  assign p5_prod__991_comb = {{7{p5_concat_147448_comb[24]}}, p5_concat_147448_comb};
  assign p5_prod__532_comb = {{7{p5_concat_147451_comb[24]}}, p5_concat_147451_comb};
  assign p5_prod__570_comb = {{7{p5_concat_147456_comb[24]}}, p5_concat_147456_comb};
  assign p5_prod__788_comb = {{7{p5_concat_147475_comb[24]}}, p5_concat_147475_comb};
  assign p5_prod__826_comb = {{7{p5_concat_147480_comb[24]}}, p5_concat_147480_comb};
  assign p5_prod__539_comb = {{8{p5_concat_147499_comb[23]}}, p5_concat_147499_comb};
  assign p5_prod__546_comb = {{7{p5_concat_147500_comb[24]}}, p5_concat_147500_comb};
  assign p5_prod__553_comb = {{8{p5_concat_147501_comb[23]}}, p5_concat_147501_comb};
  assign p5_prod__559_comb = {{7{p5_concat_147502_comb[24]}}, p5_concat_147502_comb};
  assign p5_prod__564_comb = {{7{p5_concat_147503_comb[24]}}, p5_concat_147503_comb};
  assign p5_prod__568_comb = {{8{p5_concat_147504_comb[23]}}, p5_concat_147504_comb};
  assign p5_prod__571_comb = {{7{p5_concat_147505_comb[24]}}, p5_concat_147505_comb};
  assign p5_prod__573_comb = {{8{p5_concat_147506_comb[23]}}, p5_concat_147506_comb};
  assign p5_prod__623_comb = {{7{p5_concat_147510_comb[24]}}, p5_concat_147510_comb};
  assign p5_prod__628_comb = {{7{p5_concat_147511_comb[24]}}, p5_concat_147511_comb};
  assign p5_prod__751_comb = {{7{p5_concat_147526_comb[24]}}, p5_concat_147526_comb};
  assign p5_prod__756_comb = {{7{p5_concat_147527_comb[24]}}, p5_concat_147527_comb};
  assign p5_prod__795_comb = {{8{p5_concat_147531_comb[23]}}, p5_concat_147531_comb};
  assign p5_prod__802_comb = {{7{p5_concat_147532_comb[24]}}, p5_concat_147532_comb};
  assign p5_prod__809_comb = {{8{p5_concat_147533_comb[23]}}, p5_concat_147533_comb};
  assign p5_prod__815_comb = {{7{p5_concat_147534_comb[24]}}, p5_concat_147534_comb};
  assign p5_prod__820_comb = {{7{p5_concat_147535_comb[24]}}, p5_concat_147535_comb};
  assign p5_prod__824_comb = {{8{p5_concat_147536_comb[23]}}, p5_concat_147536_comb};
  assign p5_prod__827_comb = {{7{p5_concat_147537_comb[24]}}, p5_concat_147537_comb};
  assign p5_prod__829_comb = {{8{p5_concat_147538_comb[23]}}, p5_concat_147538_comb};
  assign p5_prod__879_comb = {{7{p5_concat_147542_comb[24]}}, p5_concat_147542_comb};
  assign p5_prod__884_comb = {{7{p5_concat_147543_comb[24]}}, p5_concat_147543_comb};
  assign p5_prod__1007_comb = {{7{p5_concat_147558_comb[24]}}, p5_concat_147558_comb};
  assign p5_prod__1012_comb = {{7{p5_concat_147559_comb[24]}}, p5_concat_147559_comb};
  assign p5_prod__554_comb = {{7{p5_concat_147565_comb[24]}}, p5_concat_147565_comb};
  assign p5_prod__574_comb = {{7{p5_concat_147566_comb[24]}}, p5_concat_147566_comb};
  assign p5_prod__810_comb = {{7{p5_concat_147589_comb[24]}}, p5_concat_147589_comb};
  assign p5_prod__830_comb = {{7{p5_concat_147590_comb[24]}}, p5_concat_147590_comb};
  assign p5_prod__523_comb = {{9{p5_concat_147805_comb[22]}}, p5_concat_147805_comb};
  assign p5_prod__528_comb = {{9{p5_concat_147806_comb[22]}}, p5_concat_147806_comb};
  assign p5_prod__587_comb = {{9{p5_concat_147811_comb[22]}}, p5_concat_147811_comb};
  assign p5_prod__592_comb = {{9{p5_concat_147812_comb[22]}}, p5_concat_147812_comb};
  assign p5_prod__715_comb = {{9{p5_concat_147823_comb[22]}}, p5_concat_147823_comb};
  assign p5_prod__720_comb = {{9{p5_concat_147824_comb[22]}}, p5_concat_147824_comb};
  assign p5_prod__843_comb = {{9{p5_concat_147835_comb[22]}}, p5_concat_147835_comb};
  assign p5_prod__848_comb = {{9{p5_concat_147836_comb[22]}}, p5_concat_147836_comb};
  assign p5_prod__971_comb = {{9{p5_concat_147847_comb[22]}}, p5_concat_147847_comb};
  assign p5_prod__976_comb = {{9{p5_concat_147848_comb[22]}}, p5_concat_147848_comb};
  assign p5_prod__525_comb = {{9{p5_concat_147947_comb[22]}}, p5_concat_147947_comb};
  assign p5_prod__556_comb = {{9{p5_concat_147952_comb[22]}}, p5_concat_147952_comb};
  assign p5_prod__545_comb = {{9{p5_concat_147997_comb[22]}}, p5_concat_147997_comb};
  assign p5_prod__563_comb = {{9{p5_concat_147998_comb[22]}}, p5_concat_147998_comb};
  assign p5_prod__547_comb = {{9{p5_concat_148139_comb[22]}}, p5_concat_148139_comb};
  assign p5_prod__575_comb = {{9{p5_concat_148144_comb[22]}}, p5_concat_148144_comb};
  assign p5_or_149154_comb = p5_prod__779_comb | 32'h0000_0080;
  assign p5_or_149155_comb = p5_prod__784_comb | 32'h0000_0080;
  assign p5_or_149319_comb = p5_prod__781_comb | 32'h0000_0080;
  assign p5_or_149326_comb = p5_prod__812_comb | 32'h0000_0080;
  assign p5_or_149370_comb = p5_prod__801_comb | 32'h0000_0080;
  assign p5_or_149371_comb = p5_prod__819_comb | 32'h0000_0080;
  assign p5_or_149527_comb = p5_prod__803_comb | 32'h0000_0080;
  assign p5_or_149534_comb = p5_prod__831_comb | 32'h0000_0080;
  assign p5_smul_57326_TrailingBits___200_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___201_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___202_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___203_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___204_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___205_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___206_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___207_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___208_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___209_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___210_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___211_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___212_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___213_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___214_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___215_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___216_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___217_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___218_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___219_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___220_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___221_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___222_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___223_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___232_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___233_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___234_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___235_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___236_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___237_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___238_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___239_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___240_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___241_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___242_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___243_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___244_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___245_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___246_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___247_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___248_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___249_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___250_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___251_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___252_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___253_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___254_comb = 8'h00;
  assign p5_smul_57326_TrailingBits___255_comb = 8'h00;
  assign p5_prod__583_comb = {{7{p5_concat_147297_comb[24]}}, p5_concat_147297_comb};
  assign p5_prod__598_comb = {{7{p5_concat_147302_comb[24]}}, p5_concat_147302_comb};
  assign p5_prod__647_comb = {{7{p5_concat_147303_comb[24]}}, p5_concat_147303_comb};
  assign p5_concat_147817_comb = {p5_smul_58260_NarrowedMult__comb, p5_smul_57330_TrailingBits___201_comb};
  assign p5_concat_147818_comb = {p5_smul_58262_NarrowedMult__comb, p5_smul_57330_TrailingBits___202_comb};
  assign p5_prod__662_comb = {{7{p5_concat_147308_comb[24]}}, p5_concat_147308_comb};
  assign p5_prod__711_comb = {{7{p5_concat_147309_comb[24]}}, p5_concat_147309_comb};
  assign p5_prod__726_comb = {{7{p5_concat_147314_comb[24]}}, p5_concat_147314_comb};
  assign p5_prod__839_comb = {{7{p5_concat_147321_comb[24]}}, p5_concat_147321_comb};
  assign p5_prod__854_comb = {{7{p5_concat_147326_comb[24]}}, p5_concat_147326_comb};
  assign p5_prod__903_comb = {{7{p5_concat_147327_comb[24]}}, p5_concat_147327_comb};
  assign p5_concat_147841_comb = {p5_smul_58324_NarrowedMult__comb, p5_smul_57330_TrailingBits___217_comb};
  assign p5_concat_147842_comb = {p5_smul_58326_NarrowedMult__comb, p5_smul_57330_TrailingBits___218_comb};
  assign p5_prod__918_comb = {{7{p5_concat_147332_comb[24]}}, p5_concat_147332_comb};
  assign p5_prod__967_comb = {{7{p5_concat_147333_comb[24]}}, p5_concat_147333_comb};
  assign p5_prod__982_comb = {{7{p5_concat_147338_comb[24]}}, p5_concat_147338_comb};
  assign p5_prod__581_comb = {{7{p5_concat_147347_comb[24]}}, p5_concat_147347_comb};
  assign p5_prod__584_comb = {{8{p5_concat_147348_comb[23]}}, p5_concat_147348_comb};
  assign p5_prod__588_comb = {{8{p5_concat_147349_comb[23]}}, p5_concat_147349_comb};
  assign p5_prod__606_comb = {{8{p5_concat_147352_comb[23]}}, p5_concat_147352_comb};
  assign p5_prod__613_comb = {{8{p5_concat_147353_comb[23]}}, p5_concat_147353_comb};
  assign p5_prod__619_comb = {{7{p5_concat_147354_comb[24]}}, p5_concat_147354_comb};
  assign p5_prod__645_comb = {{7{p5_concat_147355_comb[24]}}, p5_concat_147355_comb};
  assign p5_prod__648_comb = {{8{p5_concat_147356_comb[23]}}, p5_concat_147356_comb};
  assign p5_prod__652_comb = {{8{p5_concat_147357_comb[23]}}, p5_concat_147357_comb};
  assign p5_prod__657_comb = {{7{p5_concat_147358_comb[24]}}, p5_concat_147358_comb};
  assign p5_prod__663_comb = {{7{p5_concat_147359_comb[24]}}, p5_concat_147359_comb};
  assign p5_prod__670_comb = {{8{p5_concat_147360_comb[23]}}, p5_concat_147360_comb};
  assign p5_prod__677_comb = {{8{p5_concat_147361_comb[23]}}, p5_concat_147361_comb};
  assign p5_prod__683_comb = {{7{p5_concat_147362_comb[24]}}, p5_concat_147362_comb};
  assign p5_prod__709_comb = {{7{p5_concat_147363_comb[24]}}, p5_concat_147363_comb};
  assign p5_prod__712_comb = {{8{p5_concat_147364_comb[23]}}, p5_concat_147364_comb};
  assign p5_prod__716_comb = {{8{p5_concat_147365_comb[23]}}, p5_concat_147365_comb};
  assign p5_prod__734_comb = {{8{p5_concat_147368_comb[23]}}, p5_concat_147368_comb};
  assign p5_prod__741_comb = {{8{p5_concat_147369_comb[23]}}, p5_concat_147369_comb};
  assign p5_prod__747_comb = {{7{p5_concat_147370_comb[24]}}, p5_concat_147370_comb};
  assign p5_prod__837_comb = {{7{p5_concat_147379_comb[24]}}, p5_concat_147379_comb};
  assign p5_prod__840_comb = {{8{p5_concat_147380_comb[23]}}, p5_concat_147380_comb};
  assign p5_prod__844_comb = {{8{p5_concat_147381_comb[23]}}, p5_concat_147381_comb};
  assign p5_prod__862_comb = {{8{p5_concat_147384_comb[23]}}, p5_concat_147384_comb};
  assign p5_prod__869_comb = {{8{p5_concat_147385_comb[23]}}, p5_concat_147385_comb};
  assign p5_prod__875_comb = {{7{p5_concat_147386_comb[24]}}, p5_concat_147386_comb};
  assign p5_prod__901_comb = {{7{p5_concat_147387_comb[24]}}, p5_concat_147387_comb};
  assign p5_prod__904_comb = {{8{p5_concat_147388_comb[23]}}, p5_concat_147388_comb};
  assign p5_prod__908_comb = {{8{p5_concat_147389_comb[23]}}, p5_concat_147389_comb};
  assign p5_prod__913_comb = {{7{p5_concat_147390_comb[24]}}, p5_concat_147390_comb};
  assign p5_prod__919_comb = {{7{p5_concat_147391_comb[24]}}, p5_concat_147391_comb};
  assign p5_prod__926_comb = {{8{p5_concat_147392_comb[23]}}, p5_concat_147392_comb};
  assign p5_prod__933_comb = {{8{p5_concat_147393_comb[23]}}, p5_concat_147393_comb};
  assign p5_prod__939_comb = {{7{p5_concat_147394_comb[24]}}, p5_concat_147394_comb};
  assign p5_prod__965_comb = {{7{p5_concat_147395_comb[24]}}, p5_concat_147395_comb};
  assign p5_prod__968_comb = {{8{p5_concat_147396_comb[23]}}, p5_concat_147396_comb};
  assign p5_prod__972_comb = {{8{p5_concat_147397_comb[23]}}, p5_concat_147397_comb};
  assign p5_prod__990_comb = {{8{p5_concat_147400_comb[23]}}, p5_concat_147400_comb};
  assign p5_prod__997_comb = {{8{p5_concat_147401_comb[23]}}, p5_concat_147401_comb};
  assign p5_prod__1003_comb = {{7{p5_concat_147402_comb[24]}}, p5_concat_147402_comb};
  assign p5_concat_147953_comb = {p5_smul_58496_NarrowedMult__comb, p5_smul_57330_TrailingBits___260_comb};
  assign p5_concat_147958_comb = {p5_smul_58506_NarrowedMult__comb, p5_smul_57330_TrailingBits___263_comb};
  assign p5_concat_147959_comb = {p5_smul_58512_NarrowedMult__comb, p5_smul_57330_TrailingBits___264_comb};
  assign p5_prod__664_comb = {{7{p5_concat_147417_comb[24]}}, p5_concat_147417_comb};
  assign p5_prod__671_comb = {{7{p5_concat_147418_comb[24]}}, p5_concat_147418_comb};
  assign p5_concat_147964_comb = {p5_smul_58522_NarrowedMult__comb, p5_smul_57330_TrailingBits___267_comb};
  assign p5_concat_147965_comb = {p5_smul_58528_NarrowedMult__comb, p5_smul_57330_TrailingBits___268_comb};
  assign p5_concat_147970_comb = {p5_smul_58538_NarrowedMult__comb, p5_smul_57330_TrailingBits___271_comb};
  assign p5_concat_147977_comb = {p5_smul_58560_NarrowedMult__comb, p5_smul_57330_TrailingBits___276_comb};
  assign p5_concat_147982_comb = {p5_smul_58570_NarrowedMult__comb, p5_smul_57330_TrailingBits___279_comb};
  assign p5_concat_147983_comb = {p5_smul_58576_NarrowedMult__comb, p5_smul_57330_TrailingBits___280_comb};
  assign p5_prod__920_comb = {{7{p5_concat_147441_comb[24]}}, p5_concat_147441_comb};
  assign p5_prod__927_comb = {{7{p5_concat_147442_comb[24]}}, p5_concat_147442_comb};
  assign p5_concat_147988_comb = {p5_smul_58586_NarrowedMult__comb, p5_smul_57330_TrailingBits___283_comb};
  assign p5_concat_147989_comb = {p5_smul_58592_NarrowedMult__comb, p5_smul_57330_TrailingBits___284_comb};
  assign p5_concat_147994_comb = {p5_smul_58602_NarrowedMult__comb, p5_smul_57330_TrailingBits___287_comb};
  assign p5_prod__596_comb = {{7{p5_concat_147457_comb[24]}}, p5_concat_147457_comb};
  assign p5_concat_148003_comb = {p5_smul_58754_NarrowedMult__comb, p5_smul_57330_TrailingBits___293_comb};
  assign p5_concat_148004_comb = {p5_smul_58760_NarrowedMult__comb, p5_smul_57330_TrailingBits___294_comb};
  assign p5_prod__634_comb = {{7{p5_concat_147462_comb[24]}}, p5_concat_147462_comb};
  assign p5_prod__660_comb = {{7{p5_concat_147463_comb[24]}}, p5_concat_147463_comb};
  assign p5_concat_148009_comb = {p5_smul_58770_NarrowedMult__comb, p5_smul_57330_TrailingBits___297_comb};
  assign p5_concat_148010_comb = {p5_smul_58776_NarrowedMult__comb, p5_smul_57330_TrailingBits___298_comb};
  assign p5_prod__698_comb = {{7{p5_concat_147468_comb[24]}}, p5_concat_147468_comb};
  assign p5_prod__724_comb = {{7{p5_concat_147469_comb[24]}}, p5_concat_147469_comb};
  assign p5_concat_148015_comb = {p5_smul_58786_NarrowedMult__comb, p5_smul_57330_TrailingBits___301_comb};
  assign p5_concat_148016_comb = {p5_smul_58792_NarrowedMult__comb, p5_smul_57330_TrailingBits___302_comb};
  assign p5_prod__762_comb = {{7{p5_concat_147474_comb[24]}}, p5_concat_147474_comb};
  assign p5_prod__852_comb = {{7{p5_concat_147481_comb[24]}}, p5_concat_147481_comb};
  assign p5_concat_148027_comb = {p5_smul_58818_NarrowedMult__comb, p5_smul_57330_TrailingBits___309_comb};
  assign p5_concat_148028_comb = {p5_smul_58824_NarrowedMult__comb, p5_smul_57330_TrailingBits___310_comb};
  assign p5_prod__890_comb = {{7{p5_concat_147486_comb[24]}}, p5_concat_147486_comb};
  assign p5_prod__916_comb = {{7{p5_concat_147487_comb[24]}}, p5_concat_147487_comb};
  assign p5_concat_148033_comb = {p5_smul_58834_NarrowedMult__comb, p5_smul_57330_TrailingBits___313_comb};
  assign p5_concat_148034_comb = {p5_smul_58840_NarrowedMult__comb, p5_smul_57330_TrailingBits___314_comb};
  assign p5_prod__954_comb = {{7{p5_concat_147492_comb[24]}}, p5_concat_147492_comb};
  assign p5_prod__980_comb = {{7{p5_concat_147493_comb[24]}}, p5_concat_147493_comb};
  assign p5_concat_148039_comb = {p5_smul_58850_NarrowedMult__comb, p5_smul_57330_TrailingBits___317_comb};
  assign p5_concat_148040_comb = {p5_smul_58856_NarrowedMult__comb, p5_smul_57330_TrailingBits___318_comb};
  assign p5_prod__1018_comb = {{7{p5_concat_147498_comb[24]}}, p5_concat_147498_comb};
  assign p5_prod__603_comb = {{8{p5_concat_147507_comb[23]}}, p5_concat_147507_comb};
  assign p5_prod__610_comb = {{7{p5_concat_147508_comb[24]}}, p5_concat_147508_comb};
  assign p5_prod__617_comb = {{8{p5_concat_147509_comb[23]}}, p5_concat_147509_comb};
  assign p5_prod__632_comb = {{8{p5_concat_147512_comb[23]}}, p5_concat_147512_comb};
  assign p5_prod__635_comb = {{7{p5_concat_147513_comb[24]}}, p5_concat_147513_comb};
  assign p5_prod__637_comb = {{8{p5_concat_147514_comb[23]}}, p5_concat_147514_comb};
  assign p5_prod__667_comb = {{8{p5_concat_147515_comb[23]}}, p5_concat_147515_comb};
  assign p5_prod__674_comb = {{7{p5_concat_147516_comb[24]}}, p5_concat_147516_comb};
  assign p5_prod__681_comb = {{8{p5_concat_147517_comb[23]}}, p5_concat_147517_comb};
  assign p5_prod__687_comb = {{7{p5_concat_147518_comb[24]}}, p5_concat_147518_comb};
  assign p5_prod__692_comb = {{7{p5_concat_147519_comb[24]}}, p5_concat_147519_comb};
  assign p5_prod__696_comb = {{8{p5_concat_147520_comb[23]}}, p5_concat_147520_comb};
  assign p5_prod__699_comb = {{7{p5_concat_147521_comb[24]}}, p5_concat_147521_comb};
  assign p5_prod__701_comb = {{8{p5_concat_147522_comb[23]}}, p5_concat_147522_comb};
  assign p5_prod__731_comb = {{8{p5_concat_147523_comb[23]}}, p5_concat_147523_comb};
  assign p5_prod__738_comb = {{7{p5_concat_147524_comb[24]}}, p5_concat_147524_comb};
  assign p5_prod__745_comb = {{8{p5_concat_147525_comb[23]}}, p5_concat_147525_comb};
  assign p5_prod__760_comb = {{8{p5_concat_147528_comb[23]}}, p5_concat_147528_comb};
  assign p5_prod__763_comb = {{7{p5_concat_147529_comb[24]}}, p5_concat_147529_comb};
  assign p5_prod__765_comb = {{8{p5_concat_147530_comb[23]}}, p5_concat_147530_comb};
  assign p5_prod__859_comb = {{8{p5_concat_147539_comb[23]}}, p5_concat_147539_comb};
  assign p5_prod__866_comb = {{7{p5_concat_147540_comb[24]}}, p5_concat_147540_comb};
  assign p5_prod__873_comb = {{8{p5_concat_147541_comb[23]}}, p5_concat_147541_comb};
  assign p5_prod__888_comb = {{8{p5_concat_147544_comb[23]}}, p5_concat_147544_comb};
  assign p5_prod__891_comb = {{7{p5_concat_147545_comb[24]}}, p5_concat_147545_comb};
  assign p5_prod__893_comb = {{8{p5_concat_147546_comb[23]}}, p5_concat_147546_comb};
  assign p5_prod__923_comb = {{8{p5_concat_147547_comb[23]}}, p5_concat_147547_comb};
  assign p5_prod__930_comb = {{7{p5_concat_147548_comb[24]}}, p5_concat_147548_comb};
  assign p5_prod__937_comb = {{8{p5_concat_147549_comb[23]}}, p5_concat_147549_comb};
  assign p5_prod__943_comb = {{7{p5_concat_147550_comb[24]}}, p5_concat_147550_comb};
  assign p5_prod__948_comb = {{7{p5_concat_147551_comb[24]}}, p5_concat_147551_comb};
  assign p5_prod__952_comb = {{8{p5_concat_147552_comb[23]}}, p5_concat_147552_comb};
  assign p5_prod__955_comb = {{7{p5_concat_147553_comb[24]}}, p5_concat_147553_comb};
  assign p5_prod__957_comb = {{8{p5_concat_147554_comb[23]}}, p5_concat_147554_comb};
  assign p5_prod__987_comb = {{8{p5_concat_147555_comb[23]}}, p5_concat_147555_comb};
  assign p5_prod__994_comb = {{7{p5_concat_147556_comb[24]}}, p5_concat_147556_comb};
  assign p5_prod__1001_comb = {{8{p5_concat_147557_comb[23]}}, p5_concat_147557_comb};
  assign p5_prod__1016_comb = {{8{p5_concat_147560_comb[23]}}, p5_concat_147560_comb};
  assign p5_prod__1019_comb = {{7{p5_concat_147561_comb[24]}}, p5_concat_147561_comb};
  assign p5_prod__1021_comb = {{8{p5_concat_147562_comb[23]}}, p5_concat_147562_comb};
  assign p5_concat_148145_comb = {p5_smul_59006_NarrowedMult__comb, p5_smul_57330_TrailingBits___356_comb};
  assign p5_prod__618_comb = {{7{p5_concat_147571_comb[24]}}, p5_concat_147571_comb};
  assign p5_prod__638_comb = {{7{p5_concat_147572_comb[24]}}, p5_concat_147572_comb};
  assign p5_concat_148150_comb = {p5_smul_59020_NarrowedMult__comb, p5_smul_57330_TrailingBits___359_comb};
  assign p5_concat_148151_comb = {p5_smul_59022_NarrowedMult__comb, p5_smul_57330_TrailingBits___360_comb};
  assign p5_prod__682_comb = {{7{p5_concat_147577_comb[24]}}, p5_concat_147577_comb};
  assign p5_prod__702_comb = {{7{p5_concat_147578_comb[24]}}, p5_concat_147578_comb};
  assign p5_concat_148156_comb = {p5_smul_59036_NarrowedMult__comb, p5_smul_57330_TrailingBits___363_comb};
  assign p5_concat_148157_comb = {p5_smul_59038_NarrowedMult__comb, p5_smul_57330_TrailingBits___364_comb};
  assign p5_prod__746_comb = {{7{p5_concat_147583_comb[24]}}, p5_concat_147583_comb};
  assign p5_prod__766_comb = {{7{p5_concat_147584_comb[24]}}, p5_concat_147584_comb};
  assign p5_concat_148162_comb = {p5_smul_59052_NarrowedMult__comb, p5_smul_57330_TrailingBits___367_comb};
  assign p5_concat_148169_comb = {p5_smul_59070_NarrowedMult__comb, p5_smul_57330_TrailingBits___372_comb};
  assign p5_prod__874_comb = {{7{p5_concat_147595_comb[24]}}, p5_concat_147595_comb};
  assign p5_prod__894_comb = {{7{p5_concat_147596_comb[24]}}, p5_concat_147596_comb};
  assign p5_concat_148174_comb = {p5_smul_59084_NarrowedMult__comb, p5_smul_57330_TrailingBits___375_comb};
  assign p5_concat_148175_comb = {p5_smul_59086_NarrowedMult__comb, p5_smul_57330_TrailingBits___376_comb};
  assign p5_prod__938_comb = {{7{p5_concat_147601_comb[24]}}, p5_concat_147601_comb};
  assign p5_prod__958_comb = {{7{p5_concat_147602_comb[24]}}, p5_concat_147602_comb};
  assign p5_concat_148180_comb = {p5_smul_59100_NarrowedMult__comb, p5_smul_57330_TrailingBits___379_comb};
  assign p5_concat_148181_comb = {p5_smul_59102_NarrowedMult__comb, p5_smul_57330_TrailingBits___380_comb};
  assign p5_prod__1002_comb = {{7{p5_concat_147607_comb[24]}}, p5_concat_147607_comb};
  assign p5_prod__1022_comb = {{7{p5_concat_147608_comb[24]}}, p5_concat_147608_comb};
  assign p5_concat_148186_comb = {p5_smul_59116_NarrowedMult__comb, p5_smul_57330_TrailingBits___383_comb};
  assign p5_or_148397_comb = p5_prod__519_comb | 32'h0000_0080;
  assign p5_or_148404_comb = p5_prod__534_comb | 32'h0000_0080;
  assign p5_or_148437_comb = p5_prod__775_comb | 32'h0000_0080;
  assign p5_or_148444_comb = p5_prod__790_comb | 32'h0000_0080;
  assign p5_or_148477_comb = p5_prod__517_comb | 32'h0000_0080;
  assign p5_or_148484_comb = p5_prod__529_comb | 32'h0000_0080;
  assign p5_or_148487_comb = p5_prod__535_comb | 32'h0000_0080;
  assign p5_or_148494_comb = p5_prod__555_comb | 32'h0000_0080;
  assign p5_or_148504_comb = p5_prod__593_comb | 32'h0000_0080;
  assign p5_or_148507_comb = p5_prod__599_comb | 32'h0000_0080;
  assign p5_or_148544_comb = p5_prod__721_comb | 32'h0000_0080;
  assign p5_or_148547_comb = p5_prod__727_comb | 32'h0000_0080;
  assign p5_or_148557_comb = p5_prod__773_comb | 32'h0000_0080;
  assign p5_or_148564_comb = p5_prod__785_comb | 32'h0000_0080;
  assign p5_or_148567_comb = p5_prod__791_comb | 32'h0000_0080;
  assign p5_or_148574_comb = p5_prod__811_comb | 32'h0000_0080;
  assign p5_or_148584_comb = p5_prod__849_comb | 32'h0000_0080;
  assign p5_or_148587_comb = p5_prod__855_comb | 32'h0000_0080;
  assign p5_or_148624_comb = p5_prod__977_comb | 32'h0000_0080;
  assign p5_or_148627_comb = p5_prod__983_comb | 32'h0000_0080;
  assign p5_or_148639_comb = p5_prod__536_comb | 32'h0000_0080;
  assign p5_or_148642_comb = p5_prod__543_comb | 32'h0000_0080;
  assign p5_or_148649_comb = p5_prod__600_comb | 32'h0000_0080;
  assign p5_or_148652_comb = p5_prod__607_comb | 32'h0000_0080;
  assign p5_or_148669_comb = p5_prod__728_comb | 32'h0000_0080;
  assign p5_or_148672_comb = p5_prod__735_comb | 32'h0000_0080;
  assign p5_or_148679_comb = p5_prod__792_comb | 32'h0000_0080;
  assign p5_or_148682_comb = p5_prod__799_comb | 32'h0000_0080;
  assign p5_or_148689_comb = p5_prod__856_comb | 32'h0000_0080;
  assign p5_or_148692_comb = p5_prod__863_comb | 32'h0000_0080;
  assign p5_or_148709_comb = p5_prod__984_comb | 32'h0000_0080;
  assign p5_or_148712_comb = p5_prod__991_comb | 32'h0000_0080;
  assign p5_or_148717_comb = p5_prod__532_comb | 32'h0000_0080;
  assign p5_or_148724_comb = p5_prod__570_comb | 32'h0000_0080;
  assign p5_or_148757_comb = p5_prod__788_comb | 32'h0000_0080;
  assign p5_or_148764_comb = p5_prod__826_comb | 32'h0000_0080;
  assign p5_or_148799_comb = p5_prod__546_comb | 32'h0000_0080;
  assign p5_or_148804_comb = p5_prod__559_comb | 32'h0000_0080;
  assign p5_or_148807_comb = p5_prod__564_comb | 32'h0000_0080;
  assign p5_or_148812_comb = p5_prod__571_comb | 32'h0000_0080;
  assign p5_or_148824_comb = p5_prod__623_comb | 32'h0000_0080;
  assign p5_or_148827_comb = p5_prod__628_comb | 32'h0000_0080;
  assign p5_or_148864_comb = p5_prod__751_comb | 32'h0000_0080;
  assign p5_or_148867_comb = p5_prod__756_comb | 32'h0000_0080;
  assign p5_or_148879_comb = p5_prod__802_comb | 32'h0000_0080;
  assign p5_or_148884_comb = p5_prod__815_comb | 32'h0000_0080;
  assign p5_or_148887_comb = p5_prod__820_comb | 32'h0000_0080;
  assign p5_or_148892_comb = p5_prod__827_comb | 32'h0000_0080;
  assign p5_or_148904_comb = p5_prod__879_comb | 32'h0000_0080;
  assign p5_or_148907_comb = p5_prod__884_comb | 32'h0000_0080;
  assign p5_or_148944_comb = p5_prod__1007_comb | 32'h0000_0080;
  assign p5_or_148947_comb = p5_prod__1012_comb | 32'h0000_0080;
  assign p5_or_148959_comb = p5_prod__554_comb | 32'h0000_0080;
  assign p5_or_148962_comb = p5_prod__574_comb | 32'h0000_0080;
  assign p5_or_148999_comb = p5_prod__810_comb | 32'h0000_0080;
  assign p5_or_149002_comb = p5_prod__830_comb | 32'h0000_0080;
  assign p5_or_149134_comb = p5_prod__523_comb | 32'h0000_0080;
  assign p5_or_149135_comb = p5_prod__528_comb | 32'h0000_0080;
  assign p5_or_149140_comb = p5_prod__587_comb | 32'h0000_0080;
  assign p5_or_149141_comb = p5_prod__592_comb | 32'h0000_0080;
  assign p5_or_149148_comb = p5_prod__715_comb | 32'h0000_0080;
  assign p5_or_149149_comb = p5_prod__720_comb | 32'h0000_0080;
  assign p5_or_149160_comb = p5_prod__843_comb | 32'h0000_0080;
  assign p5_or_149161_comb = p5_prod__848_comb | 32'h0000_0080;
  assign p5_or_149168_comb = p5_prod__971_comb | 32'h0000_0080;
  assign p5_or_149169_comb = p5_prod__976_comb | 32'h0000_0080;
  assign p5_or_149291_comb = p5_prod__525_comb | 32'h0000_0080;
  assign p5_or_149298_comb = p5_prod__556_comb | 32'h0000_0080;
  assign p5_or_149350_comb = p5_prod__545_comb | 32'h0000_0080;
  assign p5_or_149351_comb = p5_prod__563_comb | 32'h0000_0080;
  assign p5_or_149507_comb = p5_prod__547_comb | 32'h0000_0080;
  assign p5_or_149514_comb = p5_prod__575_comb | 32'h0000_0080;
  assign p5_sel_149547_comb = $signed(p5_shifted__64_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__64_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__64_squeezed_comb, p5_smul_57326_TrailingBits___64_comb};
  assign p5_sel_149548_comb = $signed(p5_shifted__65_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__65_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__65_squeezed_comb, p5_smul_57326_TrailingBits___65_comb};
  assign p5_sel_149549_comb = $signed(p5_shifted__66_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__66_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__66_squeezed_comb, p5_smul_57326_TrailingBits___66_comb};
  assign p5_sel_149550_comb = $signed(p5_shifted__67_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__67_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__67_squeezed_comb, p5_smul_57326_TrailingBits___67_comb};
  assign p5_sel_149551_comb = $signed(p5_shifted__68_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__68_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__68_squeezed_comb, p5_smul_57326_TrailingBits___68_comb};
  assign p5_sel_149552_comb = $signed(p5_shifted__69_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__69_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__69_squeezed_comb, p5_smul_57326_TrailingBits___69_comb};
  assign p5_sel_149553_comb = $signed(p5_shifted__70_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__70_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__70_squeezed_comb, p5_smul_57326_TrailingBits___70_comb};
  assign p5_sel_149554_comb = $signed(p5_shifted__71_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__71_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__71_squeezed_comb, p5_smul_57326_TrailingBits___71_comb};
  assign p5_sel_149555_comb = $signed(p5_shifted__96_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__96_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__96_squeezed_comb, p5_smul_57326_TrailingBits___96_comb};
  assign p5_sel_149556_comb = $signed(p5_shifted__97_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__97_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__97_squeezed_comb, p5_smul_57326_TrailingBits___97_comb};
  assign p5_sel_149557_comb = $signed(p5_shifted__98_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__98_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__98_squeezed_comb, p5_smul_57326_TrailingBits___98_comb};
  assign p5_sel_149558_comb = $signed(p5_shifted__99_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__99_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__99_squeezed_comb, p5_smul_57326_TrailingBits___99_comb};
  assign p5_sel_149559_comb = $signed(p5_shifted__100_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__100_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__100_squeezed_comb, p5_smul_57326_TrailingBits___100_comb};
  assign p5_sel_149560_comb = $signed(p5_shifted__101_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__101_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__101_squeezed_comb, p5_smul_57326_TrailingBits___101_comb};
  assign p5_sel_149561_comb = $signed(p5_shifted__102_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__102_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__102_squeezed_comb, p5_smul_57326_TrailingBits___102_comb};
  assign p5_sel_149562_comb = $signed(p5_shifted__103_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p5_shifted__103_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__103_squeezed_comb, p5_smul_57326_TrailingBits___103_comb};
  assign p5_shifted__72_comb = {~p4_clipped__9[7], p4_clipped__9[6:0], p5_smul_57326_TrailingBits___200_comb};
  assign p5_shifted__73_comb = {~p4_clipped__25[7], p4_clipped__25[6:0], p5_smul_57326_TrailingBits___201_comb};
  assign p5_shifted__74_comb = {~p4_clipped__41[7], p4_clipped__41[6:0], p5_smul_57326_TrailingBits___202_comb};
  assign p5_shifted__75_comb = {~p4_bit_slice_146165, p4_bit_slice_146191, p5_smul_57326_TrailingBits___203_comb};
  assign p5_shifted__76_comb = {~p4_bit_slice_146166, p4_bit_slice_146192, p5_smul_57326_TrailingBits___204_comb};
  assign p5_shifted__77_comb = {~p4_clipped__89[7], p4_clipped__89[6:0], p5_smul_57326_TrailingBits___205_comb};
  assign p5_shifted__78_comb = {~p4_clipped__105[7], p4_clipped__105[6:0], p5_smul_57326_TrailingBits___206_comb};
  assign p5_shifted__79_comb = {~p4_clipped__121[7], p4_clipped__121[6:0], p5_smul_57326_TrailingBits___207_comb};
  assign p5_shifted__80_comb = {~p4_clipped__10[7], p4_clipped__10[6:0], p5_smul_57326_TrailingBits___208_comb};
  assign p5_shifted__81_comb = {~p4_clipped__26[7], p4_clipped__26[6:0], p5_smul_57326_TrailingBits___209_comb};
  assign p5_shifted__82_comb = {~p4_clipped__42[7], p4_clipped__42[6:0], p5_smul_57326_TrailingBits___210_comb};
  assign p5_shifted__83_comb = {~p4_clipped__58[7], p4_clipped__58[6:0], p5_smul_57326_TrailingBits___211_comb};
  assign p5_shifted__84_comb = {~p4_clipped__74[7], p4_clipped__74[6:0], p5_smul_57326_TrailingBits___212_comb};
  assign p5_shifted__85_comb = {~p4_clipped__90[7], p4_clipped__90[6:0], p5_smul_57326_TrailingBits___213_comb};
  assign p5_shifted__86_comb = {~p4_clipped__106[7], p4_clipped__106[6:0], p5_smul_57326_TrailingBits___214_comb};
  assign p5_shifted__87_comb = {~p4_clipped__122[7], p4_clipped__122[6:0], p5_smul_57326_TrailingBits___215_comb};
  assign p5_shifted__88_comb = {~p4_clipped__11[7], p4_clipped__11[6:0], p5_smul_57326_TrailingBits___216_comb};
  assign p5_shifted__89_comb = {~p4_clipped__27[7], p4_clipped__27[6:0], p5_smul_57326_TrailingBits___217_comb};
  assign p5_shifted__90_comb = {~p4_clipped__43[7], p4_clipped__43[6:0], p5_smul_57326_TrailingBits___218_comb};
  assign p5_shifted__91_comb = {~p4_bit_slice_146167, p4_bit_slice_146193, p5_smul_57326_TrailingBits___219_comb};
  assign p5_shifted__92_comb = {~p4_bit_slice_146168, p4_bit_slice_146194, p5_smul_57326_TrailingBits___220_comb};
  assign p5_shifted__93_comb = {~p4_clipped__91[7], p4_clipped__91[6:0], p5_smul_57326_TrailingBits___221_comb};
  assign p5_shifted__94_comb = {~p4_clipped__107[7], p4_clipped__107[6:0], p5_smul_57326_TrailingBits___222_comb};
  assign p5_shifted__95_comb = {~p4_clipped__123[7], p4_clipped__123[6:0], p5_smul_57326_TrailingBits___223_comb};
  assign p5_shifted__104_comb = {~p4_clipped__13[7], p4_clipped__13[6:0], p5_smul_57326_TrailingBits___232_comb};
  assign p5_shifted__105_comb = {~p4_clipped__29[7], p4_clipped__29[6:0], p5_smul_57326_TrailingBits___233_comb};
  assign p5_shifted__106_comb = {~p4_clipped__45[7], p4_clipped__45[6:0], p5_smul_57326_TrailingBits___234_comb};
  assign p5_shifted__107_comb = {~p4_bit_slice_146175, p4_bit_slice_146207, p5_smul_57326_TrailingBits___235_comb};
  assign p5_shifted__108_comb = {~p4_bit_slice_146176, p4_bit_slice_146208, p5_smul_57326_TrailingBits___236_comb};
  assign p5_shifted__109_comb = {~p4_clipped__93[7], p4_clipped__93[6:0], p5_smul_57326_TrailingBits___237_comb};
  assign p5_shifted__110_comb = {~p4_clipped__109[7], p4_clipped__109[6:0], p5_smul_57326_TrailingBits___238_comb};
  assign p5_shifted__111_comb = {~p4_clipped__125[7], p4_clipped__125[6:0], p5_smul_57326_TrailingBits___239_comb};
  assign p5_shifted__112_comb = {~p4_clipped__14[7], p4_clipped__14[6:0], p5_smul_57326_TrailingBits___240_comb};
  assign p5_shifted__113_comb = {~p4_clipped__30[7], p4_clipped__30[6:0], p5_smul_57326_TrailingBits___241_comb};
  assign p5_shifted__114_comb = {~p4_clipped__46[7], p4_clipped__46[6:0], p5_smul_57326_TrailingBits___242_comb};
  assign p5_shifted__115_comb = {~p4_clipped__62[7], p4_clipped__62[6:0], p5_smul_57326_TrailingBits___243_comb};
  assign p5_shifted__116_comb = {~p4_clipped__78[7], p4_clipped__78[6:0], p5_smul_57326_TrailingBits___244_comb};
  assign p5_shifted__117_comb = {~p4_clipped__94[7], p4_clipped__94[6:0], p5_smul_57326_TrailingBits___245_comb};
  assign p5_shifted__118_comb = {~p4_clipped__110[7], p4_clipped__110[6:0], p5_smul_57326_TrailingBits___246_comb};
  assign p5_shifted__119_comb = {~p4_clipped__126[7], p4_clipped__126[6:0], p5_smul_57326_TrailingBits___247_comb};
  assign p5_shifted__120_comb = {~p4_clipped__15[7], p4_clipped__15[6:0], p5_smul_57326_TrailingBits___248_comb};
  assign p5_shifted__121_comb = {~p4_clipped__31[7], p4_clipped__31[6:0], p5_smul_57326_TrailingBits___249_comb};
  assign p5_shifted__122_comb = {~p4_clipped__47[7], p4_clipped__47[6:0], p5_smul_57326_TrailingBits___250_comb};
  assign p5_shifted__123_comb = {~p4_bit_slice_146177, p4_bit_slice_146209, p5_smul_57326_TrailingBits___251_comb};
  assign p5_shifted__124_comb = {~p4_bit_slice_146178, p4_bit_slice_146210, p5_smul_57326_TrailingBits___252_comb};
  assign p5_shifted__125_comb = {~p4_clipped__95[7], p4_clipped__95[6:0], p5_smul_57326_TrailingBits___253_comb};
  assign p5_shifted__126_comb = {~p4_clipped__111[7], p4_clipped__111[6:0], p5_smul_57326_TrailingBits___254_comb};
  assign p5_shifted__127_comb = {~p4_clipped__127[7], p4_clipped__127[6:0], p5_smul_57326_TrailingBits___255_comb};
  assign p5_prod__651_comb = {{9{p5_concat_147817_comb[22]}}, p5_concat_147817_comb};
  assign p5_prod__656_comb = {{9{p5_concat_147818_comb[22]}}, p5_concat_147818_comb};
  assign p5_prod__907_comb = {{9{p5_concat_147841_comb[22]}}, p5_concat_147841_comb};
  assign p5_prod__912_comb = {{9{p5_concat_147842_comb[22]}}, p5_concat_147842_comb};
  assign p5_or_148497_comb = p5_prod__581_comb | 32'h0000_0080;
  assign p5_or_148514_comb = p5_prod__619_comb | 32'h0000_0080;
  assign p5_or_148517_comb = p5_prod__645_comb | 32'h0000_0080;
  assign p5_or_148524_comb = p5_prod__657_comb | 32'h0000_0080;
  assign p5_or_148527_comb = p5_prod__663_comb | 32'h0000_0080;
  assign p5_or_148534_comb = p5_prod__683_comb | 32'h0000_0080;
  assign p5_or_148537_comb = p5_prod__709_comb | 32'h0000_0080;
  assign p5_or_148554_comb = p5_prod__747_comb | 32'h0000_0080;
  assign p5_or_148577_comb = p5_prod__837_comb | 32'h0000_0080;
  assign p5_or_148594_comb = p5_prod__875_comb | 32'h0000_0080;
  assign p5_or_148597_comb = p5_prod__901_comb | 32'h0000_0080;
  assign p5_or_148604_comb = p5_prod__913_comb | 32'h0000_0080;
  assign p5_or_148607_comb = p5_prod__919_comb | 32'h0000_0080;
  assign p5_or_148614_comb = p5_prod__939_comb | 32'h0000_0080;
  assign p5_or_148617_comb = p5_prod__965_comb | 32'h0000_0080;
  assign p5_or_148634_comb = p5_prod__1003_comb | 32'h0000_0080;
  assign p5_prod__589_comb = {{9{p5_concat_147953_comb[22]}}, p5_concat_147953_comb};
  assign p5_prod__620_comb = {{9{p5_concat_147958_comb[22]}}, p5_concat_147958_comb};
  assign p5_prod__653_comb = {{9{p5_concat_147959_comb[22]}}, p5_concat_147959_comb};
  assign p5_prod__684_comb = {{9{p5_concat_147964_comb[22]}}, p5_concat_147964_comb};
  assign p5_prod__717_comb = {{9{p5_concat_147965_comb[22]}}, p5_concat_147965_comb};
  assign p5_prod__748_comb = {{9{p5_concat_147970_comb[22]}}, p5_concat_147970_comb};
  assign p5_prod__845_comb = {{9{p5_concat_147977_comb[22]}}, p5_concat_147977_comb};
  assign p5_prod__876_comb = {{9{p5_concat_147982_comb[22]}}, p5_concat_147982_comb};
  assign p5_prod__909_comb = {{9{p5_concat_147983_comb[22]}}, p5_concat_147983_comb};
  assign p5_prod__940_comb = {{9{p5_concat_147988_comb[22]}}, p5_concat_147988_comb};
  assign p5_prod__973_comb = {{9{p5_concat_147989_comb[22]}}, p5_concat_147989_comb};
  assign p5_prod__1004_comb = {{9{p5_concat_147994_comb[22]}}, p5_concat_147994_comb};
  assign p5_prod__609_comb = {{9{p5_concat_148003_comb[22]}}, p5_concat_148003_comb};
  assign p5_prod__627_comb = {{9{p5_concat_148004_comb[22]}}, p5_concat_148004_comb};
  assign p5_prod__673_comb = {{9{p5_concat_148009_comb[22]}}, p5_concat_148009_comb};
  assign p5_prod__691_comb = {{9{p5_concat_148010_comb[22]}}, p5_concat_148010_comb};
  assign p5_prod__737_comb = {{9{p5_concat_148015_comb[22]}}, p5_concat_148015_comb};
  assign p5_prod__755_comb = {{9{p5_concat_148016_comb[22]}}, p5_concat_148016_comb};
  assign p5_prod__865_comb = {{9{p5_concat_148027_comb[22]}}, p5_concat_148027_comb};
  assign p5_prod__883_comb = {{9{p5_concat_148028_comb[22]}}, p5_concat_148028_comb};
  assign p5_prod__929_comb = {{9{p5_concat_148033_comb[22]}}, p5_concat_148033_comb};
  assign p5_prod__947_comb = {{9{p5_concat_148034_comb[22]}}, p5_concat_148034_comb};
  assign p5_prod__993_comb = {{9{p5_concat_148039_comb[22]}}, p5_concat_148039_comb};
  assign p5_prod__1011_comb = {{9{p5_concat_148040_comb[22]}}, p5_concat_148040_comb};
  assign p5_or_148819_comb = p5_prod__610_comb | 32'h0000_0080;
  assign p5_or_148832_comb = p5_prod__635_comb | 32'h0000_0080;
  assign p5_or_148839_comb = p5_prod__674_comb | 32'h0000_0080;
  assign p5_or_148844_comb = p5_prod__687_comb | 32'h0000_0080;
  assign p5_or_148847_comb = p5_prod__692_comb | 32'h0000_0080;
  assign p5_or_148852_comb = p5_prod__699_comb | 32'h0000_0080;
  assign p5_or_148859_comb = p5_prod__738_comb | 32'h0000_0080;
  assign p5_or_148872_comb = p5_prod__763_comb | 32'h0000_0080;
  assign p5_or_148899_comb = p5_prod__866_comb | 32'h0000_0080;
  assign p5_or_148912_comb = p5_prod__891_comb | 32'h0000_0080;
  assign p5_or_148919_comb = p5_prod__930_comb | 32'h0000_0080;
  assign p5_or_148924_comb = p5_prod__943_comb | 32'h0000_0080;
  assign p5_or_148927_comb = p5_prod__948_comb | 32'h0000_0080;
  assign p5_or_148932_comb = p5_prod__955_comb | 32'h0000_0080;
  assign p5_or_148939_comb = p5_prod__994_comb | 32'h0000_0080;
  assign p5_or_148952_comb = p5_prod__1019_comb | 32'h0000_0080;
  assign p5_prod__611_comb = {{9{p5_concat_148145_comb[22]}}, p5_concat_148145_comb};
  assign p5_prod__639_comb = {{9{p5_concat_148150_comb[22]}}, p5_concat_148150_comb};
  assign p5_prod__675_comb = {{9{p5_concat_148151_comb[22]}}, p5_concat_148151_comb};
  assign p5_prod__703_comb = {{9{p5_concat_148156_comb[22]}}, p5_concat_148156_comb};
  assign p5_prod__739_comb = {{9{p5_concat_148157_comb[22]}}, p5_concat_148157_comb};
  assign p5_prod__767_comb = {{9{p5_concat_148162_comb[22]}}, p5_concat_148162_comb};
  assign p5_prod__867_comb = {{9{p5_concat_148169_comb[22]}}, p5_concat_148169_comb};
  assign p5_prod__895_comb = {{9{p5_concat_148174_comb[22]}}, p5_concat_148174_comb};
  assign p5_prod__931_comb = {{9{p5_concat_148175_comb[22]}}, p5_concat_148175_comb};
  assign p5_prod__959_comb = {{9{p5_concat_148180_comb[22]}}, p5_concat_148180_comb};
  assign p5_prod__995_comb = {{9{p5_concat_148181_comb[22]}}, p5_concat_148181_comb};
  assign p5_prod__1023_comb = {{9{p5_concat_148186_comb[22]}}, p5_concat_148186_comb};
  assign p5_sel_148221_comb = $signed(p5_shifted__72_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__72_squeezed_comb;
  assign p5_sel_148224_comb = $signed(p5_shifted__73_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__73_squeezed_comb;
  assign p5_sel_148227_comb = $signed(p5_shifted__74_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__74_squeezed_comb;
  assign p5_sel_148230_comb = $signed(p5_shifted__75_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__75_squeezed_comb;
  assign p5_sel_148233_comb = $signed(p5_shifted__76_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__76_squeezed_comb;
  assign p5_sel_148236_comb = $signed(p5_shifted__77_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__77_squeezed_comb;
  assign p5_sel_148239_comb = $signed(p5_shifted__78_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__78_squeezed_comb;
  assign p5_sel_148242_comb = $signed(p5_shifted__79_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__79_squeezed_comb;
  assign p5_sel_148245_comb = $signed(p5_shifted__80_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__80_squeezed_comb;
  assign p5_sel_148248_comb = $signed(p5_shifted__81_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__81_squeezed_comb;
  assign p5_sel_148251_comb = $signed(p5_shifted__82_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__82_squeezed_comb;
  assign p5_sel_148254_comb = $signed(p5_shifted__83_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__83_squeezed_comb;
  assign p5_sel_148257_comb = $signed(p5_shifted__84_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__84_squeezed_comb;
  assign p5_sel_148260_comb = $signed(p5_shifted__85_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__85_squeezed_comb;
  assign p5_sel_148263_comb = $signed(p5_shifted__86_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__86_squeezed_comb;
  assign p5_sel_148266_comb = $signed(p5_shifted__87_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__87_squeezed_comb;
  assign p5_sel_148269_comb = $signed(p5_shifted__88_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__88_squeezed_comb;
  assign p5_sel_148272_comb = $signed(p5_shifted__89_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__89_squeezed_comb;
  assign p5_sel_148275_comb = $signed(p5_shifted__90_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__90_squeezed_comb;
  assign p5_sel_148278_comb = $signed(p5_shifted__91_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__91_squeezed_comb;
  assign p5_sel_148281_comb = $signed(p5_shifted__92_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__92_squeezed_comb;
  assign p5_sel_148284_comb = $signed(p5_shifted__93_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__93_squeezed_comb;
  assign p5_sel_148287_comb = $signed(p5_shifted__94_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__94_squeezed_comb;
  assign p5_sel_148290_comb = $signed(p5_shifted__95_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__95_squeezed_comb;
  assign p5_sel_148325_comb = $signed(p5_shifted__104_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__104_squeezed_comb;
  assign p5_sel_148328_comb = $signed(p5_shifted__105_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__105_squeezed_comb;
  assign p5_sel_148331_comb = $signed(p5_shifted__106_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__106_squeezed_comb;
  assign p5_sel_148334_comb = $signed(p5_shifted__107_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__107_squeezed_comb;
  assign p5_sel_148337_comb = $signed(p5_shifted__108_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__108_squeezed_comb;
  assign p5_sel_148340_comb = $signed(p5_shifted__109_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__109_squeezed_comb;
  assign p5_sel_148343_comb = $signed(p5_shifted__110_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__110_squeezed_comb;
  assign p5_sel_148346_comb = $signed(p5_shifted__111_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__111_squeezed_comb;
  assign p5_sel_148349_comb = $signed(p5_shifted__112_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__112_squeezed_comb;
  assign p5_sel_148352_comb = $signed(p5_shifted__113_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__113_squeezed_comb;
  assign p5_sel_148355_comb = $signed(p5_shifted__114_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__114_squeezed_comb;
  assign p5_sel_148358_comb = $signed(p5_shifted__115_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__115_squeezed_comb;
  assign p5_sel_148361_comb = $signed(p5_shifted__116_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__116_squeezed_comb;
  assign p5_sel_148364_comb = $signed(p5_shifted__117_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__117_squeezed_comb;
  assign p5_sel_148367_comb = $signed(p5_shifted__118_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__118_squeezed_comb;
  assign p5_sel_148370_comb = $signed(p5_shifted__119_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__119_squeezed_comb;
  assign p5_sel_148373_comb = $signed(p5_shifted__120_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__120_squeezed_comb;
  assign p5_sel_148376_comb = $signed(p5_shifted__121_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__121_squeezed_comb;
  assign p5_sel_148379_comb = $signed(p5_shifted__122_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__122_squeezed_comb;
  assign p5_sel_148382_comb = $signed(p5_shifted__123_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__123_squeezed_comb;
  assign p5_sel_148385_comb = $signed(p5_shifted__124_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__124_squeezed_comb;
  assign p5_sel_148388_comb = $signed(p5_shifted__125_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__125_squeezed_comb;
  assign p5_sel_148391_comb = $signed(p5_shifted__126_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__126_squeezed_comb;
  assign p5_sel_148394_comb = $signed(p5_shifted__127_squeezed_comb) < $signed(8'h80) ? 8'h80 : p5_shifted__127_squeezed_comb;
  assign p5_or_148407_comb = p5_prod__583_comb | 32'h0000_0080;
  assign p5_or_148414_comb = p5_prod__598_comb | 32'h0000_0080;
  assign p5_or_148417_comb = p5_prod__647_comb | 32'h0000_0080;
  assign p5_or_148424_comb = p5_prod__662_comb | 32'h0000_0080;
  assign p5_or_148427_comb = p5_prod__711_comb | 32'h0000_0080;
  assign p5_or_148434_comb = p5_prod__726_comb | 32'h0000_0080;
  assign p5_or_148447_comb = p5_prod__839_comb | 32'h0000_0080;
  assign p5_or_148454_comb = p5_prod__854_comb | 32'h0000_0080;
  assign p5_or_148457_comb = p5_prod__903_comb | 32'h0000_0080;
  assign p5_or_148464_comb = p5_prod__918_comb | 32'h0000_0080;
  assign p5_or_148467_comb = p5_prod__967_comb | 32'h0000_0080;
  assign p5_or_148474_comb = p5_prod__982_comb | 32'h0000_0080;
  assign p5_or_148659_comb = p5_prod__664_comb | 32'h0000_0080;
  assign p5_or_148662_comb = p5_prod__671_comb | 32'h0000_0080;
  assign p5_or_148699_comb = p5_prod__920_comb | 32'h0000_0080;
  assign p5_or_148702_comb = p5_prod__927_comb | 32'h0000_0080;
  assign p5_or_148727_comb = p5_prod__596_comb | 32'h0000_0080;
  assign p5_or_148734_comb = p5_prod__634_comb | 32'h0000_0080;
  assign p5_or_148737_comb = p5_prod__660_comb | 32'h0000_0080;
  assign p5_or_148744_comb = p5_prod__698_comb | 32'h0000_0080;
  assign p5_or_148747_comb = p5_prod__724_comb | 32'h0000_0080;
  assign p5_or_148754_comb = p5_prod__762_comb | 32'h0000_0080;
  assign p5_or_148767_comb = p5_prod__852_comb | 32'h0000_0080;
  assign p5_or_148774_comb = p5_prod__890_comb | 32'h0000_0080;
  assign p5_or_148777_comb = p5_prod__916_comb | 32'h0000_0080;
  assign p5_or_148784_comb = p5_prod__954_comb | 32'h0000_0080;
  assign p5_or_148787_comb = p5_prod__980_comb | 32'h0000_0080;
  assign p5_or_148794_comb = p5_prod__1018_comb | 32'h0000_0080;
  assign p5_or_148969_comb = p5_prod__618_comb | 32'h0000_0080;
  assign p5_or_148972_comb = p5_prod__638_comb | 32'h0000_0080;
  assign p5_or_148979_comb = p5_prod__682_comb | 32'h0000_0080;
  assign p5_or_148982_comb = p5_prod__702_comb | 32'h0000_0080;
  assign p5_or_148989_comb = p5_prod__746_comb | 32'h0000_0080;
  assign p5_or_148992_comb = p5_prod__766_comb | 32'h0000_0080;
  assign p5_or_149009_comb = p5_prod__874_comb | 32'h0000_0080;
  assign p5_or_149012_comb = p5_prod__894_comb | 32'h0000_0080;
  assign p5_or_149019_comb = p5_prod__938_comb | 32'h0000_0080;
  assign p5_or_149022_comb = p5_prod__958_comb | 32'h0000_0080;
  assign p5_or_149029_comb = p5_prod__1002_comb | 32'h0000_0080;
  assign p5_or_149032_comb = p5_prod__1022_comb | 32'h0000_0080;
  assign p5_sgt_149059_comb = $signed(p5_shifted__72_comb) > $signed(16'h7fff);
  assign p5_sgt_149060_comb = $signed(p5_shifted__73_comb) > $signed(16'h7fff);
  assign p5_sgt_149061_comb = $signed(p5_shifted__74_comb) > $signed(16'h7fff);
  assign p5_sgt_149062_comb = $signed(p5_shifted__75_comb) > $signed(16'h7fff);
  assign p5_sgt_149063_comb = $signed(p5_shifted__76_comb) > $signed(16'h7fff);
  assign p5_sgt_149064_comb = $signed(p5_shifted__77_comb) > $signed(16'h7fff);
  assign p5_sgt_149065_comb = $signed(p5_shifted__78_comb) > $signed(16'h7fff);
  assign p5_sgt_149066_comb = $signed(p5_shifted__79_comb) > $signed(16'h7fff);
  assign p5_sgt_149067_comb = $signed(p5_shifted__80_comb) > $signed(16'h7fff);
  assign p5_sgt_149068_comb = $signed(p5_shifted__81_comb) > $signed(16'h7fff);
  assign p5_sgt_149069_comb = $signed(p5_shifted__82_comb) > $signed(16'h7fff);
  assign p5_sgt_149070_comb = $signed(p5_shifted__83_comb) > $signed(16'h7fff);
  assign p5_sgt_149071_comb = $signed(p5_shifted__84_comb) > $signed(16'h7fff);
  assign p5_sgt_149072_comb = $signed(p5_shifted__85_comb) > $signed(16'h7fff);
  assign p5_sgt_149073_comb = $signed(p5_shifted__86_comb) > $signed(16'h7fff);
  assign p5_sgt_149074_comb = $signed(p5_shifted__87_comb) > $signed(16'h7fff);
  assign p5_sgt_149075_comb = $signed(p5_shifted__88_comb) > $signed(16'h7fff);
  assign p5_sgt_149076_comb = $signed(p5_shifted__89_comb) > $signed(16'h7fff);
  assign p5_sgt_149077_comb = $signed(p5_shifted__90_comb) > $signed(16'h7fff);
  assign p5_sgt_149078_comb = $signed(p5_shifted__91_comb) > $signed(16'h7fff);
  assign p5_sgt_149079_comb = $signed(p5_shifted__92_comb) > $signed(16'h7fff);
  assign p5_sgt_149080_comb = $signed(p5_shifted__93_comb) > $signed(16'h7fff);
  assign p5_sgt_149081_comb = $signed(p5_shifted__94_comb) > $signed(16'h7fff);
  assign p5_sgt_149082_comb = $signed(p5_shifted__95_comb) > $signed(16'h7fff);
  assign p5_sgt_149107_comb = $signed(p5_shifted__104_comb) > $signed(16'h7fff);
  assign p5_sgt_149108_comb = $signed(p5_shifted__105_comb) > $signed(16'h7fff);
  assign p5_sgt_149109_comb = $signed(p5_shifted__106_comb) > $signed(16'h7fff);
  assign p5_sgt_149110_comb = $signed(p5_shifted__107_comb) > $signed(16'h7fff);
  assign p5_sgt_149111_comb = $signed(p5_shifted__108_comb) > $signed(16'h7fff);
  assign p5_sgt_149112_comb = $signed(p5_shifted__109_comb) > $signed(16'h7fff);
  assign p5_sgt_149113_comb = $signed(p5_shifted__110_comb) > $signed(16'h7fff);
  assign p5_sgt_149114_comb = $signed(p5_shifted__111_comb) > $signed(16'h7fff);
  assign p5_sgt_149115_comb = $signed(p5_shifted__112_comb) > $signed(16'h7fff);
  assign p5_sgt_149116_comb = $signed(p5_shifted__113_comb) > $signed(16'h7fff);
  assign p5_sgt_149117_comb = $signed(p5_shifted__114_comb) > $signed(16'h7fff);
  assign p5_sgt_149118_comb = $signed(p5_shifted__115_comb) > $signed(16'h7fff);
  assign p5_sgt_149119_comb = $signed(p5_shifted__116_comb) > $signed(16'h7fff);
  assign p5_sgt_149120_comb = $signed(p5_shifted__117_comb) > $signed(16'h7fff);
  assign p5_sgt_149121_comb = $signed(p5_shifted__118_comb) > $signed(16'h7fff);
  assign p5_sgt_149122_comb = $signed(p5_shifted__119_comb) > $signed(16'h7fff);
  assign p5_sgt_149123_comb = $signed(p5_shifted__120_comb) > $signed(16'h7fff);
  assign p5_sgt_149124_comb = $signed(p5_shifted__121_comb) > $signed(16'h7fff);
  assign p5_sgt_149125_comb = $signed(p5_shifted__122_comb) > $signed(16'h7fff);
  assign p5_sgt_149126_comb = $signed(p5_shifted__123_comb) > $signed(16'h7fff);
  assign p5_sgt_149127_comb = $signed(p5_shifted__124_comb) > $signed(16'h7fff);
  assign p5_sgt_149128_comb = $signed(p5_shifted__125_comb) > $signed(16'h7fff);
  assign p5_sgt_149129_comb = $signed(p5_shifted__126_comb) > $signed(16'h7fff);
  assign p5_sgt_149130_comb = $signed(p5_shifted__127_comb) > $signed(16'h7fff);
  assign p5_slt_149139_comb = $signed(p5_prod__583_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149142_comb = $signed(p5_prod__598_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149143_comb = $signed(p5_prod__647_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149144_comb = p5_prod__651_comb | 32'h0000_0080;
  assign p5_or_149145_comb = p5_prod__656_comb | 32'h0000_0080;
  assign p5_slt_149146_comb = $signed(p5_prod__662_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149147_comb = $signed(p5_prod__711_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149150_comb = $signed(p5_prod__726_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149159_comb = $signed(p5_prod__839_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149162_comb = $signed(p5_prod__854_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149163_comb = $signed(p5_prod__903_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149164_comb = p5_prod__907_comb | 32'h0000_0080;
  assign p5_or_149165_comb = p5_prod__912_comb | 32'h0000_0080;
  assign p5_slt_149166_comb = $signed(p5_prod__918_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149167_comb = $signed(p5_prod__967_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149170_comb = $signed(p5_prod__982_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149191_comb = $signed(p5_prod__581_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149192_comb = p5_or_148497_comb[23:10];
  assign p5_slt_149193_comb = $signed(p5_prod__584_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149194_comb = $signed(p5_prod__588_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149201_comb = $signed(p5_prod__606_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149202_comb = $signed(p5_prod__613_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149203_comb = $signed(p5_prod__619_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149204_comb = p5_or_148514_comb[23:10];
  assign p5_slt_149205_comb = $signed(p5_prod__645_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149206_comb = p5_or_148517_comb[23:10];
  assign p5_slt_149207_comb = $signed(p5_prod__648_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149208_comb = $signed(p5_prod__652_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149209_comb = $signed(p5_prod__657_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149210_comb = p5_or_148524_comb[23:10];
  assign p5_slt_149211_comb = $signed(p5_prod__663_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149212_comb = p5_or_148527_comb[23:10];
  assign p5_slt_149213_comb = $signed(p5_prod__670_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149214_comb = $signed(p5_prod__677_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149215_comb = $signed(p5_prod__683_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149216_comb = p5_or_148534_comb[23:10];
  assign p5_slt_149217_comb = $signed(p5_prod__709_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149218_comb = p5_or_148537_comb[23:10];
  assign p5_slt_149219_comb = $signed(p5_prod__712_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149220_comb = $signed(p5_prod__716_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149227_comb = $signed(p5_prod__734_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149228_comb = $signed(p5_prod__741_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149229_comb = $signed(p5_prod__747_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149230_comb = p5_or_148554_comb[23:10];
  assign p5_slt_149251_comb = $signed(p5_prod__837_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149252_comb = p5_or_148577_comb[23:10];
  assign p5_slt_149253_comb = $signed(p5_prod__840_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149254_comb = $signed(p5_prod__844_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149261_comb = $signed(p5_prod__862_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149262_comb = $signed(p5_prod__869_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149263_comb = $signed(p5_prod__875_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149264_comb = p5_or_148594_comb[23:10];
  assign p5_slt_149265_comb = $signed(p5_prod__901_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149266_comb = p5_or_148597_comb[23:10];
  assign p5_slt_149267_comb = $signed(p5_prod__904_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149268_comb = $signed(p5_prod__908_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149269_comb = $signed(p5_prod__913_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149270_comb = p5_or_148604_comb[23:10];
  assign p5_slt_149271_comb = $signed(p5_prod__919_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149272_comb = p5_or_148607_comb[23:10];
  assign p5_slt_149273_comb = $signed(p5_prod__926_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149274_comb = $signed(p5_prod__933_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149275_comb = $signed(p5_prod__939_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149276_comb = p5_or_148614_comb[23:10];
  assign p5_slt_149277_comb = $signed(p5_prod__965_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149278_comb = p5_or_148617_comb[23:10];
  assign p5_slt_149279_comb = $signed(p5_prod__968_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149280_comb = $signed(p5_prod__972_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149287_comb = $signed(p5_prod__990_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149288_comb = $signed(p5_prod__997_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149289_comb = $signed(p5_prod__1003_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149290_comb = p5_or_148634_comb[23:10];
  assign p5_or_149299_comb = p5_prod__589_comb | 32'h0000_0080;
  assign p5_or_149306_comb = p5_prod__620_comb | 32'h0000_0080;
  assign p5_or_149307_comb = p5_prod__653_comb | 32'h0000_0080;
  assign p5_slt_149308_comb = $signed(p5_prod__664_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149309_comb = $signed(p5_prod__671_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149310_comb = p5_prod__684_comb | 32'h0000_0080;
  assign p5_or_149311_comb = p5_prod__717_comb | 32'h0000_0080;
  assign p5_or_149318_comb = p5_prod__748_comb | 32'h0000_0080;
  assign p5_or_149327_comb = p5_prod__845_comb | 32'h0000_0080;
  assign p5_or_149334_comb = p5_prod__876_comb | 32'h0000_0080;
  assign p5_or_149335_comb = p5_prod__909_comb | 32'h0000_0080;
  assign p5_slt_149336_comb = $signed(p5_prod__920_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149337_comb = $signed(p5_prod__927_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149338_comb = p5_prod__940_comb | 32'h0000_0080;
  assign p5_or_149339_comb = p5_prod__973_comb | 32'h0000_0080;
  assign p5_or_149346_comb = p5_prod__1004_comb | 32'h0000_0080;
  assign p5_slt_149355_comb = $signed(p5_prod__596_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149356_comb = p5_prod__609_comb | 32'h0000_0080;
  assign p5_or_149357_comb = p5_prod__627_comb | 32'h0000_0080;
  assign p5_slt_149358_comb = $signed(p5_prod__634_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149359_comb = $signed(p5_prod__660_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149360_comb = p5_prod__673_comb | 32'h0000_0080;
  assign p5_or_149361_comb = p5_prod__691_comb | 32'h0000_0080;
  assign p5_slt_149362_comb = $signed(p5_prod__698_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149363_comb = $signed(p5_prod__724_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149364_comb = p5_prod__737_comb | 32'h0000_0080;
  assign p5_or_149365_comb = p5_prod__755_comb | 32'h0000_0080;
  assign p5_slt_149366_comb = $signed(p5_prod__762_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149375_comb = $signed(p5_prod__852_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149376_comb = p5_prod__865_comb | 32'h0000_0080;
  assign p5_or_149377_comb = p5_prod__883_comb | 32'h0000_0080;
  assign p5_slt_149378_comb = $signed(p5_prod__890_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149379_comb = $signed(p5_prod__916_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149380_comb = p5_prod__929_comb | 32'h0000_0080;
  assign p5_or_149381_comb = p5_prod__947_comb | 32'h0000_0080;
  assign p5_slt_149382_comb = $signed(p5_prod__954_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149383_comb = $signed(p5_prod__980_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149384_comb = p5_prod__993_comb | 32'h0000_0080;
  assign p5_or_149385_comb = p5_prod__1011_comb | 32'h0000_0080;
  assign p5_slt_149386_comb = $signed(p5_prod__1018_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149407_comb = $signed(p5_prod__603_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149408_comb = $signed(p5_prod__610_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149409_comb = p5_or_148819_comb[23:10];
  assign p5_slt_149410_comb = $signed(p5_prod__617_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149417_comb = $signed(p5_prod__632_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149418_comb = $signed(p5_prod__635_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149419_comb = p5_or_148832_comb[23:10];
  assign p5_slt_149420_comb = $signed(p5_prod__637_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149421_comb = $signed(p5_prod__667_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149422_comb = $signed(p5_prod__674_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149423_comb = p5_or_148839_comb[23:10];
  assign p5_slt_149424_comb = $signed(p5_prod__681_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149425_comb = $signed(p5_prod__687_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149426_comb = p5_or_148844_comb[23:10];
  assign p5_slt_149427_comb = $signed(p5_prod__692_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149428_comb = p5_or_148847_comb[23:10];
  assign p5_slt_149429_comb = $signed(p5_prod__696_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149430_comb = $signed(p5_prod__699_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149431_comb = p5_or_148852_comb[23:10];
  assign p5_slt_149432_comb = $signed(p5_prod__701_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149433_comb = $signed(p5_prod__731_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149434_comb = $signed(p5_prod__738_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149435_comb = p5_or_148859_comb[23:10];
  assign p5_slt_149436_comb = $signed(p5_prod__745_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149443_comb = $signed(p5_prod__760_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149444_comb = $signed(p5_prod__763_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149445_comb = p5_or_148872_comb[23:10];
  assign p5_slt_149446_comb = $signed(p5_prod__765_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149467_comb = $signed(p5_prod__859_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149468_comb = $signed(p5_prod__866_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149469_comb = p5_or_148899_comb[23:10];
  assign p5_slt_149470_comb = $signed(p5_prod__873_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149477_comb = $signed(p5_prod__888_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149478_comb = $signed(p5_prod__891_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149479_comb = p5_or_148912_comb[23:10];
  assign p5_slt_149480_comb = $signed(p5_prod__893_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149481_comb = $signed(p5_prod__923_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149482_comb = $signed(p5_prod__930_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149483_comb = p5_or_148919_comb[23:10];
  assign p5_slt_149484_comb = $signed(p5_prod__937_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149485_comb = $signed(p5_prod__943_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149486_comb = p5_or_148924_comb[23:10];
  assign p5_slt_149487_comb = $signed(p5_prod__948_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149488_comb = p5_or_148927_comb[23:10];
  assign p5_slt_149489_comb = $signed(p5_prod__952_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149490_comb = $signed(p5_prod__955_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149491_comb = p5_or_148932_comb[23:10];
  assign p5_slt_149492_comb = $signed(p5_prod__957_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149493_comb = $signed(p5_prod__987_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149494_comb = $signed(p5_prod__994_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149495_comb = p5_or_148939_comb[23:10];
  assign p5_slt_149496_comb = $signed(p5_prod__1001_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149503_comb = $signed(p5_prod__1016_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149504_comb = $signed(p5_prod__1019_comb[31:10]) < $signed(22'h3f_e000);
  assign p5_bit_slice_149505_comb = p5_or_148952_comb[23:10];
  assign p5_slt_149506_comb = $signed(p5_prod__1021_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149515_comb = p5_prod__611_comb | 32'h0000_0080;
  assign p5_slt_149516_comb = $signed(p5_prod__618_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149517_comb = $signed(p5_prod__638_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149518_comb = p5_prod__639_comb | 32'h0000_0080;
  assign p5_or_149519_comb = p5_prod__675_comb | 32'h0000_0080;
  assign p5_slt_149520_comb = $signed(p5_prod__682_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149521_comb = $signed(p5_prod__702_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149522_comb = p5_prod__703_comb | 32'h0000_0080;
  assign p5_or_149523_comb = p5_prod__739_comb | 32'h0000_0080;
  assign p5_slt_149524_comb = $signed(p5_prod__746_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149525_comb = $signed(p5_prod__766_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149526_comb = p5_prod__767_comb | 32'h0000_0080;
  assign p5_or_149535_comb = p5_prod__867_comb | 32'h0000_0080;
  assign p5_slt_149536_comb = $signed(p5_prod__874_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149537_comb = $signed(p5_prod__894_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149538_comb = p5_prod__895_comb | 32'h0000_0080;
  assign p5_or_149539_comb = p5_prod__931_comb | 32'h0000_0080;
  assign p5_slt_149540_comb = $signed(p5_prod__938_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149541_comb = $signed(p5_prod__958_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149542_comb = p5_prod__959_comb | 32'h0000_0080;
  assign p5_or_149543_comb = p5_prod__995_comb | 32'h0000_0080;
  assign p5_slt_149544_comb = $signed(p5_prod__1002_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_slt_149545_comb = $signed(p5_prod__1022_comb[31:9]) < $signed(23'h7f_c000);
  assign p5_or_149546_comb = p5_prod__1023_comb | 32'h0000_0080;
  assign p5_sel_149565_comb = $signed(p5_prod__519_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148397_comb[23:9];
  assign p5_bit_slice_149568_comb = p5_or_149134_comb[23:9];
  assign p5_bit_slice_149571_comb = p5_or_149135_comb[23:9];
  assign p5_sel_149574_comb = $signed(p5_prod__534_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148404_comb[23:9];
  assign p5_bit_slice_149577_comb = p5_or_149140_comb[23:9];
  assign p5_bit_slice_149580_comb = p5_or_149141_comb[23:9];
  assign p5_bit_slice_149583_comb = p5_or_149148_comb[23:9];
  assign p5_bit_slice_149586_comb = p5_or_149149_comb[23:9];
  assign p5_sel_149589_comb = $signed(p5_prod__775_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148437_comb[23:9];
  assign p5_sel_149600_comb = $signed(p5_prod__790_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148444_comb[23:9];
  assign p5_bit_slice_149603_comb = p5_or_149160_comb[23:9];
  assign p5_bit_slice_149606_comb = p5_or_149161_comb[23:9];
  assign p5_bit_slice_149609_comb = p5_or_149168_comb[23:9];
  assign p5_bit_slice_149612_comb = p5_or_149169_comb[23:9];
  assign p5_sel_149615_comb = $signed(p5_prod__517_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148477_comb[23:10];
  assign p5_sel_149618_comb = $signed(p5_prod__520_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58352_NarrowedMult__comb;
  assign p5_sel_149621_comb = $signed(p5_prod__524_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58354_NarrowedMult__comb;
  assign p5_sel_149624_comb = $signed(p5_prod__529_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148484_comb[23:10];
  assign p5_sel_149627_comb = $signed(p5_prod__535_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148487_comb[23:10];
  assign p5_sel_149630_comb = $signed(p5_prod__542_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58360_NarrowedMult__comb;
  assign p5_sel_149633_comb = $signed(p5_prod__549_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58362_NarrowedMult__comb;
  assign p5_sel_149636_comb = $signed(p5_prod__555_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148494_comb[23:10];
  assign p5_bit_slice_149637_comb = p5_or_148497_comb[31:8];
  assign p5_sel_149644_comb = $signed(p5_prod__593_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148504_comb[23:10];
  assign p5_sel_149647_comb = $signed(p5_prod__599_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148507_comb[23:10];
  assign p5_bit_slice_149652_comb = p5_or_148514_comb[31:8];
  assign p5_bit_slice_149653_comb = p5_or_148517_comb[31:8];
  assign p5_bit_slice_149658_comb = p5_or_148524_comb[31:8];
  assign p5_bit_slice_149659_comb = p5_or_148527_comb[31:8];
  assign p5_bit_slice_149664_comb = p5_or_148534_comb[31:8];
  assign p5_bit_slice_149665_comb = p5_or_148537_comb[31:8];
  assign p5_sel_149672_comb = $signed(p5_prod__721_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148544_comb[23:10];
  assign p5_sel_149675_comb = $signed(p5_prod__727_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148547_comb[23:10];
  assign p5_bit_slice_149680_comb = p5_or_148554_comb[31:8];
  assign p5_sel_149683_comb = $signed(p5_prod__773_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148557_comb[23:10];
  assign p5_sel_149686_comb = $signed(p5_prod__776_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58416_NarrowedMult__comb;
  assign p5_sel_149689_comb = $signed(p5_prod__780_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58418_NarrowedMult__comb;
  assign p5_sel_149692_comb = $signed(p5_prod__785_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148564_comb[23:10];
  assign p5_sel_149695_comb = $signed(p5_prod__791_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148567_comb[23:10];
  assign p5_sel_149698_comb = $signed(p5_prod__798_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58424_NarrowedMult__comb;
  assign p5_sel_149701_comb = $signed(p5_prod__805_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58426_NarrowedMult__comb;
  assign p5_sel_149704_comb = $signed(p5_prod__811_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148574_comb[23:10];
  assign p5_bit_slice_149705_comb = p5_or_148577_comb[31:8];
  assign p5_sel_149712_comb = $signed(p5_prod__849_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148584_comb[23:10];
  assign p5_sel_149715_comb = $signed(p5_prod__855_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148587_comb[23:10];
  assign p5_bit_slice_149720_comb = p5_or_148594_comb[31:8];
  assign p5_bit_slice_149721_comb = p5_or_148597_comb[31:8];
  assign p5_bit_slice_149726_comb = p5_or_148604_comb[31:8];
  assign p5_bit_slice_149727_comb = p5_or_148607_comb[31:8];
  assign p5_bit_slice_149732_comb = p5_or_148614_comb[31:8];
  assign p5_bit_slice_149733_comb = p5_or_148617_comb[31:8];
  assign p5_sel_149740_comb = $signed(p5_prod__977_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148624_comb[23:10];
  assign p5_sel_149743_comb = $signed(p5_prod__983_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148627_comb[23:10];
  assign p5_bit_slice_149748_comb = p5_or_148634_comb[31:8];
  assign p5_bit_slice_149751_comb = p5_or_149291_comb[23:9];
  assign p5_sel_149754_comb = $signed(p5_prod__536_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148639_comb[23:9];
  assign p5_sel_149757_comb = $signed(p5_prod__543_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148642_comb[23:9];
  assign p5_bit_slice_149760_comb = p5_or_149298_comb[23:9];
  assign p5_sel_149763_comb = $signed(p5_prod__600_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148649_comb[23:9];
  assign p5_sel_149766_comb = $signed(p5_prod__607_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148652_comb[23:9];
  assign p5_sel_149769_comb = $signed(p5_prod__728_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148669_comb[23:9];
  assign p5_sel_149772_comb = $signed(p5_prod__735_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148672_comb[23:9];
  assign p5_sel_149779_comb = $signed(p5_prod__792_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148679_comb[23:9];
  assign p5_sel_149782_comb = $signed(p5_prod__799_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148682_comb[23:9];
  assign p5_sel_149789_comb = $signed(p5_prod__856_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148689_comb[23:9];
  assign p5_sel_149792_comb = $signed(p5_prod__863_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148692_comb[23:9];
  assign p5_sel_149795_comb = $signed(p5_prod__984_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148709_comb[23:9];
  assign p5_sel_149798_comb = $signed(p5_prod__991_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148712_comb[23:9];
  assign p5_sel_149801_comb = $signed(p5_prod__532_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148717_comb[23:9];
  assign p5_bit_slice_149804_comb = p5_or_149350_comb[23:9];
  assign p5_bit_slice_149807_comb = p5_or_149351_comb[23:9];
  assign p5_sel_149810_comb = $signed(p5_prod__570_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148724_comb[23:9];
  assign p5_sel_149813_comb = $signed(p5_prod__788_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148757_comb[23:9];
  assign p5_sel_149824_comb = $signed(p5_prod__826_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148764_comb[23:9];
  assign p5_sel_149827_comb = $signed(p5_prod__539_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58862_NarrowedMult__comb;
  assign p5_sel_149830_comb = $signed(p5_prod__546_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148799_comb[23:10];
  assign p5_sel_149833_comb = $signed(p5_prod__553_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58866_NarrowedMult__comb;
  assign p5_sel_149836_comb = $signed(p5_prod__559_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148804_comb[23:10];
  assign p5_sel_149839_comb = $signed(p5_prod__564_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148807_comb[23:10];
  assign p5_sel_149842_comb = $signed(p5_prod__568_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58872_NarrowedMult__comb;
  assign p5_sel_149845_comb = $signed(p5_prod__571_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148812_comb[23:10];
  assign p5_sel_149848_comb = $signed(p5_prod__573_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58876_NarrowedMult__comb;
  assign p5_bit_slice_149851_comb = p5_or_148819_comb[31:8];
  assign p5_sel_149856_comb = $signed(p5_prod__623_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148824_comb[23:10];
  assign p5_sel_149859_comb = $signed(p5_prod__628_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148827_comb[23:10];
  assign p5_bit_slice_149862_comb = p5_or_148832_comb[31:8];
  assign p5_bit_slice_149867_comb = p5_or_148839_comb[31:8];
  assign p5_bit_slice_149870_comb = p5_or_148844_comb[31:8];
  assign p5_bit_slice_149871_comb = p5_or_148847_comb[31:8];
  assign p5_bit_slice_149874_comb = p5_or_148852_comb[31:8];
  assign p5_bit_slice_149879_comb = p5_or_148859_comb[31:8];
  assign p5_sel_149884_comb = $signed(p5_prod__751_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148864_comb[23:10];
  assign p5_sel_149887_comb = $signed(p5_prod__756_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148867_comb[23:10];
  assign p5_bit_slice_149890_comb = p5_or_148872_comb[31:8];
  assign p5_sel_149895_comb = $signed(p5_prod__795_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58926_NarrowedMult__comb;
  assign p5_sel_149898_comb = $signed(p5_prod__802_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148879_comb[23:10];
  assign p5_sel_149901_comb = $signed(p5_prod__809_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58930_NarrowedMult__comb;
  assign p5_sel_149904_comb = $signed(p5_prod__815_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148884_comb[23:10];
  assign p5_sel_149907_comb = $signed(p5_prod__820_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148887_comb[23:10];
  assign p5_sel_149910_comb = $signed(p5_prod__824_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58936_NarrowedMult__comb;
  assign p5_sel_149913_comb = $signed(p5_prod__827_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148892_comb[23:10];
  assign p5_sel_149916_comb = $signed(p5_prod__829_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_smul_58940_NarrowedMult__comb;
  assign p5_bit_slice_149919_comb = p5_or_148899_comb[31:8];
  assign p5_sel_149924_comb = $signed(p5_prod__879_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148904_comb[23:10];
  assign p5_sel_149927_comb = $signed(p5_prod__884_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148907_comb[23:10];
  assign p5_bit_slice_149930_comb = p5_or_148912_comb[31:8];
  assign p5_bit_slice_149935_comb = p5_or_148919_comb[31:8];
  assign p5_bit_slice_149938_comb = p5_or_148924_comb[31:8];
  assign p5_bit_slice_149939_comb = p5_or_148927_comb[31:8];
  assign p5_bit_slice_149942_comb = p5_or_148932_comb[31:8];
  assign p5_bit_slice_149947_comb = p5_or_148939_comb[31:8];
  assign p5_sel_149952_comb = $signed(p5_prod__1007_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148944_comb[23:10];
  assign p5_sel_149955_comb = $signed(p5_prod__1012_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p5_or_148947_comb[23:10];
  assign p5_bit_slice_149958_comb = p5_or_148952_comb[31:8];
  assign p5_bit_slice_149963_comb = p5_or_149507_comb[23:9];
  assign p5_sel_149966_comb = $signed(p5_prod__554_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148959_comb[23:9];
  assign p5_sel_149969_comb = $signed(p5_prod__574_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148962_comb[23:9];
  assign p5_bit_slice_149972_comb = p5_or_149514_comb[23:9];
  assign p5_sel_149979_comb = $signed(p5_prod__810_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_148999_comb[23:9];
  assign p5_sel_149982_comb = $signed(p5_prod__830_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p5_or_149002_comb[23:9];
  assign p5_sgt_150003_comb = $signed(p5_or_148397_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150004_comb = $signed(p5_or_149134_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150005_comb = $signed(p5_or_149135_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150006_comb = $signed(p5_or_148404_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150007_comb = $signed(p5_or_149140_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150008_comb = $signed(p5_or_149141_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150009_comb = $signed(p5_or_149148_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150010_comb = $signed(p5_or_149149_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150011_comb = $signed(p5_or_148437_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150018_comb = $signed(p5_or_148444_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150019_comb = $signed(p5_or_149160_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150020_comb = $signed(p5_or_149161_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150021_comb = $signed(p5_or_149168_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150022_comb = $signed(p5_or_149169_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150023_comb = $signed(p5_or_148477_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150024_comb = $signed(p5_prod__520_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150025_comb = $signed(p5_prod__524_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150026_comb = $signed(p5_or_148484_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150027_comb = $signed(p5_or_148487_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150028_comb = $signed(p5_prod__542_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150029_comb = $signed(p5_prod__549_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150030_comb = $signed(p5_or_148494_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150031_comb = $signed(p5_prod__584_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150032_comb = $signed(p5_prod__588_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150033_comb = $signed(p5_or_148504_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150034_comb = $signed(p5_or_148507_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150035_comb = $signed(p5_prod__606_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150036_comb = $signed(p5_prod__613_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150037_comb = $signed(p5_prod__648_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150038_comb = $signed(p5_prod__652_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150039_comb = $signed(p5_prod__670_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150040_comb = $signed(p5_prod__677_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150041_comb = $signed(p5_prod__712_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150042_comb = $signed(p5_prod__716_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150043_comb = $signed(p5_or_148544_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150044_comb = $signed(p5_or_148547_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150045_comb = $signed(p5_prod__734_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150046_comb = $signed(p5_prod__741_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150047_comb = $signed(p5_or_148557_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150048_comb = $signed(p5_prod__776_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150049_comb = $signed(p5_prod__780_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150050_comb = $signed(p5_or_148564_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150051_comb = $signed(p5_or_148567_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150052_comb = $signed(p5_prod__798_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150053_comb = $signed(p5_prod__805_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150054_comb = $signed(p5_or_148574_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150055_comb = $signed(p5_prod__840_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150056_comb = $signed(p5_prod__844_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150057_comb = $signed(p5_or_148584_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150058_comb = $signed(p5_or_148587_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150059_comb = $signed(p5_prod__862_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150060_comb = $signed(p5_prod__869_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150061_comb = $signed(p5_prod__904_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150062_comb = $signed(p5_prod__908_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150063_comb = $signed(p5_prod__926_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150064_comb = $signed(p5_prod__933_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150065_comb = $signed(p5_prod__968_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150066_comb = $signed(p5_prod__972_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150067_comb = $signed(p5_or_148624_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150068_comb = $signed(p5_or_148627_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150069_comb = $signed(p5_prod__990_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150070_comb = $signed(p5_prod__997_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150071_comb = $signed(p5_or_149291_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150072_comb = $signed(p5_or_148639_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150073_comb = $signed(p5_or_148642_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150074_comb = $signed(p5_or_149298_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150075_comb = $signed(p5_or_148649_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150076_comb = $signed(p5_or_148652_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150077_comb = $signed(p5_or_148669_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150078_comb = $signed(p5_or_148672_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150082_comb = $signed(p5_or_148679_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150083_comb = $signed(p5_or_148682_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150087_comb = $signed(p5_or_148689_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150088_comb = $signed(p5_or_148692_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150089_comb = $signed(p5_or_148709_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150090_comb = $signed(p5_or_148712_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150091_comb = $signed(p5_or_148717_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150092_comb = $signed(p5_or_149350_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150093_comb = $signed(p5_or_149351_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150094_comb = $signed(p5_or_148724_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150095_comb = $signed(p5_or_148757_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150102_comb = $signed(p5_or_148764_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150103_comb = $signed(p5_prod__539_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150104_comb = $signed(p5_or_148799_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150105_comb = $signed(p5_prod__553_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150106_comb = $signed(p5_or_148804_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150107_comb = $signed(p5_or_148807_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150108_comb = $signed(p5_prod__568_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150109_comb = $signed(p5_or_148812_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150110_comb = $signed(p5_prod__573_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150111_comb = $signed(p5_prod__603_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150112_comb = $signed(p5_prod__617_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150113_comb = $signed(p5_or_148824_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150114_comb = $signed(p5_or_148827_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150115_comb = $signed(p5_prod__632_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150116_comb = $signed(p5_prod__637_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150117_comb = $signed(p5_prod__667_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150118_comb = $signed(p5_prod__681_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150119_comb = $signed(p5_prod__696_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150120_comb = $signed(p5_prod__701_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150121_comb = $signed(p5_prod__731_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150122_comb = $signed(p5_prod__745_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150123_comb = $signed(p5_or_148864_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150124_comb = $signed(p5_or_148867_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150125_comb = $signed(p5_prod__760_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150126_comb = $signed(p5_prod__765_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150127_comb = $signed(p5_prod__795_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150128_comb = $signed(p5_or_148879_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150129_comb = $signed(p5_prod__809_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150130_comb = $signed(p5_or_148884_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150131_comb = $signed(p5_or_148887_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150132_comb = $signed(p5_prod__824_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150133_comb = $signed(p5_or_148892_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150134_comb = $signed(p5_prod__829_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150135_comb = $signed(p5_prod__859_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150136_comb = $signed(p5_prod__873_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150137_comb = $signed(p5_or_148904_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150138_comb = $signed(p5_or_148907_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150139_comb = $signed(p5_prod__888_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150140_comb = $signed(p5_prod__893_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150141_comb = $signed(p5_prod__923_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150142_comb = $signed(p5_prod__937_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150143_comb = $signed(p5_prod__952_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150144_comb = $signed(p5_prod__957_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150145_comb = $signed(p5_prod__987_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150146_comb = $signed(p5_prod__1001_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150147_comb = $signed(p5_or_148944_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150148_comb = $signed(p5_or_148947_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150149_comb = $signed(p5_prod__1016_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150150_comb = $signed(p5_prod__1021_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150151_comb = $signed(p5_or_149507_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150152_comb = $signed(p5_or_148959_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150153_comb = $signed(p5_or_148962_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150154_comb = $signed(p5_or_149514_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150158_comb = $signed(p5_or_148999_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_sgt_150159_comb = $signed(p5_or_149002_comb[31:8]) > $signed(24'h00_7fff);
  assign p5_add_150163_comb = {{1{p5_sel_149547_comb[15]}}, p5_sel_149547_comb} + {{1{p5_sel_149548_comb[15]}}, p5_sel_149548_comb};
  assign p5_add_150164_comb = {{1{p5_sel_149549_comb[15]}}, p5_sel_149549_comb} + {{1{p5_sel_149550_comb[15]}}, p5_sel_149550_comb};
  assign p5_add_150165_comb = {{1{p5_sel_149551_comb[15]}}, p5_sel_149551_comb} + {{1{p5_sel_149552_comb[15]}}, p5_sel_149552_comb};
  assign p5_add_150166_comb = {{1{p5_sel_149553_comb[15]}}, p5_sel_149553_comb} + {{1{p5_sel_149554_comb[15]}}, p5_sel_149554_comb};
  assign p5_add_150167_comb = {{1{p5_sel_149555_comb[15]}}, p5_sel_149555_comb} + {{1{p5_sel_149556_comb[15]}}, p5_sel_149556_comb};
  assign p5_add_150168_comb = {{1{p5_sel_149557_comb[15]}}, p5_sel_149557_comb} + {{1{p5_sel_149558_comb[15]}}, p5_sel_149558_comb};
  assign p5_add_150169_comb = {{1{p5_sel_149559_comb[15]}}, p5_sel_149559_comb} + {{1{p5_sel_149560_comb[15]}}, p5_sel_149560_comb};
  assign p5_add_150170_comb = {{1{p5_sel_149561_comb[15]}}, p5_sel_149561_comb} + {{1{p5_sel_149562_comb[15]}}, p5_sel_149562_comb};
  assign p5_sel_150171_comb = $signed(p5_or_149154_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149154_comb[23:9], 1'h0};
  assign p5_sel_150172_comb = $signed(p5_or_149155_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149155_comb[23:9], 1'h0};
  assign p5_sel_150173_comb = $signed(p5_or_149319_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149319_comb[23:9], 1'h0};
  assign p5_sel_150174_comb = $signed(p5_or_149326_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149326_comb[23:9], 1'h0};
  assign p5_sel_150175_comb = $signed(p5_or_149370_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149370_comb[23:9], 1'h0};
  assign p5_sel_150176_comb = $signed(p5_or_149371_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149371_comb[23:9], 1'h0};
  assign p5_sel_150177_comb = $signed(p5_or_149527_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149527_comb[23:9], 1'h0};
  assign p5_sel_150178_comb = $signed(p5_or_149534_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149534_comb[23:9], 1'h0};

  // Registers for pipe stage 5:
  reg [7:0] p5_shifted__66_squeezed;
  reg [7:0] p5_shifted__69_squeezed;
  reg [7:0] p5_shifted__74_squeezed;
  reg [7:0] p5_shifted__77_squeezed;
  reg [7:0] p5_shifted__82_squeezed;
  reg [7:0] p5_shifted__85_squeezed;
  reg [7:0] p5_shifted__90_squeezed;
  reg [7:0] p5_shifted__93_squeezed;
  reg [7:0] p5_shifted__98_squeezed;
  reg [7:0] p5_shifted__101_squeezed;
  reg [7:0] p5_shifted__106_squeezed;
  reg [7:0] p5_shifted__109_squeezed;
  reg [7:0] p5_shifted__114_squeezed;
  reg [7:0] p5_shifted__117_squeezed;
  reg [7:0] p5_shifted__122_squeezed;
  reg [7:0] p5_shifted__125_squeezed;
  reg [7:0] p5_shifted__64_squeezed;
  reg [7:0] p5_shifted__65_squeezed;
  reg [7:0] p5_shifted__67_squeezed;
  reg [7:0] p5_shifted__68_squeezed;
  reg [7:0] p5_shifted__70_squeezed;
  reg [7:0] p5_shifted__71_squeezed;
  reg [7:0] p5_shifted__72_squeezed;
  reg [7:0] p5_shifted__73_squeezed;
  reg [7:0] p5_shifted__75_squeezed;
  reg [7:0] p5_shifted__76_squeezed;
  reg [7:0] p5_shifted__78_squeezed;
  reg [7:0] p5_shifted__79_squeezed;
  reg [7:0] p5_shifted__80_squeezed;
  reg [7:0] p5_shifted__81_squeezed;
  reg [7:0] p5_shifted__83_squeezed;
  reg [7:0] p5_shifted__84_squeezed;
  reg [7:0] p5_shifted__86_squeezed;
  reg [7:0] p5_shifted__87_squeezed;
  reg [7:0] p5_shifted__88_squeezed;
  reg [7:0] p5_shifted__89_squeezed;
  reg [7:0] p5_shifted__91_squeezed;
  reg [7:0] p5_shifted__92_squeezed;
  reg [7:0] p5_shifted__94_squeezed;
  reg [7:0] p5_shifted__95_squeezed;
  reg [7:0] p5_shifted__96_squeezed;
  reg [7:0] p5_shifted__97_squeezed;
  reg [7:0] p5_shifted__99_squeezed;
  reg [7:0] p5_shifted__100_squeezed;
  reg [7:0] p5_shifted__102_squeezed;
  reg [7:0] p5_shifted__103_squeezed;
  reg [7:0] p5_shifted__104_squeezed;
  reg [7:0] p5_shifted__105_squeezed;
  reg [7:0] p5_shifted__107_squeezed;
  reg [7:0] p5_shifted__108_squeezed;
  reg [7:0] p5_shifted__110_squeezed;
  reg [7:0] p5_shifted__111_squeezed;
  reg [7:0] p5_shifted__112_squeezed;
  reg [7:0] p5_shifted__113_squeezed;
  reg [7:0] p5_shifted__115_squeezed;
  reg [7:0] p5_shifted__116_squeezed;
  reg [7:0] p5_shifted__118_squeezed;
  reg [7:0] p5_shifted__119_squeezed;
  reg [7:0] p5_shifted__120_squeezed;
  reg [7:0] p5_shifted__121_squeezed;
  reg [7:0] p5_shifted__123_squeezed;
  reg [7:0] p5_shifted__124_squeezed;
  reg [7:0] p5_shifted__126_squeezed;
  reg [7:0] p5_shifted__127_squeezed;
  reg [14:0] p5_smul_58368_NarrowedMult_;
  reg [14:0] p5_smul_58370_NarrowedMult_;
  reg [14:0] p5_smul_58376_NarrowedMult_;
  reg [14:0] p5_smul_58378_NarrowedMult_;
  reg [14:0] p5_smul_58384_NarrowedMult_;
  reg [14:0] p5_smul_58386_NarrowedMult_;
  reg [14:0] p5_smul_58392_NarrowedMult_;
  reg [14:0] p5_smul_58394_NarrowedMult_;
  reg [14:0] p5_smul_58400_NarrowedMult_;
  reg [14:0] p5_smul_58402_NarrowedMult_;
  reg [14:0] p5_smul_58408_NarrowedMult_;
  reg [14:0] p5_smul_58410_NarrowedMult_;
  reg [14:0] p5_smul_58432_NarrowedMult_;
  reg [14:0] p5_smul_58434_NarrowedMult_;
  reg [14:0] p5_smul_58440_NarrowedMult_;
  reg [14:0] p5_smul_58442_NarrowedMult_;
  reg [14:0] p5_smul_58448_NarrowedMult_;
  reg [14:0] p5_smul_58450_NarrowedMult_;
  reg [14:0] p5_smul_58456_NarrowedMult_;
  reg [14:0] p5_smul_58458_NarrowedMult_;
  reg [14:0] p5_smul_58464_NarrowedMult_;
  reg [14:0] p5_smul_58466_NarrowedMult_;
  reg [14:0] p5_smul_58472_NarrowedMult_;
  reg [14:0] p5_smul_58474_NarrowedMult_;
  reg [14:0] p5_smul_58878_NarrowedMult_;
  reg [14:0] p5_smul_58882_NarrowedMult_;
  reg [14:0] p5_smul_58888_NarrowedMult_;
  reg [14:0] p5_smul_58892_NarrowedMult_;
  reg [14:0] p5_smul_58894_NarrowedMult_;
  reg [14:0] p5_smul_58898_NarrowedMult_;
  reg [14:0] p5_smul_58904_NarrowedMult_;
  reg [14:0] p5_smul_58908_NarrowedMult_;
  reg [14:0] p5_smul_58910_NarrowedMult_;
  reg [14:0] p5_smul_58914_NarrowedMult_;
  reg [14:0] p5_smul_58920_NarrowedMult_;
  reg [14:0] p5_smul_58924_NarrowedMult_;
  reg [14:0] p5_smul_58942_NarrowedMult_;
  reg [14:0] p5_smul_58946_NarrowedMult_;
  reg [14:0] p5_smul_58952_NarrowedMult_;
  reg [14:0] p5_smul_58956_NarrowedMult_;
  reg [14:0] p5_smul_58958_NarrowedMult_;
  reg [14:0] p5_smul_58962_NarrowedMult_;
  reg [14:0] p5_smul_58968_NarrowedMult_;
  reg [14:0] p5_smul_58972_NarrowedMult_;
  reg [14:0] p5_smul_58974_NarrowedMult_;
  reg [14:0] p5_smul_58978_NarrowedMult_;
  reg [14:0] p5_smul_58984_NarrowedMult_;
  reg [14:0] p5_smul_58988_NarrowedMult_;
  reg [7:0] p5_sel_148221;
  reg [7:0] p5_sel_148224;
  reg [7:0] p5_sel_148227;
  reg [7:0] p5_sel_148230;
  reg [7:0] p5_sel_148233;
  reg [7:0] p5_sel_148236;
  reg [7:0] p5_sel_148239;
  reg [7:0] p5_sel_148242;
  reg [7:0] p5_sel_148245;
  reg [7:0] p5_sel_148248;
  reg [7:0] p5_sel_148251;
  reg [7:0] p5_sel_148254;
  reg [7:0] p5_sel_148257;
  reg [7:0] p5_sel_148260;
  reg [7:0] p5_sel_148263;
  reg [7:0] p5_sel_148266;
  reg [7:0] p5_sel_148269;
  reg [7:0] p5_sel_148272;
  reg [7:0] p5_sel_148275;
  reg [7:0] p5_sel_148278;
  reg [7:0] p5_sel_148281;
  reg [7:0] p5_sel_148284;
  reg [7:0] p5_sel_148287;
  reg [7:0] p5_sel_148290;
  reg [7:0] p5_sel_148325;
  reg [7:0] p5_sel_148328;
  reg [7:0] p5_sel_148331;
  reg [7:0] p5_sel_148334;
  reg [7:0] p5_sel_148337;
  reg [7:0] p5_sel_148340;
  reg [7:0] p5_sel_148343;
  reg [7:0] p5_sel_148346;
  reg [7:0] p5_sel_148349;
  reg [7:0] p5_sel_148352;
  reg [7:0] p5_sel_148355;
  reg [7:0] p5_sel_148358;
  reg [7:0] p5_sel_148361;
  reg [7:0] p5_sel_148364;
  reg [7:0] p5_sel_148367;
  reg [7:0] p5_sel_148370;
  reg [7:0] p5_sel_148373;
  reg [7:0] p5_sel_148376;
  reg [7:0] p5_sel_148379;
  reg [7:0] p5_sel_148382;
  reg [7:0] p5_sel_148385;
  reg [7:0] p5_sel_148388;
  reg [7:0] p5_sel_148391;
  reg [7:0] p5_sel_148394;
  reg [31:0] p5_or_148407;
  reg [31:0] p5_or_148414;
  reg [31:0] p5_or_148417;
  reg [31:0] p5_or_148424;
  reg [31:0] p5_or_148427;
  reg [31:0] p5_or_148434;
  reg [31:0] p5_or_148447;
  reg [31:0] p5_or_148454;
  reg [31:0] p5_or_148457;
  reg [31:0] p5_or_148464;
  reg [31:0] p5_or_148467;
  reg [31:0] p5_or_148474;
  reg [31:0] p5_or_148659;
  reg [31:0] p5_or_148662;
  reg [31:0] p5_or_148699;
  reg [31:0] p5_or_148702;
  reg [31:0] p5_or_148727;
  reg [31:0] p5_or_148734;
  reg [31:0] p5_or_148737;
  reg [31:0] p5_or_148744;
  reg [31:0] p5_or_148747;
  reg [31:0] p5_or_148754;
  reg [31:0] p5_or_148767;
  reg [31:0] p5_or_148774;
  reg [31:0] p5_or_148777;
  reg [31:0] p5_or_148784;
  reg [31:0] p5_or_148787;
  reg [31:0] p5_or_148794;
  reg [31:0] p5_or_148969;
  reg [31:0] p5_or_148972;
  reg [31:0] p5_or_148979;
  reg [31:0] p5_or_148982;
  reg [31:0] p5_or_148989;
  reg [31:0] p5_or_148992;
  reg [31:0] p5_or_149009;
  reg [31:0] p5_or_149012;
  reg [31:0] p5_or_149019;
  reg [31:0] p5_or_149022;
  reg [31:0] p5_or_149029;
  reg [31:0] p5_or_149032;
  reg p5_sgt_149059;
  reg p5_sgt_149060;
  reg p5_sgt_149061;
  reg p5_sgt_149062;
  reg p5_sgt_149063;
  reg p5_sgt_149064;
  reg p5_sgt_149065;
  reg p5_sgt_149066;
  reg p5_sgt_149067;
  reg p5_sgt_149068;
  reg p5_sgt_149069;
  reg p5_sgt_149070;
  reg p5_sgt_149071;
  reg p5_sgt_149072;
  reg p5_sgt_149073;
  reg p5_sgt_149074;
  reg p5_sgt_149075;
  reg p5_sgt_149076;
  reg p5_sgt_149077;
  reg p5_sgt_149078;
  reg p5_sgt_149079;
  reg p5_sgt_149080;
  reg p5_sgt_149081;
  reg p5_sgt_149082;
  reg p5_sgt_149107;
  reg p5_sgt_149108;
  reg p5_sgt_149109;
  reg p5_sgt_149110;
  reg p5_sgt_149111;
  reg p5_sgt_149112;
  reg p5_sgt_149113;
  reg p5_sgt_149114;
  reg p5_sgt_149115;
  reg p5_sgt_149116;
  reg p5_sgt_149117;
  reg p5_sgt_149118;
  reg p5_sgt_149119;
  reg p5_sgt_149120;
  reg p5_sgt_149121;
  reg p5_sgt_149122;
  reg p5_sgt_149123;
  reg p5_sgt_149124;
  reg p5_sgt_149125;
  reg p5_sgt_149126;
  reg p5_sgt_149127;
  reg p5_sgt_149128;
  reg p5_sgt_149129;
  reg p5_sgt_149130;
  reg p5_slt_149139;
  reg p5_slt_149142;
  reg p5_slt_149143;
  reg [31:0] p5_or_149144;
  reg [31:0] p5_or_149145;
  reg p5_slt_149146;
  reg p5_slt_149147;
  reg p5_slt_149150;
  reg p5_slt_149159;
  reg p5_slt_149162;
  reg p5_slt_149163;
  reg [31:0] p5_or_149164;
  reg [31:0] p5_or_149165;
  reg p5_slt_149166;
  reg p5_slt_149167;
  reg p5_slt_149170;
  reg p5_slt_149191;
  reg [13:0] p5_bit_slice_149192;
  reg p5_slt_149193;
  reg p5_slt_149194;
  reg p5_slt_149201;
  reg p5_slt_149202;
  reg p5_slt_149203;
  reg [13:0] p5_bit_slice_149204;
  reg p5_slt_149205;
  reg [13:0] p5_bit_slice_149206;
  reg p5_slt_149207;
  reg p5_slt_149208;
  reg p5_slt_149209;
  reg [13:0] p5_bit_slice_149210;
  reg p5_slt_149211;
  reg [13:0] p5_bit_slice_149212;
  reg p5_slt_149213;
  reg p5_slt_149214;
  reg p5_slt_149215;
  reg [13:0] p5_bit_slice_149216;
  reg p5_slt_149217;
  reg [13:0] p5_bit_slice_149218;
  reg p5_slt_149219;
  reg p5_slt_149220;
  reg p5_slt_149227;
  reg p5_slt_149228;
  reg p5_slt_149229;
  reg [13:0] p5_bit_slice_149230;
  reg p5_slt_149251;
  reg [13:0] p5_bit_slice_149252;
  reg p5_slt_149253;
  reg p5_slt_149254;
  reg p5_slt_149261;
  reg p5_slt_149262;
  reg p5_slt_149263;
  reg [13:0] p5_bit_slice_149264;
  reg p5_slt_149265;
  reg [13:0] p5_bit_slice_149266;
  reg p5_slt_149267;
  reg p5_slt_149268;
  reg p5_slt_149269;
  reg [13:0] p5_bit_slice_149270;
  reg p5_slt_149271;
  reg [13:0] p5_bit_slice_149272;
  reg p5_slt_149273;
  reg p5_slt_149274;
  reg p5_slt_149275;
  reg [13:0] p5_bit_slice_149276;
  reg p5_slt_149277;
  reg [13:0] p5_bit_slice_149278;
  reg p5_slt_149279;
  reg p5_slt_149280;
  reg p5_slt_149287;
  reg p5_slt_149288;
  reg p5_slt_149289;
  reg [13:0] p5_bit_slice_149290;
  reg [31:0] p5_or_149299;
  reg [31:0] p5_or_149306;
  reg [31:0] p5_or_149307;
  reg p5_slt_149308;
  reg p5_slt_149309;
  reg [31:0] p5_or_149310;
  reg [31:0] p5_or_149311;
  reg [31:0] p5_or_149318;
  reg [31:0] p5_or_149327;
  reg [31:0] p5_or_149334;
  reg [31:0] p5_or_149335;
  reg p5_slt_149336;
  reg p5_slt_149337;
  reg [31:0] p5_or_149338;
  reg [31:0] p5_or_149339;
  reg [31:0] p5_or_149346;
  reg p5_slt_149355;
  reg [31:0] p5_or_149356;
  reg [31:0] p5_or_149357;
  reg p5_slt_149358;
  reg p5_slt_149359;
  reg [31:0] p5_or_149360;
  reg [31:0] p5_or_149361;
  reg p5_slt_149362;
  reg p5_slt_149363;
  reg [31:0] p5_or_149364;
  reg [31:0] p5_or_149365;
  reg p5_slt_149366;
  reg p5_slt_149375;
  reg [31:0] p5_or_149376;
  reg [31:0] p5_or_149377;
  reg p5_slt_149378;
  reg p5_slt_149379;
  reg [31:0] p5_or_149380;
  reg [31:0] p5_or_149381;
  reg p5_slt_149382;
  reg p5_slt_149383;
  reg [31:0] p5_or_149384;
  reg [31:0] p5_or_149385;
  reg p5_slt_149386;
  reg p5_slt_149407;
  reg p5_slt_149408;
  reg [13:0] p5_bit_slice_149409;
  reg p5_slt_149410;
  reg p5_slt_149417;
  reg p5_slt_149418;
  reg [13:0] p5_bit_slice_149419;
  reg p5_slt_149420;
  reg p5_slt_149421;
  reg p5_slt_149422;
  reg [13:0] p5_bit_slice_149423;
  reg p5_slt_149424;
  reg p5_slt_149425;
  reg [13:0] p5_bit_slice_149426;
  reg p5_slt_149427;
  reg [13:0] p5_bit_slice_149428;
  reg p5_slt_149429;
  reg p5_slt_149430;
  reg [13:0] p5_bit_slice_149431;
  reg p5_slt_149432;
  reg p5_slt_149433;
  reg p5_slt_149434;
  reg [13:0] p5_bit_slice_149435;
  reg p5_slt_149436;
  reg p5_slt_149443;
  reg p5_slt_149444;
  reg [13:0] p5_bit_slice_149445;
  reg p5_slt_149446;
  reg p5_slt_149467;
  reg p5_slt_149468;
  reg [13:0] p5_bit_slice_149469;
  reg p5_slt_149470;
  reg p5_slt_149477;
  reg p5_slt_149478;
  reg [13:0] p5_bit_slice_149479;
  reg p5_slt_149480;
  reg p5_slt_149481;
  reg p5_slt_149482;
  reg [13:0] p5_bit_slice_149483;
  reg p5_slt_149484;
  reg p5_slt_149485;
  reg [13:0] p5_bit_slice_149486;
  reg p5_slt_149487;
  reg [13:0] p5_bit_slice_149488;
  reg p5_slt_149489;
  reg p5_slt_149490;
  reg [13:0] p5_bit_slice_149491;
  reg p5_slt_149492;
  reg p5_slt_149493;
  reg p5_slt_149494;
  reg [13:0] p5_bit_slice_149495;
  reg p5_slt_149496;
  reg p5_slt_149503;
  reg p5_slt_149504;
  reg [13:0] p5_bit_slice_149505;
  reg p5_slt_149506;
  reg [31:0] p5_or_149515;
  reg p5_slt_149516;
  reg p5_slt_149517;
  reg [31:0] p5_or_149518;
  reg [31:0] p5_or_149519;
  reg p5_slt_149520;
  reg p5_slt_149521;
  reg [31:0] p5_or_149522;
  reg [31:0] p5_or_149523;
  reg p5_slt_149524;
  reg p5_slt_149525;
  reg [31:0] p5_or_149526;
  reg [31:0] p5_or_149535;
  reg p5_slt_149536;
  reg p5_slt_149537;
  reg [31:0] p5_or_149538;
  reg [31:0] p5_or_149539;
  reg p5_slt_149540;
  reg p5_slt_149541;
  reg [31:0] p5_or_149542;
  reg [31:0] p5_or_149543;
  reg p5_slt_149544;
  reg p5_slt_149545;
  reg [31:0] p5_or_149546;
  reg [14:0] p5_sel_149565;
  reg [14:0] p5_bit_slice_149568;
  reg [14:0] p5_bit_slice_149571;
  reg [14:0] p5_sel_149574;
  reg [14:0] p5_bit_slice_149577;
  reg [14:0] p5_bit_slice_149580;
  reg [14:0] p5_bit_slice_149583;
  reg [14:0] p5_bit_slice_149586;
  reg [14:0] p5_sel_149589;
  reg [14:0] p5_sel_149600;
  reg [14:0] p5_bit_slice_149603;
  reg [14:0] p5_bit_slice_149606;
  reg [14:0] p5_bit_slice_149609;
  reg [14:0] p5_bit_slice_149612;
  reg [13:0] p5_sel_149615;
  reg [14:0] p5_sel_149618;
  reg [14:0] p5_sel_149621;
  reg [13:0] p5_sel_149624;
  reg [13:0] p5_sel_149627;
  reg [14:0] p5_sel_149630;
  reg [14:0] p5_sel_149633;
  reg [13:0] p5_sel_149636;
  reg [23:0] p5_bit_slice_149637;
  reg [13:0] p5_sel_149644;
  reg [13:0] p5_sel_149647;
  reg [23:0] p5_bit_slice_149652;
  reg [23:0] p5_bit_slice_149653;
  reg [23:0] p5_bit_slice_149658;
  reg [23:0] p5_bit_slice_149659;
  reg [23:0] p5_bit_slice_149664;
  reg [23:0] p5_bit_slice_149665;
  reg [13:0] p5_sel_149672;
  reg [13:0] p5_sel_149675;
  reg [23:0] p5_bit_slice_149680;
  reg [13:0] p5_sel_149683;
  reg [14:0] p5_sel_149686;
  reg [14:0] p5_sel_149689;
  reg [13:0] p5_sel_149692;
  reg [13:0] p5_sel_149695;
  reg [14:0] p5_sel_149698;
  reg [14:0] p5_sel_149701;
  reg [13:0] p5_sel_149704;
  reg [23:0] p5_bit_slice_149705;
  reg [13:0] p5_sel_149712;
  reg [13:0] p5_sel_149715;
  reg [23:0] p5_bit_slice_149720;
  reg [23:0] p5_bit_slice_149721;
  reg [23:0] p5_bit_slice_149726;
  reg [23:0] p5_bit_slice_149727;
  reg [23:0] p5_bit_slice_149732;
  reg [23:0] p5_bit_slice_149733;
  reg [13:0] p5_sel_149740;
  reg [13:0] p5_sel_149743;
  reg [23:0] p5_bit_slice_149748;
  reg [14:0] p5_bit_slice_149751;
  reg [14:0] p5_sel_149754;
  reg [14:0] p5_sel_149757;
  reg [14:0] p5_bit_slice_149760;
  reg [14:0] p5_sel_149763;
  reg [14:0] p5_sel_149766;
  reg [14:0] p5_sel_149769;
  reg [14:0] p5_sel_149772;
  reg [14:0] p5_sel_149779;
  reg [14:0] p5_sel_149782;
  reg [14:0] p5_sel_149789;
  reg [14:0] p5_sel_149792;
  reg [14:0] p5_sel_149795;
  reg [14:0] p5_sel_149798;
  reg [14:0] p5_sel_149801;
  reg [14:0] p5_bit_slice_149804;
  reg [14:0] p5_bit_slice_149807;
  reg [14:0] p5_sel_149810;
  reg [14:0] p5_sel_149813;
  reg [14:0] p5_sel_149824;
  reg [14:0] p5_sel_149827;
  reg [13:0] p5_sel_149830;
  reg [14:0] p5_sel_149833;
  reg [13:0] p5_sel_149836;
  reg [13:0] p5_sel_149839;
  reg [14:0] p5_sel_149842;
  reg [13:0] p5_sel_149845;
  reg [14:0] p5_sel_149848;
  reg [23:0] p5_bit_slice_149851;
  reg [13:0] p5_sel_149856;
  reg [13:0] p5_sel_149859;
  reg [23:0] p5_bit_slice_149862;
  reg [23:0] p5_bit_slice_149867;
  reg [23:0] p5_bit_slice_149870;
  reg [23:0] p5_bit_slice_149871;
  reg [23:0] p5_bit_slice_149874;
  reg [23:0] p5_bit_slice_149879;
  reg [13:0] p5_sel_149884;
  reg [13:0] p5_sel_149887;
  reg [23:0] p5_bit_slice_149890;
  reg [14:0] p5_sel_149895;
  reg [13:0] p5_sel_149898;
  reg [14:0] p5_sel_149901;
  reg [13:0] p5_sel_149904;
  reg [13:0] p5_sel_149907;
  reg [14:0] p5_sel_149910;
  reg [13:0] p5_sel_149913;
  reg [14:0] p5_sel_149916;
  reg [23:0] p5_bit_slice_149919;
  reg [13:0] p5_sel_149924;
  reg [13:0] p5_sel_149927;
  reg [23:0] p5_bit_slice_149930;
  reg [23:0] p5_bit_slice_149935;
  reg [23:0] p5_bit_slice_149938;
  reg [23:0] p5_bit_slice_149939;
  reg [23:0] p5_bit_slice_149942;
  reg [23:0] p5_bit_slice_149947;
  reg [13:0] p5_sel_149952;
  reg [13:0] p5_sel_149955;
  reg [23:0] p5_bit_slice_149958;
  reg [14:0] p5_bit_slice_149963;
  reg [14:0] p5_sel_149966;
  reg [14:0] p5_sel_149969;
  reg [14:0] p5_bit_slice_149972;
  reg [14:0] p5_sel_149979;
  reg [14:0] p5_sel_149982;
  reg p5_sgt_150003;
  reg p5_sgt_150004;
  reg p5_sgt_150005;
  reg p5_sgt_150006;
  reg p5_sgt_150007;
  reg p5_sgt_150008;
  reg p5_sgt_150009;
  reg p5_sgt_150010;
  reg p5_sgt_150011;
  reg p5_sgt_150018;
  reg p5_sgt_150019;
  reg p5_sgt_150020;
  reg p5_sgt_150021;
  reg p5_sgt_150022;
  reg p5_sgt_150023;
  reg p5_sgt_150024;
  reg p5_sgt_150025;
  reg p5_sgt_150026;
  reg p5_sgt_150027;
  reg p5_sgt_150028;
  reg p5_sgt_150029;
  reg p5_sgt_150030;
  reg p5_sgt_150031;
  reg p5_sgt_150032;
  reg p5_sgt_150033;
  reg p5_sgt_150034;
  reg p5_sgt_150035;
  reg p5_sgt_150036;
  reg p5_sgt_150037;
  reg p5_sgt_150038;
  reg p5_sgt_150039;
  reg p5_sgt_150040;
  reg p5_sgt_150041;
  reg p5_sgt_150042;
  reg p5_sgt_150043;
  reg p5_sgt_150044;
  reg p5_sgt_150045;
  reg p5_sgt_150046;
  reg p5_sgt_150047;
  reg p5_sgt_150048;
  reg p5_sgt_150049;
  reg p5_sgt_150050;
  reg p5_sgt_150051;
  reg p5_sgt_150052;
  reg p5_sgt_150053;
  reg p5_sgt_150054;
  reg p5_sgt_150055;
  reg p5_sgt_150056;
  reg p5_sgt_150057;
  reg p5_sgt_150058;
  reg p5_sgt_150059;
  reg p5_sgt_150060;
  reg p5_sgt_150061;
  reg p5_sgt_150062;
  reg p5_sgt_150063;
  reg p5_sgt_150064;
  reg p5_sgt_150065;
  reg p5_sgt_150066;
  reg p5_sgt_150067;
  reg p5_sgt_150068;
  reg p5_sgt_150069;
  reg p5_sgt_150070;
  reg p5_sgt_150071;
  reg p5_sgt_150072;
  reg p5_sgt_150073;
  reg p5_sgt_150074;
  reg p5_sgt_150075;
  reg p5_sgt_150076;
  reg p5_sgt_150077;
  reg p5_sgt_150078;
  reg p5_sgt_150082;
  reg p5_sgt_150083;
  reg p5_sgt_150087;
  reg p5_sgt_150088;
  reg p5_sgt_150089;
  reg p5_sgt_150090;
  reg p5_sgt_150091;
  reg p5_sgt_150092;
  reg p5_sgt_150093;
  reg p5_sgt_150094;
  reg p5_sgt_150095;
  reg p5_sgt_150102;
  reg p5_sgt_150103;
  reg p5_sgt_150104;
  reg p5_sgt_150105;
  reg p5_sgt_150106;
  reg p5_sgt_150107;
  reg p5_sgt_150108;
  reg p5_sgt_150109;
  reg p5_sgt_150110;
  reg p5_sgt_150111;
  reg p5_sgt_150112;
  reg p5_sgt_150113;
  reg p5_sgt_150114;
  reg p5_sgt_150115;
  reg p5_sgt_150116;
  reg p5_sgt_150117;
  reg p5_sgt_150118;
  reg p5_sgt_150119;
  reg p5_sgt_150120;
  reg p5_sgt_150121;
  reg p5_sgt_150122;
  reg p5_sgt_150123;
  reg p5_sgt_150124;
  reg p5_sgt_150125;
  reg p5_sgt_150126;
  reg p5_sgt_150127;
  reg p5_sgt_150128;
  reg p5_sgt_150129;
  reg p5_sgt_150130;
  reg p5_sgt_150131;
  reg p5_sgt_150132;
  reg p5_sgt_150133;
  reg p5_sgt_150134;
  reg p5_sgt_150135;
  reg p5_sgt_150136;
  reg p5_sgt_150137;
  reg p5_sgt_150138;
  reg p5_sgt_150139;
  reg p5_sgt_150140;
  reg p5_sgt_150141;
  reg p5_sgt_150142;
  reg p5_sgt_150143;
  reg p5_sgt_150144;
  reg p5_sgt_150145;
  reg p5_sgt_150146;
  reg p5_sgt_150147;
  reg p5_sgt_150148;
  reg p5_sgt_150149;
  reg p5_sgt_150150;
  reg p5_sgt_150151;
  reg p5_sgt_150152;
  reg p5_sgt_150153;
  reg p5_sgt_150154;
  reg p5_sgt_150158;
  reg p5_sgt_150159;
  reg [16:0] p5_add_150163;
  reg [16:0] p5_add_150164;
  reg [16:0] p5_add_150165;
  reg [16:0] p5_add_150166;
  reg [16:0] p5_add_150167;
  reg [16:0] p5_add_150168;
  reg [16:0] p5_add_150169;
  reg [16:0] p5_add_150170;
  reg [15:0] p5_sel_150171;
  reg [15:0] p5_sel_150172;
  reg [15:0] p5_sel_150173;
  reg [15:0] p5_sel_150174;
  reg [15:0] p5_sel_150175;
  reg [15:0] p5_sel_150176;
  reg [15:0] p5_sel_150177;
  reg [15:0] p5_sel_150178;
  always @ (posedge clk) begin
    p5_shifted__66_squeezed <= p5_shifted__66_squeezed_comb;
    p5_shifted__69_squeezed <= p5_shifted__69_squeezed_comb;
    p5_shifted__74_squeezed <= p5_shifted__74_squeezed_comb;
    p5_shifted__77_squeezed <= p5_shifted__77_squeezed_comb;
    p5_shifted__82_squeezed <= p5_shifted__82_squeezed_comb;
    p5_shifted__85_squeezed <= p5_shifted__85_squeezed_comb;
    p5_shifted__90_squeezed <= p5_shifted__90_squeezed_comb;
    p5_shifted__93_squeezed <= p5_shifted__93_squeezed_comb;
    p5_shifted__98_squeezed <= p5_shifted__98_squeezed_comb;
    p5_shifted__101_squeezed <= p5_shifted__101_squeezed_comb;
    p5_shifted__106_squeezed <= p5_shifted__106_squeezed_comb;
    p5_shifted__109_squeezed <= p5_shifted__109_squeezed_comb;
    p5_shifted__114_squeezed <= p5_shifted__114_squeezed_comb;
    p5_shifted__117_squeezed <= p5_shifted__117_squeezed_comb;
    p5_shifted__122_squeezed <= p5_shifted__122_squeezed_comb;
    p5_shifted__125_squeezed <= p5_shifted__125_squeezed_comb;
    p5_shifted__64_squeezed <= p5_shifted__64_squeezed_comb;
    p5_shifted__65_squeezed <= p5_shifted__65_squeezed_comb;
    p5_shifted__67_squeezed <= p5_shifted__67_squeezed_comb;
    p5_shifted__68_squeezed <= p5_shifted__68_squeezed_comb;
    p5_shifted__70_squeezed <= p5_shifted__70_squeezed_comb;
    p5_shifted__71_squeezed <= p5_shifted__71_squeezed_comb;
    p5_shifted__72_squeezed <= p5_shifted__72_squeezed_comb;
    p5_shifted__73_squeezed <= p5_shifted__73_squeezed_comb;
    p5_shifted__75_squeezed <= p5_shifted__75_squeezed_comb;
    p5_shifted__76_squeezed <= p5_shifted__76_squeezed_comb;
    p5_shifted__78_squeezed <= p5_shifted__78_squeezed_comb;
    p5_shifted__79_squeezed <= p5_shifted__79_squeezed_comb;
    p5_shifted__80_squeezed <= p5_shifted__80_squeezed_comb;
    p5_shifted__81_squeezed <= p5_shifted__81_squeezed_comb;
    p5_shifted__83_squeezed <= p5_shifted__83_squeezed_comb;
    p5_shifted__84_squeezed <= p5_shifted__84_squeezed_comb;
    p5_shifted__86_squeezed <= p5_shifted__86_squeezed_comb;
    p5_shifted__87_squeezed <= p5_shifted__87_squeezed_comb;
    p5_shifted__88_squeezed <= p5_shifted__88_squeezed_comb;
    p5_shifted__89_squeezed <= p5_shifted__89_squeezed_comb;
    p5_shifted__91_squeezed <= p5_shifted__91_squeezed_comb;
    p5_shifted__92_squeezed <= p5_shifted__92_squeezed_comb;
    p5_shifted__94_squeezed <= p5_shifted__94_squeezed_comb;
    p5_shifted__95_squeezed <= p5_shifted__95_squeezed_comb;
    p5_shifted__96_squeezed <= p5_shifted__96_squeezed_comb;
    p5_shifted__97_squeezed <= p5_shifted__97_squeezed_comb;
    p5_shifted__99_squeezed <= p5_shifted__99_squeezed_comb;
    p5_shifted__100_squeezed <= p5_shifted__100_squeezed_comb;
    p5_shifted__102_squeezed <= p5_shifted__102_squeezed_comb;
    p5_shifted__103_squeezed <= p5_shifted__103_squeezed_comb;
    p5_shifted__104_squeezed <= p5_shifted__104_squeezed_comb;
    p5_shifted__105_squeezed <= p5_shifted__105_squeezed_comb;
    p5_shifted__107_squeezed <= p5_shifted__107_squeezed_comb;
    p5_shifted__108_squeezed <= p5_shifted__108_squeezed_comb;
    p5_shifted__110_squeezed <= p5_shifted__110_squeezed_comb;
    p5_shifted__111_squeezed <= p5_shifted__111_squeezed_comb;
    p5_shifted__112_squeezed <= p5_shifted__112_squeezed_comb;
    p5_shifted__113_squeezed <= p5_shifted__113_squeezed_comb;
    p5_shifted__115_squeezed <= p5_shifted__115_squeezed_comb;
    p5_shifted__116_squeezed <= p5_shifted__116_squeezed_comb;
    p5_shifted__118_squeezed <= p5_shifted__118_squeezed_comb;
    p5_shifted__119_squeezed <= p5_shifted__119_squeezed_comb;
    p5_shifted__120_squeezed <= p5_shifted__120_squeezed_comb;
    p5_shifted__121_squeezed <= p5_shifted__121_squeezed_comb;
    p5_shifted__123_squeezed <= p5_shifted__123_squeezed_comb;
    p5_shifted__124_squeezed <= p5_shifted__124_squeezed_comb;
    p5_shifted__126_squeezed <= p5_shifted__126_squeezed_comb;
    p5_shifted__127_squeezed <= p5_shifted__127_squeezed_comb;
    p5_smul_58368_NarrowedMult_ <= p5_smul_58368_NarrowedMult__comb;
    p5_smul_58370_NarrowedMult_ <= p5_smul_58370_NarrowedMult__comb;
    p5_smul_58376_NarrowedMult_ <= p5_smul_58376_NarrowedMult__comb;
    p5_smul_58378_NarrowedMult_ <= p5_smul_58378_NarrowedMult__comb;
    p5_smul_58384_NarrowedMult_ <= p5_smul_58384_NarrowedMult__comb;
    p5_smul_58386_NarrowedMult_ <= p5_smul_58386_NarrowedMult__comb;
    p5_smul_58392_NarrowedMult_ <= p5_smul_58392_NarrowedMult__comb;
    p5_smul_58394_NarrowedMult_ <= p5_smul_58394_NarrowedMult__comb;
    p5_smul_58400_NarrowedMult_ <= p5_smul_58400_NarrowedMult__comb;
    p5_smul_58402_NarrowedMult_ <= p5_smul_58402_NarrowedMult__comb;
    p5_smul_58408_NarrowedMult_ <= p5_smul_58408_NarrowedMult__comb;
    p5_smul_58410_NarrowedMult_ <= p5_smul_58410_NarrowedMult__comb;
    p5_smul_58432_NarrowedMult_ <= p5_smul_58432_NarrowedMult__comb;
    p5_smul_58434_NarrowedMult_ <= p5_smul_58434_NarrowedMult__comb;
    p5_smul_58440_NarrowedMult_ <= p5_smul_58440_NarrowedMult__comb;
    p5_smul_58442_NarrowedMult_ <= p5_smul_58442_NarrowedMult__comb;
    p5_smul_58448_NarrowedMult_ <= p5_smul_58448_NarrowedMult__comb;
    p5_smul_58450_NarrowedMult_ <= p5_smul_58450_NarrowedMult__comb;
    p5_smul_58456_NarrowedMult_ <= p5_smul_58456_NarrowedMult__comb;
    p5_smul_58458_NarrowedMult_ <= p5_smul_58458_NarrowedMult__comb;
    p5_smul_58464_NarrowedMult_ <= p5_smul_58464_NarrowedMult__comb;
    p5_smul_58466_NarrowedMult_ <= p5_smul_58466_NarrowedMult__comb;
    p5_smul_58472_NarrowedMult_ <= p5_smul_58472_NarrowedMult__comb;
    p5_smul_58474_NarrowedMult_ <= p5_smul_58474_NarrowedMult__comb;
    p5_smul_58878_NarrowedMult_ <= p5_smul_58878_NarrowedMult__comb;
    p5_smul_58882_NarrowedMult_ <= p5_smul_58882_NarrowedMult__comb;
    p5_smul_58888_NarrowedMult_ <= p5_smul_58888_NarrowedMult__comb;
    p5_smul_58892_NarrowedMult_ <= p5_smul_58892_NarrowedMult__comb;
    p5_smul_58894_NarrowedMult_ <= p5_smul_58894_NarrowedMult__comb;
    p5_smul_58898_NarrowedMult_ <= p5_smul_58898_NarrowedMult__comb;
    p5_smul_58904_NarrowedMult_ <= p5_smul_58904_NarrowedMult__comb;
    p5_smul_58908_NarrowedMult_ <= p5_smul_58908_NarrowedMult__comb;
    p5_smul_58910_NarrowedMult_ <= p5_smul_58910_NarrowedMult__comb;
    p5_smul_58914_NarrowedMult_ <= p5_smul_58914_NarrowedMult__comb;
    p5_smul_58920_NarrowedMult_ <= p5_smul_58920_NarrowedMult__comb;
    p5_smul_58924_NarrowedMult_ <= p5_smul_58924_NarrowedMult__comb;
    p5_smul_58942_NarrowedMult_ <= p5_smul_58942_NarrowedMult__comb;
    p5_smul_58946_NarrowedMult_ <= p5_smul_58946_NarrowedMult__comb;
    p5_smul_58952_NarrowedMult_ <= p5_smul_58952_NarrowedMult__comb;
    p5_smul_58956_NarrowedMult_ <= p5_smul_58956_NarrowedMult__comb;
    p5_smul_58958_NarrowedMult_ <= p5_smul_58958_NarrowedMult__comb;
    p5_smul_58962_NarrowedMult_ <= p5_smul_58962_NarrowedMult__comb;
    p5_smul_58968_NarrowedMult_ <= p5_smul_58968_NarrowedMult__comb;
    p5_smul_58972_NarrowedMult_ <= p5_smul_58972_NarrowedMult__comb;
    p5_smul_58974_NarrowedMult_ <= p5_smul_58974_NarrowedMult__comb;
    p5_smul_58978_NarrowedMult_ <= p5_smul_58978_NarrowedMult__comb;
    p5_smul_58984_NarrowedMult_ <= p5_smul_58984_NarrowedMult__comb;
    p5_smul_58988_NarrowedMult_ <= p5_smul_58988_NarrowedMult__comb;
    p5_sel_148221 <= p5_sel_148221_comb;
    p5_sel_148224 <= p5_sel_148224_comb;
    p5_sel_148227 <= p5_sel_148227_comb;
    p5_sel_148230 <= p5_sel_148230_comb;
    p5_sel_148233 <= p5_sel_148233_comb;
    p5_sel_148236 <= p5_sel_148236_comb;
    p5_sel_148239 <= p5_sel_148239_comb;
    p5_sel_148242 <= p5_sel_148242_comb;
    p5_sel_148245 <= p5_sel_148245_comb;
    p5_sel_148248 <= p5_sel_148248_comb;
    p5_sel_148251 <= p5_sel_148251_comb;
    p5_sel_148254 <= p5_sel_148254_comb;
    p5_sel_148257 <= p5_sel_148257_comb;
    p5_sel_148260 <= p5_sel_148260_comb;
    p5_sel_148263 <= p5_sel_148263_comb;
    p5_sel_148266 <= p5_sel_148266_comb;
    p5_sel_148269 <= p5_sel_148269_comb;
    p5_sel_148272 <= p5_sel_148272_comb;
    p5_sel_148275 <= p5_sel_148275_comb;
    p5_sel_148278 <= p5_sel_148278_comb;
    p5_sel_148281 <= p5_sel_148281_comb;
    p5_sel_148284 <= p5_sel_148284_comb;
    p5_sel_148287 <= p5_sel_148287_comb;
    p5_sel_148290 <= p5_sel_148290_comb;
    p5_sel_148325 <= p5_sel_148325_comb;
    p5_sel_148328 <= p5_sel_148328_comb;
    p5_sel_148331 <= p5_sel_148331_comb;
    p5_sel_148334 <= p5_sel_148334_comb;
    p5_sel_148337 <= p5_sel_148337_comb;
    p5_sel_148340 <= p5_sel_148340_comb;
    p5_sel_148343 <= p5_sel_148343_comb;
    p5_sel_148346 <= p5_sel_148346_comb;
    p5_sel_148349 <= p5_sel_148349_comb;
    p5_sel_148352 <= p5_sel_148352_comb;
    p5_sel_148355 <= p5_sel_148355_comb;
    p5_sel_148358 <= p5_sel_148358_comb;
    p5_sel_148361 <= p5_sel_148361_comb;
    p5_sel_148364 <= p5_sel_148364_comb;
    p5_sel_148367 <= p5_sel_148367_comb;
    p5_sel_148370 <= p5_sel_148370_comb;
    p5_sel_148373 <= p5_sel_148373_comb;
    p5_sel_148376 <= p5_sel_148376_comb;
    p5_sel_148379 <= p5_sel_148379_comb;
    p5_sel_148382 <= p5_sel_148382_comb;
    p5_sel_148385 <= p5_sel_148385_comb;
    p5_sel_148388 <= p5_sel_148388_comb;
    p5_sel_148391 <= p5_sel_148391_comb;
    p5_sel_148394 <= p5_sel_148394_comb;
    p5_or_148407 <= p5_or_148407_comb;
    p5_or_148414 <= p5_or_148414_comb;
    p5_or_148417 <= p5_or_148417_comb;
    p5_or_148424 <= p5_or_148424_comb;
    p5_or_148427 <= p5_or_148427_comb;
    p5_or_148434 <= p5_or_148434_comb;
    p5_or_148447 <= p5_or_148447_comb;
    p5_or_148454 <= p5_or_148454_comb;
    p5_or_148457 <= p5_or_148457_comb;
    p5_or_148464 <= p5_or_148464_comb;
    p5_or_148467 <= p5_or_148467_comb;
    p5_or_148474 <= p5_or_148474_comb;
    p5_or_148659 <= p5_or_148659_comb;
    p5_or_148662 <= p5_or_148662_comb;
    p5_or_148699 <= p5_or_148699_comb;
    p5_or_148702 <= p5_or_148702_comb;
    p5_or_148727 <= p5_or_148727_comb;
    p5_or_148734 <= p5_or_148734_comb;
    p5_or_148737 <= p5_or_148737_comb;
    p5_or_148744 <= p5_or_148744_comb;
    p5_or_148747 <= p5_or_148747_comb;
    p5_or_148754 <= p5_or_148754_comb;
    p5_or_148767 <= p5_or_148767_comb;
    p5_or_148774 <= p5_or_148774_comb;
    p5_or_148777 <= p5_or_148777_comb;
    p5_or_148784 <= p5_or_148784_comb;
    p5_or_148787 <= p5_or_148787_comb;
    p5_or_148794 <= p5_or_148794_comb;
    p5_or_148969 <= p5_or_148969_comb;
    p5_or_148972 <= p5_or_148972_comb;
    p5_or_148979 <= p5_or_148979_comb;
    p5_or_148982 <= p5_or_148982_comb;
    p5_or_148989 <= p5_or_148989_comb;
    p5_or_148992 <= p5_or_148992_comb;
    p5_or_149009 <= p5_or_149009_comb;
    p5_or_149012 <= p5_or_149012_comb;
    p5_or_149019 <= p5_or_149019_comb;
    p5_or_149022 <= p5_or_149022_comb;
    p5_or_149029 <= p5_or_149029_comb;
    p5_or_149032 <= p5_or_149032_comb;
    p5_sgt_149059 <= p5_sgt_149059_comb;
    p5_sgt_149060 <= p5_sgt_149060_comb;
    p5_sgt_149061 <= p5_sgt_149061_comb;
    p5_sgt_149062 <= p5_sgt_149062_comb;
    p5_sgt_149063 <= p5_sgt_149063_comb;
    p5_sgt_149064 <= p5_sgt_149064_comb;
    p5_sgt_149065 <= p5_sgt_149065_comb;
    p5_sgt_149066 <= p5_sgt_149066_comb;
    p5_sgt_149067 <= p5_sgt_149067_comb;
    p5_sgt_149068 <= p5_sgt_149068_comb;
    p5_sgt_149069 <= p5_sgt_149069_comb;
    p5_sgt_149070 <= p5_sgt_149070_comb;
    p5_sgt_149071 <= p5_sgt_149071_comb;
    p5_sgt_149072 <= p5_sgt_149072_comb;
    p5_sgt_149073 <= p5_sgt_149073_comb;
    p5_sgt_149074 <= p5_sgt_149074_comb;
    p5_sgt_149075 <= p5_sgt_149075_comb;
    p5_sgt_149076 <= p5_sgt_149076_comb;
    p5_sgt_149077 <= p5_sgt_149077_comb;
    p5_sgt_149078 <= p5_sgt_149078_comb;
    p5_sgt_149079 <= p5_sgt_149079_comb;
    p5_sgt_149080 <= p5_sgt_149080_comb;
    p5_sgt_149081 <= p5_sgt_149081_comb;
    p5_sgt_149082 <= p5_sgt_149082_comb;
    p5_sgt_149107 <= p5_sgt_149107_comb;
    p5_sgt_149108 <= p5_sgt_149108_comb;
    p5_sgt_149109 <= p5_sgt_149109_comb;
    p5_sgt_149110 <= p5_sgt_149110_comb;
    p5_sgt_149111 <= p5_sgt_149111_comb;
    p5_sgt_149112 <= p5_sgt_149112_comb;
    p5_sgt_149113 <= p5_sgt_149113_comb;
    p5_sgt_149114 <= p5_sgt_149114_comb;
    p5_sgt_149115 <= p5_sgt_149115_comb;
    p5_sgt_149116 <= p5_sgt_149116_comb;
    p5_sgt_149117 <= p5_sgt_149117_comb;
    p5_sgt_149118 <= p5_sgt_149118_comb;
    p5_sgt_149119 <= p5_sgt_149119_comb;
    p5_sgt_149120 <= p5_sgt_149120_comb;
    p5_sgt_149121 <= p5_sgt_149121_comb;
    p5_sgt_149122 <= p5_sgt_149122_comb;
    p5_sgt_149123 <= p5_sgt_149123_comb;
    p5_sgt_149124 <= p5_sgt_149124_comb;
    p5_sgt_149125 <= p5_sgt_149125_comb;
    p5_sgt_149126 <= p5_sgt_149126_comb;
    p5_sgt_149127 <= p5_sgt_149127_comb;
    p5_sgt_149128 <= p5_sgt_149128_comb;
    p5_sgt_149129 <= p5_sgt_149129_comb;
    p5_sgt_149130 <= p5_sgt_149130_comb;
    p5_slt_149139 <= p5_slt_149139_comb;
    p5_slt_149142 <= p5_slt_149142_comb;
    p5_slt_149143 <= p5_slt_149143_comb;
    p5_or_149144 <= p5_or_149144_comb;
    p5_or_149145 <= p5_or_149145_comb;
    p5_slt_149146 <= p5_slt_149146_comb;
    p5_slt_149147 <= p5_slt_149147_comb;
    p5_slt_149150 <= p5_slt_149150_comb;
    p5_slt_149159 <= p5_slt_149159_comb;
    p5_slt_149162 <= p5_slt_149162_comb;
    p5_slt_149163 <= p5_slt_149163_comb;
    p5_or_149164 <= p5_or_149164_comb;
    p5_or_149165 <= p5_or_149165_comb;
    p5_slt_149166 <= p5_slt_149166_comb;
    p5_slt_149167 <= p5_slt_149167_comb;
    p5_slt_149170 <= p5_slt_149170_comb;
    p5_slt_149191 <= p5_slt_149191_comb;
    p5_bit_slice_149192 <= p5_bit_slice_149192_comb;
    p5_slt_149193 <= p5_slt_149193_comb;
    p5_slt_149194 <= p5_slt_149194_comb;
    p5_slt_149201 <= p5_slt_149201_comb;
    p5_slt_149202 <= p5_slt_149202_comb;
    p5_slt_149203 <= p5_slt_149203_comb;
    p5_bit_slice_149204 <= p5_bit_slice_149204_comb;
    p5_slt_149205 <= p5_slt_149205_comb;
    p5_bit_slice_149206 <= p5_bit_slice_149206_comb;
    p5_slt_149207 <= p5_slt_149207_comb;
    p5_slt_149208 <= p5_slt_149208_comb;
    p5_slt_149209 <= p5_slt_149209_comb;
    p5_bit_slice_149210 <= p5_bit_slice_149210_comb;
    p5_slt_149211 <= p5_slt_149211_comb;
    p5_bit_slice_149212 <= p5_bit_slice_149212_comb;
    p5_slt_149213 <= p5_slt_149213_comb;
    p5_slt_149214 <= p5_slt_149214_comb;
    p5_slt_149215 <= p5_slt_149215_comb;
    p5_bit_slice_149216 <= p5_bit_slice_149216_comb;
    p5_slt_149217 <= p5_slt_149217_comb;
    p5_bit_slice_149218 <= p5_bit_slice_149218_comb;
    p5_slt_149219 <= p5_slt_149219_comb;
    p5_slt_149220 <= p5_slt_149220_comb;
    p5_slt_149227 <= p5_slt_149227_comb;
    p5_slt_149228 <= p5_slt_149228_comb;
    p5_slt_149229 <= p5_slt_149229_comb;
    p5_bit_slice_149230 <= p5_bit_slice_149230_comb;
    p5_slt_149251 <= p5_slt_149251_comb;
    p5_bit_slice_149252 <= p5_bit_slice_149252_comb;
    p5_slt_149253 <= p5_slt_149253_comb;
    p5_slt_149254 <= p5_slt_149254_comb;
    p5_slt_149261 <= p5_slt_149261_comb;
    p5_slt_149262 <= p5_slt_149262_comb;
    p5_slt_149263 <= p5_slt_149263_comb;
    p5_bit_slice_149264 <= p5_bit_slice_149264_comb;
    p5_slt_149265 <= p5_slt_149265_comb;
    p5_bit_slice_149266 <= p5_bit_slice_149266_comb;
    p5_slt_149267 <= p5_slt_149267_comb;
    p5_slt_149268 <= p5_slt_149268_comb;
    p5_slt_149269 <= p5_slt_149269_comb;
    p5_bit_slice_149270 <= p5_bit_slice_149270_comb;
    p5_slt_149271 <= p5_slt_149271_comb;
    p5_bit_slice_149272 <= p5_bit_slice_149272_comb;
    p5_slt_149273 <= p5_slt_149273_comb;
    p5_slt_149274 <= p5_slt_149274_comb;
    p5_slt_149275 <= p5_slt_149275_comb;
    p5_bit_slice_149276 <= p5_bit_slice_149276_comb;
    p5_slt_149277 <= p5_slt_149277_comb;
    p5_bit_slice_149278 <= p5_bit_slice_149278_comb;
    p5_slt_149279 <= p5_slt_149279_comb;
    p5_slt_149280 <= p5_slt_149280_comb;
    p5_slt_149287 <= p5_slt_149287_comb;
    p5_slt_149288 <= p5_slt_149288_comb;
    p5_slt_149289 <= p5_slt_149289_comb;
    p5_bit_slice_149290 <= p5_bit_slice_149290_comb;
    p5_or_149299 <= p5_or_149299_comb;
    p5_or_149306 <= p5_or_149306_comb;
    p5_or_149307 <= p5_or_149307_comb;
    p5_slt_149308 <= p5_slt_149308_comb;
    p5_slt_149309 <= p5_slt_149309_comb;
    p5_or_149310 <= p5_or_149310_comb;
    p5_or_149311 <= p5_or_149311_comb;
    p5_or_149318 <= p5_or_149318_comb;
    p5_or_149327 <= p5_or_149327_comb;
    p5_or_149334 <= p5_or_149334_comb;
    p5_or_149335 <= p5_or_149335_comb;
    p5_slt_149336 <= p5_slt_149336_comb;
    p5_slt_149337 <= p5_slt_149337_comb;
    p5_or_149338 <= p5_or_149338_comb;
    p5_or_149339 <= p5_or_149339_comb;
    p5_or_149346 <= p5_or_149346_comb;
    p5_slt_149355 <= p5_slt_149355_comb;
    p5_or_149356 <= p5_or_149356_comb;
    p5_or_149357 <= p5_or_149357_comb;
    p5_slt_149358 <= p5_slt_149358_comb;
    p5_slt_149359 <= p5_slt_149359_comb;
    p5_or_149360 <= p5_or_149360_comb;
    p5_or_149361 <= p5_or_149361_comb;
    p5_slt_149362 <= p5_slt_149362_comb;
    p5_slt_149363 <= p5_slt_149363_comb;
    p5_or_149364 <= p5_or_149364_comb;
    p5_or_149365 <= p5_or_149365_comb;
    p5_slt_149366 <= p5_slt_149366_comb;
    p5_slt_149375 <= p5_slt_149375_comb;
    p5_or_149376 <= p5_or_149376_comb;
    p5_or_149377 <= p5_or_149377_comb;
    p5_slt_149378 <= p5_slt_149378_comb;
    p5_slt_149379 <= p5_slt_149379_comb;
    p5_or_149380 <= p5_or_149380_comb;
    p5_or_149381 <= p5_or_149381_comb;
    p5_slt_149382 <= p5_slt_149382_comb;
    p5_slt_149383 <= p5_slt_149383_comb;
    p5_or_149384 <= p5_or_149384_comb;
    p5_or_149385 <= p5_or_149385_comb;
    p5_slt_149386 <= p5_slt_149386_comb;
    p5_slt_149407 <= p5_slt_149407_comb;
    p5_slt_149408 <= p5_slt_149408_comb;
    p5_bit_slice_149409 <= p5_bit_slice_149409_comb;
    p5_slt_149410 <= p5_slt_149410_comb;
    p5_slt_149417 <= p5_slt_149417_comb;
    p5_slt_149418 <= p5_slt_149418_comb;
    p5_bit_slice_149419 <= p5_bit_slice_149419_comb;
    p5_slt_149420 <= p5_slt_149420_comb;
    p5_slt_149421 <= p5_slt_149421_comb;
    p5_slt_149422 <= p5_slt_149422_comb;
    p5_bit_slice_149423 <= p5_bit_slice_149423_comb;
    p5_slt_149424 <= p5_slt_149424_comb;
    p5_slt_149425 <= p5_slt_149425_comb;
    p5_bit_slice_149426 <= p5_bit_slice_149426_comb;
    p5_slt_149427 <= p5_slt_149427_comb;
    p5_bit_slice_149428 <= p5_bit_slice_149428_comb;
    p5_slt_149429 <= p5_slt_149429_comb;
    p5_slt_149430 <= p5_slt_149430_comb;
    p5_bit_slice_149431 <= p5_bit_slice_149431_comb;
    p5_slt_149432 <= p5_slt_149432_comb;
    p5_slt_149433 <= p5_slt_149433_comb;
    p5_slt_149434 <= p5_slt_149434_comb;
    p5_bit_slice_149435 <= p5_bit_slice_149435_comb;
    p5_slt_149436 <= p5_slt_149436_comb;
    p5_slt_149443 <= p5_slt_149443_comb;
    p5_slt_149444 <= p5_slt_149444_comb;
    p5_bit_slice_149445 <= p5_bit_slice_149445_comb;
    p5_slt_149446 <= p5_slt_149446_comb;
    p5_slt_149467 <= p5_slt_149467_comb;
    p5_slt_149468 <= p5_slt_149468_comb;
    p5_bit_slice_149469 <= p5_bit_slice_149469_comb;
    p5_slt_149470 <= p5_slt_149470_comb;
    p5_slt_149477 <= p5_slt_149477_comb;
    p5_slt_149478 <= p5_slt_149478_comb;
    p5_bit_slice_149479 <= p5_bit_slice_149479_comb;
    p5_slt_149480 <= p5_slt_149480_comb;
    p5_slt_149481 <= p5_slt_149481_comb;
    p5_slt_149482 <= p5_slt_149482_comb;
    p5_bit_slice_149483 <= p5_bit_slice_149483_comb;
    p5_slt_149484 <= p5_slt_149484_comb;
    p5_slt_149485 <= p5_slt_149485_comb;
    p5_bit_slice_149486 <= p5_bit_slice_149486_comb;
    p5_slt_149487 <= p5_slt_149487_comb;
    p5_bit_slice_149488 <= p5_bit_slice_149488_comb;
    p5_slt_149489 <= p5_slt_149489_comb;
    p5_slt_149490 <= p5_slt_149490_comb;
    p5_bit_slice_149491 <= p5_bit_slice_149491_comb;
    p5_slt_149492 <= p5_slt_149492_comb;
    p5_slt_149493 <= p5_slt_149493_comb;
    p5_slt_149494 <= p5_slt_149494_comb;
    p5_bit_slice_149495 <= p5_bit_slice_149495_comb;
    p5_slt_149496 <= p5_slt_149496_comb;
    p5_slt_149503 <= p5_slt_149503_comb;
    p5_slt_149504 <= p5_slt_149504_comb;
    p5_bit_slice_149505 <= p5_bit_slice_149505_comb;
    p5_slt_149506 <= p5_slt_149506_comb;
    p5_or_149515 <= p5_or_149515_comb;
    p5_slt_149516 <= p5_slt_149516_comb;
    p5_slt_149517 <= p5_slt_149517_comb;
    p5_or_149518 <= p5_or_149518_comb;
    p5_or_149519 <= p5_or_149519_comb;
    p5_slt_149520 <= p5_slt_149520_comb;
    p5_slt_149521 <= p5_slt_149521_comb;
    p5_or_149522 <= p5_or_149522_comb;
    p5_or_149523 <= p5_or_149523_comb;
    p5_slt_149524 <= p5_slt_149524_comb;
    p5_slt_149525 <= p5_slt_149525_comb;
    p5_or_149526 <= p5_or_149526_comb;
    p5_or_149535 <= p5_or_149535_comb;
    p5_slt_149536 <= p5_slt_149536_comb;
    p5_slt_149537 <= p5_slt_149537_comb;
    p5_or_149538 <= p5_or_149538_comb;
    p5_or_149539 <= p5_or_149539_comb;
    p5_slt_149540 <= p5_slt_149540_comb;
    p5_slt_149541 <= p5_slt_149541_comb;
    p5_or_149542 <= p5_or_149542_comb;
    p5_or_149543 <= p5_or_149543_comb;
    p5_slt_149544 <= p5_slt_149544_comb;
    p5_slt_149545 <= p5_slt_149545_comb;
    p5_or_149546 <= p5_or_149546_comb;
    p5_sel_149565 <= p5_sel_149565_comb;
    p5_bit_slice_149568 <= p5_bit_slice_149568_comb;
    p5_bit_slice_149571 <= p5_bit_slice_149571_comb;
    p5_sel_149574 <= p5_sel_149574_comb;
    p5_bit_slice_149577 <= p5_bit_slice_149577_comb;
    p5_bit_slice_149580 <= p5_bit_slice_149580_comb;
    p5_bit_slice_149583 <= p5_bit_slice_149583_comb;
    p5_bit_slice_149586 <= p5_bit_slice_149586_comb;
    p5_sel_149589 <= p5_sel_149589_comb;
    p5_sel_149600 <= p5_sel_149600_comb;
    p5_bit_slice_149603 <= p5_bit_slice_149603_comb;
    p5_bit_slice_149606 <= p5_bit_slice_149606_comb;
    p5_bit_slice_149609 <= p5_bit_slice_149609_comb;
    p5_bit_slice_149612 <= p5_bit_slice_149612_comb;
    p5_sel_149615 <= p5_sel_149615_comb;
    p5_sel_149618 <= p5_sel_149618_comb;
    p5_sel_149621 <= p5_sel_149621_comb;
    p5_sel_149624 <= p5_sel_149624_comb;
    p5_sel_149627 <= p5_sel_149627_comb;
    p5_sel_149630 <= p5_sel_149630_comb;
    p5_sel_149633 <= p5_sel_149633_comb;
    p5_sel_149636 <= p5_sel_149636_comb;
    p5_bit_slice_149637 <= p5_bit_slice_149637_comb;
    p5_sel_149644 <= p5_sel_149644_comb;
    p5_sel_149647 <= p5_sel_149647_comb;
    p5_bit_slice_149652 <= p5_bit_slice_149652_comb;
    p5_bit_slice_149653 <= p5_bit_slice_149653_comb;
    p5_bit_slice_149658 <= p5_bit_slice_149658_comb;
    p5_bit_slice_149659 <= p5_bit_slice_149659_comb;
    p5_bit_slice_149664 <= p5_bit_slice_149664_comb;
    p5_bit_slice_149665 <= p5_bit_slice_149665_comb;
    p5_sel_149672 <= p5_sel_149672_comb;
    p5_sel_149675 <= p5_sel_149675_comb;
    p5_bit_slice_149680 <= p5_bit_slice_149680_comb;
    p5_sel_149683 <= p5_sel_149683_comb;
    p5_sel_149686 <= p5_sel_149686_comb;
    p5_sel_149689 <= p5_sel_149689_comb;
    p5_sel_149692 <= p5_sel_149692_comb;
    p5_sel_149695 <= p5_sel_149695_comb;
    p5_sel_149698 <= p5_sel_149698_comb;
    p5_sel_149701 <= p5_sel_149701_comb;
    p5_sel_149704 <= p5_sel_149704_comb;
    p5_bit_slice_149705 <= p5_bit_slice_149705_comb;
    p5_sel_149712 <= p5_sel_149712_comb;
    p5_sel_149715 <= p5_sel_149715_comb;
    p5_bit_slice_149720 <= p5_bit_slice_149720_comb;
    p5_bit_slice_149721 <= p5_bit_slice_149721_comb;
    p5_bit_slice_149726 <= p5_bit_slice_149726_comb;
    p5_bit_slice_149727 <= p5_bit_slice_149727_comb;
    p5_bit_slice_149732 <= p5_bit_slice_149732_comb;
    p5_bit_slice_149733 <= p5_bit_slice_149733_comb;
    p5_sel_149740 <= p5_sel_149740_comb;
    p5_sel_149743 <= p5_sel_149743_comb;
    p5_bit_slice_149748 <= p5_bit_slice_149748_comb;
    p5_bit_slice_149751 <= p5_bit_slice_149751_comb;
    p5_sel_149754 <= p5_sel_149754_comb;
    p5_sel_149757 <= p5_sel_149757_comb;
    p5_bit_slice_149760 <= p5_bit_slice_149760_comb;
    p5_sel_149763 <= p5_sel_149763_comb;
    p5_sel_149766 <= p5_sel_149766_comb;
    p5_sel_149769 <= p5_sel_149769_comb;
    p5_sel_149772 <= p5_sel_149772_comb;
    p5_sel_149779 <= p5_sel_149779_comb;
    p5_sel_149782 <= p5_sel_149782_comb;
    p5_sel_149789 <= p5_sel_149789_comb;
    p5_sel_149792 <= p5_sel_149792_comb;
    p5_sel_149795 <= p5_sel_149795_comb;
    p5_sel_149798 <= p5_sel_149798_comb;
    p5_sel_149801 <= p5_sel_149801_comb;
    p5_bit_slice_149804 <= p5_bit_slice_149804_comb;
    p5_bit_slice_149807 <= p5_bit_slice_149807_comb;
    p5_sel_149810 <= p5_sel_149810_comb;
    p5_sel_149813 <= p5_sel_149813_comb;
    p5_sel_149824 <= p5_sel_149824_comb;
    p5_sel_149827 <= p5_sel_149827_comb;
    p5_sel_149830 <= p5_sel_149830_comb;
    p5_sel_149833 <= p5_sel_149833_comb;
    p5_sel_149836 <= p5_sel_149836_comb;
    p5_sel_149839 <= p5_sel_149839_comb;
    p5_sel_149842 <= p5_sel_149842_comb;
    p5_sel_149845 <= p5_sel_149845_comb;
    p5_sel_149848 <= p5_sel_149848_comb;
    p5_bit_slice_149851 <= p5_bit_slice_149851_comb;
    p5_sel_149856 <= p5_sel_149856_comb;
    p5_sel_149859 <= p5_sel_149859_comb;
    p5_bit_slice_149862 <= p5_bit_slice_149862_comb;
    p5_bit_slice_149867 <= p5_bit_slice_149867_comb;
    p5_bit_slice_149870 <= p5_bit_slice_149870_comb;
    p5_bit_slice_149871 <= p5_bit_slice_149871_comb;
    p5_bit_slice_149874 <= p5_bit_slice_149874_comb;
    p5_bit_slice_149879 <= p5_bit_slice_149879_comb;
    p5_sel_149884 <= p5_sel_149884_comb;
    p5_sel_149887 <= p5_sel_149887_comb;
    p5_bit_slice_149890 <= p5_bit_slice_149890_comb;
    p5_sel_149895 <= p5_sel_149895_comb;
    p5_sel_149898 <= p5_sel_149898_comb;
    p5_sel_149901 <= p5_sel_149901_comb;
    p5_sel_149904 <= p5_sel_149904_comb;
    p5_sel_149907 <= p5_sel_149907_comb;
    p5_sel_149910 <= p5_sel_149910_comb;
    p5_sel_149913 <= p5_sel_149913_comb;
    p5_sel_149916 <= p5_sel_149916_comb;
    p5_bit_slice_149919 <= p5_bit_slice_149919_comb;
    p5_sel_149924 <= p5_sel_149924_comb;
    p5_sel_149927 <= p5_sel_149927_comb;
    p5_bit_slice_149930 <= p5_bit_slice_149930_comb;
    p5_bit_slice_149935 <= p5_bit_slice_149935_comb;
    p5_bit_slice_149938 <= p5_bit_slice_149938_comb;
    p5_bit_slice_149939 <= p5_bit_slice_149939_comb;
    p5_bit_slice_149942 <= p5_bit_slice_149942_comb;
    p5_bit_slice_149947 <= p5_bit_slice_149947_comb;
    p5_sel_149952 <= p5_sel_149952_comb;
    p5_sel_149955 <= p5_sel_149955_comb;
    p5_bit_slice_149958 <= p5_bit_slice_149958_comb;
    p5_bit_slice_149963 <= p5_bit_slice_149963_comb;
    p5_sel_149966 <= p5_sel_149966_comb;
    p5_sel_149969 <= p5_sel_149969_comb;
    p5_bit_slice_149972 <= p5_bit_slice_149972_comb;
    p5_sel_149979 <= p5_sel_149979_comb;
    p5_sel_149982 <= p5_sel_149982_comb;
    p5_sgt_150003 <= p5_sgt_150003_comb;
    p5_sgt_150004 <= p5_sgt_150004_comb;
    p5_sgt_150005 <= p5_sgt_150005_comb;
    p5_sgt_150006 <= p5_sgt_150006_comb;
    p5_sgt_150007 <= p5_sgt_150007_comb;
    p5_sgt_150008 <= p5_sgt_150008_comb;
    p5_sgt_150009 <= p5_sgt_150009_comb;
    p5_sgt_150010 <= p5_sgt_150010_comb;
    p5_sgt_150011 <= p5_sgt_150011_comb;
    p5_sgt_150018 <= p5_sgt_150018_comb;
    p5_sgt_150019 <= p5_sgt_150019_comb;
    p5_sgt_150020 <= p5_sgt_150020_comb;
    p5_sgt_150021 <= p5_sgt_150021_comb;
    p5_sgt_150022 <= p5_sgt_150022_comb;
    p5_sgt_150023 <= p5_sgt_150023_comb;
    p5_sgt_150024 <= p5_sgt_150024_comb;
    p5_sgt_150025 <= p5_sgt_150025_comb;
    p5_sgt_150026 <= p5_sgt_150026_comb;
    p5_sgt_150027 <= p5_sgt_150027_comb;
    p5_sgt_150028 <= p5_sgt_150028_comb;
    p5_sgt_150029 <= p5_sgt_150029_comb;
    p5_sgt_150030 <= p5_sgt_150030_comb;
    p5_sgt_150031 <= p5_sgt_150031_comb;
    p5_sgt_150032 <= p5_sgt_150032_comb;
    p5_sgt_150033 <= p5_sgt_150033_comb;
    p5_sgt_150034 <= p5_sgt_150034_comb;
    p5_sgt_150035 <= p5_sgt_150035_comb;
    p5_sgt_150036 <= p5_sgt_150036_comb;
    p5_sgt_150037 <= p5_sgt_150037_comb;
    p5_sgt_150038 <= p5_sgt_150038_comb;
    p5_sgt_150039 <= p5_sgt_150039_comb;
    p5_sgt_150040 <= p5_sgt_150040_comb;
    p5_sgt_150041 <= p5_sgt_150041_comb;
    p5_sgt_150042 <= p5_sgt_150042_comb;
    p5_sgt_150043 <= p5_sgt_150043_comb;
    p5_sgt_150044 <= p5_sgt_150044_comb;
    p5_sgt_150045 <= p5_sgt_150045_comb;
    p5_sgt_150046 <= p5_sgt_150046_comb;
    p5_sgt_150047 <= p5_sgt_150047_comb;
    p5_sgt_150048 <= p5_sgt_150048_comb;
    p5_sgt_150049 <= p5_sgt_150049_comb;
    p5_sgt_150050 <= p5_sgt_150050_comb;
    p5_sgt_150051 <= p5_sgt_150051_comb;
    p5_sgt_150052 <= p5_sgt_150052_comb;
    p5_sgt_150053 <= p5_sgt_150053_comb;
    p5_sgt_150054 <= p5_sgt_150054_comb;
    p5_sgt_150055 <= p5_sgt_150055_comb;
    p5_sgt_150056 <= p5_sgt_150056_comb;
    p5_sgt_150057 <= p5_sgt_150057_comb;
    p5_sgt_150058 <= p5_sgt_150058_comb;
    p5_sgt_150059 <= p5_sgt_150059_comb;
    p5_sgt_150060 <= p5_sgt_150060_comb;
    p5_sgt_150061 <= p5_sgt_150061_comb;
    p5_sgt_150062 <= p5_sgt_150062_comb;
    p5_sgt_150063 <= p5_sgt_150063_comb;
    p5_sgt_150064 <= p5_sgt_150064_comb;
    p5_sgt_150065 <= p5_sgt_150065_comb;
    p5_sgt_150066 <= p5_sgt_150066_comb;
    p5_sgt_150067 <= p5_sgt_150067_comb;
    p5_sgt_150068 <= p5_sgt_150068_comb;
    p5_sgt_150069 <= p5_sgt_150069_comb;
    p5_sgt_150070 <= p5_sgt_150070_comb;
    p5_sgt_150071 <= p5_sgt_150071_comb;
    p5_sgt_150072 <= p5_sgt_150072_comb;
    p5_sgt_150073 <= p5_sgt_150073_comb;
    p5_sgt_150074 <= p5_sgt_150074_comb;
    p5_sgt_150075 <= p5_sgt_150075_comb;
    p5_sgt_150076 <= p5_sgt_150076_comb;
    p5_sgt_150077 <= p5_sgt_150077_comb;
    p5_sgt_150078 <= p5_sgt_150078_comb;
    p5_sgt_150082 <= p5_sgt_150082_comb;
    p5_sgt_150083 <= p5_sgt_150083_comb;
    p5_sgt_150087 <= p5_sgt_150087_comb;
    p5_sgt_150088 <= p5_sgt_150088_comb;
    p5_sgt_150089 <= p5_sgt_150089_comb;
    p5_sgt_150090 <= p5_sgt_150090_comb;
    p5_sgt_150091 <= p5_sgt_150091_comb;
    p5_sgt_150092 <= p5_sgt_150092_comb;
    p5_sgt_150093 <= p5_sgt_150093_comb;
    p5_sgt_150094 <= p5_sgt_150094_comb;
    p5_sgt_150095 <= p5_sgt_150095_comb;
    p5_sgt_150102 <= p5_sgt_150102_comb;
    p5_sgt_150103 <= p5_sgt_150103_comb;
    p5_sgt_150104 <= p5_sgt_150104_comb;
    p5_sgt_150105 <= p5_sgt_150105_comb;
    p5_sgt_150106 <= p5_sgt_150106_comb;
    p5_sgt_150107 <= p5_sgt_150107_comb;
    p5_sgt_150108 <= p5_sgt_150108_comb;
    p5_sgt_150109 <= p5_sgt_150109_comb;
    p5_sgt_150110 <= p5_sgt_150110_comb;
    p5_sgt_150111 <= p5_sgt_150111_comb;
    p5_sgt_150112 <= p5_sgt_150112_comb;
    p5_sgt_150113 <= p5_sgt_150113_comb;
    p5_sgt_150114 <= p5_sgt_150114_comb;
    p5_sgt_150115 <= p5_sgt_150115_comb;
    p5_sgt_150116 <= p5_sgt_150116_comb;
    p5_sgt_150117 <= p5_sgt_150117_comb;
    p5_sgt_150118 <= p5_sgt_150118_comb;
    p5_sgt_150119 <= p5_sgt_150119_comb;
    p5_sgt_150120 <= p5_sgt_150120_comb;
    p5_sgt_150121 <= p5_sgt_150121_comb;
    p5_sgt_150122 <= p5_sgt_150122_comb;
    p5_sgt_150123 <= p5_sgt_150123_comb;
    p5_sgt_150124 <= p5_sgt_150124_comb;
    p5_sgt_150125 <= p5_sgt_150125_comb;
    p5_sgt_150126 <= p5_sgt_150126_comb;
    p5_sgt_150127 <= p5_sgt_150127_comb;
    p5_sgt_150128 <= p5_sgt_150128_comb;
    p5_sgt_150129 <= p5_sgt_150129_comb;
    p5_sgt_150130 <= p5_sgt_150130_comb;
    p5_sgt_150131 <= p5_sgt_150131_comb;
    p5_sgt_150132 <= p5_sgt_150132_comb;
    p5_sgt_150133 <= p5_sgt_150133_comb;
    p5_sgt_150134 <= p5_sgt_150134_comb;
    p5_sgt_150135 <= p5_sgt_150135_comb;
    p5_sgt_150136 <= p5_sgt_150136_comb;
    p5_sgt_150137 <= p5_sgt_150137_comb;
    p5_sgt_150138 <= p5_sgt_150138_comb;
    p5_sgt_150139 <= p5_sgt_150139_comb;
    p5_sgt_150140 <= p5_sgt_150140_comb;
    p5_sgt_150141 <= p5_sgt_150141_comb;
    p5_sgt_150142 <= p5_sgt_150142_comb;
    p5_sgt_150143 <= p5_sgt_150143_comb;
    p5_sgt_150144 <= p5_sgt_150144_comb;
    p5_sgt_150145 <= p5_sgt_150145_comb;
    p5_sgt_150146 <= p5_sgt_150146_comb;
    p5_sgt_150147 <= p5_sgt_150147_comb;
    p5_sgt_150148 <= p5_sgt_150148_comb;
    p5_sgt_150149 <= p5_sgt_150149_comb;
    p5_sgt_150150 <= p5_sgt_150150_comb;
    p5_sgt_150151 <= p5_sgt_150151_comb;
    p5_sgt_150152 <= p5_sgt_150152_comb;
    p5_sgt_150153 <= p5_sgt_150153_comb;
    p5_sgt_150154 <= p5_sgt_150154_comb;
    p5_sgt_150158 <= p5_sgt_150158_comb;
    p5_sgt_150159 <= p5_sgt_150159_comb;
    p5_add_150163 <= p5_add_150163_comb;
    p5_add_150164 <= p5_add_150164_comb;
    p5_add_150165 <= p5_add_150165_comb;
    p5_add_150166 <= p5_add_150166_comb;
    p5_add_150167 <= p5_add_150167_comb;
    p5_add_150168 <= p5_add_150168_comb;
    p5_add_150169 <= p5_add_150169_comb;
    p5_add_150170 <= p5_add_150170_comb;
    p5_sel_150171 <= p5_sel_150171_comb;
    p5_sel_150172 <= p5_sel_150172_comb;
    p5_sel_150173 <= p5_sel_150173_comb;
    p5_sel_150174 <= p5_sel_150174_comb;
    p5_sel_150175 <= p5_sel_150175_comb;
    p5_sel_150176 <= p5_sel_150176_comb;
    p5_sel_150177 <= p5_sel_150177_comb;
    p5_sel_150178 <= p5_sel_150178_comb;
  end

  // ===== Pipe stage 6:
  wire [7:0] p6_smul_57326_TrailingBits___72_comb;
  wire [7:0] p6_smul_57326_TrailingBits___73_comb;
  wire [7:0] p6_smul_57326_TrailingBits___74_comb;
  wire [7:0] p6_smul_57326_TrailingBits___75_comb;
  wire [7:0] p6_smul_57326_TrailingBits___76_comb;
  wire [7:0] p6_smul_57326_TrailingBits___77_comb;
  wire [7:0] p6_smul_57326_TrailingBits___78_comb;
  wire [7:0] p6_smul_57326_TrailingBits___79_comb;
  wire [7:0] p6_smul_57326_TrailingBits___80_comb;
  wire [7:0] p6_smul_57326_TrailingBits___81_comb;
  wire [7:0] p6_smul_57326_TrailingBits___82_comb;
  wire [7:0] p6_smul_57326_TrailingBits___83_comb;
  wire [7:0] p6_smul_57326_TrailingBits___84_comb;
  wire [7:0] p6_smul_57326_TrailingBits___85_comb;
  wire [7:0] p6_smul_57326_TrailingBits___86_comb;
  wire [7:0] p6_smul_57326_TrailingBits___87_comb;
  wire [7:0] p6_smul_57326_TrailingBits___88_comb;
  wire [7:0] p6_smul_57326_TrailingBits___89_comb;
  wire [7:0] p6_smul_57326_TrailingBits___90_comb;
  wire [7:0] p6_smul_57326_TrailingBits___91_comb;
  wire [7:0] p6_smul_57326_TrailingBits___92_comb;
  wire [7:0] p6_smul_57326_TrailingBits___93_comb;
  wire [7:0] p6_smul_57326_TrailingBits___94_comb;
  wire [7:0] p6_smul_57326_TrailingBits___95_comb;
  wire [7:0] p6_smul_57326_TrailingBits___104_comb;
  wire [7:0] p6_smul_57326_TrailingBits___105_comb;
  wire [7:0] p6_smul_57326_TrailingBits___106_comb;
  wire [7:0] p6_smul_57326_TrailingBits___107_comb;
  wire [7:0] p6_smul_57326_TrailingBits___108_comb;
  wire [7:0] p6_smul_57326_TrailingBits___109_comb;
  wire [7:0] p6_smul_57326_TrailingBits___110_comb;
  wire [7:0] p6_smul_57326_TrailingBits___111_comb;
  wire [7:0] p6_smul_57326_TrailingBits___112_comb;
  wire [7:0] p6_smul_57326_TrailingBits___113_comb;
  wire [7:0] p6_smul_57326_TrailingBits___114_comb;
  wire [7:0] p6_smul_57326_TrailingBits___115_comb;
  wire [7:0] p6_smul_57326_TrailingBits___116_comb;
  wire [7:0] p6_smul_57326_TrailingBits___117_comb;
  wire [7:0] p6_smul_57326_TrailingBits___118_comb;
  wire [7:0] p6_smul_57326_TrailingBits___119_comb;
  wire [7:0] p6_smul_57326_TrailingBits___120_comb;
  wire [7:0] p6_smul_57326_TrailingBits___121_comb;
  wire [7:0] p6_smul_57326_TrailingBits___122_comb;
  wire [7:0] p6_smul_57326_TrailingBits___123_comb;
  wire [7:0] p6_smul_57326_TrailingBits___124_comb;
  wire [7:0] p6_smul_57326_TrailingBits___125_comb;
  wire [7:0] p6_smul_57326_TrailingBits___126_comb;
  wire [7:0] p6_smul_57326_TrailingBits___127_comb;
  wire [16:0] p6_smul_58222_NarrowedMult__comb;
  wire [16:0] p6_smul_58224_NarrowedMult__comb;
  wire [16:0] p6_smul_58234_NarrowedMult__comb;
  wire [16:0] p6_smul_58236_NarrowedMult__comb;
  wire [16:0] p6_smul_58238_NarrowedMult__comb;
  wire [16:0] p6_smul_58240_NarrowedMult__comb;
  wire [16:0] p6_smul_58250_NarrowedMult__comb;
  wire [16:0] p6_smul_58252_NarrowedMult__comb;
  wire [16:0] p6_smul_58254_NarrowedMult__comb;
  wire [16:0] p6_smul_58256_NarrowedMult__comb;
  wire [16:0] p6_smul_58266_NarrowedMult__comb;
  wire [16:0] p6_smul_58268_NarrowedMult__comb;
  wire [16:0] p6_smul_58270_NarrowedMult__comb;
  wire [16:0] p6_smul_58272_NarrowedMult__comb;
  wire [16:0] p6_smul_58282_NarrowedMult__comb;
  wire [16:0] p6_smul_58284_NarrowedMult__comb;
  wire [16:0] p6_smul_58286_NarrowedMult__comb;
  wire [16:0] p6_smul_58288_NarrowedMult__comb;
  wire [16:0] p6_smul_58298_NarrowedMult__comb;
  wire [16:0] p6_smul_58300_NarrowedMult__comb;
  wire [16:0] p6_smul_58302_NarrowedMult__comb;
  wire [16:0] p6_smul_58304_NarrowedMult__comb;
  wire [16:0] p6_smul_58314_NarrowedMult__comb;
  wire [16:0] p6_smul_58316_NarrowedMult__comb;
  wire [16:0] p6_smul_58318_NarrowedMult__comb;
  wire [16:0] p6_smul_58320_NarrowedMult__comb;
  wire [16:0] p6_smul_58330_NarrowedMult__comb;
  wire [16:0] p6_smul_58332_NarrowedMult__comb;
  wire [16:0] p6_smul_58334_NarrowedMult__comb;
  wire [16:0] p6_smul_58336_NarrowedMult__comb;
  wire [16:0] p6_smul_58346_NarrowedMult__comb;
  wire [16:0] p6_smul_58348_NarrowedMult__comb;
  wire [16:0] p6_smul_58478_NarrowedMult__comb;
  wire [16:0] p6_smul_58482_NarrowedMult__comb;
  wire [16:0] p6_smul_58488_NarrowedMult__comb;
  wire [16:0] p6_smul_58492_NarrowedMult__comb;
  wire [16:0] p6_smul_58494_NarrowedMult__comb;
  wire [16:0] p6_smul_58498_NarrowedMult__comb;
  wire [16:0] p6_smul_58504_NarrowedMult__comb;
  wire [16:0] p6_smul_58508_NarrowedMult__comb;
  wire [16:0] p6_smul_58510_NarrowedMult__comb;
  wire [16:0] p6_smul_58514_NarrowedMult__comb;
  wire [16:0] p6_smul_58520_NarrowedMult__comb;
  wire [16:0] p6_smul_58524_NarrowedMult__comb;
  wire [16:0] p6_smul_58526_NarrowedMult__comb;
  wire [16:0] p6_smul_58530_NarrowedMult__comb;
  wire [16:0] p6_smul_58536_NarrowedMult__comb;
  wire [16:0] p6_smul_58540_NarrowedMult__comb;
  wire [16:0] p6_smul_58542_NarrowedMult__comb;
  wire [16:0] p6_smul_58546_NarrowedMult__comb;
  wire [16:0] p6_smul_58552_NarrowedMult__comb;
  wire [16:0] p6_smul_58556_NarrowedMult__comb;
  wire [16:0] p6_smul_58558_NarrowedMult__comb;
  wire [16:0] p6_smul_58562_NarrowedMult__comb;
  wire [16:0] p6_smul_58568_NarrowedMult__comb;
  wire [16:0] p6_smul_58572_NarrowedMult__comb;
  wire [16:0] p6_smul_58574_NarrowedMult__comb;
  wire [16:0] p6_smul_58578_NarrowedMult__comb;
  wire [16:0] p6_smul_58584_NarrowedMult__comb;
  wire [16:0] p6_smul_58588_NarrowedMult__comb;
  wire [16:0] p6_smul_58590_NarrowedMult__comb;
  wire [16:0] p6_smul_58594_NarrowedMult__comb;
  wire [16:0] p6_smul_58600_NarrowedMult__comb;
  wire [16:0] p6_smul_58604_NarrowedMult__comb;
  wire [16:0] p6_smul_58606_NarrowedMult__comb;
  wire [16:0] p6_smul_58608_NarrowedMult__comb;
  wire [16:0] p6_smul_58610_NarrowedMult__comb;
  wire [16:0] p6_smul_58612_NarrowedMult__comb;
  wire [16:0] p6_smul_58614_NarrowedMult__comb;
  wire [16:0] p6_smul_58616_NarrowedMult__comb;
  wire [16:0] p6_smul_58618_NarrowedMult__comb;
  wire [16:0] p6_smul_58620_NarrowedMult__comb;
  wire [16:0] p6_smul_58622_NarrowedMult__comb;
  wire [16:0] p6_smul_58624_NarrowedMult__comb;
  wire [16:0] p6_smul_58626_NarrowedMult__comb;
  wire [16:0] p6_smul_58628_NarrowedMult__comb;
  wire [16:0] p6_smul_58630_NarrowedMult__comb;
  wire [16:0] p6_smul_58632_NarrowedMult__comb;
  wire [16:0] p6_smul_58634_NarrowedMult__comb;
  wire [16:0] p6_smul_58636_NarrowedMult__comb;
  wire [16:0] p6_smul_58638_NarrowedMult__comb;
  wire [16:0] p6_smul_58640_NarrowedMult__comb;
  wire [16:0] p6_smul_58642_NarrowedMult__comb;
  wire [16:0] p6_smul_58644_NarrowedMult__comb;
  wire [16:0] p6_smul_58646_NarrowedMult__comb;
  wire [16:0] p6_smul_58648_NarrowedMult__comb;
  wire [16:0] p6_smul_58650_NarrowedMult__comb;
  wire [16:0] p6_smul_58652_NarrowedMult__comb;
  wire [16:0] p6_smul_58654_NarrowedMult__comb;
  wire [16:0] p6_smul_58656_NarrowedMult__comb;
  wire [16:0] p6_smul_58658_NarrowedMult__comb;
  wire [16:0] p6_smul_58660_NarrowedMult__comb;
  wire [16:0] p6_smul_58662_NarrowedMult__comb;
  wire [16:0] p6_smul_58664_NarrowedMult__comb;
  wire [16:0] p6_smul_58666_NarrowedMult__comb;
  wire [16:0] p6_smul_58668_NarrowedMult__comb;
  wire [16:0] p6_smul_58670_NarrowedMult__comb;
  wire [16:0] p6_smul_58672_NarrowedMult__comb;
  wire [16:0] p6_smul_58674_NarrowedMult__comb;
  wire [16:0] p6_smul_58676_NarrowedMult__comb;
  wire [16:0] p6_smul_58678_NarrowedMult__comb;
  wire [16:0] p6_smul_58680_NarrowedMult__comb;
  wire [16:0] p6_smul_58682_NarrowedMult__comb;
  wire [16:0] p6_smul_58684_NarrowedMult__comb;
  wire [16:0] p6_smul_58686_NarrowedMult__comb;
  wire [16:0] p6_smul_58688_NarrowedMult__comb;
  wire [16:0] p6_smul_58690_NarrowedMult__comb;
  wire [16:0] p6_smul_58692_NarrowedMult__comb;
  wire [16:0] p6_smul_58694_NarrowedMult__comb;
  wire [16:0] p6_smul_58696_NarrowedMult__comb;
  wire [16:0] p6_smul_58698_NarrowedMult__comb;
  wire [16:0] p6_smul_58700_NarrowedMult__comb;
  wire [16:0] p6_smul_58702_NarrowedMult__comb;
  wire [16:0] p6_smul_58704_NarrowedMult__comb;
  wire [16:0] p6_smul_58706_NarrowedMult__comb;
  wire [16:0] p6_smul_58708_NarrowedMult__comb;
  wire [16:0] p6_smul_58710_NarrowedMult__comb;
  wire [16:0] p6_smul_58712_NarrowedMult__comb;
  wire [16:0] p6_smul_58714_NarrowedMult__comb;
  wire [16:0] p6_smul_58716_NarrowedMult__comb;
  wire [16:0] p6_smul_58718_NarrowedMult__comb;
  wire [16:0] p6_smul_58720_NarrowedMult__comb;
  wire [16:0] p6_smul_58722_NarrowedMult__comb;
  wire [16:0] p6_smul_58724_NarrowedMult__comb;
  wire [16:0] p6_smul_58726_NarrowedMult__comb;
  wire [16:0] p6_smul_58728_NarrowedMult__comb;
  wire [16:0] p6_smul_58730_NarrowedMult__comb;
  wire [16:0] p6_smul_58732_NarrowedMult__comb;
  wire [16:0] p6_smul_58736_NarrowedMult__comb;
  wire [16:0] p6_smul_58740_NarrowedMult__comb;
  wire [16:0] p6_smul_58742_NarrowedMult__comb;
  wire [16:0] p6_smul_58746_NarrowedMult__comb;
  wire [16:0] p6_smul_58752_NarrowedMult__comb;
  wire [16:0] p6_smul_58756_NarrowedMult__comb;
  wire [16:0] p6_smul_58758_NarrowedMult__comb;
  wire [16:0] p6_smul_58762_NarrowedMult__comb;
  wire [16:0] p6_smul_58768_NarrowedMult__comb;
  wire [16:0] p6_smul_58772_NarrowedMult__comb;
  wire [16:0] p6_smul_58774_NarrowedMult__comb;
  wire [16:0] p6_smul_58778_NarrowedMult__comb;
  wire [16:0] p6_smul_58784_NarrowedMult__comb;
  wire [16:0] p6_smul_58788_NarrowedMult__comb;
  wire [16:0] p6_smul_58790_NarrowedMult__comb;
  wire [16:0] p6_smul_58794_NarrowedMult__comb;
  wire [16:0] p6_smul_58800_NarrowedMult__comb;
  wire [16:0] p6_smul_58804_NarrowedMult__comb;
  wire [16:0] p6_smul_58806_NarrowedMult__comb;
  wire [16:0] p6_smul_58810_NarrowedMult__comb;
  wire [16:0] p6_smul_58816_NarrowedMult__comb;
  wire [16:0] p6_smul_58820_NarrowedMult__comb;
  wire [16:0] p6_smul_58822_NarrowedMult__comb;
  wire [16:0] p6_smul_58826_NarrowedMult__comb;
  wire [16:0] p6_smul_58832_NarrowedMult__comb;
  wire [16:0] p6_smul_58836_NarrowedMult__comb;
  wire [16:0] p6_smul_58838_NarrowedMult__comb;
  wire [16:0] p6_smul_58842_NarrowedMult__comb;
  wire [16:0] p6_smul_58848_NarrowedMult__comb;
  wire [16:0] p6_smul_58852_NarrowedMult__comb;
  wire [16:0] p6_smul_58854_NarrowedMult__comb;
  wire [16:0] p6_smul_58858_NarrowedMult__comb;
  wire [16:0] p6_smul_58994_NarrowedMult__comb;
  wire [16:0] p6_smul_58996_NarrowedMult__comb;
  wire [16:0] p6_smul_58998_NarrowedMult__comb;
  wire [16:0] p6_smul_59000_NarrowedMult__comb;
  wire [16:0] p6_smul_59010_NarrowedMult__comb;
  wire [16:0] p6_smul_59012_NarrowedMult__comb;
  wire [16:0] p6_smul_59014_NarrowedMult__comb;
  wire [16:0] p6_smul_59016_NarrowedMult__comb;
  wire [16:0] p6_smul_59026_NarrowedMult__comb;
  wire [16:0] p6_smul_59028_NarrowedMult__comb;
  wire [16:0] p6_smul_59030_NarrowedMult__comb;
  wire [16:0] p6_smul_59032_NarrowedMult__comb;
  wire [16:0] p6_smul_59042_NarrowedMult__comb;
  wire [16:0] p6_smul_59044_NarrowedMult__comb;
  wire [16:0] p6_smul_59046_NarrowedMult__comb;
  wire [16:0] p6_smul_59048_NarrowedMult__comb;
  wire [16:0] p6_smul_59058_NarrowedMult__comb;
  wire [16:0] p6_smul_59060_NarrowedMult__comb;
  wire [16:0] p6_smul_59062_NarrowedMult__comb;
  wire [16:0] p6_smul_59064_NarrowedMult__comb;
  wire [16:0] p6_smul_59074_NarrowedMult__comb;
  wire [16:0] p6_smul_59076_NarrowedMult__comb;
  wire [16:0] p6_smul_59078_NarrowedMult__comb;
  wire [16:0] p6_smul_59080_NarrowedMult__comb;
  wire [16:0] p6_smul_59090_NarrowedMult__comb;
  wire [16:0] p6_smul_59092_NarrowedMult__comb;
  wire [16:0] p6_smul_59094_NarrowedMult__comb;
  wire [16:0] p6_smul_59096_NarrowedMult__comb;
  wire [16:0] p6_smul_59106_NarrowedMult__comb;
  wire [16:0] p6_smul_59108_NarrowedMult__comb;
  wire [16:0] p6_smul_59110_NarrowedMult__comb;
  wire [16:0] p6_smul_59112_NarrowedMult__comb;
  wire [31:0] p6_sum__520_comb;
  wire [31:0] p6_sum__521_comb;
  wire [31:0] p6_sum__522_comb;
  wire [31:0] p6_sum__523_comb;
  wire [31:0] p6_sum__296_comb;
  wire [31:0] p6_sum__297_comb;
  wire [31:0] p6_sum__298_comb;
  wire [31:0] p6_sum__299_comb;
  wire [15:0] p6_sel_152483_comb;
  wire [15:0] p6_sel_152484_comb;
  wire [15:0] p6_sel_152485_comb;
  wire [15:0] p6_sel_152486_comb;
  wire [15:0] p6_sel_152487_comb;
  wire [15:0] p6_sel_152488_comb;
  wire [15:0] p6_sel_152489_comb;
  wire [15:0] p6_sel_152490_comb;
  wire [15:0] p6_sel_152491_comb;
  wire [15:0] p6_sel_152492_comb;
  wire [15:0] p6_sel_152493_comb;
  wire [15:0] p6_sel_152494_comb;
  wire [15:0] p6_sel_152495_comb;
  wire [15:0] p6_sel_152496_comb;
  wire [15:0] p6_sel_152497_comb;
  wire [15:0] p6_sel_152498_comb;
  wire [15:0] p6_sel_152499_comb;
  wire [15:0] p6_sel_152500_comb;
  wire [15:0] p6_sel_152501_comb;
  wire [15:0] p6_sel_152502_comb;
  wire [15:0] p6_sel_152503_comb;
  wire [15:0] p6_sel_152504_comb;
  wire [15:0] p6_sel_152505_comb;
  wire [15:0] p6_sel_152506_comb;
  wire [15:0] p6_sel_152507_comb;
  wire [15:0] p6_sel_152508_comb;
  wire [15:0] p6_sel_152509_comb;
  wire [15:0] p6_sel_152510_comb;
  wire [15:0] p6_sel_152511_comb;
  wire [15:0] p6_sel_152512_comb;
  wire [15:0] p6_sel_152513_comb;
  wire [15:0] p6_sel_152514_comb;
  wire [15:0] p6_sel_152515_comb;
  wire [15:0] p6_sel_152516_comb;
  wire [15:0] p6_sel_152517_comb;
  wire [15:0] p6_sel_152518_comb;
  wire [15:0] p6_sel_152519_comb;
  wire [15:0] p6_sel_152520_comb;
  wire [15:0] p6_sel_152521_comb;
  wire [15:0] p6_sel_152522_comb;
  wire [15:0] p6_sel_152523_comb;
  wire [15:0] p6_sel_152524_comb;
  wire [15:0] p6_sel_152525_comb;
  wire [15:0] p6_sel_152526_comb;
  wire [15:0] p6_sel_152527_comb;
  wire [15:0] p6_sel_152528_comb;
  wire [15:0] p6_sel_152529_comb;
  wire [15:0] p6_sel_152530_comb;
  wire [15:0] p6_sel_155217_comb;
  wire [15:0] p6_sel_155218_comb;
  wire [15:0] p6_sel_155219_comb;
  wire [15:0] p6_sel_155220_comb;
  wire [15:0] p6_sel_155221_comb;
  wire [15:0] p6_sel_155222_comb;
  wire [15:0] p6_sel_155223_comb;
  wire [15:0] p6_sel_155224_comb;
  wire [15:0] p6_sel_155249_comb;
  wire [15:0] p6_sel_155250_comb;
  wire [15:0] p6_sel_155251_comb;
  wire [15:0] p6_sel_155252_comb;
  wire [15:0] p6_sel_155253_comb;
  wire [15:0] p6_sel_155254_comb;
  wire [15:0] p6_sel_155255_comb;
  wire [15:0] p6_sel_155256_comb;
  wire [15:0] p6_sel_155469_comb;
  wire [15:0] p6_sel_155470_comb;
  wire [15:0] p6_sel_155471_comb;
  wire [15:0] p6_sel_155472_comb;
  wire [15:0] p6_sel_155473_comb;
  wire [15:0] p6_sel_155474_comb;
  wire [15:0] p6_sel_155475_comb;
  wire [15:0] p6_sel_155476_comb;
  wire [15:0] p6_sel_155501_comb;
  wire [15:0] p6_sel_155502_comb;
  wire [15:0] p6_sel_155503_comb;
  wire [15:0] p6_sel_155504_comb;
  wire [15:0] p6_sel_155505_comb;
  wire [15:0] p6_sel_155506_comb;
  wire [15:0] p6_sel_155507_comb;
  wire [15:0] p6_sel_155508_comb;
  wire [31:0] p6_sum__524_comb;
  wire [31:0] p6_sum__525_comb;
  wire [31:0] p6_sum__300_comb;
  wire [31:0] p6_sum__301_comb;
  wire [15:0] p6_sel_155225_comb;
  wire [15:0] p6_sel_155226_comb;
  wire [15:0] p6_sel_155227_comb;
  wire [15:0] p6_sel_155228_comb;
  wire [15:0] p6_sel_155229_comb;
  wire [15:0] p6_sel_155230_comb;
  wire [15:0] p6_sel_155231_comb;
  wire [15:0] p6_sel_155232_comb;
  wire [15:0] p6_sel_155233_comb;
  wire [15:0] p6_sel_155234_comb;
  wire [15:0] p6_sel_155235_comb;
  wire [15:0] p6_sel_155236_comb;
  wire [15:0] p6_sel_155237_comb;
  wire [15:0] p6_sel_155238_comb;
  wire [15:0] p6_sel_155239_comb;
  wire [15:0] p6_sel_155240_comb;
  wire [15:0] p6_sel_155241_comb;
  wire [15:0] p6_sel_155242_comb;
  wire [15:0] p6_sel_155243_comb;
  wire [15:0] p6_sel_155244_comb;
  wire [15:0] p6_sel_155245_comb;
  wire [15:0] p6_sel_155246_comb;
  wire [15:0] p6_sel_155247_comb;
  wire [15:0] p6_sel_155248_comb;
  wire [15:0] p6_sel_155257_comb;
  wire [15:0] p6_sel_155258_comb;
  wire [15:0] p6_sel_155259_comb;
  wire [15:0] p6_sel_155260_comb;
  wire [15:0] p6_sel_155261_comb;
  wire [15:0] p6_sel_155262_comb;
  wire [15:0] p6_sel_155263_comb;
  wire [15:0] p6_sel_155264_comb;
  wire [15:0] p6_sel_155265_comb;
  wire [15:0] p6_sel_155266_comb;
  wire [15:0] p6_sel_155267_comb;
  wire [15:0] p6_sel_155268_comb;
  wire [15:0] p6_sel_155269_comb;
  wire [15:0] p6_sel_155270_comb;
  wire [15:0] p6_sel_155271_comb;
  wire [15:0] p6_sel_155272_comb;
  wire [15:0] p6_sel_155273_comb;
  wire [15:0] p6_sel_155274_comb;
  wire [15:0] p6_sel_155275_comb;
  wire [15:0] p6_sel_155276_comb;
  wire [15:0] p6_sel_155277_comb;
  wire [15:0] p6_sel_155278_comb;
  wire [15:0] p6_sel_155279_comb;
  wire [15:0] p6_sel_155280_comb;
  wire [15:0] p6_sel_155477_comb;
  wire [15:0] p6_sel_155478_comb;
  wire [15:0] p6_sel_155479_comb;
  wire [15:0] p6_sel_155480_comb;
  wire [15:0] p6_sel_155481_comb;
  wire [15:0] p6_sel_155482_comb;
  wire [15:0] p6_sel_155483_comb;
  wire [15:0] p6_sel_155484_comb;
  wire [15:0] p6_sel_155485_comb;
  wire [15:0] p6_sel_155486_comb;
  wire [15:0] p6_sel_155487_comb;
  wire [15:0] p6_sel_155488_comb;
  wire [15:0] p6_sel_155489_comb;
  wire [15:0] p6_sel_155490_comb;
  wire [15:0] p6_sel_155491_comb;
  wire [15:0] p6_sel_155492_comb;
  wire [15:0] p6_sel_155493_comb;
  wire [15:0] p6_sel_155494_comb;
  wire [15:0] p6_sel_155495_comb;
  wire [15:0] p6_sel_155496_comb;
  wire [15:0] p6_sel_155497_comb;
  wire [15:0] p6_sel_155498_comb;
  wire [15:0] p6_sel_155499_comb;
  wire [15:0] p6_sel_155500_comb;
  wire [15:0] p6_sel_155509_comb;
  wire [15:0] p6_sel_155510_comb;
  wire [15:0] p6_sel_155511_comb;
  wire [15:0] p6_sel_155512_comb;
  wire [15:0] p6_sel_155513_comb;
  wire [15:0] p6_sel_155514_comb;
  wire [15:0] p6_sel_155515_comb;
  wire [15:0] p6_sel_155516_comb;
  wire [15:0] p6_sel_155517_comb;
  wire [15:0] p6_sel_155518_comb;
  wire [15:0] p6_sel_155519_comb;
  wire [15:0] p6_sel_155520_comb;
  wire [15:0] p6_sel_155521_comb;
  wire [15:0] p6_sel_155522_comb;
  wire [15:0] p6_sel_155523_comb;
  wire [15:0] p6_sel_155524_comb;
  wire [15:0] p6_sel_155525_comb;
  wire [15:0] p6_sel_155526_comb;
  wire [15:0] p6_sel_155527_comb;
  wire [15:0] p6_sel_155528_comb;
  wire [15:0] p6_sel_155529_comb;
  wire [15:0] p6_sel_155530_comb;
  wire [15:0] p6_sel_155531_comb;
  wire [15:0] p6_sel_155532_comb;
  wire [31:0] p6_sum__526_comb;
  wire [31:0] p6_sum__302_comb;
  wire [16:0] p6_add_155131_comb;
  wire [16:0] p6_add_155132_comb;
  wire [16:0] p6_add_155133_comb;
  wire [16:0] p6_add_155134_comb;
  wire [16:0] p6_add_155135_comb;
  wire [16:0] p6_add_155136_comb;
  wire [16:0] p6_add_155137_comb;
  wire [16:0] p6_add_155138_comb;
  wire [16:0] p6_add_155139_comb;
  wire [16:0] p6_add_155140_comb;
  wire [16:0] p6_add_155141_comb;
  wire [16:0] p6_add_155142_comb;
  wire [16:0] p6_add_155143_comb;
  wire [16:0] p6_add_155144_comb;
  wire [16:0] p6_add_155145_comb;
  wire [16:0] p6_add_155146_comb;
  wire [16:0] p6_add_155147_comb;
  wire [16:0] p6_add_155148_comb;
  wire [16:0] p6_add_155149_comb;
  wire [16:0] p6_add_155150_comb;
  wire [16:0] p6_add_155151_comb;
  wire [16:0] p6_add_155152_comb;
  wire [16:0] p6_add_155153_comb;
  wire [16:0] p6_add_155154_comb;
  wire [15:0] p6_sel_155155_comb;
  wire [15:0] p6_sel_155156_comb;
  wire [15:0] p6_sel_155157_comb;
  wire [15:0] p6_sel_155158_comb;
  wire [15:0] p6_sel_155159_comb;
  wire [15:0] p6_sel_155160_comb;
  wire [15:0] p6_sel_155161_comb;
  wire [15:0] p6_sel_155162_comb;
  wire [15:0] p6_sel_155163_comb;
  wire [15:0] p6_sel_155164_comb;
  wire [15:0] p6_sel_155165_comb;
  wire [15:0] p6_sel_155166_comb;
  wire [15:0] p6_sel_155167_comb;
  wire [15:0] p6_sel_155168_comb;
  wire [15:0] p6_sel_155169_comb;
  wire [15:0] p6_sel_155170_comb;
  wire [15:0] p6_sel_155171_comb;
  wire [15:0] p6_sel_155172_comb;
  wire [15:0] p6_sel_155173_comb;
  wire [15:0] p6_sel_155174_comb;
  wire [15:0] p6_sel_155175_comb;
  wire [15:0] p6_sel_155176_comb;
  wire [15:0] p6_sel_155177_comb;
  wire [15:0] p6_sel_155178_comb;
  wire [15:0] p6_sel_155179_comb;
  wire [15:0] p6_sel_155180_comb;
  wire [15:0] p6_sel_155181_comb;
  wire [15:0] p6_sel_155182_comb;
  wire [15:0] p6_sel_155183_comb;
  wire [15:0] p6_sel_155184_comb;
  wire [15:0] p6_sel_155185_comb;
  wire [15:0] p6_sel_155186_comb;
  wire [15:0] p6_sel_155187_comb;
  wire [15:0] p6_sel_155188_comb;
  wire [15:0] p6_sel_155189_comb;
  wire [15:0] p6_sel_155190_comb;
  wire [15:0] p6_sel_155191_comb;
  wire [15:0] p6_sel_155192_comb;
  wire [15:0] p6_sel_155193_comb;
  wire [15:0] p6_sel_155194_comb;
  wire [15:0] p6_sel_155195_comb;
  wire [15:0] p6_sel_155196_comb;
  wire [15:0] p6_sel_155197_comb;
  wire [15:0] p6_sel_155198_comb;
  wire [15:0] p6_sel_155199_comb;
  wire [15:0] p6_sel_155200_comb;
  wire [15:0] p6_sel_155201_comb;
  wire [15:0] p6_sel_155202_comb;
  wire [15:0] p6_sel_155203_comb;
  wire [15:0] p6_sel_155204_comb;
  wire [15:0] p6_sel_155205_comb;
  wire [15:0] p6_sel_155206_comb;
  wire [15:0] p6_sel_155207_comb;
  wire [15:0] p6_sel_155208_comb;
  wire [15:0] p6_sel_155209_comb;
  wire [15:0] p6_sel_155210_comb;
  wire [15:0] p6_sel_155211_comb;
  wire [15:0] p6_sel_155212_comb;
  wire [15:0] p6_sel_155213_comb;
  wire [15:0] p6_sel_155214_comb;
  wire [15:0] p6_sel_155215_comb;
  wire [15:0] p6_sel_155216_comb;
  wire [15:0] p6_sel_155281_comb;
  wire [15:0] p6_sel_155282_comb;
  wire [15:0] p6_sel_155283_comb;
  wire [15:0] p6_sel_155284_comb;
  wire [15:0] p6_sel_155285_comb;
  wire [15:0] p6_sel_155286_comb;
  wire [15:0] p6_sel_155287_comb;
  wire [15:0] p6_sel_155288_comb;
  wire [15:0] p6_sel_155289_comb;
  wire [15:0] p6_sel_155290_comb;
  wire [15:0] p6_sel_155291_comb;
  wire [15:0] p6_sel_155292_comb;
  wire [15:0] p6_sel_155293_comb;
  wire [15:0] p6_sel_155294_comb;
  wire [15:0] p6_sel_155295_comb;
  wire [15:0] p6_sel_155296_comb;
  wire [15:0] p6_sel_155297_comb;
  wire [15:0] p6_sel_155298_comb;
  wire [15:0] p6_sel_155299_comb;
  wire [15:0] p6_sel_155300_comb;
  wire [15:0] p6_sel_155301_comb;
  wire [15:0] p6_sel_155302_comb;
  wire [15:0] p6_sel_155303_comb;
  wire [15:0] p6_sel_155304_comb;
  wire [15:0] p6_sel_155305_comb;
  wire [15:0] p6_sel_155306_comb;
  wire [15:0] p6_sel_155307_comb;
  wire [15:0] p6_sel_155308_comb;
  wire [15:0] p6_sel_155309_comb;
  wire [15:0] p6_sel_155310_comb;
  wire [15:0] p6_sel_155311_comb;
  wire [15:0] p6_sel_155312_comb;
  wire [15:0] p6_sel_155313_comb;
  wire [15:0] p6_sel_155314_comb;
  wire [15:0] p6_sel_155315_comb;
  wire [15:0] p6_sel_155316_comb;
  wire [15:0] p6_sel_155317_comb;
  wire [15:0] p6_sel_155318_comb;
  wire [15:0] p6_sel_155319_comb;
  wire [15:0] p6_sel_155320_comb;
  wire [15:0] p6_sel_155321_comb;
  wire [15:0] p6_sel_155322_comb;
  wire [15:0] p6_sel_155323_comb;
  wire [15:0] p6_sel_155324_comb;
  wire [15:0] p6_sel_155325_comb;
  wire [15:0] p6_sel_155326_comb;
  wire [15:0] p6_sel_155327_comb;
  wire [15:0] p6_sel_155328_comb;
  wire [15:0] p6_sel_155329_comb;
  wire [15:0] p6_sel_155330_comb;
  wire [15:0] p6_sel_155331_comb;
  wire [15:0] p6_sel_155332_comb;
  wire [15:0] p6_sel_155333_comb;
  wire [15:0] p6_sel_155334_comb;
  wire [15:0] p6_sel_155335_comb;
  wire [15:0] p6_sel_155336_comb;
  wire [15:0] p6_sel_155337_comb;
  wire [15:0] p6_sel_155338_comb;
  wire [15:0] p6_sel_155339_comb;
  wire [15:0] p6_sel_155340_comb;
  wire [15:0] p6_sel_155341_comb;
  wire [15:0] p6_sel_155342_comb;
  wire [15:0] p6_sel_155343_comb;
  wire [15:0] p6_sel_155344_comb;
  wire [15:0] p6_sel_155345_comb;
  wire [15:0] p6_sel_155346_comb;
  wire [15:0] p6_sel_155347_comb;
  wire [15:0] p6_sel_155348_comb;
  wire [15:0] p6_sel_155349_comb;
  wire [15:0] p6_sel_155350_comb;
  wire [15:0] p6_sel_155351_comb;
  wire [15:0] p6_sel_155352_comb;
  wire [15:0] p6_sel_155353_comb;
  wire [15:0] p6_sel_155354_comb;
  wire [15:0] p6_sel_155355_comb;
  wire [15:0] p6_sel_155356_comb;
  wire [15:0] p6_sel_155357_comb;
  wire [15:0] p6_sel_155358_comb;
  wire [15:0] p6_sel_155359_comb;
  wire [15:0] p6_sel_155360_comb;
  wire [15:0] p6_sel_155361_comb;
  wire [15:0] p6_sel_155362_comb;
  wire [15:0] p6_sel_155363_comb;
  wire [15:0] p6_sel_155364_comb;
  wire [15:0] p6_sel_155365_comb;
  wire [15:0] p6_sel_155366_comb;
  wire [15:0] p6_sel_155367_comb;
  wire [15:0] p6_sel_155368_comb;
  wire [15:0] p6_sel_155369_comb;
  wire [15:0] p6_sel_155370_comb;
  wire [15:0] p6_sel_155371_comb;
  wire [15:0] p6_sel_155372_comb;
  wire [15:0] p6_sel_155373_comb;
  wire [15:0] p6_sel_155374_comb;
  wire [15:0] p6_sel_155375_comb;
  wire [15:0] p6_sel_155376_comb;
  wire [15:0] p6_sel_155377_comb;
  wire [15:0] p6_sel_155378_comb;
  wire [15:0] p6_sel_155379_comb;
  wire [15:0] p6_sel_155380_comb;
  wire [15:0] p6_sel_155381_comb;
  wire [15:0] p6_sel_155382_comb;
  wire [15:0] p6_sel_155383_comb;
  wire [15:0] p6_sel_155384_comb;
  wire [15:0] p6_sel_155385_comb;
  wire [15:0] p6_sel_155386_comb;
  wire [15:0] p6_sel_155387_comb;
  wire [15:0] p6_sel_155388_comb;
  wire [15:0] p6_sel_155389_comb;
  wire [15:0] p6_sel_155390_comb;
  wire [15:0] p6_sel_155391_comb;
  wire [15:0] p6_sel_155392_comb;
  wire [15:0] p6_sel_155393_comb;
  wire [15:0] p6_sel_155394_comb;
  wire [15:0] p6_sel_155395_comb;
  wire [15:0] p6_sel_155396_comb;
  wire [15:0] p6_sel_155397_comb;
  wire [15:0] p6_sel_155398_comb;
  wire [15:0] p6_sel_155399_comb;
  wire [15:0] p6_sel_155400_comb;
  wire [15:0] p6_sel_155401_comb;
  wire [15:0] p6_sel_155402_comb;
  wire [15:0] p6_sel_155403_comb;
  wire [15:0] p6_sel_155404_comb;
  wire [15:0] p6_sel_155405_comb;
  wire [15:0] p6_sel_155406_comb;
  wire [15:0] p6_sel_155407_comb;
  wire [15:0] p6_sel_155408_comb;
  wire [15:0] p6_sel_155409_comb;
  wire [15:0] p6_sel_155410_comb;
  wire [15:0] p6_sel_155411_comb;
  wire [15:0] p6_sel_155412_comb;
  wire [15:0] p6_sel_155413_comb;
  wire [15:0] p6_sel_155414_comb;
  wire [15:0] p6_sel_155415_comb;
  wire [15:0] p6_sel_155416_comb;
  wire [15:0] p6_sel_155417_comb;
  wire [15:0] p6_sel_155418_comb;
  wire [15:0] p6_sel_155419_comb;
  wire [15:0] p6_sel_155420_comb;
  wire [15:0] p6_sel_155421_comb;
  wire [15:0] p6_sel_155422_comb;
  wire [15:0] p6_sel_155423_comb;
  wire [15:0] p6_sel_155424_comb;
  wire [15:0] p6_sel_155425_comb;
  wire [15:0] p6_sel_155426_comb;
  wire [15:0] p6_sel_155427_comb;
  wire [15:0] p6_sel_155428_comb;
  wire [15:0] p6_sel_155429_comb;
  wire [15:0] p6_sel_155430_comb;
  wire [15:0] p6_sel_155431_comb;
  wire [15:0] p6_sel_155432_comb;
  wire [15:0] p6_sel_155433_comb;
  wire [15:0] p6_sel_155434_comb;
  wire [15:0] p6_sel_155435_comb;
  wire [15:0] p6_sel_155436_comb;
  wire [15:0] p6_sel_155437_comb;
  wire [15:0] p6_sel_155438_comb;
  wire [15:0] p6_sel_155439_comb;
  wire [15:0] p6_sel_155440_comb;
  wire [15:0] p6_sel_155441_comb;
  wire [15:0] p6_sel_155442_comb;
  wire [15:0] p6_sel_155443_comb;
  wire [15:0] p6_sel_155444_comb;
  wire [15:0] p6_sel_155445_comb;
  wire [15:0] p6_sel_155446_comb;
  wire [15:0] p6_sel_155447_comb;
  wire [15:0] p6_sel_155448_comb;
  wire [15:0] p6_sel_155449_comb;
  wire [15:0] p6_sel_155450_comb;
  wire [15:0] p6_sel_155451_comb;
  wire [15:0] p6_sel_155452_comb;
  wire [15:0] p6_sel_155453_comb;
  wire [15:0] p6_sel_155454_comb;
  wire [15:0] p6_sel_155455_comb;
  wire [15:0] p6_sel_155456_comb;
  wire [15:0] p6_sel_155457_comb;
  wire [15:0] p6_sel_155458_comb;
  wire [15:0] p6_sel_155459_comb;
  wire [15:0] p6_sel_155460_comb;
  wire [15:0] p6_sel_155461_comb;
  wire [15:0] p6_sel_155462_comb;
  wire [15:0] p6_sel_155463_comb;
  wire [15:0] p6_sel_155464_comb;
  wire [15:0] p6_sel_155465_comb;
  wire [15:0] p6_sel_155466_comb;
  wire [15:0] p6_sel_155467_comb;
  wire [15:0] p6_sel_155468_comb;
  wire [15:0] p6_sel_155533_comb;
  wire [15:0] p6_sel_155534_comb;
  wire [15:0] p6_sel_155535_comb;
  wire [15:0] p6_sel_155536_comb;
  wire [15:0] p6_sel_155537_comb;
  wire [15:0] p6_sel_155538_comb;
  wire [15:0] p6_sel_155539_comb;
  wire [15:0] p6_sel_155540_comb;
  wire [15:0] p6_sel_155541_comb;
  wire [15:0] p6_sel_155542_comb;
  wire [15:0] p6_sel_155543_comb;
  wire [15:0] p6_sel_155544_comb;
  wire [15:0] p6_sel_155545_comb;
  wire [15:0] p6_sel_155546_comb;
  wire [15:0] p6_sel_155547_comb;
  wire [15:0] p6_sel_155548_comb;
  wire [15:0] p6_sel_155549_comb;
  wire [15:0] p6_sel_155550_comb;
  wire [15:0] p6_sel_155551_comb;
  wire [15:0] p6_sel_155552_comb;
  wire [15:0] p6_sel_155553_comb;
  wire [15:0] p6_sel_155554_comb;
  wire [15:0] p6_sel_155555_comb;
  wire [15:0] p6_sel_155556_comb;
  wire [15:0] p6_sel_155557_comb;
  wire [15:0] p6_sel_155558_comb;
  wire [15:0] p6_sel_155559_comb;
  wire [15:0] p6_sel_155560_comb;
  wire [15:0] p6_sel_155561_comb;
  wire [15:0] p6_sel_155562_comb;
  wire [15:0] p6_sel_155563_comb;
  wire [15:0] p6_sel_155564_comb;
  wire [15:0] p6_sel_155565_comb;
  wire [15:0] p6_sel_155566_comb;
  wire [15:0] p6_sel_155567_comb;
  wire [15:0] p6_sel_155568_comb;
  wire [15:0] p6_sel_155569_comb;
  wire [15:0] p6_sel_155570_comb;
  wire [15:0] p6_sel_155571_comb;
  wire [15:0] p6_sel_155572_comb;
  wire [15:0] p6_sel_155573_comb;
  wire [15:0] p6_sel_155574_comb;
  wire [15:0] p6_sel_155575_comb;
  wire [15:0] p6_sel_155576_comb;
  wire [15:0] p6_sel_155577_comb;
  wire [15:0] p6_sel_155578_comb;
  wire [15:0] p6_sel_155579_comb;
  wire [15:0] p6_sel_155580_comb;
  wire [15:0] p6_sel_155581_comb;
  wire [15:0] p6_sel_155582_comb;
  wire [15:0] p6_sel_155583_comb;
  wire [15:0] p6_sel_155584_comb;
  wire [15:0] p6_sel_155585_comb;
  wire [15:0] p6_sel_155586_comb;
  wire [15:0] p6_sel_155587_comb;
  wire [15:0] p6_sel_155588_comb;
  wire [15:0] p6_sel_155589_comb;
  wire [15:0] p6_sel_155590_comb;
  wire [15:0] p6_sel_155591_comb;
  wire [15:0] p6_sel_155592_comb;
  wire [15:0] p6_sel_155593_comb;
  wire [15:0] p6_sel_155594_comb;
  wire [16:0] p6_add_156123_comb;
  wire [16:0] p6_add_156124_comb;
  wire [16:0] p6_add_156125_comb;
  wire [16:0] p6_add_156126_comb;
  wire [16:0] p6_add_156139_comb;
  wire [16:0] p6_add_156140_comb;
  wire [16:0] p6_add_156141_comb;
  wire [16:0] p6_add_156142_comb;
  wire [16:0] p6_add_156251_comb;
  wire [16:0] p6_add_156252_comb;
  wire [16:0] p6_add_156253_comb;
  wire [16:0] p6_add_156254_comb;
  wire [16:0] p6_add_156267_comb;
  wire [16:0] p6_add_156268_comb;
  wire [16:0] p6_add_156269_comb;
  wire [16:0] p6_add_156270_comb;
  wire [31:0] p6_umul_156555_comb;
  wire [31:0] p6_umul_156559_comb;
  wire [31:0] p6_sum__464_comb;
  wire [31:0] p6_sum__465_comb;
  wire [31:0] p6_sum__466_comb;
  wire [31:0] p6_sum__467_comb;
  wire [31:0] p6_sum__408_comb;
  wire [31:0] p6_sum__409_comb;
  wire [31:0] p6_sum__410_comb;
  wire [31:0] p6_sum__411_comb;
  wire [31:0] p6_sum__352_comb;
  wire [31:0] p6_sum__353_comb;
  wire [31:0] p6_sum__354_comb;
  wire [31:0] p6_sum__355_comb;
  wire [31:0] p6_sum__240_comb;
  wire [31:0] p6_sum__241_comb;
  wire [31:0] p6_sum__242_comb;
  wire [31:0] p6_sum__243_comb;
  wire [31:0] p6_sum__184_comb;
  wire [31:0] p6_sum__185_comb;
  wire [31:0] p6_sum__186_comb;
  wire [31:0] p6_sum__187_comb;
  wire [31:0] p6_sum__128_comb;
  wire [31:0] p6_sum__129_comb;
  wire [31:0] p6_sum__130_comb;
  wire [31:0] p6_sum__131_comb;
  wire [16:0] p6_add_156127_comb;
  wire [16:0] p6_add_156128_comb;
  wire [16:0] p6_add_156129_comb;
  wire [16:0] p6_add_156130_comb;
  wire [16:0] p6_add_156131_comb;
  wire [16:0] p6_add_156132_comb;
  wire [16:0] p6_add_156133_comb;
  wire [16:0] p6_add_156134_comb;
  wire [16:0] p6_add_156135_comb;
  wire [16:0] p6_add_156136_comb;
  wire [16:0] p6_add_156137_comb;
  wire [16:0] p6_add_156138_comb;
  wire [16:0] p6_add_156143_comb;
  wire [16:0] p6_add_156144_comb;
  wire [16:0] p6_add_156145_comb;
  wire [16:0] p6_add_156146_comb;
  wire [16:0] p6_add_156147_comb;
  wire [16:0] p6_add_156148_comb;
  wire [16:0] p6_add_156149_comb;
  wire [16:0] p6_add_156150_comb;
  wire [16:0] p6_add_156151_comb;
  wire [16:0] p6_add_156152_comb;
  wire [16:0] p6_add_156153_comb;
  wire [16:0] p6_add_156154_comb;
  wire [16:0] p6_add_156255_comb;
  wire [16:0] p6_add_156256_comb;
  wire [16:0] p6_add_156257_comb;
  wire [16:0] p6_add_156258_comb;
  wire [16:0] p6_add_156259_comb;
  wire [16:0] p6_add_156260_comb;
  wire [16:0] p6_add_156261_comb;
  wire [16:0] p6_add_156262_comb;
  wire [16:0] p6_add_156263_comb;
  wire [16:0] p6_add_156264_comb;
  wire [16:0] p6_add_156265_comb;
  wire [16:0] p6_add_156266_comb;
  wire [16:0] p6_add_156271_comb;
  wire [16:0] p6_add_156272_comb;
  wire [16:0] p6_add_156273_comb;
  wire [16:0] p6_add_156274_comb;
  wire [16:0] p6_add_156275_comb;
  wire [16:0] p6_add_156276_comb;
  wire [16:0] p6_add_156277_comb;
  wire [16:0] p6_add_156278_comb;
  wire [16:0] p6_add_156279_comb;
  wire [16:0] p6_add_156280_comb;
  wire [16:0] p6_add_156281_comb;
  wire [16:0] p6_add_156282_comb;
  wire [24:0] p6_sum__1576_comb;
  wire [24:0] p6_sum__1577_comb;
  wire [24:0] p6_sum__1578_comb;
  wire [24:0] p6_sum__1579_comb;
  wire [24:0] p6_sum__1464_comb;
  wire [24:0] p6_sum__1465_comb;
  wire [24:0] p6_sum__1466_comb;
  wire [24:0] p6_sum__1467_comb;
  wire [24:0] p6_sum__1560_comb;
  wire [24:0] p6_sum__1561_comb;
  wire [24:0] p6_sum__1562_comb;
  wire [24:0] p6_sum__1563_comb;
  wire [24:0] p6_sum__1448_comb;
  wire [24:0] p6_sum__1449_comb;
  wire [24:0] p6_sum__1450_comb;
  wire [24:0] p6_sum__1451_comb;
  wire [31:0] p6_sum__468_comb;
  wire [31:0] p6_sum__469_comb;
  wire [31:0] p6_sum__412_comb;
  wire [31:0] p6_sum__413_comb;
  wire [31:0] p6_sum__356_comb;
  wire [31:0] p6_sum__357_comb;
  wire [31:0] p6_sum__244_comb;
  wire [31:0] p6_sum__245_comb;
  wire [31:0] p6_sum__188_comb;
  wire [31:0] p6_sum__189_comb;
  wire [31:0] p6_sum__132_comb;
  wire [31:0] p6_sum__133_comb;
  wire [16:0] p6_add_156091_comb;
  wire [16:0] p6_add_156092_comb;
  wire [16:0] p6_add_156093_comb;
  wire [16:0] p6_add_156094_comb;
  wire [16:0] p6_add_156095_comb;
  wire [16:0] p6_add_156096_comb;
  wire [16:0] p6_add_156097_comb;
  wire [16:0] p6_add_156098_comb;
  wire [16:0] p6_add_156099_comb;
  wire [16:0] p6_add_156100_comb;
  wire [16:0] p6_add_156101_comb;
  wire [16:0] p6_add_156102_comb;
  wire [16:0] p6_add_156103_comb;
  wire [16:0] p6_add_156104_comb;
  wire [16:0] p6_add_156105_comb;
  wire [16:0] p6_add_156106_comb;
  wire [16:0] p6_add_156107_comb;
  wire [16:0] p6_add_156108_comb;
  wire [16:0] p6_add_156109_comb;
  wire [16:0] p6_add_156110_comb;
  wire [16:0] p6_add_156111_comb;
  wire [16:0] p6_add_156112_comb;
  wire [16:0] p6_add_156113_comb;
  wire [16:0] p6_add_156114_comb;
  wire [16:0] p6_add_156115_comb;
  wire [16:0] p6_add_156116_comb;
  wire [16:0] p6_add_156117_comb;
  wire [16:0] p6_add_156118_comb;
  wire [16:0] p6_add_156119_comb;
  wire [16:0] p6_add_156120_comb;
  wire [16:0] p6_add_156121_comb;
  wire [16:0] p6_add_156122_comb;
  wire [16:0] p6_add_156155_comb;
  wire [16:0] p6_add_156156_comb;
  wire [16:0] p6_add_156157_comb;
  wire [16:0] p6_add_156158_comb;
  wire [16:0] p6_add_156159_comb;
  wire [16:0] p6_add_156160_comb;
  wire [16:0] p6_add_156161_comb;
  wire [16:0] p6_add_156162_comb;
  wire [16:0] p6_add_156163_comb;
  wire [16:0] p6_add_156164_comb;
  wire [16:0] p6_add_156165_comb;
  wire [16:0] p6_add_156166_comb;
  wire [16:0] p6_add_156167_comb;
  wire [16:0] p6_add_156168_comb;
  wire [16:0] p6_add_156169_comb;
  wire [16:0] p6_add_156170_comb;
  wire [16:0] p6_add_156171_comb;
  wire [16:0] p6_add_156172_comb;
  wire [16:0] p6_add_156173_comb;
  wire [16:0] p6_add_156174_comb;
  wire [16:0] p6_add_156175_comb;
  wire [16:0] p6_add_156176_comb;
  wire [16:0] p6_add_156177_comb;
  wire [16:0] p6_add_156178_comb;
  wire [16:0] p6_add_156179_comb;
  wire [16:0] p6_add_156180_comb;
  wire [16:0] p6_add_156181_comb;
  wire [16:0] p6_add_156182_comb;
  wire [16:0] p6_add_156183_comb;
  wire [16:0] p6_add_156184_comb;
  wire [16:0] p6_add_156185_comb;
  wire [16:0] p6_add_156186_comb;
  wire [16:0] p6_add_156187_comb;
  wire [16:0] p6_add_156188_comb;
  wire [16:0] p6_add_156189_comb;
  wire [16:0] p6_add_156190_comb;
  wire [16:0] p6_add_156191_comb;
  wire [16:0] p6_add_156192_comb;
  wire [16:0] p6_add_156193_comb;
  wire [16:0] p6_add_156194_comb;
  wire [16:0] p6_add_156195_comb;
  wire [16:0] p6_add_156196_comb;
  wire [16:0] p6_add_156197_comb;
  wire [16:0] p6_add_156198_comb;
  wire [16:0] p6_add_156199_comb;
  wire [16:0] p6_add_156200_comb;
  wire [16:0] p6_add_156201_comb;
  wire [16:0] p6_add_156202_comb;
  wire [16:0] p6_add_156203_comb;
  wire [16:0] p6_add_156204_comb;
  wire [16:0] p6_add_156205_comb;
  wire [16:0] p6_add_156206_comb;
  wire [16:0] p6_add_156207_comb;
  wire [16:0] p6_add_156208_comb;
  wire [16:0] p6_add_156209_comb;
  wire [16:0] p6_add_156210_comb;
  wire [16:0] p6_add_156211_comb;
  wire [16:0] p6_add_156212_comb;
  wire [16:0] p6_add_156213_comb;
  wire [16:0] p6_add_156214_comb;
  wire [16:0] p6_add_156215_comb;
  wire [16:0] p6_add_156216_comb;
  wire [16:0] p6_add_156217_comb;
  wire [16:0] p6_add_156218_comb;
  wire [16:0] p6_add_156219_comb;
  wire [16:0] p6_add_156220_comb;
  wire [16:0] p6_add_156221_comb;
  wire [16:0] p6_add_156222_comb;
  wire [16:0] p6_add_156223_comb;
  wire [16:0] p6_add_156224_comb;
  wire [16:0] p6_add_156225_comb;
  wire [16:0] p6_add_156226_comb;
  wire [16:0] p6_add_156227_comb;
  wire [16:0] p6_add_156228_comb;
  wire [16:0] p6_add_156229_comb;
  wire [16:0] p6_add_156230_comb;
  wire [16:0] p6_add_156231_comb;
  wire [16:0] p6_add_156232_comb;
  wire [16:0] p6_add_156233_comb;
  wire [16:0] p6_add_156234_comb;
  wire [16:0] p6_add_156235_comb;
  wire [16:0] p6_add_156236_comb;
  wire [16:0] p6_add_156237_comb;
  wire [16:0] p6_add_156238_comb;
  wire [16:0] p6_add_156239_comb;
  wire [16:0] p6_add_156240_comb;
  wire [16:0] p6_add_156241_comb;
  wire [16:0] p6_add_156242_comb;
  wire [16:0] p6_add_156243_comb;
  wire [16:0] p6_add_156244_comb;
  wire [16:0] p6_add_156245_comb;
  wire [16:0] p6_add_156246_comb;
  wire [16:0] p6_add_156247_comb;
  wire [16:0] p6_add_156248_comb;
  wire [16:0] p6_add_156249_comb;
  wire [16:0] p6_add_156250_comb;
  wire [16:0] p6_add_156283_comb;
  wire [16:0] p6_add_156284_comb;
  wire [16:0] p6_add_156285_comb;
  wire [16:0] p6_add_156286_comb;
  wire [16:0] p6_add_156287_comb;
  wire [16:0] p6_add_156288_comb;
  wire [16:0] p6_add_156289_comb;
  wire [16:0] p6_add_156290_comb;
  wire [16:0] p6_add_156291_comb;
  wire [16:0] p6_add_156292_comb;
  wire [16:0] p6_add_156293_comb;
  wire [16:0] p6_add_156294_comb;
  wire [16:0] p6_add_156295_comb;
  wire [16:0] p6_add_156296_comb;
  wire [16:0] p6_add_156297_comb;
  wire [16:0] p6_add_156298_comb;
  wire [16:0] p6_add_156299_comb;
  wire [16:0] p6_add_156300_comb;
  wire [16:0] p6_add_156301_comb;
  wire [16:0] p6_add_156302_comb;
  wire [16:0] p6_add_156303_comb;
  wire [16:0] p6_add_156304_comb;
  wire [16:0] p6_add_156305_comb;
  wire [16:0] p6_add_156306_comb;
  wire [16:0] p6_add_156307_comb;
  wire [16:0] p6_add_156308_comb;
  wire [16:0] p6_add_156309_comb;
  wire [16:0] p6_add_156310_comb;
  wire [16:0] p6_add_156311_comb;
  wire [16:0] p6_add_156312_comb;
  wire [16:0] p6_add_156313_comb;
  wire [16:0] p6_add_156314_comb;
  wire [24:0] p6_sum__1548_comb;
  wire [24:0] p6_sum__1549_comb;
  wire [24:0] p6_sum__1550_comb;
  wire [24:0] p6_sum__1551_comb;
  wire [24:0] p6_sum__1520_comb;
  wire [24:0] p6_sum__1521_comb;
  wire [24:0] p6_sum__1522_comb;
  wire [24:0] p6_sum__1523_comb;
  wire [24:0] p6_sum__1492_comb;
  wire [24:0] p6_sum__1493_comb;
  wire [24:0] p6_sum__1494_comb;
  wire [24:0] p6_sum__1495_comb;
  wire [24:0] p6_sum__1436_comb;
  wire [24:0] p6_sum__1437_comb;
  wire [24:0] p6_sum__1438_comb;
  wire [24:0] p6_sum__1439_comb;
  wire [24:0] p6_sum__1408_comb;
  wire [24:0] p6_sum__1409_comb;
  wire [24:0] p6_sum__1410_comb;
  wire [24:0] p6_sum__1411_comb;
  wire [24:0] p6_sum__1380_comb;
  wire [24:0] p6_sum__1381_comb;
  wire [24:0] p6_sum__1382_comb;
  wire [24:0] p6_sum__1383_comb;
  wire [24:0] p6_sum__1532_comb;
  wire [24:0] p6_sum__1533_comb;
  wire [24:0] p6_sum__1534_comb;
  wire [24:0] p6_sum__1535_comb;
  wire [24:0] p6_sum__1504_comb;
  wire [24:0] p6_sum__1505_comb;
  wire [24:0] p6_sum__1506_comb;
  wire [24:0] p6_sum__1507_comb;
  wire [24:0] p6_sum__1476_comb;
  wire [24:0] p6_sum__1477_comb;
  wire [24:0] p6_sum__1478_comb;
  wire [24:0] p6_sum__1479_comb;
  wire [24:0] p6_sum__1420_comb;
  wire [24:0] p6_sum__1421_comb;
  wire [24:0] p6_sum__1422_comb;
  wire [24:0] p6_sum__1423_comb;
  wire [24:0] p6_sum__1392_comb;
  wire [24:0] p6_sum__1393_comb;
  wire [24:0] p6_sum__1394_comb;
  wire [24:0] p6_sum__1395_comb;
  wire [24:0] p6_sum__1364_comb;
  wire [24:0] p6_sum__1365_comb;
  wire [24:0] p6_sum__1366_comb;
  wire [24:0] p6_sum__1367_comb;
  wire [24:0] p6_sum__1244_comb;
  wire [24:0] p6_sum__1245_comb;
  wire [24:0] p6_sum__1188_comb;
  wire [24:0] p6_sum__1189_comb;
  wire [24:0] p6_sum__1236_comb;
  wire [24:0] p6_sum__1237_comb;
  wire [24:0] p6_sum__1180_comb;
  wire [24:0] p6_sum__1181_comb;
  wire [24:0] p6_add_156699_comb;
  wire [24:0] p6_add_156700_comb;
  wire [31:0] p6_sum__470_comb;
  wire [31:0] p6_sum__414_comb;
  wire [31:0] p6_sum__358_comb;
  wire [31:0] p6_sum__246_comb;
  wire [31:0] p6_sum__190_comb;
  wire [31:0] p6_sum__134_comb;
  wire [24:0] p6_sum__1580_comb;
  wire [24:0] p6_sum__1581_comb;
  wire [24:0] p6_sum__1582_comb;
  wire [24:0] p6_sum__1583_comb;
  wire [24:0] p6_sum__1552_comb;
  wire [24:0] p6_sum__1553_comb;
  wire [24:0] p6_sum__1554_comb;
  wire [24:0] p6_sum__1555_comb;
  wire [24:0] p6_sum__1524_comb;
  wire [24:0] p6_sum__1525_comb;
  wire [24:0] p6_sum__1526_comb;
  wire [24:0] p6_sum__1527_comb;
  wire [24:0] p6_sum__1496_comb;
  wire [24:0] p6_sum__1497_comb;
  wire [24:0] p6_sum__1498_comb;
  wire [24:0] p6_sum__1499_comb;
  wire [24:0] p6_sum__1468_comb;
  wire [24:0] p6_sum__1469_comb;
  wire [24:0] p6_sum__1470_comb;
  wire [24:0] p6_sum__1471_comb;
  wire [24:0] p6_sum__1440_comb;
  wire [24:0] p6_sum__1441_comb;
  wire [24:0] p6_sum__1442_comb;
  wire [24:0] p6_sum__1443_comb;
  wire [24:0] p6_sum__1412_comb;
  wire [24:0] p6_sum__1413_comb;
  wire [24:0] p6_sum__1414_comb;
  wire [24:0] p6_sum__1415_comb;
  wire [24:0] p6_sum__1384_comb;
  wire [24:0] p6_sum__1385_comb;
  wire [24:0] p6_sum__1386_comb;
  wire [24:0] p6_sum__1387_comb;
  wire [24:0] p6_sum__1572_comb;
  wire [24:0] p6_sum__1573_comb;
  wire [24:0] p6_sum__1574_comb;
  wire [24:0] p6_sum__1575_comb;
  wire [24:0] p6_sum__1544_comb;
  wire [24:0] p6_sum__1545_comb;
  wire [24:0] p6_sum__1546_comb;
  wire [24:0] p6_sum__1547_comb;
  wire [24:0] p6_sum__1516_comb;
  wire [24:0] p6_sum__1517_comb;
  wire [24:0] p6_sum__1518_comb;
  wire [24:0] p6_sum__1519_comb;
  wire [24:0] p6_sum__1488_comb;
  wire [24:0] p6_sum__1489_comb;
  wire [24:0] p6_sum__1490_comb;
  wire [24:0] p6_sum__1491_comb;
  wire [24:0] p6_sum__1460_comb;
  wire [24:0] p6_sum__1461_comb;
  wire [24:0] p6_sum__1462_comb;
  wire [24:0] p6_sum__1463_comb;
  wire [24:0] p6_sum__1432_comb;
  wire [24:0] p6_sum__1433_comb;
  wire [24:0] p6_sum__1434_comb;
  wire [24:0] p6_sum__1435_comb;
  wire [24:0] p6_sum__1404_comb;
  wire [24:0] p6_sum__1405_comb;
  wire [24:0] p6_sum__1406_comb;
  wire [24:0] p6_sum__1407_comb;
  wire [24:0] p6_sum__1376_comb;
  wire [24:0] p6_sum__1377_comb;
  wire [24:0] p6_sum__1378_comb;
  wire [24:0] p6_sum__1379_comb;
  wire [24:0] p6_sum__1568_comb;
  wire [24:0] p6_sum__1569_comb;
  wire [24:0] p6_sum__1570_comb;
  wire [24:0] p6_sum__1571_comb;
  wire [24:0] p6_sum__1540_comb;
  wire [24:0] p6_sum__1541_comb;
  wire [24:0] p6_sum__1542_comb;
  wire [24:0] p6_sum__1543_comb;
  wire [24:0] p6_sum__1512_comb;
  wire [24:0] p6_sum__1513_comb;
  wire [24:0] p6_sum__1514_comb;
  wire [24:0] p6_sum__1515_comb;
  wire [24:0] p6_sum__1484_comb;
  wire [24:0] p6_sum__1485_comb;
  wire [24:0] p6_sum__1486_comb;
  wire [24:0] p6_sum__1487_comb;
  wire [24:0] p6_sum__1456_comb;
  wire [24:0] p6_sum__1457_comb;
  wire [24:0] p6_sum__1458_comb;
  wire [24:0] p6_sum__1459_comb;
  wire [24:0] p6_sum__1428_comb;
  wire [24:0] p6_sum__1429_comb;
  wire [24:0] p6_sum__1430_comb;
  wire [24:0] p6_sum__1431_comb;
  wire [24:0] p6_sum__1400_comb;
  wire [24:0] p6_sum__1401_comb;
  wire [24:0] p6_sum__1402_comb;
  wire [24:0] p6_sum__1403_comb;
  wire [24:0] p6_sum__1372_comb;
  wire [24:0] p6_sum__1373_comb;
  wire [24:0] p6_sum__1374_comb;
  wire [24:0] p6_sum__1375_comb;
  wire [24:0] p6_sum__1564_comb;
  wire [24:0] p6_sum__1565_comb;
  wire [24:0] p6_sum__1566_comb;
  wire [24:0] p6_sum__1567_comb;
  wire [24:0] p6_sum__1536_comb;
  wire [24:0] p6_sum__1537_comb;
  wire [24:0] p6_sum__1538_comb;
  wire [24:0] p6_sum__1539_comb;
  wire [24:0] p6_sum__1508_comb;
  wire [24:0] p6_sum__1509_comb;
  wire [24:0] p6_sum__1510_comb;
  wire [24:0] p6_sum__1511_comb;
  wire [24:0] p6_sum__1480_comb;
  wire [24:0] p6_sum__1481_comb;
  wire [24:0] p6_sum__1482_comb;
  wire [24:0] p6_sum__1483_comb;
  wire [24:0] p6_sum__1452_comb;
  wire [24:0] p6_sum__1453_comb;
  wire [24:0] p6_sum__1454_comb;
  wire [24:0] p6_sum__1455_comb;
  wire [24:0] p6_sum__1424_comb;
  wire [24:0] p6_sum__1425_comb;
  wire [24:0] p6_sum__1426_comb;
  wire [24:0] p6_sum__1427_comb;
  wire [24:0] p6_sum__1396_comb;
  wire [24:0] p6_sum__1397_comb;
  wire [24:0] p6_sum__1398_comb;
  wire [24:0] p6_sum__1399_comb;
  wire [24:0] p6_sum__1368_comb;
  wire [24:0] p6_sum__1369_comb;
  wire [24:0] p6_sum__1370_comb;
  wire [24:0] p6_sum__1371_comb;
  wire [24:0] p6_sum__1556_comb;
  wire [24:0] p6_sum__1557_comb;
  wire [24:0] p6_sum__1558_comb;
  wire [24:0] p6_sum__1559_comb;
  wire [24:0] p6_sum__1528_comb;
  wire [24:0] p6_sum__1529_comb;
  wire [24:0] p6_sum__1530_comb;
  wire [24:0] p6_sum__1531_comb;
  wire [24:0] p6_sum__1500_comb;
  wire [24:0] p6_sum__1501_comb;
  wire [24:0] p6_sum__1502_comb;
  wire [24:0] p6_sum__1503_comb;
  wire [24:0] p6_sum__1472_comb;
  wire [24:0] p6_sum__1473_comb;
  wire [24:0] p6_sum__1474_comb;
  wire [24:0] p6_sum__1475_comb;
  wire [24:0] p6_sum__1444_comb;
  wire [24:0] p6_sum__1445_comb;
  wire [24:0] p6_sum__1446_comb;
  wire [24:0] p6_sum__1447_comb;
  wire [24:0] p6_sum__1416_comb;
  wire [24:0] p6_sum__1417_comb;
  wire [24:0] p6_sum__1418_comb;
  wire [24:0] p6_sum__1419_comb;
  wire [24:0] p6_sum__1388_comb;
  wire [24:0] p6_sum__1389_comb;
  wire [24:0] p6_sum__1390_comb;
  wire [24:0] p6_sum__1391_comb;
  wire [24:0] p6_sum__1360_comb;
  wire [24:0] p6_sum__1361_comb;
  wire [24:0] p6_sum__1362_comb;
  wire [24:0] p6_sum__1363_comb;
  wire [24:0] p6_sum__1230_comb;
  wire [24:0] p6_sum__1231_comb;
  wire [24:0] p6_sum__1216_comb;
  wire [24:0] p6_sum__1217_comb;
  wire [24:0] p6_sum__1202_comb;
  wire [24:0] p6_sum__1203_comb;
  wire [24:0] p6_sum__1174_comb;
  wire [24:0] p6_sum__1175_comb;
  wire [24:0] p6_sum__1160_comb;
  wire [24:0] p6_sum__1161_comb;
  wire [24:0] p6_sum__1146_comb;
  wire [24:0] p6_sum__1147_comb;
  wire [24:0] p6_sum__1222_comb;
  wire [24:0] p6_sum__1223_comb;
  wire [24:0] p6_sum__1208_comb;
  wire [24:0] p6_sum__1209_comb;
  wire [24:0] p6_sum__1194_comb;
  wire [24:0] p6_sum__1195_comb;
  wire [24:0] p6_sum__1166_comb;
  wire [24:0] p6_sum__1167_comb;
  wire [24:0] p6_sum__1152_comb;
  wire [24:0] p6_sum__1153_comb;
  wire [24:0] p6_sum__1138_comb;
  wire [24:0] p6_sum__1139_comb;
  wire [24:0] p6_sum__1078_comb;
  wire [24:0] p6_sum__1050_comb;
  wire [24:0] p6_sum__1074_comb;
  wire [24:0] p6_sum__1046_comb;
  wire [31:0] p6_umul_156556_comb;
  wire [31:0] p6_umul_156557_comb;
  wire [31:0] p6_umul_156558_comb;
  wire [31:0] p6_umul_156560_comb;
  wire [31:0] p6_umul_156561_comb;
  wire [31:0] p6_umul_156562_comb;
  wire [24:0] p6_sum__1246_comb;
  wire [24:0] p6_sum__1247_comb;
  wire [24:0] p6_sum__1232_comb;
  wire [24:0] p6_sum__1233_comb;
  wire [24:0] p6_sum__1218_comb;
  wire [24:0] p6_sum__1219_comb;
  wire [24:0] p6_sum__1204_comb;
  wire [24:0] p6_sum__1205_comb;
  wire [24:0] p6_sum__1190_comb;
  wire [24:0] p6_sum__1191_comb;
  wire [24:0] p6_sum__1176_comb;
  wire [24:0] p6_sum__1177_comb;
  wire [24:0] p6_sum__1162_comb;
  wire [24:0] p6_sum__1163_comb;
  wire [24:0] p6_sum__1148_comb;
  wire [24:0] p6_sum__1149_comb;
  wire [24:0] p6_sum__1242_comb;
  wire [24:0] p6_sum__1243_comb;
  wire [24:0] p6_sum__1228_comb;
  wire [24:0] p6_sum__1229_comb;
  wire [24:0] p6_sum__1214_comb;
  wire [24:0] p6_sum__1215_comb;
  wire [24:0] p6_sum__1200_comb;
  wire [24:0] p6_sum__1201_comb;
  wire [24:0] p6_sum__1186_comb;
  wire [24:0] p6_sum__1187_comb;
  wire [24:0] p6_sum__1172_comb;
  wire [24:0] p6_sum__1173_comb;
  wire [24:0] p6_sum__1158_comb;
  wire [24:0] p6_sum__1159_comb;
  wire [24:0] p6_sum__1144_comb;
  wire [24:0] p6_sum__1145_comb;
  wire [24:0] p6_sum__1240_comb;
  wire [24:0] p6_sum__1241_comb;
  wire [24:0] p6_sum__1226_comb;
  wire [24:0] p6_sum__1227_comb;
  wire [24:0] p6_sum__1212_comb;
  wire [24:0] p6_sum__1213_comb;
  wire [24:0] p6_sum__1198_comb;
  wire [24:0] p6_sum__1199_comb;
  wire [24:0] p6_sum__1184_comb;
  wire [24:0] p6_sum__1185_comb;
  wire [24:0] p6_sum__1170_comb;
  wire [24:0] p6_sum__1171_comb;
  wire [24:0] p6_sum__1156_comb;
  wire [24:0] p6_sum__1157_comb;
  wire [24:0] p6_sum__1142_comb;
  wire [24:0] p6_sum__1143_comb;
  wire [24:0] p6_sum__1238_comb;
  wire [24:0] p6_sum__1239_comb;
  wire [24:0] p6_sum__1224_comb;
  wire [24:0] p6_sum__1225_comb;
  wire [24:0] p6_sum__1210_comb;
  wire [24:0] p6_sum__1211_comb;
  wire [24:0] p6_sum__1196_comb;
  wire [24:0] p6_sum__1197_comb;
  wire [24:0] p6_sum__1182_comb;
  wire [24:0] p6_sum__1183_comb;
  wire [24:0] p6_sum__1168_comb;
  wire [24:0] p6_sum__1169_comb;
  wire [24:0] p6_sum__1154_comb;
  wire [24:0] p6_sum__1155_comb;
  wire [24:0] p6_sum__1140_comb;
  wire [24:0] p6_sum__1141_comb;
  wire [24:0] p6_sum__1234_comb;
  wire [24:0] p6_sum__1235_comb;
  wire [24:0] p6_sum__1220_comb;
  wire [24:0] p6_sum__1221_comb;
  wire [24:0] p6_sum__1206_comb;
  wire [24:0] p6_sum__1207_comb;
  wire [24:0] p6_sum__1192_comb;
  wire [24:0] p6_sum__1193_comb;
  wire [24:0] p6_sum__1178_comb;
  wire [24:0] p6_sum__1179_comb;
  wire [24:0] p6_sum__1164_comb;
  wire [24:0] p6_sum__1165_comb;
  wire [24:0] p6_sum__1150_comb;
  wire [24:0] p6_sum__1151_comb;
  wire [24:0] p6_sum__1136_comb;
  wire [24:0] p6_sum__1137_comb;
  wire [24:0] p6_sum__1071_comb;
  wire [24:0] p6_sum__1064_comb;
  wire [24:0] p6_sum__1057_comb;
  wire [24:0] p6_sum__1043_comb;
  wire [24:0] p6_sum__1036_comb;
  wire [24:0] p6_sum__1029_comb;
  wire [24:0] p6_sum__1067_comb;
  wire [24:0] p6_sum__1060_comb;
  wire [24:0] p6_sum__1053_comb;
  wire [24:0] p6_sum__1039_comb;
  wire [24:0] p6_sum__1032_comb;
  wire [24:0] p6_sum__1025_comb;
  wire [24:0] p6_add_156701_comb;
  wire [24:0] p6_add_156702_comb;
  wire [24:0] p6_add_156703_comb;
  wire [24:0] p6_add_156704_comb;
  wire p6_sgt_156710_comb;
  wire [8:0] p6_bit_slice_156711_comb;
  wire p6_sgt_156713_comb;
  wire [8:0] p6_bit_slice_156714_comb;
  wire p6_slt_156715_comb;
  wire p6_slt_156716_comb;
  assign p6_smul_57326_TrailingBits___72_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___73_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___74_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___75_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___76_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___77_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___78_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___79_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___80_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___81_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___82_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___83_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___84_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___85_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___86_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___87_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___88_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___89_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___90_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___91_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___92_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___93_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___94_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___95_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___104_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___105_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___106_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___107_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___108_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___109_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___110_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___111_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___112_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___113_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___114_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___115_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___116_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___117_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___118_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___119_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___120_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___121_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___122_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___123_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___124_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___125_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___126_comb = 8'h00;
  assign p6_smul_57326_TrailingBits___127_comb = 8'h00;
  assign p6_smul_58222_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__64_squeezed, 9'h0fb);
  assign p6_smul_58224_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__65_squeezed, 9'h0d5);
  assign p6_smul_58234_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__70_squeezed, 9'h12b);
  assign p6_smul_58236_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__71_squeezed, 9'h105);
  assign p6_smul_58238_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__72_squeezed, 9'h0fb);
  assign p6_smul_58240_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__73_squeezed, 9'h0d5);
  assign p6_smul_58250_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__78_squeezed, 9'h12b);
  assign p6_smul_58252_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__79_squeezed, 9'h105);
  assign p6_smul_58254_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__80_squeezed, 9'h0fb);
  assign p6_smul_58256_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__81_squeezed, 9'h0d5);
  assign p6_smul_58266_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__86_squeezed, 9'h12b);
  assign p6_smul_58268_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__87_squeezed, 9'h105);
  assign p6_smul_58270_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__88_squeezed, 9'h0fb);
  assign p6_smul_58272_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__89_squeezed, 9'h0d5);
  assign p6_smul_58282_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__94_squeezed, 9'h12b);
  assign p6_smul_58284_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__95_squeezed, 9'h105);
  assign p6_smul_58286_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__96_squeezed, 9'h0fb);
  assign p6_smul_58288_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__97_squeezed, 9'h0d5);
  assign p6_smul_58298_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__102_squeezed, 9'h12b);
  assign p6_smul_58300_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__103_squeezed, 9'h105);
  assign p6_smul_58302_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__104_squeezed, 9'h0fb);
  assign p6_smul_58304_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__105_squeezed, 9'h0d5);
  assign p6_smul_58314_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__110_squeezed, 9'h12b);
  assign p6_smul_58316_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__111_squeezed, 9'h105);
  assign p6_smul_58318_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__112_squeezed, 9'h0fb);
  assign p6_smul_58320_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__113_squeezed, 9'h0d5);
  assign p6_smul_58330_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__118_squeezed, 9'h12b);
  assign p6_smul_58332_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__119_squeezed, 9'h105);
  assign p6_smul_58334_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__120_squeezed, 9'h0fb);
  assign p6_smul_58336_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__121_squeezed, 9'h0d5);
  assign p6_smul_58346_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__126_squeezed, 9'h12b);
  assign p6_smul_58348_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__127_squeezed, 9'h105);
  assign p6_smul_58478_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__64_squeezed, 9'h0d5);
  assign p6_smul_58482_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__66_squeezed, 9'h105);
  assign p6_smul_58488_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__69_squeezed, 9'h0fb);
  assign p6_smul_58492_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__71_squeezed, 9'h12b);
  assign p6_smul_58494_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__72_squeezed, 9'h0d5);
  assign p6_smul_58498_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__74_squeezed, 9'h105);
  assign p6_smul_58504_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__77_squeezed, 9'h0fb);
  assign p6_smul_58508_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__79_squeezed, 9'h12b);
  assign p6_smul_58510_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__80_squeezed, 9'h0d5);
  assign p6_smul_58514_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__82_squeezed, 9'h105);
  assign p6_smul_58520_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__85_squeezed, 9'h0fb);
  assign p6_smul_58524_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__87_squeezed, 9'h12b);
  assign p6_smul_58526_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__88_squeezed, 9'h0d5);
  assign p6_smul_58530_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__90_squeezed, 9'h105);
  assign p6_smul_58536_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__93_squeezed, 9'h0fb);
  assign p6_smul_58540_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__95_squeezed, 9'h12b);
  assign p6_smul_58542_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__96_squeezed, 9'h0d5);
  assign p6_smul_58546_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__98_squeezed, 9'h105);
  assign p6_smul_58552_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__101_squeezed, 9'h0fb);
  assign p6_smul_58556_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__103_squeezed, 9'h12b);
  assign p6_smul_58558_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__104_squeezed, 9'h0d5);
  assign p6_smul_58562_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__106_squeezed, 9'h105);
  assign p6_smul_58568_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__109_squeezed, 9'h0fb);
  assign p6_smul_58572_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__111_squeezed, 9'h12b);
  assign p6_smul_58574_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__112_squeezed, 9'h0d5);
  assign p6_smul_58578_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__114_squeezed, 9'h105);
  assign p6_smul_58584_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__117_squeezed, 9'h0fb);
  assign p6_smul_58588_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__119_squeezed, 9'h12b);
  assign p6_smul_58590_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__120_squeezed, 9'h0d5);
  assign p6_smul_58594_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__122_squeezed, 9'h105);
  assign p6_smul_58600_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__125_squeezed, 9'h0fb);
  assign p6_smul_58604_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__127_squeezed, 9'h12b);
  assign p6_smul_58606_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__64_squeezed, 9'h0b5);
  assign p6_smul_58608_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__65_squeezed, 9'h14b);
  assign p6_smul_58610_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__66_squeezed, 9'h14b);
  assign p6_smul_58612_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__67_squeezed, 9'h0b5);
  assign p6_smul_58614_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__68_squeezed, 9'h0b5);
  assign p6_smul_58616_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__69_squeezed, 9'h14b);
  assign p6_smul_58618_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__70_squeezed, 9'h14b);
  assign p6_smul_58620_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__71_squeezed, 9'h0b5);
  assign p6_smul_58622_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__72_squeezed, 9'h0b5);
  assign p6_smul_58624_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__73_squeezed, 9'h14b);
  assign p6_smul_58626_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__74_squeezed, 9'h14b);
  assign p6_smul_58628_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__75_squeezed, 9'h0b5);
  assign p6_smul_58630_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__76_squeezed, 9'h0b5);
  assign p6_smul_58632_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__77_squeezed, 9'h14b);
  assign p6_smul_58634_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__78_squeezed, 9'h14b);
  assign p6_smul_58636_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__79_squeezed, 9'h0b5);
  assign p6_smul_58638_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__80_squeezed, 9'h0b5);
  assign p6_smul_58640_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__81_squeezed, 9'h14b);
  assign p6_smul_58642_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__82_squeezed, 9'h14b);
  assign p6_smul_58644_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__83_squeezed, 9'h0b5);
  assign p6_smul_58646_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__84_squeezed, 9'h0b5);
  assign p6_smul_58648_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__85_squeezed, 9'h14b);
  assign p6_smul_58650_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__86_squeezed, 9'h14b);
  assign p6_smul_58652_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__87_squeezed, 9'h0b5);
  assign p6_smul_58654_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__88_squeezed, 9'h0b5);
  assign p6_smul_58656_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__89_squeezed, 9'h14b);
  assign p6_smul_58658_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__90_squeezed, 9'h14b);
  assign p6_smul_58660_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__91_squeezed, 9'h0b5);
  assign p6_smul_58662_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__92_squeezed, 9'h0b5);
  assign p6_smul_58664_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__93_squeezed, 9'h14b);
  assign p6_smul_58666_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__94_squeezed, 9'h14b);
  assign p6_smul_58668_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__95_squeezed, 9'h0b5);
  assign p6_smul_58670_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__96_squeezed, 9'h0b5);
  assign p6_smul_58672_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__97_squeezed, 9'h14b);
  assign p6_smul_58674_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__98_squeezed, 9'h14b);
  assign p6_smul_58676_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__99_squeezed, 9'h0b5);
  assign p6_smul_58678_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__100_squeezed, 9'h0b5);
  assign p6_smul_58680_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__101_squeezed, 9'h14b);
  assign p6_smul_58682_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__102_squeezed, 9'h14b);
  assign p6_smul_58684_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__103_squeezed, 9'h0b5);
  assign p6_smul_58686_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__104_squeezed, 9'h0b5);
  assign p6_smul_58688_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__105_squeezed, 9'h14b);
  assign p6_smul_58690_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__106_squeezed, 9'h14b);
  assign p6_smul_58692_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__107_squeezed, 9'h0b5);
  assign p6_smul_58694_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__108_squeezed, 9'h0b5);
  assign p6_smul_58696_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__109_squeezed, 9'h14b);
  assign p6_smul_58698_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__110_squeezed, 9'h14b);
  assign p6_smul_58700_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__111_squeezed, 9'h0b5);
  assign p6_smul_58702_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__112_squeezed, 9'h0b5);
  assign p6_smul_58704_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__113_squeezed, 9'h14b);
  assign p6_smul_58706_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__114_squeezed, 9'h14b);
  assign p6_smul_58708_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__115_squeezed, 9'h0b5);
  assign p6_smul_58710_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__116_squeezed, 9'h0b5);
  assign p6_smul_58712_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__117_squeezed, 9'h14b);
  assign p6_smul_58714_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__118_squeezed, 9'h14b);
  assign p6_smul_58716_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__119_squeezed, 9'h0b5);
  assign p6_smul_58718_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__120_squeezed, 9'h0b5);
  assign p6_smul_58720_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__121_squeezed, 9'h14b);
  assign p6_smul_58722_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__122_squeezed, 9'h14b);
  assign p6_smul_58724_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__123_squeezed, 9'h0b5);
  assign p6_smul_58726_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__124_squeezed, 9'h0b5);
  assign p6_smul_58728_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__125_squeezed, 9'h14b);
  assign p6_smul_58730_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__126_squeezed, 9'h14b);
  assign p6_smul_58732_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__127_squeezed, 9'h0b5);
  assign p6_smul_58736_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__65_squeezed, 9'h105);
  assign p6_smul_58740_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__67_squeezed, 9'h0d5);
  assign p6_smul_58742_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__68_squeezed, 9'h0d5);
  assign p6_smul_58746_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__70_squeezed, 9'h105);
  assign p6_smul_58752_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__73_squeezed, 9'h105);
  assign p6_smul_58756_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__75_squeezed, 9'h0d5);
  assign p6_smul_58758_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__76_squeezed, 9'h0d5);
  assign p6_smul_58762_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__78_squeezed, 9'h105);
  assign p6_smul_58768_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__81_squeezed, 9'h105);
  assign p6_smul_58772_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__83_squeezed, 9'h0d5);
  assign p6_smul_58774_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__84_squeezed, 9'h0d5);
  assign p6_smul_58778_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__86_squeezed, 9'h105);
  assign p6_smul_58784_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__89_squeezed, 9'h105);
  assign p6_smul_58788_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__91_squeezed, 9'h0d5);
  assign p6_smul_58790_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__92_squeezed, 9'h0d5);
  assign p6_smul_58794_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__94_squeezed, 9'h105);
  assign p6_smul_58800_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__97_squeezed, 9'h105);
  assign p6_smul_58804_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__99_squeezed, 9'h0d5);
  assign p6_smul_58806_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__100_squeezed, 9'h0d5);
  assign p6_smul_58810_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__102_squeezed, 9'h105);
  assign p6_smul_58816_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__105_squeezed, 9'h105);
  assign p6_smul_58820_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__107_squeezed, 9'h0d5);
  assign p6_smul_58822_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__108_squeezed, 9'h0d5);
  assign p6_smul_58826_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__110_squeezed, 9'h105);
  assign p6_smul_58832_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__113_squeezed, 9'h105);
  assign p6_smul_58836_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__115_squeezed, 9'h0d5);
  assign p6_smul_58838_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__116_squeezed, 9'h0d5);
  assign p6_smul_58842_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__118_squeezed, 9'h105);
  assign p6_smul_58848_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__121_squeezed, 9'h105);
  assign p6_smul_58852_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__123_squeezed, 9'h0d5);
  assign p6_smul_58854_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__124_squeezed, 9'h0d5);
  assign p6_smul_58858_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__126_squeezed, 9'h105);
  assign p6_smul_58994_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__66_squeezed, 9'h0d5);
  assign p6_smul_58996_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__67_squeezed, 9'h105);
  assign p6_smul_58998_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__68_squeezed, 9'h105);
  assign p6_smul_59000_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__69_squeezed, 9'h0d5);
  assign p6_smul_59010_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__74_squeezed, 9'h0d5);
  assign p6_smul_59012_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__75_squeezed, 9'h105);
  assign p6_smul_59014_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__76_squeezed, 9'h105);
  assign p6_smul_59016_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__77_squeezed, 9'h0d5);
  assign p6_smul_59026_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__82_squeezed, 9'h0d5);
  assign p6_smul_59028_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__83_squeezed, 9'h105);
  assign p6_smul_59030_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__84_squeezed, 9'h105);
  assign p6_smul_59032_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__85_squeezed, 9'h0d5);
  assign p6_smul_59042_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__90_squeezed, 9'h0d5);
  assign p6_smul_59044_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__91_squeezed, 9'h105);
  assign p6_smul_59046_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__92_squeezed, 9'h105);
  assign p6_smul_59048_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__93_squeezed, 9'h0d5);
  assign p6_smul_59058_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__98_squeezed, 9'h0d5);
  assign p6_smul_59060_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__99_squeezed, 9'h105);
  assign p6_smul_59062_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__100_squeezed, 9'h105);
  assign p6_smul_59064_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__101_squeezed, 9'h0d5);
  assign p6_smul_59074_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__106_squeezed, 9'h0d5);
  assign p6_smul_59076_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__107_squeezed, 9'h105);
  assign p6_smul_59078_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__108_squeezed, 9'h105);
  assign p6_smul_59080_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__109_squeezed, 9'h0d5);
  assign p6_smul_59090_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__114_squeezed, 9'h0d5);
  assign p6_smul_59092_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__115_squeezed, 9'h105);
  assign p6_smul_59094_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__116_squeezed, 9'h105);
  assign p6_smul_59096_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__117_squeezed, 9'h0d5);
  assign p6_smul_59106_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__122_squeezed, 9'h0d5);
  assign p6_smul_59108_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__123_squeezed, 9'h105);
  assign p6_smul_59110_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__124_squeezed, 9'h105);
  assign p6_smul_59112_NarrowedMult__comb = smul17b_8b_x_9b(p5_shifted__125_squeezed, 9'h0d5);
  assign p6_sum__520_comb = {{15{p5_add_150163[16]}}, p5_add_150163};
  assign p6_sum__521_comb = {{15{p5_add_150164[16]}}, p5_add_150164};
  assign p6_sum__522_comb = {{15{p5_add_150165[16]}}, p5_add_150165};
  assign p6_sum__523_comb = {{15{p5_add_150166[16]}}, p5_add_150166};
  assign p6_sum__296_comb = {{15{p5_add_150167[16]}}, p5_add_150167};
  assign p6_sum__297_comb = {{15{p5_add_150168[16]}}, p5_add_150168};
  assign p6_sum__298_comb = {{15{p5_add_150169[16]}}, p5_add_150169};
  assign p6_sum__299_comb = {{15{p5_add_150170[16]}}, p5_add_150170};
  assign p6_sel_152483_comb = p5_sgt_149059 ? 16'h7fff : {p5_sel_148221, p6_smul_57326_TrailingBits___72_comb};
  assign p6_sel_152484_comb = p5_sgt_149060 ? 16'h7fff : {p5_sel_148224, p6_smul_57326_TrailingBits___73_comb};
  assign p6_sel_152485_comb = p5_sgt_149061 ? 16'h7fff : {p5_sel_148227, p6_smul_57326_TrailingBits___74_comb};
  assign p6_sel_152486_comb = p5_sgt_149062 ? 16'h7fff : {p5_sel_148230, p6_smul_57326_TrailingBits___75_comb};
  assign p6_sel_152487_comb = p5_sgt_149063 ? 16'h7fff : {p5_sel_148233, p6_smul_57326_TrailingBits___76_comb};
  assign p6_sel_152488_comb = p5_sgt_149064 ? 16'h7fff : {p5_sel_148236, p6_smul_57326_TrailingBits___77_comb};
  assign p6_sel_152489_comb = p5_sgt_149065 ? 16'h7fff : {p5_sel_148239, p6_smul_57326_TrailingBits___78_comb};
  assign p6_sel_152490_comb = p5_sgt_149066 ? 16'h7fff : {p5_sel_148242, p6_smul_57326_TrailingBits___79_comb};
  assign p6_sel_152491_comb = p5_sgt_149067 ? 16'h7fff : {p5_sel_148245, p6_smul_57326_TrailingBits___80_comb};
  assign p6_sel_152492_comb = p5_sgt_149068 ? 16'h7fff : {p5_sel_148248, p6_smul_57326_TrailingBits___81_comb};
  assign p6_sel_152493_comb = p5_sgt_149069 ? 16'h7fff : {p5_sel_148251, p6_smul_57326_TrailingBits___82_comb};
  assign p6_sel_152494_comb = p5_sgt_149070 ? 16'h7fff : {p5_sel_148254, p6_smul_57326_TrailingBits___83_comb};
  assign p6_sel_152495_comb = p5_sgt_149071 ? 16'h7fff : {p5_sel_148257, p6_smul_57326_TrailingBits___84_comb};
  assign p6_sel_152496_comb = p5_sgt_149072 ? 16'h7fff : {p5_sel_148260, p6_smul_57326_TrailingBits___85_comb};
  assign p6_sel_152497_comb = p5_sgt_149073 ? 16'h7fff : {p5_sel_148263, p6_smul_57326_TrailingBits___86_comb};
  assign p6_sel_152498_comb = p5_sgt_149074 ? 16'h7fff : {p5_sel_148266, p6_smul_57326_TrailingBits___87_comb};
  assign p6_sel_152499_comb = p5_sgt_149075 ? 16'h7fff : {p5_sel_148269, p6_smul_57326_TrailingBits___88_comb};
  assign p6_sel_152500_comb = p5_sgt_149076 ? 16'h7fff : {p5_sel_148272, p6_smul_57326_TrailingBits___89_comb};
  assign p6_sel_152501_comb = p5_sgt_149077 ? 16'h7fff : {p5_sel_148275, p6_smul_57326_TrailingBits___90_comb};
  assign p6_sel_152502_comb = p5_sgt_149078 ? 16'h7fff : {p5_sel_148278, p6_smul_57326_TrailingBits___91_comb};
  assign p6_sel_152503_comb = p5_sgt_149079 ? 16'h7fff : {p5_sel_148281, p6_smul_57326_TrailingBits___92_comb};
  assign p6_sel_152504_comb = p5_sgt_149080 ? 16'h7fff : {p5_sel_148284, p6_smul_57326_TrailingBits___93_comb};
  assign p6_sel_152505_comb = p5_sgt_149081 ? 16'h7fff : {p5_sel_148287, p6_smul_57326_TrailingBits___94_comb};
  assign p6_sel_152506_comb = p5_sgt_149082 ? 16'h7fff : {p5_sel_148290, p6_smul_57326_TrailingBits___95_comb};
  assign p6_sel_152507_comb = p5_sgt_149107 ? 16'h7fff : {p5_sel_148325, p6_smul_57326_TrailingBits___104_comb};
  assign p6_sel_152508_comb = p5_sgt_149108 ? 16'h7fff : {p5_sel_148328, p6_smul_57326_TrailingBits___105_comb};
  assign p6_sel_152509_comb = p5_sgt_149109 ? 16'h7fff : {p5_sel_148331, p6_smul_57326_TrailingBits___106_comb};
  assign p6_sel_152510_comb = p5_sgt_149110 ? 16'h7fff : {p5_sel_148334, p6_smul_57326_TrailingBits___107_comb};
  assign p6_sel_152511_comb = p5_sgt_149111 ? 16'h7fff : {p5_sel_148337, p6_smul_57326_TrailingBits___108_comb};
  assign p6_sel_152512_comb = p5_sgt_149112 ? 16'h7fff : {p5_sel_148340, p6_smul_57326_TrailingBits___109_comb};
  assign p6_sel_152513_comb = p5_sgt_149113 ? 16'h7fff : {p5_sel_148343, p6_smul_57326_TrailingBits___110_comb};
  assign p6_sel_152514_comb = p5_sgt_149114 ? 16'h7fff : {p5_sel_148346, p6_smul_57326_TrailingBits___111_comb};
  assign p6_sel_152515_comb = p5_sgt_149115 ? 16'h7fff : {p5_sel_148349, p6_smul_57326_TrailingBits___112_comb};
  assign p6_sel_152516_comb = p5_sgt_149116 ? 16'h7fff : {p5_sel_148352, p6_smul_57326_TrailingBits___113_comb};
  assign p6_sel_152517_comb = p5_sgt_149117 ? 16'h7fff : {p5_sel_148355, p6_smul_57326_TrailingBits___114_comb};
  assign p6_sel_152518_comb = p5_sgt_149118 ? 16'h7fff : {p5_sel_148358, p6_smul_57326_TrailingBits___115_comb};
  assign p6_sel_152519_comb = p5_sgt_149119 ? 16'h7fff : {p5_sel_148361, p6_smul_57326_TrailingBits___116_comb};
  assign p6_sel_152520_comb = p5_sgt_149120 ? 16'h7fff : {p5_sel_148364, p6_smul_57326_TrailingBits___117_comb};
  assign p6_sel_152521_comb = p5_sgt_149121 ? 16'h7fff : {p5_sel_148367, p6_smul_57326_TrailingBits___118_comb};
  assign p6_sel_152522_comb = p5_sgt_149122 ? 16'h7fff : {p5_sel_148370, p6_smul_57326_TrailingBits___119_comb};
  assign p6_sel_152523_comb = p5_sgt_149123 ? 16'h7fff : {p5_sel_148373, p6_smul_57326_TrailingBits___120_comb};
  assign p6_sel_152524_comb = p5_sgt_149124 ? 16'h7fff : {p5_sel_148376, p6_smul_57326_TrailingBits___121_comb};
  assign p6_sel_152525_comb = p5_sgt_149125 ? 16'h7fff : {p5_sel_148379, p6_smul_57326_TrailingBits___122_comb};
  assign p6_sel_152526_comb = p5_sgt_149126 ? 16'h7fff : {p5_sel_148382, p6_smul_57326_TrailingBits___123_comb};
  assign p6_sel_152527_comb = p5_sgt_149127 ? 16'h7fff : {p5_sel_148385, p6_smul_57326_TrailingBits___124_comb};
  assign p6_sel_152528_comb = p5_sgt_149128 ? 16'h7fff : {p5_sel_148388, p6_smul_57326_TrailingBits___125_comb};
  assign p6_sel_152529_comb = p5_sgt_149129 ? 16'h7fff : {p5_sel_148391, p6_smul_57326_TrailingBits___126_comb};
  assign p6_sel_152530_comb = p5_sgt_149130 ? 16'h7fff : {p5_sel_148394, p6_smul_57326_TrailingBits___127_comb};
  assign p6_sel_155217_comb = p5_sgt_150023 ? 16'h7fff : {p5_sel_149615, 2'h0};
  assign p6_sel_155218_comb = p5_sgt_150024 ? 16'h7fff : {p5_sel_149618, 1'h0};
  assign p6_sel_155219_comb = p5_sgt_150025 ? 16'h7fff : {p5_sel_149621, 1'h0};
  assign p6_sel_155220_comb = p5_sgt_150026 ? 16'h7fff : {p5_sel_149624, 2'h0};
  assign p6_sel_155221_comb = p5_sgt_150027 ? 16'h7fff : {p5_sel_149627, 2'h0};
  assign p6_sel_155222_comb = p5_sgt_150028 ? 16'h7fff : {p5_sel_149630, 1'h0};
  assign p6_sel_155223_comb = p5_sgt_150029 ? 16'h7fff : {p5_sel_149633, 1'h0};
  assign p6_sel_155224_comb = p5_sgt_150030 ? 16'h7fff : {p5_sel_149636, 2'h0};
  assign p6_sel_155249_comb = p5_sgt_150047 ? 16'h7fff : {p5_sel_149683, 2'h0};
  assign p6_sel_155250_comb = p5_sgt_150048 ? 16'h7fff : {p5_sel_149686, 1'h0};
  assign p6_sel_155251_comb = p5_sgt_150049 ? 16'h7fff : {p5_sel_149689, 1'h0};
  assign p6_sel_155252_comb = p5_sgt_150050 ? 16'h7fff : {p5_sel_149692, 2'h0};
  assign p6_sel_155253_comb = p5_sgt_150051 ? 16'h7fff : {p5_sel_149695, 2'h0};
  assign p6_sel_155254_comb = p5_sgt_150052 ? 16'h7fff : {p5_sel_149698, 1'h0};
  assign p6_sel_155255_comb = p5_sgt_150053 ? 16'h7fff : {p5_sel_149701, 1'h0};
  assign p6_sel_155256_comb = p5_sgt_150054 ? 16'h7fff : {p5_sel_149704, 2'h0};
  assign p6_sel_155469_comb = p5_sgt_150103 ? 16'h7fff : {p5_sel_149827, 1'h0};
  assign p6_sel_155470_comb = p5_sgt_150104 ? 16'h7fff : {p5_sel_149830, 2'h0};
  assign p6_sel_155471_comb = p5_sgt_150105 ? 16'h7fff : {p5_sel_149833, 1'h0};
  assign p6_sel_155472_comb = p5_sgt_150106 ? 16'h7fff : {p5_sel_149836, 2'h0};
  assign p6_sel_155473_comb = p5_sgt_150107 ? 16'h7fff : {p5_sel_149839, 2'h0};
  assign p6_sel_155474_comb = p5_sgt_150108 ? 16'h7fff : {p5_sel_149842, 1'h0};
  assign p6_sel_155475_comb = p5_sgt_150109 ? 16'h7fff : {p5_sel_149845, 2'h0};
  assign p6_sel_155476_comb = p5_sgt_150110 ? 16'h7fff : {p5_sel_149848, 1'h0};
  assign p6_sel_155501_comb = p5_sgt_150127 ? 16'h7fff : {p5_sel_149895, 1'h0};
  assign p6_sel_155502_comb = p5_sgt_150128 ? 16'h7fff : {p5_sel_149898, 2'h0};
  assign p6_sel_155503_comb = p5_sgt_150129 ? 16'h7fff : {p5_sel_149901, 1'h0};
  assign p6_sel_155504_comb = p5_sgt_150130 ? 16'h7fff : {p5_sel_149904, 2'h0};
  assign p6_sel_155505_comb = p5_sgt_150131 ? 16'h7fff : {p5_sel_149907, 2'h0};
  assign p6_sel_155506_comb = p5_sgt_150132 ? 16'h7fff : {p5_sel_149910, 1'h0};
  assign p6_sel_155507_comb = p5_sgt_150133 ? 16'h7fff : {p5_sel_149913, 2'h0};
  assign p6_sel_155508_comb = p5_sgt_150134 ? 16'h7fff : {p5_sel_149916, 1'h0};
  assign p6_sum__524_comb = p6_sum__520_comb + p6_sum__521_comb;
  assign p6_sum__525_comb = p6_sum__522_comb + p6_sum__523_comb;
  assign p6_sum__300_comb = p6_sum__296_comb + p6_sum__297_comb;
  assign p6_sum__301_comb = p6_sum__298_comb + p6_sum__299_comb;
  assign p6_sel_155225_comb = $signed(p5_bit_slice_149637) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149191 ? 14'h2000 : p5_bit_slice_149192, 2'h0};
  assign p6_sel_155226_comb = p5_sgt_150031 ? 16'h7fff : {p5_slt_149193 ? 15'h4000 : p5_smul_58368_NarrowedMult_, 1'h0};
  assign p6_sel_155227_comb = p5_sgt_150032 ? 16'h7fff : {p5_slt_149194 ? 15'h4000 : p5_smul_58370_NarrowedMult_, 1'h0};
  assign p6_sel_155228_comb = p5_sgt_150033 ? 16'h7fff : {p5_sel_149644, 2'h0};
  assign p6_sel_155229_comb = p5_sgt_150034 ? 16'h7fff : {p5_sel_149647, 2'h0};
  assign p6_sel_155230_comb = p5_sgt_150035 ? 16'h7fff : {p5_slt_149201 ? 15'h4000 : p5_smul_58376_NarrowedMult_, 1'h0};
  assign p6_sel_155231_comb = p5_sgt_150036 ? 16'h7fff : {p5_slt_149202 ? 15'h4000 : p5_smul_58378_NarrowedMult_, 1'h0};
  assign p6_sel_155232_comb = $signed(p5_bit_slice_149652) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149203 ? 14'h2000 : p5_bit_slice_149204, 2'h0};
  assign p6_sel_155233_comb = $signed(p5_bit_slice_149653) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149205 ? 14'h2000 : p5_bit_slice_149206, 2'h0};
  assign p6_sel_155234_comb = p5_sgt_150037 ? 16'h7fff : {p5_slt_149207 ? 15'h4000 : p5_smul_58384_NarrowedMult_, 1'h0};
  assign p6_sel_155235_comb = p5_sgt_150038 ? 16'h7fff : {p5_slt_149208 ? 15'h4000 : p5_smul_58386_NarrowedMult_, 1'h0};
  assign p6_sel_155236_comb = $signed(p5_bit_slice_149658) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149209 ? 14'h2000 : p5_bit_slice_149210, 2'h0};
  assign p6_sel_155237_comb = $signed(p5_bit_slice_149659) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149211 ? 14'h2000 : p5_bit_slice_149212, 2'h0};
  assign p6_sel_155238_comb = p5_sgt_150039 ? 16'h7fff : {p5_slt_149213 ? 15'h4000 : p5_smul_58392_NarrowedMult_, 1'h0};
  assign p6_sel_155239_comb = p5_sgt_150040 ? 16'h7fff : {p5_slt_149214 ? 15'h4000 : p5_smul_58394_NarrowedMult_, 1'h0};
  assign p6_sel_155240_comb = $signed(p5_bit_slice_149664) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149215 ? 14'h2000 : p5_bit_slice_149216, 2'h0};
  assign p6_sel_155241_comb = $signed(p5_bit_slice_149665) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149217 ? 14'h2000 : p5_bit_slice_149218, 2'h0};
  assign p6_sel_155242_comb = p5_sgt_150041 ? 16'h7fff : {p5_slt_149219 ? 15'h4000 : p5_smul_58400_NarrowedMult_, 1'h0};
  assign p6_sel_155243_comb = p5_sgt_150042 ? 16'h7fff : {p5_slt_149220 ? 15'h4000 : p5_smul_58402_NarrowedMult_, 1'h0};
  assign p6_sel_155244_comb = p5_sgt_150043 ? 16'h7fff : {p5_sel_149672, 2'h0};
  assign p6_sel_155245_comb = p5_sgt_150044 ? 16'h7fff : {p5_sel_149675, 2'h0};
  assign p6_sel_155246_comb = p5_sgt_150045 ? 16'h7fff : {p5_slt_149227 ? 15'h4000 : p5_smul_58408_NarrowedMult_, 1'h0};
  assign p6_sel_155247_comb = p5_sgt_150046 ? 16'h7fff : {p5_slt_149228 ? 15'h4000 : p5_smul_58410_NarrowedMult_, 1'h0};
  assign p6_sel_155248_comb = $signed(p5_bit_slice_149680) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149229 ? 14'h2000 : p5_bit_slice_149230, 2'h0};
  assign p6_sel_155257_comb = $signed(p5_bit_slice_149705) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149251 ? 14'h2000 : p5_bit_slice_149252, 2'h0};
  assign p6_sel_155258_comb = p5_sgt_150055 ? 16'h7fff : {p5_slt_149253 ? 15'h4000 : p5_smul_58432_NarrowedMult_, 1'h0};
  assign p6_sel_155259_comb = p5_sgt_150056 ? 16'h7fff : {p5_slt_149254 ? 15'h4000 : p5_smul_58434_NarrowedMult_, 1'h0};
  assign p6_sel_155260_comb = p5_sgt_150057 ? 16'h7fff : {p5_sel_149712, 2'h0};
  assign p6_sel_155261_comb = p5_sgt_150058 ? 16'h7fff : {p5_sel_149715, 2'h0};
  assign p6_sel_155262_comb = p5_sgt_150059 ? 16'h7fff : {p5_slt_149261 ? 15'h4000 : p5_smul_58440_NarrowedMult_, 1'h0};
  assign p6_sel_155263_comb = p5_sgt_150060 ? 16'h7fff : {p5_slt_149262 ? 15'h4000 : p5_smul_58442_NarrowedMult_, 1'h0};
  assign p6_sel_155264_comb = $signed(p5_bit_slice_149720) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149263 ? 14'h2000 : p5_bit_slice_149264, 2'h0};
  assign p6_sel_155265_comb = $signed(p5_bit_slice_149721) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149265 ? 14'h2000 : p5_bit_slice_149266, 2'h0};
  assign p6_sel_155266_comb = p5_sgt_150061 ? 16'h7fff : {p5_slt_149267 ? 15'h4000 : p5_smul_58448_NarrowedMult_, 1'h0};
  assign p6_sel_155267_comb = p5_sgt_150062 ? 16'h7fff : {p5_slt_149268 ? 15'h4000 : p5_smul_58450_NarrowedMult_, 1'h0};
  assign p6_sel_155268_comb = $signed(p5_bit_slice_149726) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149269 ? 14'h2000 : p5_bit_slice_149270, 2'h0};
  assign p6_sel_155269_comb = $signed(p5_bit_slice_149727) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149271 ? 14'h2000 : p5_bit_slice_149272, 2'h0};
  assign p6_sel_155270_comb = p5_sgt_150063 ? 16'h7fff : {p5_slt_149273 ? 15'h4000 : p5_smul_58456_NarrowedMult_, 1'h0};
  assign p6_sel_155271_comb = p5_sgt_150064 ? 16'h7fff : {p5_slt_149274 ? 15'h4000 : p5_smul_58458_NarrowedMult_, 1'h0};
  assign p6_sel_155272_comb = $signed(p5_bit_slice_149732) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149275 ? 14'h2000 : p5_bit_slice_149276, 2'h0};
  assign p6_sel_155273_comb = $signed(p5_bit_slice_149733) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149277 ? 14'h2000 : p5_bit_slice_149278, 2'h0};
  assign p6_sel_155274_comb = p5_sgt_150065 ? 16'h7fff : {p5_slt_149279 ? 15'h4000 : p5_smul_58464_NarrowedMult_, 1'h0};
  assign p6_sel_155275_comb = p5_sgt_150066 ? 16'h7fff : {p5_slt_149280 ? 15'h4000 : p5_smul_58466_NarrowedMult_, 1'h0};
  assign p6_sel_155276_comb = p5_sgt_150067 ? 16'h7fff : {p5_sel_149740, 2'h0};
  assign p6_sel_155277_comb = p5_sgt_150068 ? 16'h7fff : {p5_sel_149743, 2'h0};
  assign p6_sel_155278_comb = p5_sgt_150069 ? 16'h7fff : {p5_slt_149287 ? 15'h4000 : p5_smul_58472_NarrowedMult_, 1'h0};
  assign p6_sel_155279_comb = p5_sgt_150070 ? 16'h7fff : {p5_slt_149288 ? 15'h4000 : p5_smul_58474_NarrowedMult_, 1'h0};
  assign p6_sel_155280_comb = $signed(p5_bit_slice_149748) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149289 ? 14'h2000 : p5_bit_slice_149290, 2'h0};
  assign p6_sel_155477_comb = p5_sgt_150111 ? 16'h7fff : {p5_slt_149407 ? 15'h4000 : p5_smul_58878_NarrowedMult_, 1'h0};
  assign p6_sel_155478_comb = $signed(p5_bit_slice_149851) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149408 ? 14'h2000 : p5_bit_slice_149409, 2'h0};
  assign p6_sel_155479_comb = p5_sgt_150112 ? 16'h7fff : {p5_slt_149410 ? 15'h4000 : p5_smul_58882_NarrowedMult_, 1'h0};
  assign p6_sel_155480_comb = p5_sgt_150113 ? 16'h7fff : {p5_sel_149856, 2'h0};
  assign p6_sel_155481_comb = p5_sgt_150114 ? 16'h7fff : {p5_sel_149859, 2'h0};
  assign p6_sel_155482_comb = p5_sgt_150115 ? 16'h7fff : {p5_slt_149417 ? 15'h4000 : p5_smul_58888_NarrowedMult_, 1'h0};
  assign p6_sel_155483_comb = $signed(p5_bit_slice_149862) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149418 ? 14'h2000 : p5_bit_slice_149419, 2'h0};
  assign p6_sel_155484_comb = p5_sgt_150116 ? 16'h7fff : {p5_slt_149420 ? 15'h4000 : p5_smul_58892_NarrowedMult_, 1'h0};
  assign p6_sel_155485_comb = p5_sgt_150117 ? 16'h7fff : {p5_slt_149421 ? 15'h4000 : p5_smul_58894_NarrowedMult_, 1'h0};
  assign p6_sel_155486_comb = $signed(p5_bit_slice_149867) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149422 ? 14'h2000 : p5_bit_slice_149423, 2'h0};
  assign p6_sel_155487_comb = p5_sgt_150118 ? 16'h7fff : {p5_slt_149424 ? 15'h4000 : p5_smul_58898_NarrowedMult_, 1'h0};
  assign p6_sel_155488_comb = $signed(p5_bit_slice_149870) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149425 ? 14'h2000 : p5_bit_slice_149426, 2'h0};
  assign p6_sel_155489_comb = $signed(p5_bit_slice_149871) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149427 ? 14'h2000 : p5_bit_slice_149428, 2'h0};
  assign p6_sel_155490_comb = p5_sgt_150119 ? 16'h7fff : {p5_slt_149429 ? 15'h4000 : p5_smul_58904_NarrowedMult_, 1'h0};
  assign p6_sel_155491_comb = $signed(p5_bit_slice_149874) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149430 ? 14'h2000 : p5_bit_slice_149431, 2'h0};
  assign p6_sel_155492_comb = p5_sgt_150120 ? 16'h7fff : {p5_slt_149432 ? 15'h4000 : p5_smul_58908_NarrowedMult_, 1'h0};
  assign p6_sel_155493_comb = p5_sgt_150121 ? 16'h7fff : {p5_slt_149433 ? 15'h4000 : p5_smul_58910_NarrowedMult_, 1'h0};
  assign p6_sel_155494_comb = $signed(p5_bit_slice_149879) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149434 ? 14'h2000 : p5_bit_slice_149435, 2'h0};
  assign p6_sel_155495_comb = p5_sgt_150122 ? 16'h7fff : {p5_slt_149436 ? 15'h4000 : p5_smul_58914_NarrowedMult_, 1'h0};
  assign p6_sel_155496_comb = p5_sgt_150123 ? 16'h7fff : {p5_sel_149884, 2'h0};
  assign p6_sel_155497_comb = p5_sgt_150124 ? 16'h7fff : {p5_sel_149887, 2'h0};
  assign p6_sel_155498_comb = p5_sgt_150125 ? 16'h7fff : {p5_slt_149443 ? 15'h4000 : p5_smul_58920_NarrowedMult_, 1'h0};
  assign p6_sel_155499_comb = $signed(p5_bit_slice_149890) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149444 ? 14'h2000 : p5_bit_slice_149445, 2'h0};
  assign p6_sel_155500_comb = p5_sgt_150126 ? 16'h7fff : {p5_slt_149446 ? 15'h4000 : p5_smul_58924_NarrowedMult_, 1'h0};
  assign p6_sel_155509_comb = p5_sgt_150135 ? 16'h7fff : {p5_slt_149467 ? 15'h4000 : p5_smul_58942_NarrowedMult_, 1'h0};
  assign p6_sel_155510_comb = $signed(p5_bit_slice_149919) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149468 ? 14'h2000 : p5_bit_slice_149469, 2'h0};
  assign p6_sel_155511_comb = p5_sgt_150136 ? 16'h7fff : {p5_slt_149470 ? 15'h4000 : p5_smul_58946_NarrowedMult_, 1'h0};
  assign p6_sel_155512_comb = p5_sgt_150137 ? 16'h7fff : {p5_sel_149924, 2'h0};
  assign p6_sel_155513_comb = p5_sgt_150138 ? 16'h7fff : {p5_sel_149927, 2'h0};
  assign p6_sel_155514_comb = p5_sgt_150139 ? 16'h7fff : {p5_slt_149477 ? 15'h4000 : p5_smul_58952_NarrowedMult_, 1'h0};
  assign p6_sel_155515_comb = $signed(p5_bit_slice_149930) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149478 ? 14'h2000 : p5_bit_slice_149479, 2'h0};
  assign p6_sel_155516_comb = p5_sgt_150140 ? 16'h7fff : {p5_slt_149480 ? 15'h4000 : p5_smul_58956_NarrowedMult_, 1'h0};
  assign p6_sel_155517_comb = p5_sgt_150141 ? 16'h7fff : {p5_slt_149481 ? 15'h4000 : p5_smul_58958_NarrowedMult_, 1'h0};
  assign p6_sel_155518_comb = $signed(p5_bit_slice_149935) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149482 ? 14'h2000 : p5_bit_slice_149483, 2'h0};
  assign p6_sel_155519_comb = p5_sgt_150142 ? 16'h7fff : {p5_slt_149484 ? 15'h4000 : p5_smul_58962_NarrowedMult_, 1'h0};
  assign p6_sel_155520_comb = $signed(p5_bit_slice_149938) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149485 ? 14'h2000 : p5_bit_slice_149486, 2'h0};
  assign p6_sel_155521_comb = $signed(p5_bit_slice_149939) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149487 ? 14'h2000 : p5_bit_slice_149488, 2'h0};
  assign p6_sel_155522_comb = p5_sgt_150143 ? 16'h7fff : {p5_slt_149489 ? 15'h4000 : p5_smul_58968_NarrowedMult_, 1'h0};
  assign p6_sel_155523_comb = $signed(p5_bit_slice_149942) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149490 ? 14'h2000 : p5_bit_slice_149491, 2'h0};
  assign p6_sel_155524_comb = p5_sgt_150144 ? 16'h7fff : {p5_slt_149492 ? 15'h4000 : p5_smul_58972_NarrowedMult_, 1'h0};
  assign p6_sel_155525_comb = p5_sgt_150145 ? 16'h7fff : {p5_slt_149493 ? 15'h4000 : p5_smul_58974_NarrowedMult_, 1'h0};
  assign p6_sel_155526_comb = $signed(p5_bit_slice_149947) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149494 ? 14'h2000 : p5_bit_slice_149495, 2'h0};
  assign p6_sel_155527_comb = p5_sgt_150146 ? 16'h7fff : {p5_slt_149496 ? 15'h4000 : p5_smul_58978_NarrowedMult_, 1'h0};
  assign p6_sel_155528_comb = p5_sgt_150147 ? 16'h7fff : {p5_sel_149952, 2'h0};
  assign p6_sel_155529_comb = p5_sgt_150148 ? 16'h7fff : {p5_sel_149955, 2'h0};
  assign p6_sel_155530_comb = p5_sgt_150149 ? 16'h7fff : {p5_slt_149503 ? 15'h4000 : p5_smul_58984_NarrowedMult_, 1'h0};
  assign p6_sel_155531_comb = $signed(p5_bit_slice_149958) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149504 ? 14'h2000 : p5_bit_slice_149505, 2'h0};
  assign p6_sel_155532_comb = p5_sgt_150150 ? 16'h7fff : {p5_slt_149506 ? 15'h4000 : p5_smul_58988_NarrowedMult_, 1'h0};
  assign p6_sum__526_comb = p6_sum__524_comb + p6_sum__525_comb;
  assign p6_sum__302_comb = p6_sum__300_comb + p6_sum__301_comb;
  assign p6_add_155131_comb = {{1{p6_sel_152483_comb[15]}}, p6_sel_152483_comb} + {{1{p6_sel_152484_comb[15]}}, p6_sel_152484_comb};
  assign p6_add_155132_comb = {{1{p6_sel_152485_comb[15]}}, p6_sel_152485_comb} + {{1{p6_sel_152486_comb[15]}}, p6_sel_152486_comb};
  assign p6_add_155133_comb = {{1{p6_sel_152487_comb[15]}}, p6_sel_152487_comb} + {{1{p6_sel_152488_comb[15]}}, p6_sel_152488_comb};
  assign p6_add_155134_comb = {{1{p6_sel_152489_comb[15]}}, p6_sel_152489_comb} + {{1{p6_sel_152490_comb[15]}}, p6_sel_152490_comb};
  assign p6_add_155135_comb = {{1{p6_sel_152491_comb[15]}}, p6_sel_152491_comb} + {{1{p6_sel_152492_comb[15]}}, p6_sel_152492_comb};
  assign p6_add_155136_comb = {{1{p6_sel_152493_comb[15]}}, p6_sel_152493_comb} + {{1{p6_sel_152494_comb[15]}}, p6_sel_152494_comb};
  assign p6_add_155137_comb = {{1{p6_sel_152495_comb[15]}}, p6_sel_152495_comb} + {{1{p6_sel_152496_comb[15]}}, p6_sel_152496_comb};
  assign p6_add_155138_comb = {{1{p6_sel_152497_comb[15]}}, p6_sel_152497_comb} + {{1{p6_sel_152498_comb[15]}}, p6_sel_152498_comb};
  assign p6_add_155139_comb = {{1{p6_sel_152499_comb[15]}}, p6_sel_152499_comb} + {{1{p6_sel_152500_comb[15]}}, p6_sel_152500_comb};
  assign p6_add_155140_comb = {{1{p6_sel_152501_comb[15]}}, p6_sel_152501_comb} + {{1{p6_sel_152502_comb[15]}}, p6_sel_152502_comb};
  assign p6_add_155141_comb = {{1{p6_sel_152503_comb[15]}}, p6_sel_152503_comb} + {{1{p6_sel_152504_comb[15]}}, p6_sel_152504_comb};
  assign p6_add_155142_comb = {{1{p6_sel_152505_comb[15]}}, p6_sel_152505_comb} + {{1{p6_sel_152506_comb[15]}}, p6_sel_152506_comb};
  assign p6_add_155143_comb = {{1{p6_sel_152507_comb[15]}}, p6_sel_152507_comb} + {{1{p6_sel_152508_comb[15]}}, p6_sel_152508_comb};
  assign p6_add_155144_comb = {{1{p6_sel_152509_comb[15]}}, p6_sel_152509_comb} + {{1{p6_sel_152510_comb[15]}}, p6_sel_152510_comb};
  assign p6_add_155145_comb = {{1{p6_sel_152511_comb[15]}}, p6_sel_152511_comb} + {{1{p6_sel_152512_comb[15]}}, p6_sel_152512_comb};
  assign p6_add_155146_comb = {{1{p6_sel_152513_comb[15]}}, p6_sel_152513_comb} + {{1{p6_sel_152514_comb[15]}}, p6_sel_152514_comb};
  assign p6_add_155147_comb = {{1{p6_sel_152515_comb[15]}}, p6_sel_152515_comb} + {{1{p6_sel_152516_comb[15]}}, p6_sel_152516_comb};
  assign p6_add_155148_comb = {{1{p6_sel_152517_comb[15]}}, p6_sel_152517_comb} + {{1{p6_sel_152518_comb[15]}}, p6_sel_152518_comb};
  assign p6_add_155149_comb = {{1{p6_sel_152519_comb[15]}}, p6_sel_152519_comb} + {{1{p6_sel_152520_comb[15]}}, p6_sel_152520_comb};
  assign p6_add_155150_comb = {{1{p6_sel_152521_comb[15]}}, p6_sel_152521_comb} + {{1{p6_sel_152522_comb[15]}}, p6_sel_152522_comb};
  assign p6_add_155151_comb = {{1{p6_sel_152523_comb[15]}}, p6_sel_152523_comb} + {{1{p6_sel_152524_comb[15]}}, p6_sel_152524_comb};
  assign p6_add_155152_comb = {{1{p6_sel_152525_comb[15]}}, p6_sel_152525_comb} + {{1{p6_sel_152526_comb[15]}}, p6_sel_152526_comb};
  assign p6_add_155153_comb = {{1{p6_sel_152527_comb[15]}}, p6_sel_152527_comb} + {{1{p6_sel_152528_comb[15]}}, p6_sel_152528_comb};
  assign p6_add_155154_comb = {{1{p6_sel_152529_comb[15]}}, p6_sel_152529_comb} + {{1{p6_sel_152530_comb[15]}}, p6_sel_152530_comb};
  assign p6_sel_155155_comb = $signed(p6_smul_58222_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58222_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58222_NarrowedMult__comb[15:0]);
  assign p6_sel_155156_comb = $signed(p6_smul_58224_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58224_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58224_NarrowedMult__comb[15:0]);
  assign p6_sel_155157_comb = p5_sgt_150003 ? 16'h7fff : {p5_sel_149565, 1'h0};
  assign p6_sel_155158_comb = p5_sgt_150004 ? 16'h7fff : {p5_bit_slice_149568, 1'h0};
  assign p6_sel_155159_comb = p5_sgt_150005 ? 16'h7fff : {p5_bit_slice_149571, 1'h0};
  assign p6_sel_155160_comb = p5_sgt_150006 ? 16'h7fff : {p5_sel_149574, 1'h0};
  assign p6_sel_155161_comb = $signed(p6_smul_58234_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58234_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58234_NarrowedMult__comb[15:0]);
  assign p6_sel_155162_comb = $signed(p6_smul_58236_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58236_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58236_NarrowedMult__comb[15:0]);
  assign p6_sel_155163_comb = $signed(p6_smul_58238_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58238_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58238_NarrowedMult__comb[15:0]);
  assign p6_sel_155164_comb = $signed(p6_smul_58240_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58240_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58240_NarrowedMult__comb[15:0]);
  assign p6_sel_155165_comb = $signed(p5_or_148407[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149139 ? 15'h4000 : p5_or_148407[23:9], 1'h0};
  assign p6_sel_155166_comb = p5_sgt_150007 ? 16'h7fff : {p5_bit_slice_149577, 1'h0};
  assign p6_sel_155167_comb = p5_sgt_150008 ? 16'h7fff : {p5_bit_slice_149580, 1'h0};
  assign p6_sel_155168_comb = $signed(p5_or_148414[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149142 ? 15'h4000 : p5_or_148414[23:9], 1'h0};
  assign p6_sel_155169_comb = $signed(p6_smul_58250_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58250_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58250_NarrowedMult__comb[15:0]);
  assign p6_sel_155170_comb = $signed(p6_smul_58252_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58252_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58252_NarrowedMult__comb[15:0]);
  assign p6_sel_155171_comb = $signed(p6_smul_58254_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58254_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58254_NarrowedMult__comb[15:0]);
  assign p6_sel_155172_comb = $signed(p6_smul_58256_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58256_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58256_NarrowedMult__comb[15:0]);
  assign p6_sel_155173_comb = $signed(p5_or_148417[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149143 ? 15'h4000 : p5_or_148417[23:9], 1'h0};
  assign p6_sel_155174_comb = $signed(p5_or_149144[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149144[23:9], 1'h0};
  assign p6_sel_155175_comb = $signed(p5_or_149145[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149145[23:9], 1'h0};
  assign p6_sel_155176_comb = $signed(p5_or_148424[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149146 ? 15'h4000 : p5_or_148424[23:9], 1'h0};
  assign p6_sel_155177_comb = $signed(p6_smul_58266_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58266_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58266_NarrowedMult__comb[15:0]);
  assign p6_sel_155178_comb = $signed(p6_smul_58268_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58268_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58268_NarrowedMult__comb[15:0]);
  assign p6_sel_155179_comb = $signed(p6_smul_58270_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58270_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58270_NarrowedMult__comb[15:0]);
  assign p6_sel_155180_comb = $signed(p6_smul_58272_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58272_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58272_NarrowedMult__comb[15:0]);
  assign p6_sel_155181_comb = $signed(p5_or_148427[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149147 ? 15'h4000 : p5_or_148427[23:9], 1'h0};
  assign p6_sel_155182_comb = p5_sgt_150009 ? 16'h7fff : {p5_bit_slice_149583, 1'h0};
  assign p6_sel_155183_comb = p5_sgt_150010 ? 16'h7fff : {p5_bit_slice_149586, 1'h0};
  assign p6_sel_155184_comb = $signed(p5_or_148434[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149150 ? 15'h4000 : p5_or_148434[23:9], 1'h0};
  assign p6_sel_155185_comb = $signed(p6_smul_58282_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58282_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58282_NarrowedMult__comb[15:0]);
  assign p6_sel_155186_comb = $signed(p6_smul_58284_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58284_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58284_NarrowedMult__comb[15:0]);
  assign p6_sel_155187_comb = $signed(p6_smul_58286_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58286_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58286_NarrowedMult__comb[15:0]);
  assign p6_sel_155188_comb = $signed(p6_smul_58288_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58288_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58288_NarrowedMult__comb[15:0]);
  assign p6_sel_155189_comb = p5_sgt_150011 ? 16'h7fff : {p5_sel_149589, 1'h0};
  assign p6_sel_155190_comb = p5_sgt_150018 ? 16'h7fff : {p5_sel_149600, 1'h0};
  assign p6_sel_155191_comb = $signed(p6_smul_58298_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58298_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58298_NarrowedMult__comb[15:0]);
  assign p6_sel_155192_comb = $signed(p6_smul_58300_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58300_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58300_NarrowedMult__comb[15:0]);
  assign p6_sel_155193_comb = $signed(p6_smul_58302_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58302_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58302_NarrowedMult__comb[15:0]);
  assign p6_sel_155194_comb = $signed(p6_smul_58304_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58304_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58304_NarrowedMult__comb[15:0]);
  assign p6_sel_155195_comb = $signed(p5_or_148447[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149159 ? 15'h4000 : p5_or_148447[23:9], 1'h0};
  assign p6_sel_155196_comb = p5_sgt_150019 ? 16'h7fff : {p5_bit_slice_149603, 1'h0};
  assign p6_sel_155197_comb = p5_sgt_150020 ? 16'h7fff : {p5_bit_slice_149606, 1'h0};
  assign p6_sel_155198_comb = $signed(p5_or_148454[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149162 ? 15'h4000 : p5_or_148454[23:9], 1'h0};
  assign p6_sel_155199_comb = $signed(p6_smul_58314_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58314_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58314_NarrowedMult__comb[15:0]);
  assign p6_sel_155200_comb = $signed(p6_smul_58316_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58316_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58316_NarrowedMult__comb[15:0]);
  assign p6_sel_155201_comb = $signed(p6_smul_58318_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58318_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58318_NarrowedMult__comb[15:0]);
  assign p6_sel_155202_comb = $signed(p6_smul_58320_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58320_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58320_NarrowedMult__comb[15:0]);
  assign p6_sel_155203_comb = $signed(p5_or_148457[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149163 ? 15'h4000 : p5_or_148457[23:9], 1'h0};
  assign p6_sel_155204_comb = $signed(p5_or_149164[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149164[23:9], 1'h0};
  assign p6_sel_155205_comb = $signed(p5_or_149165[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149165[23:9], 1'h0};
  assign p6_sel_155206_comb = $signed(p5_or_148464[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149166 ? 15'h4000 : p5_or_148464[23:9], 1'h0};
  assign p6_sel_155207_comb = $signed(p6_smul_58330_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58330_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58330_NarrowedMult__comb[15:0]);
  assign p6_sel_155208_comb = $signed(p6_smul_58332_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58332_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58332_NarrowedMult__comb[15:0]);
  assign p6_sel_155209_comb = $signed(p6_smul_58334_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58334_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58334_NarrowedMult__comb[15:0]);
  assign p6_sel_155210_comb = $signed(p6_smul_58336_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58336_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58336_NarrowedMult__comb[15:0]);
  assign p6_sel_155211_comb = $signed(p5_or_148467[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149167 ? 15'h4000 : p5_or_148467[23:9], 1'h0};
  assign p6_sel_155212_comb = p5_sgt_150021 ? 16'h7fff : {p5_bit_slice_149609, 1'h0};
  assign p6_sel_155213_comb = p5_sgt_150022 ? 16'h7fff : {p5_bit_slice_149612, 1'h0};
  assign p6_sel_155214_comb = $signed(p5_or_148474[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149170 ? 15'h4000 : p5_or_148474[23:9], 1'h0};
  assign p6_sel_155215_comb = $signed(p6_smul_58346_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58346_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58346_NarrowedMult__comb[15:0]);
  assign p6_sel_155216_comb = $signed(p6_smul_58348_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58348_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58348_NarrowedMult__comb[15:0]);
  assign p6_sel_155281_comb = $signed(p6_smul_58478_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58478_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58478_NarrowedMult__comb[15:0]);
  assign p6_sel_155282_comb = p5_sgt_150071 ? 16'h7fff : {p5_bit_slice_149751, 1'h0};
  assign p6_sel_155283_comb = $signed(p6_smul_58482_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58482_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58482_NarrowedMult__comb[15:0]);
  assign p6_sel_155284_comb = p5_sgt_150072 ? 16'h7fff : {p5_sel_149754, 1'h0};
  assign p6_sel_155285_comb = p5_sgt_150073 ? 16'h7fff : {p5_sel_149757, 1'h0};
  assign p6_sel_155286_comb = $signed(p6_smul_58488_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58488_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58488_NarrowedMult__comb[15:0]);
  assign p6_sel_155287_comb = p5_sgt_150074 ? 16'h7fff : {p5_bit_slice_149760, 1'h0};
  assign p6_sel_155288_comb = $signed(p6_smul_58492_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58492_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58492_NarrowedMult__comb[15:0]);
  assign p6_sel_155289_comb = $signed(p6_smul_58494_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58494_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58494_NarrowedMult__comb[15:0]);
  assign p6_sel_155290_comb = $signed(p5_or_149299[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149299[23:9], 1'h0};
  assign p6_sel_155291_comb = $signed(p6_smul_58498_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58498_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58498_NarrowedMult__comb[15:0]);
  assign p6_sel_155292_comb = p5_sgt_150075 ? 16'h7fff : {p5_sel_149763, 1'h0};
  assign p6_sel_155293_comb = p5_sgt_150076 ? 16'h7fff : {p5_sel_149766, 1'h0};
  assign p6_sel_155294_comb = $signed(p6_smul_58504_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58504_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58504_NarrowedMult__comb[15:0]);
  assign p6_sel_155295_comb = $signed(p5_or_149306[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149306[23:9], 1'h0};
  assign p6_sel_155296_comb = $signed(p6_smul_58508_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58508_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58508_NarrowedMult__comb[15:0]);
  assign p6_sel_155297_comb = $signed(p6_smul_58510_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58510_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58510_NarrowedMult__comb[15:0]);
  assign p6_sel_155298_comb = $signed(p5_or_149307[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149307[23:9], 1'h0};
  assign p6_sel_155299_comb = $signed(p6_smul_58514_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58514_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58514_NarrowedMult__comb[15:0]);
  assign p6_sel_155300_comb = $signed(p5_or_148659[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149308 ? 15'h4000 : p5_or_148659[23:9], 1'h0};
  assign p6_sel_155301_comb = $signed(p5_or_148662[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149309 ? 15'h4000 : p5_or_148662[23:9], 1'h0};
  assign p6_sel_155302_comb = $signed(p6_smul_58520_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58520_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58520_NarrowedMult__comb[15:0]);
  assign p6_sel_155303_comb = $signed(p5_or_149310[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149310[23:9], 1'h0};
  assign p6_sel_155304_comb = $signed(p6_smul_58524_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58524_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58524_NarrowedMult__comb[15:0]);
  assign p6_sel_155305_comb = $signed(p6_smul_58526_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58526_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58526_NarrowedMult__comb[15:0]);
  assign p6_sel_155306_comb = $signed(p5_or_149311[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149311[23:9], 1'h0};
  assign p6_sel_155307_comb = $signed(p6_smul_58530_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58530_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58530_NarrowedMult__comb[15:0]);
  assign p6_sel_155308_comb = p5_sgt_150077 ? 16'h7fff : {p5_sel_149769, 1'h0};
  assign p6_sel_155309_comb = p5_sgt_150078 ? 16'h7fff : {p5_sel_149772, 1'h0};
  assign p6_sel_155310_comb = $signed(p6_smul_58536_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58536_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58536_NarrowedMult__comb[15:0]);
  assign p6_sel_155311_comb = $signed(p5_or_149318[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149318[23:9], 1'h0};
  assign p6_sel_155312_comb = $signed(p6_smul_58540_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58540_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58540_NarrowedMult__comb[15:0]);
  assign p6_sel_155313_comb = $signed(p6_smul_58542_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58542_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58542_NarrowedMult__comb[15:0]);
  assign p6_sel_155314_comb = $signed(p6_smul_58546_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58546_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58546_NarrowedMult__comb[15:0]);
  assign p6_sel_155315_comb = p5_sgt_150082 ? 16'h7fff : {p5_sel_149779, 1'h0};
  assign p6_sel_155316_comb = p5_sgt_150083 ? 16'h7fff : {p5_sel_149782, 1'h0};
  assign p6_sel_155317_comb = $signed(p6_smul_58552_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58552_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58552_NarrowedMult__comb[15:0]);
  assign p6_sel_155318_comb = $signed(p6_smul_58556_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58556_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58556_NarrowedMult__comb[15:0]);
  assign p6_sel_155319_comb = $signed(p6_smul_58558_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58558_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58558_NarrowedMult__comb[15:0]);
  assign p6_sel_155320_comb = $signed(p5_or_149327[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149327[23:9], 1'h0};
  assign p6_sel_155321_comb = $signed(p6_smul_58562_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58562_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58562_NarrowedMult__comb[15:0]);
  assign p6_sel_155322_comb = p5_sgt_150087 ? 16'h7fff : {p5_sel_149789, 1'h0};
  assign p6_sel_155323_comb = p5_sgt_150088 ? 16'h7fff : {p5_sel_149792, 1'h0};
  assign p6_sel_155324_comb = $signed(p6_smul_58568_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58568_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58568_NarrowedMult__comb[15:0]);
  assign p6_sel_155325_comb = $signed(p5_or_149334[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149334[23:9], 1'h0};
  assign p6_sel_155326_comb = $signed(p6_smul_58572_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58572_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58572_NarrowedMult__comb[15:0]);
  assign p6_sel_155327_comb = $signed(p6_smul_58574_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58574_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58574_NarrowedMult__comb[15:0]);
  assign p6_sel_155328_comb = $signed(p5_or_149335[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149335[23:9], 1'h0};
  assign p6_sel_155329_comb = $signed(p6_smul_58578_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58578_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58578_NarrowedMult__comb[15:0]);
  assign p6_sel_155330_comb = $signed(p5_or_148699[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149336 ? 15'h4000 : p5_or_148699[23:9], 1'h0};
  assign p6_sel_155331_comb = $signed(p5_or_148702[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149337 ? 15'h4000 : p5_or_148702[23:9], 1'h0};
  assign p6_sel_155332_comb = $signed(p6_smul_58584_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58584_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58584_NarrowedMult__comb[15:0]);
  assign p6_sel_155333_comb = $signed(p5_or_149338[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149338[23:9], 1'h0};
  assign p6_sel_155334_comb = $signed(p6_smul_58588_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58588_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58588_NarrowedMult__comb[15:0]);
  assign p6_sel_155335_comb = $signed(p6_smul_58590_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58590_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58590_NarrowedMult__comb[15:0]);
  assign p6_sel_155336_comb = $signed(p5_or_149339[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149339[23:9], 1'h0};
  assign p6_sel_155337_comb = $signed(p6_smul_58594_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58594_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58594_NarrowedMult__comb[15:0]);
  assign p6_sel_155338_comb = p5_sgt_150089 ? 16'h7fff : {p5_sel_149795, 1'h0};
  assign p6_sel_155339_comb = p5_sgt_150090 ? 16'h7fff : {p5_sel_149798, 1'h0};
  assign p6_sel_155340_comb = $signed(p6_smul_58600_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58600_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58600_NarrowedMult__comb[15:0]);
  assign p6_sel_155341_comb = $signed(p5_or_149346[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149346[23:9], 1'h0};
  assign p6_sel_155342_comb = $signed(p6_smul_58604_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58604_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58604_NarrowedMult__comb[15:0]);
  assign p6_sel_155343_comb = $signed(p6_smul_58606_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58606_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58606_NarrowedMult__comb[15:0]);
  assign p6_sel_155344_comb = $signed(p6_smul_58608_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58608_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58608_NarrowedMult__comb[15:0]);
  assign p6_sel_155345_comb = $signed(p6_smul_58610_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58610_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58610_NarrowedMult__comb[15:0]);
  assign p6_sel_155346_comb = $signed(p6_smul_58612_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58612_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58612_NarrowedMult__comb[15:0]);
  assign p6_sel_155347_comb = $signed(p6_smul_58614_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58614_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58614_NarrowedMult__comb[15:0]);
  assign p6_sel_155348_comb = $signed(p6_smul_58616_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58616_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58616_NarrowedMult__comb[15:0]);
  assign p6_sel_155349_comb = $signed(p6_smul_58618_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58618_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58618_NarrowedMult__comb[15:0]);
  assign p6_sel_155350_comb = $signed(p6_smul_58620_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58620_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58620_NarrowedMult__comb[15:0]);
  assign p6_sel_155351_comb = $signed(p6_smul_58622_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58622_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58622_NarrowedMult__comb[15:0]);
  assign p6_sel_155352_comb = $signed(p6_smul_58624_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58624_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58624_NarrowedMult__comb[15:0]);
  assign p6_sel_155353_comb = $signed(p6_smul_58626_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58626_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58626_NarrowedMult__comb[15:0]);
  assign p6_sel_155354_comb = $signed(p6_smul_58628_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58628_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58628_NarrowedMult__comb[15:0]);
  assign p6_sel_155355_comb = $signed(p6_smul_58630_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58630_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58630_NarrowedMult__comb[15:0]);
  assign p6_sel_155356_comb = $signed(p6_smul_58632_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58632_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58632_NarrowedMult__comb[15:0]);
  assign p6_sel_155357_comb = $signed(p6_smul_58634_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58634_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58634_NarrowedMult__comb[15:0]);
  assign p6_sel_155358_comb = $signed(p6_smul_58636_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58636_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58636_NarrowedMult__comb[15:0]);
  assign p6_sel_155359_comb = $signed(p6_smul_58638_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58638_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58638_NarrowedMult__comb[15:0]);
  assign p6_sel_155360_comb = $signed(p6_smul_58640_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58640_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58640_NarrowedMult__comb[15:0]);
  assign p6_sel_155361_comb = $signed(p6_smul_58642_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58642_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58642_NarrowedMult__comb[15:0]);
  assign p6_sel_155362_comb = $signed(p6_smul_58644_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58644_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58644_NarrowedMult__comb[15:0]);
  assign p6_sel_155363_comb = $signed(p6_smul_58646_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58646_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58646_NarrowedMult__comb[15:0]);
  assign p6_sel_155364_comb = $signed(p6_smul_58648_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58648_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58648_NarrowedMult__comb[15:0]);
  assign p6_sel_155365_comb = $signed(p6_smul_58650_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58650_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58650_NarrowedMult__comb[15:0]);
  assign p6_sel_155366_comb = $signed(p6_smul_58652_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58652_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58652_NarrowedMult__comb[15:0]);
  assign p6_sel_155367_comb = $signed(p6_smul_58654_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58654_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58654_NarrowedMult__comb[15:0]);
  assign p6_sel_155368_comb = $signed(p6_smul_58656_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58656_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58656_NarrowedMult__comb[15:0]);
  assign p6_sel_155369_comb = $signed(p6_smul_58658_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58658_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58658_NarrowedMult__comb[15:0]);
  assign p6_sel_155370_comb = $signed(p6_smul_58660_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58660_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58660_NarrowedMult__comb[15:0]);
  assign p6_sel_155371_comb = $signed(p6_smul_58662_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58662_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58662_NarrowedMult__comb[15:0]);
  assign p6_sel_155372_comb = $signed(p6_smul_58664_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58664_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58664_NarrowedMult__comb[15:0]);
  assign p6_sel_155373_comb = $signed(p6_smul_58666_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58666_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58666_NarrowedMult__comb[15:0]);
  assign p6_sel_155374_comb = $signed(p6_smul_58668_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58668_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58668_NarrowedMult__comb[15:0]);
  assign p6_sel_155375_comb = $signed(p6_smul_58670_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58670_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58670_NarrowedMult__comb[15:0]);
  assign p6_sel_155376_comb = $signed(p6_smul_58672_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58672_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58672_NarrowedMult__comb[15:0]);
  assign p6_sel_155377_comb = $signed(p6_smul_58674_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58674_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58674_NarrowedMult__comb[15:0]);
  assign p6_sel_155378_comb = $signed(p6_smul_58676_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58676_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58676_NarrowedMult__comb[15:0]);
  assign p6_sel_155379_comb = $signed(p6_smul_58678_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58678_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58678_NarrowedMult__comb[15:0]);
  assign p6_sel_155380_comb = $signed(p6_smul_58680_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58680_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58680_NarrowedMult__comb[15:0]);
  assign p6_sel_155381_comb = $signed(p6_smul_58682_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58682_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58682_NarrowedMult__comb[15:0]);
  assign p6_sel_155382_comb = $signed(p6_smul_58684_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58684_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58684_NarrowedMult__comb[15:0]);
  assign p6_sel_155383_comb = $signed(p6_smul_58686_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58686_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58686_NarrowedMult__comb[15:0]);
  assign p6_sel_155384_comb = $signed(p6_smul_58688_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58688_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58688_NarrowedMult__comb[15:0]);
  assign p6_sel_155385_comb = $signed(p6_smul_58690_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58690_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58690_NarrowedMult__comb[15:0]);
  assign p6_sel_155386_comb = $signed(p6_smul_58692_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58692_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58692_NarrowedMult__comb[15:0]);
  assign p6_sel_155387_comb = $signed(p6_smul_58694_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58694_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58694_NarrowedMult__comb[15:0]);
  assign p6_sel_155388_comb = $signed(p6_smul_58696_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58696_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58696_NarrowedMult__comb[15:0]);
  assign p6_sel_155389_comb = $signed(p6_smul_58698_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58698_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58698_NarrowedMult__comb[15:0]);
  assign p6_sel_155390_comb = $signed(p6_smul_58700_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58700_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58700_NarrowedMult__comb[15:0]);
  assign p6_sel_155391_comb = $signed(p6_smul_58702_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58702_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58702_NarrowedMult__comb[15:0]);
  assign p6_sel_155392_comb = $signed(p6_smul_58704_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58704_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58704_NarrowedMult__comb[15:0]);
  assign p6_sel_155393_comb = $signed(p6_smul_58706_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58706_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58706_NarrowedMult__comb[15:0]);
  assign p6_sel_155394_comb = $signed(p6_smul_58708_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58708_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58708_NarrowedMult__comb[15:0]);
  assign p6_sel_155395_comb = $signed(p6_smul_58710_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58710_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58710_NarrowedMult__comb[15:0]);
  assign p6_sel_155396_comb = $signed(p6_smul_58712_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58712_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58712_NarrowedMult__comb[15:0]);
  assign p6_sel_155397_comb = $signed(p6_smul_58714_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58714_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58714_NarrowedMult__comb[15:0]);
  assign p6_sel_155398_comb = $signed(p6_smul_58716_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58716_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58716_NarrowedMult__comb[15:0]);
  assign p6_sel_155399_comb = $signed(p6_smul_58718_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58718_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58718_NarrowedMult__comb[15:0]);
  assign p6_sel_155400_comb = $signed(p6_smul_58720_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58720_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58720_NarrowedMult__comb[15:0]);
  assign p6_sel_155401_comb = $signed(p6_smul_58722_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58722_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58722_NarrowedMult__comb[15:0]);
  assign p6_sel_155402_comb = $signed(p6_smul_58724_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58724_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58724_NarrowedMult__comb[15:0]);
  assign p6_sel_155403_comb = $signed(p6_smul_58726_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58726_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58726_NarrowedMult__comb[15:0]);
  assign p6_sel_155404_comb = $signed(p6_smul_58728_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58728_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58728_NarrowedMult__comb[15:0]);
  assign p6_sel_155405_comb = $signed(p6_smul_58730_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58730_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58730_NarrowedMult__comb[15:0]);
  assign p6_sel_155406_comb = $signed(p6_smul_58732_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58732_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58732_NarrowedMult__comb[15:0]);
  assign p6_sel_155407_comb = p5_sgt_150091 ? 16'h7fff : {p5_sel_149801, 1'h0};
  assign p6_sel_155408_comb = $signed(p6_smul_58736_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58736_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58736_NarrowedMult__comb[15:0]);
  assign p6_sel_155409_comb = p5_sgt_150092 ? 16'h7fff : {p5_bit_slice_149804, 1'h0};
  assign p6_sel_155410_comb = $signed(p6_smul_58740_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58740_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58740_NarrowedMult__comb[15:0]);
  assign p6_sel_155411_comb = $signed(p6_smul_58742_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58742_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58742_NarrowedMult__comb[15:0]);
  assign p6_sel_155412_comb = p5_sgt_150093 ? 16'h7fff : {p5_bit_slice_149807, 1'h0};
  assign p6_sel_155413_comb = $signed(p6_smul_58746_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58746_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58746_NarrowedMult__comb[15:0]);
  assign p6_sel_155414_comb = p5_sgt_150094 ? 16'h7fff : {p5_sel_149810, 1'h0};
  assign p6_sel_155415_comb = $signed(p5_or_148727[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149355 ? 15'h4000 : p5_or_148727[23:9], 1'h0};
  assign p6_sel_155416_comb = $signed(p6_smul_58752_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58752_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58752_NarrowedMult__comb[15:0]);
  assign p6_sel_155417_comb = $signed(p5_or_149356[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149356[23:9], 1'h0};
  assign p6_sel_155418_comb = $signed(p6_smul_58756_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58756_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58756_NarrowedMult__comb[15:0]);
  assign p6_sel_155419_comb = $signed(p6_smul_58758_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58758_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58758_NarrowedMult__comb[15:0]);
  assign p6_sel_155420_comb = $signed(p5_or_149357[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149357[23:9], 1'h0};
  assign p6_sel_155421_comb = $signed(p6_smul_58762_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58762_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58762_NarrowedMult__comb[15:0]);
  assign p6_sel_155422_comb = $signed(p5_or_148734[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149358 ? 15'h4000 : p5_or_148734[23:9], 1'h0};
  assign p6_sel_155423_comb = $signed(p5_or_148737[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149359 ? 15'h4000 : p5_or_148737[23:9], 1'h0};
  assign p6_sel_155424_comb = $signed(p6_smul_58768_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58768_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58768_NarrowedMult__comb[15:0]);
  assign p6_sel_155425_comb = $signed(p5_or_149360[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149360[23:9], 1'h0};
  assign p6_sel_155426_comb = $signed(p6_smul_58772_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58772_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58772_NarrowedMult__comb[15:0]);
  assign p6_sel_155427_comb = $signed(p6_smul_58774_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58774_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58774_NarrowedMult__comb[15:0]);
  assign p6_sel_155428_comb = $signed(p5_or_149361[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149361[23:9], 1'h0};
  assign p6_sel_155429_comb = $signed(p6_smul_58778_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58778_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58778_NarrowedMult__comb[15:0]);
  assign p6_sel_155430_comb = $signed(p5_or_148744[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149362 ? 15'h4000 : p5_or_148744[23:9], 1'h0};
  assign p6_sel_155431_comb = $signed(p5_or_148747[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149363 ? 15'h4000 : p5_or_148747[23:9], 1'h0};
  assign p6_sel_155432_comb = $signed(p6_smul_58784_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58784_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58784_NarrowedMult__comb[15:0]);
  assign p6_sel_155433_comb = $signed(p5_or_149364[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149364[23:9], 1'h0};
  assign p6_sel_155434_comb = $signed(p6_smul_58788_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58788_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58788_NarrowedMult__comb[15:0]);
  assign p6_sel_155435_comb = $signed(p6_smul_58790_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58790_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58790_NarrowedMult__comb[15:0]);
  assign p6_sel_155436_comb = $signed(p5_or_149365[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149365[23:9], 1'h0};
  assign p6_sel_155437_comb = $signed(p6_smul_58794_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58794_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58794_NarrowedMult__comb[15:0]);
  assign p6_sel_155438_comb = $signed(p5_or_148754[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149366 ? 15'h4000 : p5_or_148754[23:9], 1'h0};
  assign p6_sel_155439_comb = p5_sgt_150095 ? 16'h7fff : {p5_sel_149813, 1'h0};
  assign p6_sel_155440_comb = $signed(p6_smul_58800_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58800_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58800_NarrowedMult__comb[15:0]);
  assign p6_sel_155441_comb = $signed(p6_smul_58804_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58804_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58804_NarrowedMult__comb[15:0]);
  assign p6_sel_155442_comb = $signed(p6_smul_58806_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58806_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58806_NarrowedMult__comb[15:0]);
  assign p6_sel_155443_comb = $signed(p6_smul_58810_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58810_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58810_NarrowedMult__comb[15:0]);
  assign p6_sel_155444_comb = p5_sgt_150102 ? 16'h7fff : {p5_sel_149824, 1'h0};
  assign p6_sel_155445_comb = $signed(p5_or_148767[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149375 ? 15'h4000 : p5_or_148767[23:9], 1'h0};
  assign p6_sel_155446_comb = $signed(p6_smul_58816_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58816_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58816_NarrowedMult__comb[15:0]);
  assign p6_sel_155447_comb = $signed(p5_or_149376[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149376[23:9], 1'h0};
  assign p6_sel_155448_comb = $signed(p6_smul_58820_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58820_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58820_NarrowedMult__comb[15:0]);
  assign p6_sel_155449_comb = $signed(p6_smul_58822_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58822_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58822_NarrowedMult__comb[15:0]);
  assign p6_sel_155450_comb = $signed(p5_or_149377[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149377[23:9], 1'h0};
  assign p6_sel_155451_comb = $signed(p6_smul_58826_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58826_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58826_NarrowedMult__comb[15:0]);
  assign p6_sel_155452_comb = $signed(p5_or_148774[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149378 ? 15'h4000 : p5_or_148774[23:9], 1'h0};
  assign p6_sel_155453_comb = $signed(p5_or_148777[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149379 ? 15'h4000 : p5_or_148777[23:9], 1'h0};
  assign p6_sel_155454_comb = $signed(p6_smul_58832_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58832_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58832_NarrowedMult__comb[15:0]);
  assign p6_sel_155455_comb = $signed(p5_or_149380[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149380[23:9], 1'h0};
  assign p6_sel_155456_comb = $signed(p6_smul_58836_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58836_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58836_NarrowedMult__comb[15:0]);
  assign p6_sel_155457_comb = $signed(p6_smul_58838_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58838_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58838_NarrowedMult__comb[15:0]);
  assign p6_sel_155458_comb = $signed(p5_or_149381[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149381[23:9], 1'h0};
  assign p6_sel_155459_comb = $signed(p6_smul_58842_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58842_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58842_NarrowedMult__comb[15:0]);
  assign p6_sel_155460_comb = $signed(p5_or_148784[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149382 ? 15'h4000 : p5_or_148784[23:9], 1'h0};
  assign p6_sel_155461_comb = $signed(p5_or_148787[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149383 ? 15'h4000 : p5_or_148787[23:9], 1'h0};
  assign p6_sel_155462_comb = $signed(p6_smul_58848_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58848_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58848_NarrowedMult__comb[15:0]);
  assign p6_sel_155463_comb = $signed(p5_or_149384[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149384[23:9], 1'h0};
  assign p6_sel_155464_comb = $signed(p6_smul_58852_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58852_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58852_NarrowedMult__comb[15:0]);
  assign p6_sel_155465_comb = $signed(p6_smul_58854_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58854_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58854_NarrowedMult__comb[15:0]);
  assign p6_sel_155466_comb = $signed(p5_or_149385[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149385[23:9], 1'h0};
  assign p6_sel_155467_comb = $signed(p6_smul_58858_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58858_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58858_NarrowedMult__comb[15:0]);
  assign p6_sel_155468_comb = $signed(p5_or_148794[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149386 ? 15'h4000 : p5_or_148794[23:9], 1'h0};
  assign p6_sel_155533_comb = p5_sgt_150151 ? 16'h7fff : {p5_bit_slice_149963, 1'h0};
  assign p6_sel_155534_comb = p5_sgt_150152 ? 16'h7fff : {p5_sel_149966, 1'h0};
  assign p6_sel_155535_comb = $signed(p6_smul_58994_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58994_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58994_NarrowedMult__comb[15:0]);
  assign p6_sel_155536_comb = $signed(p6_smul_58996_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58996_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58996_NarrowedMult__comb[15:0]);
  assign p6_sel_155537_comb = $signed(p6_smul_58998_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_58998_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_58998_NarrowedMult__comb[15:0]);
  assign p6_sel_155538_comb = $signed(p6_smul_59000_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59000_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59000_NarrowedMult__comb[15:0]);
  assign p6_sel_155539_comb = p5_sgt_150153 ? 16'h7fff : {p5_sel_149969, 1'h0};
  assign p6_sel_155540_comb = p5_sgt_150154 ? 16'h7fff : {p5_bit_slice_149972, 1'h0};
  assign p6_sel_155541_comb = $signed(p5_or_149515[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149515[23:9], 1'h0};
  assign p6_sel_155542_comb = $signed(p5_or_148969[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149516 ? 15'h4000 : p5_or_148969[23:9], 1'h0};
  assign p6_sel_155543_comb = $signed(p6_smul_59010_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59010_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59010_NarrowedMult__comb[15:0]);
  assign p6_sel_155544_comb = $signed(p6_smul_59012_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59012_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59012_NarrowedMult__comb[15:0]);
  assign p6_sel_155545_comb = $signed(p6_smul_59014_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59014_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59014_NarrowedMult__comb[15:0]);
  assign p6_sel_155546_comb = $signed(p6_smul_59016_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59016_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59016_NarrowedMult__comb[15:0]);
  assign p6_sel_155547_comb = $signed(p5_or_148972[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149517 ? 15'h4000 : p5_or_148972[23:9], 1'h0};
  assign p6_sel_155548_comb = $signed(p5_or_149518[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149518[23:9], 1'h0};
  assign p6_sel_155549_comb = $signed(p5_or_149519[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149519[23:9], 1'h0};
  assign p6_sel_155550_comb = $signed(p5_or_148979[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149520 ? 15'h4000 : p5_or_148979[23:9], 1'h0};
  assign p6_sel_155551_comb = $signed(p6_smul_59026_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59026_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59026_NarrowedMult__comb[15:0]);
  assign p6_sel_155552_comb = $signed(p6_smul_59028_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59028_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59028_NarrowedMult__comb[15:0]);
  assign p6_sel_155553_comb = $signed(p6_smul_59030_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59030_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59030_NarrowedMult__comb[15:0]);
  assign p6_sel_155554_comb = $signed(p6_smul_59032_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59032_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59032_NarrowedMult__comb[15:0]);
  assign p6_sel_155555_comb = $signed(p5_or_148982[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149521 ? 15'h4000 : p5_or_148982[23:9], 1'h0};
  assign p6_sel_155556_comb = $signed(p5_or_149522[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149522[23:9], 1'h0};
  assign p6_sel_155557_comb = $signed(p5_or_149523[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149523[23:9], 1'h0};
  assign p6_sel_155558_comb = $signed(p5_or_148989[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149524 ? 15'h4000 : p5_or_148989[23:9], 1'h0};
  assign p6_sel_155559_comb = $signed(p6_smul_59042_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59042_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59042_NarrowedMult__comb[15:0]);
  assign p6_sel_155560_comb = $signed(p6_smul_59044_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59044_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59044_NarrowedMult__comb[15:0]);
  assign p6_sel_155561_comb = $signed(p6_smul_59046_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59046_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59046_NarrowedMult__comb[15:0]);
  assign p6_sel_155562_comb = $signed(p6_smul_59048_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59048_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59048_NarrowedMult__comb[15:0]);
  assign p6_sel_155563_comb = $signed(p5_or_148992[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149525 ? 15'h4000 : p5_or_148992[23:9], 1'h0};
  assign p6_sel_155564_comb = $signed(p5_or_149526[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149526[23:9], 1'h0};
  assign p6_sel_155565_comb = p5_sgt_150158 ? 16'h7fff : {p5_sel_149979, 1'h0};
  assign p6_sel_155566_comb = $signed(p6_smul_59058_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59058_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59058_NarrowedMult__comb[15:0]);
  assign p6_sel_155567_comb = $signed(p6_smul_59060_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59060_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59060_NarrowedMult__comb[15:0]);
  assign p6_sel_155568_comb = $signed(p6_smul_59062_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59062_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59062_NarrowedMult__comb[15:0]);
  assign p6_sel_155569_comb = $signed(p6_smul_59064_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59064_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59064_NarrowedMult__comb[15:0]);
  assign p6_sel_155570_comb = p5_sgt_150159 ? 16'h7fff : {p5_sel_149982, 1'h0};
  assign p6_sel_155571_comb = $signed(p5_or_149535[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149535[23:9], 1'h0};
  assign p6_sel_155572_comb = $signed(p5_or_149009[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149536 ? 15'h4000 : p5_or_149009[23:9], 1'h0};
  assign p6_sel_155573_comb = $signed(p6_smul_59074_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59074_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59074_NarrowedMult__comb[15:0]);
  assign p6_sel_155574_comb = $signed(p6_smul_59076_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59076_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59076_NarrowedMult__comb[15:0]);
  assign p6_sel_155575_comb = $signed(p6_smul_59078_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59078_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59078_NarrowedMult__comb[15:0]);
  assign p6_sel_155576_comb = $signed(p6_smul_59080_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59080_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59080_NarrowedMult__comb[15:0]);
  assign p6_sel_155577_comb = $signed(p5_or_149012[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149537 ? 15'h4000 : p5_or_149012[23:9], 1'h0};
  assign p6_sel_155578_comb = $signed(p5_or_149538[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149538[23:9], 1'h0};
  assign p6_sel_155579_comb = $signed(p5_or_149539[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149539[23:9], 1'h0};
  assign p6_sel_155580_comb = $signed(p5_or_149019[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149540 ? 15'h4000 : p5_or_149019[23:9], 1'h0};
  assign p6_sel_155581_comb = $signed(p6_smul_59090_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59090_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59090_NarrowedMult__comb[15:0]);
  assign p6_sel_155582_comb = $signed(p6_smul_59092_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59092_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59092_NarrowedMult__comb[15:0]);
  assign p6_sel_155583_comb = $signed(p6_smul_59094_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59094_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59094_NarrowedMult__comb[15:0]);
  assign p6_sel_155584_comb = $signed(p6_smul_59096_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59096_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59096_NarrowedMult__comb[15:0]);
  assign p6_sel_155585_comb = $signed(p5_or_149022[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149541 ? 15'h4000 : p5_or_149022[23:9], 1'h0};
  assign p6_sel_155586_comb = $signed(p5_or_149542[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149542[23:9], 1'h0};
  assign p6_sel_155587_comb = $signed(p5_or_149543[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149543[23:9], 1'h0};
  assign p6_sel_155588_comb = $signed(p5_or_149029[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149544 ? 15'h4000 : p5_or_149029[23:9], 1'h0};
  assign p6_sel_155589_comb = $signed(p6_smul_59106_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59106_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59106_NarrowedMult__comb[15:0]);
  assign p6_sel_155590_comb = $signed(p6_smul_59108_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59108_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59108_NarrowedMult__comb[15:0]);
  assign p6_sel_155591_comb = $signed(p6_smul_59110_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59110_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59110_NarrowedMult__comb[15:0]);
  assign p6_sel_155592_comb = $signed(p6_smul_59112_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p6_smul_59112_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p6_smul_59112_NarrowedMult__comb[15:0]);
  assign p6_sel_155593_comb = $signed(p5_or_149032[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_slt_149545 ? 15'h4000 : p5_or_149032[23:9], 1'h0};
  assign p6_sel_155594_comb = $signed(p5_or_149546[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p5_or_149546[23:9], 1'h0};
  assign p6_add_156123_comb = {{1{p6_sel_155217_comb[15]}}, p6_sel_155217_comb} + {{1{p6_sel_155218_comb[15]}}, p6_sel_155218_comb};
  assign p6_add_156124_comb = {{1{p6_sel_155219_comb[15]}}, p6_sel_155219_comb} + {{1{p6_sel_155220_comb[15]}}, p6_sel_155220_comb};
  assign p6_add_156125_comb = {{1{p6_sel_155221_comb[15]}}, p6_sel_155221_comb} + {{1{p6_sel_155222_comb[15]}}, p6_sel_155222_comb};
  assign p6_add_156126_comb = {{1{p6_sel_155223_comb[15]}}, p6_sel_155223_comb} + {{1{p6_sel_155224_comb[15]}}, p6_sel_155224_comb};
  assign p6_add_156139_comb = {{1{p6_sel_155249_comb[15]}}, p6_sel_155249_comb} + {{1{p6_sel_155250_comb[15]}}, p6_sel_155250_comb};
  assign p6_add_156140_comb = {{1{p6_sel_155251_comb[15]}}, p6_sel_155251_comb} + {{1{p6_sel_155252_comb[15]}}, p6_sel_155252_comb};
  assign p6_add_156141_comb = {{1{p6_sel_155253_comb[15]}}, p6_sel_155253_comb} + {{1{p6_sel_155254_comb[15]}}, p6_sel_155254_comb};
  assign p6_add_156142_comb = {{1{p6_sel_155255_comb[15]}}, p6_sel_155255_comb} + {{1{p6_sel_155256_comb[15]}}, p6_sel_155256_comb};
  assign p6_add_156251_comb = {{1{p6_sel_155469_comb[15]}}, p6_sel_155469_comb} + {{1{p6_sel_155470_comb[15]}}, p6_sel_155470_comb};
  assign p6_add_156252_comb = {{1{p6_sel_155471_comb[15]}}, p6_sel_155471_comb} + {{1{p6_sel_155472_comb[15]}}, p6_sel_155472_comb};
  assign p6_add_156253_comb = {{1{p6_sel_155473_comb[15]}}, p6_sel_155473_comb} + {{1{p6_sel_155474_comb[15]}}, p6_sel_155474_comb};
  assign p6_add_156254_comb = {{1{p6_sel_155475_comb[15]}}, p6_sel_155475_comb} + {{1{p6_sel_155476_comb[15]}}, p6_sel_155476_comb};
  assign p6_add_156267_comb = {{1{p6_sel_155501_comb[15]}}, p6_sel_155501_comb} + {{1{p6_sel_155502_comb[15]}}, p6_sel_155502_comb};
  assign p6_add_156268_comb = {{1{p6_sel_155503_comb[15]}}, p6_sel_155503_comb} + {{1{p6_sel_155504_comb[15]}}, p6_sel_155504_comb};
  assign p6_add_156269_comb = {{1{p6_sel_155505_comb[15]}}, p6_sel_155505_comb} + {{1{p6_sel_155506_comb[15]}}, p6_sel_155506_comb};
  assign p6_add_156270_comb = {{1{p6_sel_155507_comb[15]}}, p6_sel_155507_comb} + {{1{p6_sel_155508_comb[15]}}, p6_sel_155508_comb};
  assign p6_umul_156555_comb = umul32b_32b_x_7b(p6_sum__526_comb, 7'h5b);
  assign p6_umul_156559_comb = umul32b_32b_x_7b(p6_sum__302_comb, 7'h5b);
  assign p6_sum__464_comb = {{15{p6_add_155131_comb[16]}}, p6_add_155131_comb};
  assign p6_sum__465_comb = {{15{p6_add_155132_comb[16]}}, p6_add_155132_comb};
  assign p6_sum__466_comb = {{15{p6_add_155133_comb[16]}}, p6_add_155133_comb};
  assign p6_sum__467_comb = {{15{p6_add_155134_comb[16]}}, p6_add_155134_comb};
  assign p6_sum__408_comb = {{15{p6_add_155135_comb[16]}}, p6_add_155135_comb};
  assign p6_sum__409_comb = {{15{p6_add_155136_comb[16]}}, p6_add_155136_comb};
  assign p6_sum__410_comb = {{15{p6_add_155137_comb[16]}}, p6_add_155137_comb};
  assign p6_sum__411_comb = {{15{p6_add_155138_comb[16]}}, p6_add_155138_comb};
  assign p6_sum__352_comb = {{15{p6_add_155139_comb[16]}}, p6_add_155139_comb};
  assign p6_sum__353_comb = {{15{p6_add_155140_comb[16]}}, p6_add_155140_comb};
  assign p6_sum__354_comb = {{15{p6_add_155141_comb[16]}}, p6_add_155141_comb};
  assign p6_sum__355_comb = {{15{p6_add_155142_comb[16]}}, p6_add_155142_comb};
  assign p6_sum__240_comb = {{15{p6_add_155143_comb[16]}}, p6_add_155143_comb};
  assign p6_sum__241_comb = {{15{p6_add_155144_comb[16]}}, p6_add_155144_comb};
  assign p6_sum__242_comb = {{15{p6_add_155145_comb[16]}}, p6_add_155145_comb};
  assign p6_sum__243_comb = {{15{p6_add_155146_comb[16]}}, p6_add_155146_comb};
  assign p6_sum__184_comb = {{15{p6_add_155147_comb[16]}}, p6_add_155147_comb};
  assign p6_sum__185_comb = {{15{p6_add_155148_comb[16]}}, p6_add_155148_comb};
  assign p6_sum__186_comb = {{15{p6_add_155149_comb[16]}}, p6_add_155149_comb};
  assign p6_sum__187_comb = {{15{p6_add_155150_comb[16]}}, p6_add_155150_comb};
  assign p6_sum__128_comb = {{15{p6_add_155151_comb[16]}}, p6_add_155151_comb};
  assign p6_sum__129_comb = {{15{p6_add_155152_comb[16]}}, p6_add_155152_comb};
  assign p6_sum__130_comb = {{15{p6_add_155153_comb[16]}}, p6_add_155153_comb};
  assign p6_sum__131_comb = {{15{p6_add_155154_comb[16]}}, p6_add_155154_comb};
  assign p6_add_156127_comb = {{1{p6_sel_155225_comb[15]}}, p6_sel_155225_comb} + {{1{p6_sel_155226_comb[15]}}, p6_sel_155226_comb};
  assign p6_add_156128_comb = {{1{p6_sel_155227_comb[15]}}, p6_sel_155227_comb} + {{1{p6_sel_155228_comb[15]}}, p6_sel_155228_comb};
  assign p6_add_156129_comb = {{1{p6_sel_155229_comb[15]}}, p6_sel_155229_comb} + {{1{p6_sel_155230_comb[15]}}, p6_sel_155230_comb};
  assign p6_add_156130_comb = {{1{p6_sel_155231_comb[15]}}, p6_sel_155231_comb} + {{1{p6_sel_155232_comb[15]}}, p6_sel_155232_comb};
  assign p6_add_156131_comb = {{1{p6_sel_155233_comb[15]}}, p6_sel_155233_comb} + {{1{p6_sel_155234_comb[15]}}, p6_sel_155234_comb};
  assign p6_add_156132_comb = {{1{p6_sel_155235_comb[15]}}, p6_sel_155235_comb} + {{1{p6_sel_155236_comb[15]}}, p6_sel_155236_comb};
  assign p6_add_156133_comb = {{1{p6_sel_155237_comb[15]}}, p6_sel_155237_comb} + {{1{p6_sel_155238_comb[15]}}, p6_sel_155238_comb};
  assign p6_add_156134_comb = {{1{p6_sel_155239_comb[15]}}, p6_sel_155239_comb} + {{1{p6_sel_155240_comb[15]}}, p6_sel_155240_comb};
  assign p6_add_156135_comb = {{1{p6_sel_155241_comb[15]}}, p6_sel_155241_comb} + {{1{p6_sel_155242_comb[15]}}, p6_sel_155242_comb};
  assign p6_add_156136_comb = {{1{p6_sel_155243_comb[15]}}, p6_sel_155243_comb} + {{1{p6_sel_155244_comb[15]}}, p6_sel_155244_comb};
  assign p6_add_156137_comb = {{1{p6_sel_155245_comb[15]}}, p6_sel_155245_comb} + {{1{p6_sel_155246_comb[15]}}, p6_sel_155246_comb};
  assign p6_add_156138_comb = {{1{p6_sel_155247_comb[15]}}, p6_sel_155247_comb} + {{1{p6_sel_155248_comb[15]}}, p6_sel_155248_comb};
  assign p6_add_156143_comb = {{1{p6_sel_155257_comb[15]}}, p6_sel_155257_comb} + {{1{p6_sel_155258_comb[15]}}, p6_sel_155258_comb};
  assign p6_add_156144_comb = {{1{p6_sel_155259_comb[15]}}, p6_sel_155259_comb} + {{1{p6_sel_155260_comb[15]}}, p6_sel_155260_comb};
  assign p6_add_156145_comb = {{1{p6_sel_155261_comb[15]}}, p6_sel_155261_comb} + {{1{p6_sel_155262_comb[15]}}, p6_sel_155262_comb};
  assign p6_add_156146_comb = {{1{p6_sel_155263_comb[15]}}, p6_sel_155263_comb} + {{1{p6_sel_155264_comb[15]}}, p6_sel_155264_comb};
  assign p6_add_156147_comb = {{1{p6_sel_155265_comb[15]}}, p6_sel_155265_comb} + {{1{p6_sel_155266_comb[15]}}, p6_sel_155266_comb};
  assign p6_add_156148_comb = {{1{p6_sel_155267_comb[15]}}, p6_sel_155267_comb} + {{1{p6_sel_155268_comb[15]}}, p6_sel_155268_comb};
  assign p6_add_156149_comb = {{1{p6_sel_155269_comb[15]}}, p6_sel_155269_comb} + {{1{p6_sel_155270_comb[15]}}, p6_sel_155270_comb};
  assign p6_add_156150_comb = {{1{p6_sel_155271_comb[15]}}, p6_sel_155271_comb} + {{1{p6_sel_155272_comb[15]}}, p6_sel_155272_comb};
  assign p6_add_156151_comb = {{1{p6_sel_155273_comb[15]}}, p6_sel_155273_comb} + {{1{p6_sel_155274_comb[15]}}, p6_sel_155274_comb};
  assign p6_add_156152_comb = {{1{p6_sel_155275_comb[15]}}, p6_sel_155275_comb} + {{1{p6_sel_155276_comb[15]}}, p6_sel_155276_comb};
  assign p6_add_156153_comb = {{1{p6_sel_155277_comb[15]}}, p6_sel_155277_comb} + {{1{p6_sel_155278_comb[15]}}, p6_sel_155278_comb};
  assign p6_add_156154_comb = {{1{p6_sel_155279_comb[15]}}, p6_sel_155279_comb} + {{1{p6_sel_155280_comb[15]}}, p6_sel_155280_comb};
  assign p6_add_156255_comb = {{1{p6_sel_155477_comb[15]}}, p6_sel_155477_comb} + {{1{p6_sel_155478_comb[15]}}, p6_sel_155478_comb};
  assign p6_add_156256_comb = {{1{p6_sel_155479_comb[15]}}, p6_sel_155479_comb} + {{1{p6_sel_155480_comb[15]}}, p6_sel_155480_comb};
  assign p6_add_156257_comb = {{1{p6_sel_155481_comb[15]}}, p6_sel_155481_comb} + {{1{p6_sel_155482_comb[15]}}, p6_sel_155482_comb};
  assign p6_add_156258_comb = {{1{p6_sel_155483_comb[15]}}, p6_sel_155483_comb} + {{1{p6_sel_155484_comb[15]}}, p6_sel_155484_comb};
  assign p6_add_156259_comb = {{1{p6_sel_155485_comb[15]}}, p6_sel_155485_comb} + {{1{p6_sel_155486_comb[15]}}, p6_sel_155486_comb};
  assign p6_add_156260_comb = {{1{p6_sel_155487_comb[15]}}, p6_sel_155487_comb} + {{1{p6_sel_155488_comb[15]}}, p6_sel_155488_comb};
  assign p6_add_156261_comb = {{1{p6_sel_155489_comb[15]}}, p6_sel_155489_comb} + {{1{p6_sel_155490_comb[15]}}, p6_sel_155490_comb};
  assign p6_add_156262_comb = {{1{p6_sel_155491_comb[15]}}, p6_sel_155491_comb} + {{1{p6_sel_155492_comb[15]}}, p6_sel_155492_comb};
  assign p6_add_156263_comb = {{1{p6_sel_155493_comb[15]}}, p6_sel_155493_comb} + {{1{p6_sel_155494_comb[15]}}, p6_sel_155494_comb};
  assign p6_add_156264_comb = {{1{p6_sel_155495_comb[15]}}, p6_sel_155495_comb} + {{1{p6_sel_155496_comb[15]}}, p6_sel_155496_comb};
  assign p6_add_156265_comb = {{1{p6_sel_155497_comb[15]}}, p6_sel_155497_comb} + {{1{p6_sel_155498_comb[15]}}, p6_sel_155498_comb};
  assign p6_add_156266_comb = {{1{p6_sel_155499_comb[15]}}, p6_sel_155499_comb} + {{1{p6_sel_155500_comb[15]}}, p6_sel_155500_comb};
  assign p6_add_156271_comb = {{1{p6_sel_155509_comb[15]}}, p6_sel_155509_comb} + {{1{p6_sel_155510_comb[15]}}, p6_sel_155510_comb};
  assign p6_add_156272_comb = {{1{p6_sel_155511_comb[15]}}, p6_sel_155511_comb} + {{1{p6_sel_155512_comb[15]}}, p6_sel_155512_comb};
  assign p6_add_156273_comb = {{1{p6_sel_155513_comb[15]}}, p6_sel_155513_comb} + {{1{p6_sel_155514_comb[15]}}, p6_sel_155514_comb};
  assign p6_add_156274_comb = {{1{p6_sel_155515_comb[15]}}, p6_sel_155515_comb} + {{1{p6_sel_155516_comb[15]}}, p6_sel_155516_comb};
  assign p6_add_156275_comb = {{1{p6_sel_155517_comb[15]}}, p6_sel_155517_comb} + {{1{p6_sel_155518_comb[15]}}, p6_sel_155518_comb};
  assign p6_add_156276_comb = {{1{p6_sel_155519_comb[15]}}, p6_sel_155519_comb} + {{1{p6_sel_155520_comb[15]}}, p6_sel_155520_comb};
  assign p6_add_156277_comb = {{1{p6_sel_155521_comb[15]}}, p6_sel_155521_comb} + {{1{p6_sel_155522_comb[15]}}, p6_sel_155522_comb};
  assign p6_add_156278_comb = {{1{p6_sel_155523_comb[15]}}, p6_sel_155523_comb} + {{1{p6_sel_155524_comb[15]}}, p6_sel_155524_comb};
  assign p6_add_156279_comb = {{1{p6_sel_155525_comb[15]}}, p6_sel_155525_comb} + {{1{p6_sel_155526_comb[15]}}, p6_sel_155526_comb};
  assign p6_add_156280_comb = {{1{p6_sel_155527_comb[15]}}, p6_sel_155527_comb} + {{1{p6_sel_155528_comb[15]}}, p6_sel_155528_comb};
  assign p6_add_156281_comb = {{1{p6_sel_155529_comb[15]}}, p6_sel_155529_comb} + {{1{p6_sel_155530_comb[15]}}, p6_sel_155530_comb};
  assign p6_add_156282_comb = {{1{p6_sel_155531_comb[15]}}, p6_sel_155531_comb} + {{1{p6_sel_155532_comb[15]}}, p6_sel_155532_comb};
  assign p6_sum__1576_comb = {{8{p6_add_156123_comb[16]}}, p6_add_156123_comb};
  assign p6_sum__1577_comb = {{8{p6_add_156124_comb[16]}}, p6_add_156124_comb};
  assign p6_sum__1578_comb = {{8{p6_add_156125_comb[16]}}, p6_add_156125_comb};
  assign p6_sum__1579_comb = {{8{p6_add_156126_comb[16]}}, p6_add_156126_comb};
  assign p6_sum__1464_comb = {{8{p6_add_156139_comb[16]}}, p6_add_156139_comb};
  assign p6_sum__1465_comb = {{8{p6_add_156140_comb[16]}}, p6_add_156140_comb};
  assign p6_sum__1466_comb = {{8{p6_add_156141_comb[16]}}, p6_add_156141_comb};
  assign p6_sum__1467_comb = {{8{p6_add_156142_comb[16]}}, p6_add_156142_comb};
  assign p6_sum__1560_comb = {{8{p6_add_156251_comb[16]}}, p6_add_156251_comb};
  assign p6_sum__1561_comb = {{8{p6_add_156252_comb[16]}}, p6_add_156252_comb};
  assign p6_sum__1562_comb = {{8{p6_add_156253_comb[16]}}, p6_add_156253_comb};
  assign p6_sum__1563_comb = {{8{p6_add_156254_comb[16]}}, p6_add_156254_comb};
  assign p6_sum__1448_comb = {{8{p6_add_156267_comb[16]}}, p6_add_156267_comb};
  assign p6_sum__1449_comb = {{8{p6_add_156268_comb[16]}}, p6_add_156268_comb};
  assign p6_sum__1450_comb = {{8{p6_add_156269_comb[16]}}, p6_add_156269_comb};
  assign p6_sum__1451_comb = {{8{p6_add_156270_comb[16]}}, p6_add_156270_comb};
  assign p6_sum__468_comb = p6_sum__464_comb + p6_sum__465_comb;
  assign p6_sum__469_comb = p6_sum__466_comb + p6_sum__467_comb;
  assign p6_sum__412_comb = p6_sum__408_comb + p6_sum__409_comb;
  assign p6_sum__413_comb = p6_sum__410_comb + p6_sum__411_comb;
  assign p6_sum__356_comb = p6_sum__352_comb + p6_sum__353_comb;
  assign p6_sum__357_comb = p6_sum__354_comb + p6_sum__355_comb;
  assign p6_sum__244_comb = p6_sum__240_comb + p6_sum__241_comb;
  assign p6_sum__245_comb = p6_sum__242_comb + p6_sum__243_comb;
  assign p6_sum__188_comb = p6_sum__184_comb + p6_sum__185_comb;
  assign p6_sum__189_comb = p6_sum__186_comb + p6_sum__187_comb;
  assign p6_sum__132_comb = p6_sum__128_comb + p6_sum__129_comb;
  assign p6_sum__133_comb = p6_sum__130_comb + p6_sum__131_comb;
  assign p6_add_156091_comb = {{1{p6_sel_155155_comb[15]}}, p6_sel_155155_comb} + {{1{p6_sel_155156_comb[15]}}, p6_sel_155156_comb};
  assign p6_add_156092_comb = {{1{p6_sel_155157_comb[15]}}, p6_sel_155157_comb} + {{1{p6_sel_155158_comb[15]}}, p6_sel_155158_comb};
  assign p6_add_156093_comb = {{1{p6_sel_155159_comb[15]}}, p6_sel_155159_comb} + {{1{p6_sel_155160_comb[15]}}, p6_sel_155160_comb};
  assign p6_add_156094_comb = {{1{p6_sel_155161_comb[15]}}, p6_sel_155161_comb} + {{1{p6_sel_155162_comb[15]}}, p6_sel_155162_comb};
  assign p6_add_156095_comb = {{1{p6_sel_155163_comb[15]}}, p6_sel_155163_comb} + {{1{p6_sel_155164_comb[15]}}, p6_sel_155164_comb};
  assign p6_add_156096_comb = {{1{p6_sel_155165_comb[15]}}, p6_sel_155165_comb} + {{1{p6_sel_155166_comb[15]}}, p6_sel_155166_comb};
  assign p6_add_156097_comb = {{1{p6_sel_155167_comb[15]}}, p6_sel_155167_comb} + {{1{p6_sel_155168_comb[15]}}, p6_sel_155168_comb};
  assign p6_add_156098_comb = {{1{p6_sel_155169_comb[15]}}, p6_sel_155169_comb} + {{1{p6_sel_155170_comb[15]}}, p6_sel_155170_comb};
  assign p6_add_156099_comb = {{1{p6_sel_155171_comb[15]}}, p6_sel_155171_comb} + {{1{p6_sel_155172_comb[15]}}, p6_sel_155172_comb};
  assign p6_add_156100_comb = {{1{p6_sel_155173_comb[15]}}, p6_sel_155173_comb} + {{1{p6_sel_155174_comb[15]}}, p6_sel_155174_comb};
  assign p6_add_156101_comb = {{1{p6_sel_155175_comb[15]}}, p6_sel_155175_comb} + {{1{p6_sel_155176_comb[15]}}, p6_sel_155176_comb};
  assign p6_add_156102_comb = {{1{p6_sel_155177_comb[15]}}, p6_sel_155177_comb} + {{1{p6_sel_155178_comb[15]}}, p6_sel_155178_comb};
  assign p6_add_156103_comb = {{1{p6_sel_155179_comb[15]}}, p6_sel_155179_comb} + {{1{p6_sel_155180_comb[15]}}, p6_sel_155180_comb};
  assign p6_add_156104_comb = {{1{p6_sel_155181_comb[15]}}, p6_sel_155181_comb} + {{1{p6_sel_155182_comb[15]}}, p6_sel_155182_comb};
  assign p6_add_156105_comb = {{1{p6_sel_155183_comb[15]}}, p6_sel_155183_comb} + {{1{p6_sel_155184_comb[15]}}, p6_sel_155184_comb};
  assign p6_add_156106_comb = {{1{p6_sel_155185_comb[15]}}, p6_sel_155185_comb} + {{1{p6_sel_155186_comb[15]}}, p6_sel_155186_comb};
  assign p6_add_156107_comb = {{1{p6_sel_155187_comb[15]}}, p6_sel_155187_comb} + {{1{p6_sel_155188_comb[15]}}, p6_sel_155188_comb};
  assign p6_add_156108_comb = {{1{p6_sel_155189_comb[15]}}, p6_sel_155189_comb} + {{1{p5_sel_150171[15]}}, p5_sel_150171};
  assign p6_add_156109_comb = {{1{p5_sel_150172[15]}}, p5_sel_150172} + {{1{p6_sel_155190_comb[15]}}, p6_sel_155190_comb};
  assign p6_add_156110_comb = {{1{p6_sel_155191_comb[15]}}, p6_sel_155191_comb} + {{1{p6_sel_155192_comb[15]}}, p6_sel_155192_comb};
  assign p6_add_156111_comb = {{1{p6_sel_155193_comb[15]}}, p6_sel_155193_comb} + {{1{p6_sel_155194_comb[15]}}, p6_sel_155194_comb};
  assign p6_add_156112_comb = {{1{p6_sel_155195_comb[15]}}, p6_sel_155195_comb} + {{1{p6_sel_155196_comb[15]}}, p6_sel_155196_comb};
  assign p6_add_156113_comb = {{1{p6_sel_155197_comb[15]}}, p6_sel_155197_comb} + {{1{p6_sel_155198_comb[15]}}, p6_sel_155198_comb};
  assign p6_add_156114_comb = {{1{p6_sel_155199_comb[15]}}, p6_sel_155199_comb} + {{1{p6_sel_155200_comb[15]}}, p6_sel_155200_comb};
  assign p6_add_156115_comb = {{1{p6_sel_155201_comb[15]}}, p6_sel_155201_comb} + {{1{p6_sel_155202_comb[15]}}, p6_sel_155202_comb};
  assign p6_add_156116_comb = {{1{p6_sel_155203_comb[15]}}, p6_sel_155203_comb} + {{1{p6_sel_155204_comb[15]}}, p6_sel_155204_comb};
  assign p6_add_156117_comb = {{1{p6_sel_155205_comb[15]}}, p6_sel_155205_comb} + {{1{p6_sel_155206_comb[15]}}, p6_sel_155206_comb};
  assign p6_add_156118_comb = {{1{p6_sel_155207_comb[15]}}, p6_sel_155207_comb} + {{1{p6_sel_155208_comb[15]}}, p6_sel_155208_comb};
  assign p6_add_156119_comb = {{1{p6_sel_155209_comb[15]}}, p6_sel_155209_comb} + {{1{p6_sel_155210_comb[15]}}, p6_sel_155210_comb};
  assign p6_add_156120_comb = {{1{p6_sel_155211_comb[15]}}, p6_sel_155211_comb} + {{1{p6_sel_155212_comb[15]}}, p6_sel_155212_comb};
  assign p6_add_156121_comb = {{1{p6_sel_155213_comb[15]}}, p6_sel_155213_comb} + {{1{p6_sel_155214_comb[15]}}, p6_sel_155214_comb};
  assign p6_add_156122_comb = {{1{p6_sel_155215_comb[15]}}, p6_sel_155215_comb} + {{1{p6_sel_155216_comb[15]}}, p6_sel_155216_comb};
  assign p6_add_156155_comb = {{1{p6_sel_155281_comb[15]}}, p6_sel_155281_comb} + {{1{p6_sel_155282_comb[15]}}, p6_sel_155282_comb};
  assign p6_add_156156_comb = {{1{p6_sel_155283_comb[15]}}, p6_sel_155283_comb} + {{1{p6_sel_155284_comb[15]}}, p6_sel_155284_comb};
  assign p6_add_156157_comb = {{1{p6_sel_155285_comb[15]}}, p6_sel_155285_comb} + {{1{p6_sel_155286_comb[15]}}, p6_sel_155286_comb};
  assign p6_add_156158_comb = {{1{p6_sel_155287_comb[15]}}, p6_sel_155287_comb} + {{1{p6_sel_155288_comb[15]}}, p6_sel_155288_comb};
  assign p6_add_156159_comb = {{1{p6_sel_155289_comb[15]}}, p6_sel_155289_comb} + {{1{p6_sel_155290_comb[15]}}, p6_sel_155290_comb};
  assign p6_add_156160_comb = {{1{p6_sel_155291_comb[15]}}, p6_sel_155291_comb} + {{1{p6_sel_155292_comb[15]}}, p6_sel_155292_comb};
  assign p6_add_156161_comb = {{1{p6_sel_155293_comb[15]}}, p6_sel_155293_comb} + {{1{p6_sel_155294_comb[15]}}, p6_sel_155294_comb};
  assign p6_add_156162_comb = {{1{p6_sel_155295_comb[15]}}, p6_sel_155295_comb} + {{1{p6_sel_155296_comb[15]}}, p6_sel_155296_comb};
  assign p6_add_156163_comb = {{1{p6_sel_155297_comb[15]}}, p6_sel_155297_comb} + {{1{p6_sel_155298_comb[15]}}, p6_sel_155298_comb};
  assign p6_add_156164_comb = {{1{p6_sel_155299_comb[15]}}, p6_sel_155299_comb} + {{1{p6_sel_155300_comb[15]}}, p6_sel_155300_comb};
  assign p6_add_156165_comb = {{1{p6_sel_155301_comb[15]}}, p6_sel_155301_comb} + {{1{p6_sel_155302_comb[15]}}, p6_sel_155302_comb};
  assign p6_add_156166_comb = {{1{p6_sel_155303_comb[15]}}, p6_sel_155303_comb} + {{1{p6_sel_155304_comb[15]}}, p6_sel_155304_comb};
  assign p6_add_156167_comb = {{1{p6_sel_155305_comb[15]}}, p6_sel_155305_comb} + {{1{p6_sel_155306_comb[15]}}, p6_sel_155306_comb};
  assign p6_add_156168_comb = {{1{p6_sel_155307_comb[15]}}, p6_sel_155307_comb} + {{1{p6_sel_155308_comb[15]}}, p6_sel_155308_comb};
  assign p6_add_156169_comb = {{1{p6_sel_155309_comb[15]}}, p6_sel_155309_comb} + {{1{p6_sel_155310_comb[15]}}, p6_sel_155310_comb};
  assign p6_add_156170_comb = {{1{p6_sel_155311_comb[15]}}, p6_sel_155311_comb} + {{1{p6_sel_155312_comb[15]}}, p6_sel_155312_comb};
  assign p6_add_156171_comb = {{1{p6_sel_155313_comb[15]}}, p6_sel_155313_comb} + {{1{p5_sel_150173[15]}}, p5_sel_150173};
  assign p6_add_156172_comb = {{1{p6_sel_155314_comb[15]}}, p6_sel_155314_comb} + {{1{p6_sel_155315_comb[15]}}, p6_sel_155315_comb};
  assign p6_add_156173_comb = {{1{p6_sel_155316_comb[15]}}, p6_sel_155316_comb} + {{1{p6_sel_155317_comb[15]}}, p6_sel_155317_comb};
  assign p6_add_156174_comb = {{1{p5_sel_150174[15]}}, p5_sel_150174} + {{1{p6_sel_155318_comb[15]}}, p6_sel_155318_comb};
  assign p6_add_156175_comb = {{1{p6_sel_155319_comb[15]}}, p6_sel_155319_comb} + {{1{p6_sel_155320_comb[15]}}, p6_sel_155320_comb};
  assign p6_add_156176_comb = {{1{p6_sel_155321_comb[15]}}, p6_sel_155321_comb} + {{1{p6_sel_155322_comb[15]}}, p6_sel_155322_comb};
  assign p6_add_156177_comb = {{1{p6_sel_155323_comb[15]}}, p6_sel_155323_comb} + {{1{p6_sel_155324_comb[15]}}, p6_sel_155324_comb};
  assign p6_add_156178_comb = {{1{p6_sel_155325_comb[15]}}, p6_sel_155325_comb} + {{1{p6_sel_155326_comb[15]}}, p6_sel_155326_comb};
  assign p6_add_156179_comb = {{1{p6_sel_155327_comb[15]}}, p6_sel_155327_comb} + {{1{p6_sel_155328_comb[15]}}, p6_sel_155328_comb};
  assign p6_add_156180_comb = {{1{p6_sel_155329_comb[15]}}, p6_sel_155329_comb} + {{1{p6_sel_155330_comb[15]}}, p6_sel_155330_comb};
  assign p6_add_156181_comb = {{1{p6_sel_155331_comb[15]}}, p6_sel_155331_comb} + {{1{p6_sel_155332_comb[15]}}, p6_sel_155332_comb};
  assign p6_add_156182_comb = {{1{p6_sel_155333_comb[15]}}, p6_sel_155333_comb} + {{1{p6_sel_155334_comb[15]}}, p6_sel_155334_comb};
  assign p6_add_156183_comb = {{1{p6_sel_155335_comb[15]}}, p6_sel_155335_comb} + {{1{p6_sel_155336_comb[15]}}, p6_sel_155336_comb};
  assign p6_add_156184_comb = {{1{p6_sel_155337_comb[15]}}, p6_sel_155337_comb} + {{1{p6_sel_155338_comb[15]}}, p6_sel_155338_comb};
  assign p6_add_156185_comb = {{1{p6_sel_155339_comb[15]}}, p6_sel_155339_comb} + {{1{p6_sel_155340_comb[15]}}, p6_sel_155340_comb};
  assign p6_add_156186_comb = {{1{p6_sel_155341_comb[15]}}, p6_sel_155341_comb} + {{1{p6_sel_155342_comb[15]}}, p6_sel_155342_comb};
  assign p6_add_156187_comb = {{1{p6_sel_155343_comb[15]}}, p6_sel_155343_comb} + {{1{p6_sel_155344_comb[15]}}, p6_sel_155344_comb};
  assign p6_add_156188_comb = {{1{p6_sel_155345_comb[15]}}, p6_sel_155345_comb} + {{1{p6_sel_155346_comb[15]}}, p6_sel_155346_comb};
  assign p6_add_156189_comb = {{1{p6_sel_155347_comb[15]}}, p6_sel_155347_comb} + {{1{p6_sel_155348_comb[15]}}, p6_sel_155348_comb};
  assign p6_add_156190_comb = {{1{p6_sel_155349_comb[15]}}, p6_sel_155349_comb} + {{1{p6_sel_155350_comb[15]}}, p6_sel_155350_comb};
  assign p6_add_156191_comb = {{1{p6_sel_155351_comb[15]}}, p6_sel_155351_comb} + {{1{p6_sel_155352_comb[15]}}, p6_sel_155352_comb};
  assign p6_add_156192_comb = {{1{p6_sel_155353_comb[15]}}, p6_sel_155353_comb} + {{1{p6_sel_155354_comb[15]}}, p6_sel_155354_comb};
  assign p6_add_156193_comb = {{1{p6_sel_155355_comb[15]}}, p6_sel_155355_comb} + {{1{p6_sel_155356_comb[15]}}, p6_sel_155356_comb};
  assign p6_add_156194_comb = {{1{p6_sel_155357_comb[15]}}, p6_sel_155357_comb} + {{1{p6_sel_155358_comb[15]}}, p6_sel_155358_comb};
  assign p6_add_156195_comb = {{1{p6_sel_155359_comb[15]}}, p6_sel_155359_comb} + {{1{p6_sel_155360_comb[15]}}, p6_sel_155360_comb};
  assign p6_add_156196_comb = {{1{p6_sel_155361_comb[15]}}, p6_sel_155361_comb} + {{1{p6_sel_155362_comb[15]}}, p6_sel_155362_comb};
  assign p6_add_156197_comb = {{1{p6_sel_155363_comb[15]}}, p6_sel_155363_comb} + {{1{p6_sel_155364_comb[15]}}, p6_sel_155364_comb};
  assign p6_add_156198_comb = {{1{p6_sel_155365_comb[15]}}, p6_sel_155365_comb} + {{1{p6_sel_155366_comb[15]}}, p6_sel_155366_comb};
  assign p6_add_156199_comb = {{1{p6_sel_155367_comb[15]}}, p6_sel_155367_comb} + {{1{p6_sel_155368_comb[15]}}, p6_sel_155368_comb};
  assign p6_add_156200_comb = {{1{p6_sel_155369_comb[15]}}, p6_sel_155369_comb} + {{1{p6_sel_155370_comb[15]}}, p6_sel_155370_comb};
  assign p6_add_156201_comb = {{1{p6_sel_155371_comb[15]}}, p6_sel_155371_comb} + {{1{p6_sel_155372_comb[15]}}, p6_sel_155372_comb};
  assign p6_add_156202_comb = {{1{p6_sel_155373_comb[15]}}, p6_sel_155373_comb} + {{1{p6_sel_155374_comb[15]}}, p6_sel_155374_comb};
  assign p6_add_156203_comb = {{1{p6_sel_155375_comb[15]}}, p6_sel_155375_comb} + {{1{p6_sel_155376_comb[15]}}, p6_sel_155376_comb};
  assign p6_add_156204_comb = {{1{p6_sel_155377_comb[15]}}, p6_sel_155377_comb} + {{1{p6_sel_155378_comb[15]}}, p6_sel_155378_comb};
  assign p6_add_156205_comb = {{1{p6_sel_155379_comb[15]}}, p6_sel_155379_comb} + {{1{p6_sel_155380_comb[15]}}, p6_sel_155380_comb};
  assign p6_add_156206_comb = {{1{p6_sel_155381_comb[15]}}, p6_sel_155381_comb} + {{1{p6_sel_155382_comb[15]}}, p6_sel_155382_comb};
  assign p6_add_156207_comb = {{1{p6_sel_155383_comb[15]}}, p6_sel_155383_comb} + {{1{p6_sel_155384_comb[15]}}, p6_sel_155384_comb};
  assign p6_add_156208_comb = {{1{p6_sel_155385_comb[15]}}, p6_sel_155385_comb} + {{1{p6_sel_155386_comb[15]}}, p6_sel_155386_comb};
  assign p6_add_156209_comb = {{1{p6_sel_155387_comb[15]}}, p6_sel_155387_comb} + {{1{p6_sel_155388_comb[15]}}, p6_sel_155388_comb};
  assign p6_add_156210_comb = {{1{p6_sel_155389_comb[15]}}, p6_sel_155389_comb} + {{1{p6_sel_155390_comb[15]}}, p6_sel_155390_comb};
  assign p6_add_156211_comb = {{1{p6_sel_155391_comb[15]}}, p6_sel_155391_comb} + {{1{p6_sel_155392_comb[15]}}, p6_sel_155392_comb};
  assign p6_add_156212_comb = {{1{p6_sel_155393_comb[15]}}, p6_sel_155393_comb} + {{1{p6_sel_155394_comb[15]}}, p6_sel_155394_comb};
  assign p6_add_156213_comb = {{1{p6_sel_155395_comb[15]}}, p6_sel_155395_comb} + {{1{p6_sel_155396_comb[15]}}, p6_sel_155396_comb};
  assign p6_add_156214_comb = {{1{p6_sel_155397_comb[15]}}, p6_sel_155397_comb} + {{1{p6_sel_155398_comb[15]}}, p6_sel_155398_comb};
  assign p6_add_156215_comb = {{1{p6_sel_155399_comb[15]}}, p6_sel_155399_comb} + {{1{p6_sel_155400_comb[15]}}, p6_sel_155400_comb};
  assign p6_add_156216_comb = {{1{p6_sel_155401_comb[15]}}, p6_sel_155401_comb} + {{1{p6_sel_155402_comb[15]}}, p6_sel_155402_comb};
  assign p6_add_156217_comb = {{1{p6_sel_155403_comb[15]}}, p6_sel_155403_comb} + {{1{p6_sel_155404_comb[15]}}, p6_sel_155404_comb};
  assign p6_add_156218_comb = {{1{p6_sel_155405_comb[15]}}, p6_sel_155405_comb} + {{1{p6_sel_155406_comb[15]}}, p6_sel_155406_comb};
  assign p6_add_156219_comb = {{1{p6_sel_155407_comb[15]}}, p6_sel_155407_comb} + {{1{p6_sel_155408_comb[15]}}, p6_sel_155408_comb};
  assign p6_add_156220_comb = {{1{p6_sel_155409_comb[15]}}, p6_sel_155409_comb} + {{1{p6_sel_155410_comb[15]}}, p6_sel_155410_comb};
  assign p6_add_156221_comb = {{1{p6_sel_155411_comb[15]}}, p6_sel_155411_comb} + {{1{p6_sel_155412_comb[15]}}, p6_sel_155412_comb};
  assign p6_add_156222_comb = {{1{p6_sel_155413_comb[15]}}, p6_sel_155413_comb} + {{1{p6_sel_155414_comb[15]}}, p6_sel_155414_comb};
  assign p6_add_156223_comb = {{1{p6_sel_155415_comb[15]}}, p6_sel_155415_comb} + {{1{p6_sel_155416_comb[15]}}, p6_sel_155416_comb};
  assign p6_add_156224_comb = {{1{p6_sel_155417_comb[15]}}, p6_sel_155417_comb} + {{1{p6_sel_155418_comb[15]}}, p6_sel_155418_comb};
  assign p6_add_156225_comb = {{1{p6_sel_155419_comb[15]}}, p6_sel_155419_comb} + {{1{p6_sel_155420_comb[15]}}, p6_sel_155420_comb};
  assign p6_add_156226_comb = {{1{p6_sel_155421_comb[15]}}, p6_sel_155421_comb} + {{1{p6_sel_155422_comb[15]}}, p6_sel_155422_comb};
  assign p6_add_156227_comb = {{1{p6_sel_155423_comb[15]}}, p6_sel_155423_comb} + {{1{p6_sel_155424_comb[15]}}, p6_sel_155424_comb};
  assign p6_add_156228_comb = {{1{p6_sel_155425_comb[15]}}, p6_sel_155425_comb} + {{1{p6_sel_155426_comb[15]}}, p6_sel_155426_comb};
  assign p6_add_156229_comb = {{1{p6_sel_155427_comb[15]}}, p6_sel_155427_comb} + {{1{p6_sel_155428_comb[15]}}, p6_sel_155428_comb};
  assign p6_add_156230_comb = {{1{p6_sel_155429_comb[15]}}, p6_sel_155429_comb} + {{1{p6_sel_155430_comb[15]}}, p6_sel_155430_comb};
  assign p6_add_156231_comb = {{1{p6_sel_155431_comb[15]}}, p6_sel_155431_comb} + {{1{p6_sel_155432_comb[15]}}, p6_sel_155432_comb};
  assign p6_add_156232_comb = {{1{p6_sel_155433_comb[15]}}, p6_sel_155433_comb} + {{1{p6_sel_155434_comb[15]}}, p6_sel_155434_comb};
  assign p6_add_156233_comb = {{1{p6_sel_155435_comb[15]}}, p6_sel_155435_comb} + {{1{p6_sel_155436_comb[15]}}, p6_sel_155436_comb};
  assign p6_add_156234_comb = {{1{p6_sel_155437_comb[15]}}, p6_sel_155437_comb} + {{1{p6_sel_155438_comb[15]}}, p6_sel_155438_comb};
  assign p6_add_156235_comb = {{1{p6_sel_155439_comb[15]}}, p6_sel_155439_comb} + {{1{p6_sel_155440_comb[15]}}, p6_sel_155440_comb};
  assign p6_add_156236_comb = {{1{p5_sel_150175[15]}}, p5_sel_150175} + {{1{p6_sel_155441_comb[15]}}, p6_sel_155441_comb};
  assign p6_add_156237_comb = {{1{p6_sel_155442_comb[15]}}, p6_sel_155442_comb} + {{1{p5_sel_150176[15]}}, p5_sel_150176};
  assign p6_add_156238_comb = {{1{p6_sel_155443_comb[15]}}, p6_sel_155443_comb} + {{1{p6_sel_155444_comb[15]}}, p6_sel_155444_comb};
  assign p6_add_156239_comb = {{1{p6_sel_155445_comb[15]}}, p6_sel_155445_comb} + {{1{p6_sel_155446_comb[15]}}, p6_sel_155446_comb};
  assign p6_add_156240_comb = {{1{p6_sel_155447_comb[15]}}, p6_sel_155447_comb} + {{1{p6_sel_155448_comb[15]}}, p6_sel_155448_comb};
  assign p6_add_156241_comb = {{1{p6_sel_155449_comb[15]}}, p6_sel_155449_comb} + {{1{p6_sel_155450_comb[15]}}, p6_sel_155450_comb};
  assign p6_add_156242_comb = {{1{p6_sel_155451_comb[15]}}, p6_sel_155451_comb} + {{1{p6_sel_155452_comb[15]}}, p6_sel_155452_comb};
  assign p6_add_156243_comb = {{1{p6_sel_155453_comb[15]}}, p6_sel_155453_comb} + {{1{p6_sel_155454_comb[15]}}, p6_sel_155454_comb};
  assign p6_add_156244_comb = {{1{p6_sel_155455_comb[15]}}, p6_sel_155455_comb} + {{1{p6_sel_155456_comb[15]}}, p6_sel_155456_comb};
  assign p6_add_156245_comb = {{1{p6_sel_155457_comb[15]}}, p6_sel_155457_comb} + {{1{p6_sel_155458_comb[15]}}, p6_sel_155458_comb};
  assign p6_add_156246_comb = {{1{p6_sel_155459_comb[15]}}, p6_sel_155459_comb} + {{1{p6_sel_155460_comb[15]}}, p6_sel_155460_comb};
  assign p6_add_156247_comb = {{1{p6_sel_155461_comb[15]}}, p6_sel_155461_comb} + {{1{p6_sel_155462_comb[15]}}, p6_sel_155462_comb};
  assign p6_add_156248_comb = {{1{p6_sel_155463_comb[15]}}, p6_sel_155463_comb} + {{1{p6_sel_155464_comb[15]}}, p6_sel_155464_comb};
  assign p6_add_156249_comb = {{1{p6_sel_155465_comb[15]}}, p6_sel_155465_comb} + {{1{p6_sel_155466_comb[15]}}, p6_sel_155466_comb};
  assign p6_add_156250_comb = {{1{p6_sel_155467_comb[15]}}, p6_sel_155467_comb} + {{1{p6_sel_155468_comb[15]}}, p6_sel_155468_comb};
  assign p6_add_156283_comb = {{1{p6_sel_155533_comb[15]}}, p6_sel_155533_comb} + {{1{p6_sel_155534_comb[15]}}, p6_sel_155534_comb};
  assign p6_add_156284_comb = {{1{p6_sel_155535_comb[15]}}, p6_sel_155535_comb} + {{1{p6_sel_155536_comb[15]}}, p6_sel_155536_comb};
  assign p6_add_156285_comb = {{1{p6_sel_155537_comb[15]}}, p6_sel_155537_comb} + {{1{p6_sel_155538_comb[15]}}, p6_sel_155538_comb};
  assign p6_add_156286_comb = {{1{p6_sel_155539_comb[15]}}, p6_sel_155539_comb} + {{1{p6_sel_155540_comb[15]}}, p6_sel_155540_comb};
  assign p6_add_156287_comb = {{1{p6_sel_155541_comb[15]}}, p6_sel_155541_comb} + {{1{p6_sel_155542_comb[15]}}, p6_sel_155542_comb};
  assign p6_add_156288_comb = {{1{p6_sel_155543_comb[15]}}, p6_sel_155543_comb} + {{1{p6_sel_155544_comb[15]}}, p6_sel_155544_comb};
  assign p6_add_156289_comb = {{1{p6_sel_155545_comb[15]}}, p6_sel_155545_comb} + {{1{p6_sel_155546_comb[15]}}, p6_sel_155546_comb};
  assign p6_add_156290_comb = {{1{p6_sel_155547_comb[15]}}, p6_sel_155547_comb} + {{1{p6_sel_155548_comb[15]}}, p6_sel_155548_comb};
  assign p6_add_156291_comb = {{1{p6_sel_155549_comb[15]}}, p6_sel_155549_comb} + {{1{p6_sel_155550_comb[15]}}, p6_sel_155550_comb};
  assign p6_add_156292_comb = {{1{p6_sel_155551_comb[15]}}, p6_sel_155551_comb} + {{1{p6_sel_155552_comb[15]}}, p6_sel_155552_comb};
  assign p6_add_156293_comb = {{1{p6_sel_155553_comb[15]}}, p6_sel_155553_comb} + {{1{p6_sel_155554_comb[15]}}, p6_sel_155554_comb};
  assign p6_add_156294_comb = {{1{p6_sel_155555_comb[15]}}, p6_sel_155555_comb} + {{1{p6_sel_155556_comb[15]}}, p6_sel_155556_comb};
  assign p6_add_156295_comb = {{1{p6_sel_155557_comb[15]}}, p6_sel_155557_comb} + {{1{p6_sel_155558_comb[15]}}, p6_sel_155558_comb};
  assign p6_add_156296_comb = {{1{p6_sel_155559_comb[15]}}, p6_sel_155559_comb} + {{1{p6_sel_155560_comb[15]}}, p6_sel_155560_comb};
  assign p6_add_156297_comb = {{1{p6_sel_155561_comb[15]}}, p6_sel_155561_comb} + {{1{p6_sel_155562_comb[15]}}, p6_sel_155562_comb};
  assign p6_add_156298_comb = {{1{p6_sel_155563_comb[15]}}, p6_sel_155563_comb} + {{1{p6_sel_155564_comb[15]}}, p6_sel_155564_comb};
  assign p6_add_156299_comb = {{1{p5_sel_150177[15]}}, p5_sel_150177} + {{1{p6_sel_155565_comb[15]}}, p6_sel_155565_comb};
  assign p6_add_156300_comb = {{1{p6_sel_155566_comb[15]}}, p6_sel_155566_comb} + {{1{p6_sel_155567_comb[15]}}, p6_sel_155567_comb};
  assign p6_add_156301_comb = {{1{p6_sel_155568_comb[15]}}, p6_sel_155568_comb} + {{1{p6_sel_155569_comb[15]}}, p6_sel_155569_comb};
  assign p6_add_156302_comb = {{1{p6_sel_155570_comb[15]}}, p6_sel_155570_comb} + {{1{p5_sel_150178[15]}}, p5_sel_150178};
  assign p6_add_156303_comb = {{1{p6_sel_155571_comb[15]}}, p6_sel_155571_comb} + {{1{p6_sel_155572_comb[15]}}, p6_sel_155572_comb};
  assign p6_add_156304_comb = {{1{p6_sel_155573_comb[15]}}, p6_sel_155573_comb} + {{1{p6_sel_155574_comb[15]}}, p6_sel_155574_comb};
  assign p6_add_156305_comb = {{1{p6_sel_155575_comb[15]}}, p6_sel_155575_comb} + {{1{p6_sel_155576_comb[15]}}, p6_sel_155576_comb};
  assign p6_add_156306_comb = {{1{p6_sel_155577_comb[15]}}, p6_sel_155577_comb} + {{1{p6_sel_155578_comb[15]}}, p6_sel_155578_comb};
  assign p6_add_156307_comb = {{1{p6_sel_155579_comb[15]}}, p6_sel_155579_comb} + {{1{p6_sel_155580_comb[15]}}, p6_sel_155580_comb};
  assign p6_add_156308_comb = {{1{p6_sel_155581_comb[15]}}, p6_sel_155581_comb} + {{1{p6_sel_155582_comb[15]}}, p6_sel_155582_comb};
  assign p6_add_156309_comb = {{1{p6_sel_155583_comb[15]}}, p6_sel_155583_comb} + {{1{p6_sel_155584_comb[15]}}, p6_sel_155584_comb};
  assign p6_add_156310_comb = {{1{p6_sel_155585_comb[15]}}, p6_sel_155585_comb} + {{1{p6_sel_155586_comb[15]}}, p6_sel_155586_comb};
  assign p6_add_156311_comb = {{1{p6_sel_155587_comb[15]}}, p6_sel_155587_comb} + {{1{p6_sel_155588_comb[15]}}, p6_sel_155588_comb};
  assign p6_add_156312_comb = {{1{p6_sel_155589_comb[15]}}, p6_sel_155589_comb} + {{1{p6_sel_155590_comb[15]}}, p6_sel_155590_comb};
  assign p6_add_156313_comb = {{1{p6_sel_155591_comb[15]}}, p6_sel_155591_comb} + {{1{p6_sel_155592_comb[15]}}, p6_sel_155592_comb};
  assign p6_add_156314_comb = {{1{p6_sel_155593_comb[15]}}, p6_sel_155593_comb} + {{1{p6_sel_155594_comb[15]}}, p6_sel_155594_comb};
  assign p6_sum__1548_comb = {{8{p6_add_156127_comb[16]}}, p6_add_156127_comb};
  assign p6_sum__1549_comb = {{8{p6_add_156128_comb[16]}}, p6_add_156128_comb};
  assign p6_sum__1550_comb = {{8{p6_add_156129_comb[16]}}, p6_add_156129_comb};
  assign p6_sum__1551_comb = {{8{p6_add_156130_comb[16]}}, p6_add_156130_comb};
  assign p6_sum__1520_comb = {{8{p6_add_156131_comb[16]}}, p6_add_156131_comb};
  assign p6_sum__1521_comb = {{8{p6_add_156132_comb[16]}}, p6_add_156132_comb};
  assign p6_sum__1522_comb = {{8{p6_add_156133_comb[16]}}, p6_add_156133_comb};
  assign p6_sum__1523_comb = {{8{p6_add_156134_comb[16]}}, p6_add_156134_comb};
  assign p6_sum__1492_comb = {{8{p6_add_156135_comb[16]}}, p6_add_156135_comb};
  assign p6_sum__1493_comb = {{8{p6_add_156136_comb[16]}}, p6_add_156136_comb};
  assign p6_sum__1494_comb = {{8{p6_add_156137_comb[16]}}, p6_add_156137_comb};
  assign p6_sum__1495_comb = {{8{p6_add_156138_comb[16]}}, p6_add_156138_comb};
  assign p6_sum__1436_comb = {{8{p6_add_156143_comb[16]}}, p6_add_156143_comb};
  assign p6_sum__1437_comb = {{8{p6_add_156144_comb[16]}}, p6_add_156144_comb};
  assign p6_sum__1438_comb = {{8{p6_add_156145_comb[16]}}, p6_add_156145_comb};
  assign p6_sum__1439_comb = {{8{p6_add_156146_comb[16]}}, p6_add_156146_comb};
  assign p6_sum__1408_comb = {{8{p6_add_156147_comb[16]}}, p6_add_156147_comb};
  assign p6_sum__1409_comb = {{8{p6_add_156148_comb[16]}}, p6_add_156148_comb};
  assign p6_sum__1410_comb = {{8{p6_add_156149_comb[16]}}, p6_add_156149_comb};
  assign p6_sum__1411_comb = {{8{p6_add_156150_comb[16]}}, p6_add_156150_comb};
  assign p6_sum__1380_comb = {{8{p6_add_156151_comb[16]}}, p6_add_156151_comb};
  assign p6_sum__1381_comb = {{8{p6_add_156152_comb[16]}}, p6_add_156152_comb};
  assign p6_sum__1382_comb = {{8{p6_add_156153_comb[16]}}, p6_add_156153_comb};
  assign p6_sum__1383_comb = {{8{p6_add_156154_comb[16]}}, p6_add_156154_comb};
  assign p6_sum__1532_comb = {{8{p6_add_156255_comb[16]}}, p6_add_156255_comb};
  assign p6_sum__1533_comb = {{8{p6_add_156256_comb[16]}}, p6_add_156256_comb};
  assign p6_sum__1534_comb = {{8{p6_add_156257_comb[16]}}, p6_add_156257_comb};
  assign p6_sum__1535_comb = {{8{p6_add_156258_comb[16]}}, p6_add_156258_comb};
  assign p6_sum__1504_comb = {{8{p6_add_156259_comb[16]}}, p6_add_156259_comb};
  assign p6_sum__1505_comb = {{8{p6_add_156260_comb[16]}}, p6_add_156260_comb};
  assign p6_sum__1506_comb = {{8{p6_add_156261_comb[16]}}, p6_add_156261_comb};
  assign p6_sum__1507_comb = {{8{p6_add_156262_comb[16]}}, p6_add_156262_comb};
  assign p6_sum__1476_comb = {{8{p6_add_156263_comb[16]}}, p6_add_156263_comb};
  assign p6_sum__1477_comb = {{8{p6_add_156264_comb[16]}}, p6_add_156264_comb};
  assign p6_sum__1478_comb = {{8{p6_add_156265_comb[16]}}, p6_add_156265_comb};
  assign p6_sum__1479_comb = {{8{p6_add_156266_comb[16]}}, p6_add_156266_comb};
  assign p6_sum__1420_comb = {{8{p6_add_156271_comb[16]}}, p6_add_156271_comb};
  assign p6_sum__1421_comb = {{8{p6_add_156272_comb[16]}}, p6_add_156272_comb};
  assign p6_sum__1422_comb = {{8{p6_add_156273_comb[16]}}, p6_add_156273_comb};
  assign p6_sum__1423_comb = {{8{p6_add_156274_comb[16]}}, p6_add_156274_comb};
  assign p6_sum__1392_comb = {{8{p6_add_156275_comb[16]}}, p6_add_156275_comb};
  assign p6_sum__1393_comb = {{8{p6_add_156276_comb[16]}}, p6_add_156276_comb};
  assign p6_sum__1394_comb = {{8{p6_add_156277_comb[16]}}, p6_add_156277_comb};
  assign p6_sum__1395_comb = {{8{p6_add_156278_comb[16]}}, p6_add_156278_comb};
  assign p6_sum__1364_comb = {{8{p6_add_156279_comb[16]}}, p6_add_156279_comb};
  assign p6_sum__1365_comb = {{8{p6_add_156280_comb[16]}}, p6_add_156280_comb};
  assign p6_sum__1366_comb = {{8{p6_add_156281_comb[16]}}, p6_add_156281_comb};
  assign p6_sum__1367_comb = {{8{p6_add_156282_comb[16]}}, p6_add_156282_comb};
  assign p6_sum__1244_comb = p6_sum__1576_comb + p6_sum__1577_comb;
  assign p6_sum__1245_comb = p6_sum__1578_comb + p6_sum__1579_comb;
  assign p6_sum__1188_comb = p6_sum__1464_comb + p6_sum__1465_comb;
  assign p6_sum__1189_comb = p6_sum__1466_comb + p6_sum__1467_comb;
  assign p6_sum__1236_comb = p6_sum__1560_comb + p6_sum__1561_comb;
  assign p6_sum__1237_comb = p6_sum__1562_comb + p6_sum__1563_comb;
  assign p6_sum__1180_comb = p6_sum__1448_comb + p6_sum__1449_comb;
  assign p6_sum__1181_comb = p6_sum__1450_comb + p6_sum__1451_comb;
  assign p6_add_156699_comb = p6_umul_156555_comb[31:7] + 25'h000_0001;
  assign p6_add_156700_comb = p6_umul_156559_comb[31:7] + 25'h000_0001;
  assign p6_sum__470_comb = p6_sum__468_comb + p6_sum__469_comb;
  assign p6_sum__414_comb = p6_sum__412_comb + p6_sum__413_comb;
  assign p6_sum__358_comb = p6_sum__356_comb + p6_sum__357_comb;
  assign p6_sum__246_comb = p6_sum__244_comb + p6_sum__245_comb;
  assign p6_sum__190_comb = p6_sum__188_comb + p6_sum__189_comb;
  assign p6_sum__134_comb = p6_sum__132_comb + p6_sum__133_comb;
  assign p6_sum__1580_comb = {{8{p6_add_156091_comb[16]}}, p6_add_156091_comb};
  assign p6_sum__1581_comb = {{8{p6_add_156092_comb[16]}}, p6_add_156092_comb};
  assign p6_sum__1582_comb = {{8{p6_add_156093_comb[16]}}, p6_add_156093_comb};
  assign p6_sum__1583_comb = {{8{p6_add_156094_comb[16]}}, p6_add_156094_comb};
  assign p6_sum__1552_comb = {{8{p6_add_156095_comb[16]}}, p6_add_156095_comb};
  assign p6_sum__1553_comb = {{8{p6_add_156096_comb[16]}}, p6_add_156096_comb};
  assign p6_sum__1554_comb = {{8{p6_add_156097_comb[16]}}, p6_add_156097_comb};
  assign p6_sum__1555_comb = {{8{p6_add_156098_comb[16]}}, p6_add_156098_comb};
  assign p6_sum__1524_comb = {{8{p6_add_156099_comb[16]}}, p6_add_156099_comb};
  assign p6_sum__1525_comb = {{8{p6_add_156100_comb[16]}}, p6_add_156100_comb};
  assign p6_sum__1526_comb = {{8{p6_add_156101_comb[16]}}, p6_add_156101_comb};
  assign p6_sum__1527_comb = {{8{p6_add_156102_comb[16]}}, p6_add_156102_comb};
  assign p6_sum__1496_comb = {{8{p6_add_156103_comb[16]}}, p6_add_156103_comb};
  assign p6_sum__1497_comb = {{8{p6_add_156104_comb[16]}}, p6_add_156104_comb};
  assign p6_sum__1498_comb = {{8{p6_add_156105_comb[16]}}, p6_add_156105_comb};
  assign p6_sum__1499_comb = {{8{p6_add_156106_comb[16]}}, p6_add_156106_comb};
  assign p6_sum__1468_comb = {{8{p6_add_156107_comb[16]}}, p6_add_156107_comb};
  assign p6_sum__1469_comb = {{8{p6_add_156108_comb[16]}}, p6_add_156108_comb};
  assign p6_sum__1470_comb = {{8{p6_add_156109_comb[16]}}, p6_add_156109_comb};
  assign p6_sum__1471_comb = {{8{p6_add_156110_comb[16]}}, p6_add_156110_comb};
  assign p6_sum__1440_comb = {{8{p6_add_156111_comb[16]}}, p6_add_156111_comb};
  assign p6_sum__1441_comb = {{8{p6_add_156112_comb[16]}}, p6_add_156112_comb};
  assign p6_sum__1442_comb = {{8{p6_add_156113_comb[16]}}, p6_add_156113_comb};
  assign p6_sum__1443_comb = {{8{p6_add_156114_comb[16]}}, p6_add_156114_comb};
  assign p6_sum__1412_comb = {{8{p6_add_156115_comb[16]}}, p6_add_156115_comb};
  assign p6_sum__1413_comb = {{8{p6_add_156116_comb[16]}}, p6_add_156116_comb};
  assign p6_sum__1414_comb = {{8{p6_add_156117_comb[16]}}, p6_add_156117_comb};
  assign p6_sum__1415_comb = {{8{p6_add_156118_comb[16]}}, p6_add_156118_comb};
  assign p6_sum__1384_comb = {{8{p6_add_156119_comb[16]}}, p6_add_156119_comb};
  assign p6_sum__1385_comb = {{8{p6_add_156120_comb[16]}}, p6_add_156120_comb};
  assign p6_sum__1386_comb = {{8{p6_add_156121_comb[16]}}, p6_add_156121_comb};
  assign p6_sum__1387_comb = {{8{p6_add_156122_comb[16]}}, p6_add_156122_comb};
  assign p6_sum__1572_comb = {{8{p6_add_156155_comb[16]}}, p6_add_156155_comb};
  assign p6_sum__1573_comb = {{8{p6_add_156156_comb[16]}}, p6_add_156156_comb};
  assign p6_sum__1574_comb = {{8{p6_add_156157_comb[16]}}, p6_add_156157_comb};
  assign p6_sum__1575_comb = {{8{p6_add_156158_comb[16]}}, p6_add_156158_comb};
  assign p6_sum__1544_comb = {{8{p6_add_156159_comb[16]}}, p6_add_156159_comb};
  assign p6_sum__1545_comb = {{8{p6_add_156160_comb[16]}}, p6_add_156160_comb};
  assign p6_sum__1546_comb = {{8{p6_add_156161_comb[16]}}, p6_add_156161_comb};
  assign p6_sum__1547_comb = {{8{p6_add_156162_comb[16]}}, p6_add_156162_comb};
  assign p6_sum__1516_comb = {{8{p6_add_156163_comb[16]}}, p6_add_156163_comb};
  assign p6_sum__1517_comb = {{8{p6_add_156164_comb[16]}}, p6_add_156164_comb};
  assign p6_sum__1518_comb = {{8{p6_add_156165_comb[16]}}, p6_add_156165_comb};
  assign p6_sum__1519_comb = {{8{p6_add_156166_comb[16]}}, p6_add_156166_comb};
  assign p6_sum__1488_comb = {{8{p6_add_156167_comb[16]}}, p6_add_156167_comb};
  assign p6_sum__1489_comb = {{8{p6_add_156168_comb[16]}}, p6_add_156168_comb};
  assign p6_sum__1490_comb = {{8{p6_add_156169_comb[16]}}, p6_add_156169_comb};
  assign p6_sum__1491_comb = {{8{p6_add_156170_comb[16]}}, p6_add_156170_comb};
  assign p6_sum__1460_comb = {{8{p6_add_156171_comb[16]}}, p6_add_156171_comb};
  assign p6_sum__1461_comb = {{8{p6_add_156172_comb[16]}}, p6_add_156172_comb};
  assign p6_sum__1462_comb = {{8{p6_add_156173_comb[16]}}, p6_add_156173_comb};
  assign p6_sum__1463_comb = {{8{p6_add_156174_comb[16]}}, p6_add_156174_comb};
  assign p6_sum__1432_comb = {{8{p6_add_156175_comb[16]}}, p6_add_156175_comb};
  assign p6_sum__1433_comb = {{8{p6_add_156176_comb[16]}}, p6_add_156176_comb};
  assign p6_sum__1434_comb = {{8{p6_add_156177_comb[16]}}, p6_add_156177_comb};
  assign p6_sum__1435_comb = {{8{p6_add_156178_comb[16]}}, p6_add_156178_comb};
  assign p6_sum__1404_comb = {{8{p6_add_156179_comb[16]}}, p6_add_156179_comb};
  assign p6_sum__1405_comb = {{8{p6_add_156180_comb[16]}}, p6_add_156180_comb};
  assign p6_sum__1406_comb = {{8{p6_add_156181_comb[16]}}, p6_add_156181_comb};
  assign p6_sum__1407_comb = {{8{p6_add_156182_comb[16]}}, p6_add_156182_comb};
  assign p6_sum__1376_comb = {{8{p6_add_156183_comb[16]}}, p6_add_156183_comb};
  assign p6_sum__1377_comb = {{8{p6_add_156184_comb[16]}}, p6_add_156184_comb};
  assign p6_sum__1378_comb = {{8{p6_add_156185_comb[16]}}, p6_add_156185_comb};
  assign p6_sum__1379_comb = {{8{p6_add_156186_comb[16]}}, p6_add_156186_comb};
  assign p6_sum__1568_comb = {{8{p6_add_156187_comb[16]}}, p6_add_156187_comb};
  assign p6_sum__1569_comb = {{8{p6_add_156188_comb[16]}}, p6_add_156188_comb};
  assign p6_sum__1570_comb = {{8{p6_add_156189_comb[16]}}, p6_add_156189_comb};
  assign p6_sum__1571_comb = {{8{p6_add_156190_comb[16]}}, p6_add_156190_comb};
  assign p6_sum__1540_comb = {{8{p6_add_156191_comb[16]}}, p6_add_156191_comb};
  assign p6_sum__1541_comb = {{8{p6_add_156192_comb[16]}}, p6_add_156192_comb};
  assign p6_sum__1542_comb = {{8{p6_add_156193_comb[16]}}, p6_add_156193_comb};
  assign p6_sum__1543_comb = {{8{p6_add_156194_comb[16]}}, p6_add_156194_comb};
  assign p6_sum__1512_comb = {{8{p6_add_156195_comb[16]}}, p6_add_156195_comb};
  assign p6_sum__1513_comb = {{8{p6_add_156196_comb[16]}}, p6_add_156196_comb};
  assign p6_sum__1514_comb = {{8{p6_add_156197_comb[16]}}, p6_add_156197_comb};
  assign p6_sum__1515_comb = {{8{p6_add_156198_comb[16]}}, p6_add_156198_comb};
  assign p6_sum__1484_comb = {{8{p6_add_156199_comb[16]}}, p6_add_156199_comb};
  assign p6_sum__1485_comb = {{8{p6_add_156200_comb[16]}}, p6_add_156200_comb};
  assign p6_sum__1486_comb = {{8{p6_add_156201_comb[16]}}, p6_add_156201_comb};
  assign p6_sum__1487_comb = {{8{p6_add_156202_comb[16]}}, p6_add_156202_comb};
  assign p6_sum__1456_comb = {{8{p6_add_156203_comb[16]}}, p6_add_156203_comb};
  assign p6_sum__1457_comb = {{8{p6_add_156204_comb[16]}}, p6_add_156204_comb};
  assign p6_sum__1458_comb = {{8{p6_add_156205_comb[16]}}, p6_add_156205_comb};
  assign p6_sum__1459_comb = {{8{p6_add_156206_comb[16]}}, p6_add_156206_comb};
  assign p6_sum__1428_comb = {{8{p6_add_156207_comb[16]}}, p6_add_156207_comb};
  assign p6_sum__1429_comb = {{8{p6_add_156208_comb[16]}}, p6_add_156208_comb};
  assign p6_sum__1430_comb = {{8{p6_add_156209_comb[16]}}, p6_add_156209_comb};
  assign p6_sum__1431_comb = {{8{p6_add_156210_comb[16]}}, p6_add_156210_comb};
  assign p6_sum__1400_comb = {{8{p6_add_156211_comb[16]}}, p6_add_156211_comb};
  assign p6_sum__1401_comb = {{8{p6_add_156212_comb[16]}}, p6_add_156212_comb};
  assign p6_sum__1402_comb = {{8{p6_add_156213_comb[16]}}, p6_add_156213_comb};
  assign p6_sum__1403_comb = {{8{p6_add_156214_comb[16]}}, p6_add_156214_comb};
  assign p6_sum__1372_comb = {{8{p6_add_156215_comb[16]}}, p6_add_156215_comb};
  assign p6_sum__1373_comb = {{8{p6_add_156216_comb[16]}}, p6_add_156216_comb};
  assign p6_sum__1374_comb = {{8{p6_add_156217_comb[16]}}, p6_add_156217_comb};
  assign p6_sum__1375_comb = {{8{p6_add_156218_comb[16]}}, p6_add_156218_comb};
  assign p6_sum__1564_comb = {{8{p6_add_156219_comb[16]}}, p6_add_156219_comb};
  assign p6_sum__1565_comb = {{8{p6_add_156220_comb[16]}}, p6_add_156220_comb};
  assign p6_sum__1566_comb = {{8{p6_add_156221_comb[16]}}, p6_add_156221_comb};
  assign p6_sum__1567_comb = {{8{p6_add_156222_comb[16]}}, p6_add_156222_comb};
  assign p6_sum__1536_comb = {{8{p6_add_156223_comb[16]}}, p6_add_156223_comb};
  assign p6_sum__1537_comb = {{8{p6_add_156224_comb[16]}}, p6_add_156224_comb};
  assign p6_sum__1538_comb = {{8{p6_add_156225_comb[16]}}, p6_add_156225_comb};
  assign p6_sum__1539_comb = {{8{p6_add_156226_comb[16]}}, p6_add_156226_comb};
  assign p6_sum__1508_comb = {{8{p6_add_156227_comb[16]}}, p6_add_156227_comb};
  assign p6_sum__1509_comb = {{8{p6_add_156228_comb[16]}}, p6_add_156228_comb};
  assign p6_sum__1510_comb = {{8{p6_add_156229_comb[16]}}, p6_add_156229_comb};
  assign p6_sum__1511_comb = {{8{p6_add_156230_comb[16]}}, p6_add_156230_comb};
  assign p6_sum__1480_comb = {{8{p6_add_156231_comb[16]}}, p6_add_156231_comb};
  assign p6_sum__1481_comb = {{8{p6_add_156232_comb[16]}}, p6_add_156232_comb};
  assign p6_sum__1482_comb = {{8{p6_add_156233_comb[16]}}, p6_add_156233_comb};
  assign p6_sum__1483_comb = {{8{p6_add_156234_comb[16]}}, p6_add_156234_comb};
  assign p6_sum__1452_comb = {{8{p6_add_156235_comb[16]}}, p6_add_156235_comb};
  assign p6_sum__1453_comb = {{8{p6_add_156236_comb[16]}}, p6_add_156236_comb};
  assign p6_sum__1454_comb = {{8{p6_add_156237_comb[16]}}, p6_add_156237_comb};
  assign p6_sum__1455_comb = {{8{p6_add_156238_comb[16]}}, p6_add_156238_comb};
  assign p6_sum__1424_comb = {{8{p6_add_156239_comb[16]}}, p6_add_156239_comb};
  assign p6_sum__1425_comb = {{8{p6_add_156240_comb[16]}}, p6_add_156240_comb};
  assign p6_sum__1426_comb = {{8{p6_add_156241_comb[16]}}, p6_add_156241_comb};
  assign p6_sum__1427_comb = {{8{p6_add_156242_comb[16]}}, p6_add_156242_comb};
  assign p6_sum__1396_comb = {{8{p6_add_156243_comb[16]}}, p6_add_156243_comb};
  assign p6_sum__1397_comb = {{8{p6_add_156244_comb[16]}}, p6_add_156244_comb};
  assign p6_sum__1398_comb = {{8{p6_add_156245_comb[16]}}, p6_add_156245_comb};
  assign p6_sum__1399_comb = {{8{p6_add_156246_comb[16]}}, p6_add_156246_comb};
  assign p6_sum__1368_comb = {{8{p6_add_156247_comb[16]}}, p6_add_156247_comb};
  assign p6_sum__1369_comb = {{8{p6_add_156248_comb[16]}}, p6_add_156248_comb};
  assign p6_sum__1370_comb = {{8{p6_add_156249_comb[16]}}, p6_add_156249_comb};
  assign p6_sum__1371_comb = {{8{p6_add_156250_comb[16]}}, p6_add_156250_comb};
  assign p6_sum__1556_comb = {{8{p6_add_156283_comb[16]}}, p6_add_156283_comb};
  assign p6_sum__1557_comb = {{8{p6_add_156284_comb[16]}}, p6_add_156284_comb};
  assign p6_sum__1558_comb = {{8{p6_add_156285_comb[16]}}, p6_add_156285_comb};
  assign p6_sum__1559_comb = {{8{p6_add_156286_comb[16]}}, p6_add_156286_comb};
  assign p6_sum__1528_comb = {{8{p6_add_156287_comb[16]}}, p6_add_156287_comb};
  assign p6_sum__1529_comb = {{8{p6_add_156288_comb[16]}}, p6_add_156288_comb};
  assign p6_sum__1530_comb = {{8{p6_add_156289_comb[16]}}, p6_add_156289_comb};
  assign p6_sum__1531_comb = {{8{p6_add_156290_comb[16]}}, p6_add_156290_comb};
  assign p6_sum__1500_comb = {{8{p6_add_156291_comb[16]}}, p6_add_156291_comb};
  assign p6_sum__1501_comb = {{8{p6_add_156292_comb[16]}}, p6_add_156292_comb};
  assign p6_sum__1502_comb = {{8{p6_add_156293_comb[16]}}, p6_add_156293_comb};
  assign p6_sum__1503_comb = {{8{p6_add_156294_comb[16]}}, p6_add_156294_comb};
  assign p6_sum__1472_comb = {{8{p6_add_156295_comb[16]}}, p6_add_156295_comb};
  assign p6_sum__1473_comb = {{8{p6_add_156296_comb[16]}}, p6_add_156296_comb};
  assign p6_sum__1474_comb = {{8{p6_add_156297_comb[16]}}, p6_add_156297_comb};
  assign p6_sum__1475_comb = {{8{p6_add_156298_comb[16]}}, p6_add_156298_comb};
  assign p6_sum__1444_comb = {{8{p6_add_156299_comb[16]}}, p6_add_156299_comb};
  assign p6_sum__1445_comb = {{8{p6_add_156300_comb[16]}}, p6_add_156300_comb};
  assign p6_sum__1446_comb = {{8{p6_add_156301_comb[16]}}, p6_add_156301_comb};
  assign p6_sum__1447_comb = {{8{p6_add_156302_comb[16]}}, p6_add_156302_comb};
  assign p6_sum__1416_comb = {{8{p6_add_156303_comb[16]}}, p6_add_156303_comb};
  assign p6_sum__1417_comb = {{8{p6_add_156304_comb[16]}}, p6_add_156304_comb};
  assign p6_sum__1418_comb = {{8{p6_add_156305_comb[16]}}, p6_add_156305_comb};
  assign p6_sum__1419_comb = {{8{p6_add_156306_comb[16]}}, p6_add_156306_comb};
  assign p6_sum__1388_comb = {{8{p6_add_156307_comb[16]}}, p6_add_156307_comb};
  assign p6_sum__1389_comb = {{8{p6_add_156308_comb[16]}}, p6_add_156308_comb};
  assign p6_sum__1390_comb = {{8{p6_add_156309_comb[16]}}, p6_add_156309_comb};
  assign p6_sum__1391_comb = {{8{p6_add_156310_comb[16]}}, p6_add_156310_comb};
  assign p6_sum__1360_comb = {{8{p6_add_156311_comb[16]}}, p6_add_156311_comb};
  assign p6_sum__1361_comb = {{8{p6_add_156312_comb[16]}}, p6_add_156312_comb};
  assign p6_sum__1362_comb = {{8{p6_add_156313_comb[16]}}, p6_add_156313_comb};
  assign p6_sum__1363_comb = {{8{p6_add_156314_comb[16]}}, p6_add_156314_comb};
  assign p6_sum__1230_comb = p6_sum__1548_comb + p6_sum__1549_comb;
  assign p6_sum__1231_comb = p6_sum__1550_comb + p6_sum__1551_comb;
  assign p6_sum__1216_comb = p6_sum__1520_comb + p6_sum__1521_comb;
  assign p6_sum__1217_comb = p6_sum__1522_comb + p6_sum__1523_comb;
  assign p6_sum__1202_comb = p6_sum__1492_comb + p6_sum__1493_comb;
  assign p6_sum__1203_comb = p6_sum__1494_comb + p6_sum__1495_comb;
  assign p6_sum__1174_comb = p6_sum__1436_comb + p6_sum__1437_comb;
  assign p6_sum__1175_comb = p6_sum__1438_comb + p6_sum__1439_comb;
  assign p6_sum__1160_comb = p6_sum__1408_comb + p6_sum__1409_comb;
  assign p6_sum__1161_comb = p6_sum__1410_comb + p6_sum__1411_comb;
  assign p6_sum__1146_comb = p6_sum__1380_comb + p6_sum__1381_comb;
  assign p6_sum__1147_comb = p6_sum__1382_comb + p6_sum__1383_comb;
  assign p6_sum__1222_comb = p6_sum__1532_comb + p6_sum__1533_comb;
  assign p6_sum__1223_comb = p6_sum__1534_comb + p6_sum__1535_comb;
  assign p6_sum__1208_comb = p6_sum__1504_comb + p6_sum__1505_comb;
  assign p6_sum__1209_comb = p6_sum__1506_comb + p6_sum__1507_comb;
  assign p6_sum__1194_comb = p6_sum__1476_comb + p6_sum__1477_comb;
  assign p6_sum__1195_comb = p6_sum__1478_comb + p6_sum__1479_comb;
  assign p6_sum__1166_comb = p6_sum__1420_comb + p6_sum__1421_comb;
  assign p6_sum__1167_comb = p6_sum__1422_comb + p6_sum__1423_comb;
  assign p6_sum__1152_comb = p6_sum__1392_comb + p6_sum__1393_comb;
  assign p6_sum__1153_comb = p6_sum__1394_comb + p6_sum__1395_comb;
  assign p6_sum__1138_comb = p6_sum__1364_comb + p6_sum__1365_comb;
  assign p6_sum__1139_comb = p6_sum__1366_comb + p6_sum__1367_comb;
  assign p6_sum__1078_comb = p6_sum__1244_comb + p6_sum__1245_comb;
  assign p6_sum__1050_comb = p6_sum__1188_comb + p6_sum__1189_comb;
  assign p6_sum__1074_comb = p6_sum__1236_comb + p6_sum__1237_comb;
  assign p6_sum__1046_comb = p6_sum__1180_comb + p6_sum__1181_comb;
  assign p6_umul_156556_comb = umul32b_32b_x_7b(p6_sum__470_comb, 7'h5b);
  assign p6_umul_156557_comb = umul32b_32b_x_7b(p6_sum__414_comb, 7'h5b);
  assign p6_umul_156558_comb = umul32b_32b_x_7b(p6_sum__358_comb, 7'h5b);
  assign p6_umul_156560_comb = umul32b_32b_x_7b(p6_sum__246_comb, 7'h5b);
  assign p6_umul_156561_comb = umul32b_32b_x_7b(p6_sum__190_comb, 7'h5b);
  assign p6_umul_156562_comb = umul32b_32b_x_7b(p6_sum__134_comb, 7'h5b);
  assign p6_sum__1246_comb = p6_sum__1580_comb + p6_sum__1581_comb;
  assign p6_sum__1247_comb = p6_sum__1582_comb + p6_sum__1583_comb;
  assign p6_sum__1232_comb = p6_sum__1552_comb + p6_sum__1553_comb;
  assign p6_sum__1233_comb = p6_sum__1554_comb + p6_sum__1555_comb;
  assign p6_sum__1218_comb = p6_sum__1524_comb + p6_sum__1525_comb;
  assign p6_sum__1219_comb = p6_sum__1526_comb + p6_sum__1527_comb;
  assign p6_sum__1204_comb = p6_sum__1496_comb + p6_sum__1497_comb;
  assign p6_sum__1205_comb = p6_sum__1498_comb + p6_sum__1499_comb;
  assign p6_sum__1190_comb = p6_sum__1468_comb + p6_sum__1469_comb;
  assign p6_sum__1191_comb = p6_sum__1470_comb + p6_sum__1471_comb;
  assign p6_sum__1176_comb = p6_sum__1440_comb + p6_sum__1441_comb;
  assign p6_sum__1177_comb = p6_sum__1442_comb + p6_sum__1443_comb;
  assign p6_sum__1162_comb = p6_sum__1412_comb + p6_sum__1413_comb;
  assign p6_sum__1163_comb = p6_sum__1414_comb + p6_sum__1415_comb;
  assign p6_sum__1148_comb = p6_sum__1384_comb + p6_sum__1385_comb;
  assign p6_sum__1149_comb = p6_sum__1386_comb + p6_sum__1387_comb;
  assign p6_sum__1242_comb = p6_sum__1572_comb + p6_sum__1573_comb;
  assign p6_sum__1243_comb = p6_sum__1574_comb + p6_sum__1575_comb;
  assign p6_sum__1228_comb = p6_sum__1544_comb + p6_sum__1545_comb;
  assign p6_sum__1229_comb = p6_sum__1546_comb + p6_sum__1547_comb;
  assign p6_sum__1214_comb = p6_sum__1516_comb + p6_sum__1517_comb;
  assign p6_sum__1215_comb = p6_sum__1518_comb + p6_sum__1519_comb;
  assign p6_sum__1200_comb = p6_sum__1488_comb + p6_sum__1489_comb;
  assign p6_sum__1201_comb = p6_sum__1490_comb + p6_sum__1491_comb;
  assign p6_sum__1186_comb = p6_sum__1460_comb + p6_sum__1461_comb;
  assign p6_sum__1187_comb = p6_sum__1462_comb + p6_sum__1463_comb;
  assign p6_sum__1172_comb = p6_sum__1432_comb + p6_sum__1433_comb;
  assign p6_sum__1173_comb = p6_sum__1434_comb + p6_sum__1435_comb;
  assign p6_sum__1158_comb = p6_sum__1404_comb + p6_sum__1405_comb;
  assign p6_sum__1159_comb = p6_sum__1406_comb + p6_sum__1407_comb;
  assign p6_sum__1144_comb = p6_sum__1376_comb + p6_sum__1377_comb;
  assign p6_sum__1145_comb = p6_sum__1378_comb + p6_sum__1379_comb;
  assign p6_sum__1240_comb = p6_sum__1568_comb + p6_sum__1569_comb;
  assign p6_sum__1241_comb = p6_sum__1570_comb + p6_sum__1571_comb;
  assign p6_sum__1226_comb = p6_sum__1540_comb + p6_sum__1541_comb;
  assign p6_sum__1227_comb = p6_sum__1542_comb + p6_sum__1543_comb;
  assign p6_sum__1212_comb = p6_sum__1512_comb + p6_sum__1513_comb;
  assign p6_sum__1213_comb = p6_sum__1514_comb + p6_sum__1515_comb;
  assign p6_sum__1198_comb = p6_sum__1484_comb + p6_sum__1485_comb;
  assign p6_sum__1199_comb = p6_sum__1486_comb + p6_sum__1487_comb;
  assign p6_sum__1184_comb = p6_sum__1456_comb + p6_sum__1457_comb;
  assign p6_sum__1185_comb = p6_sum__1458_comb + p6_sum__1459_comb;
  assign p6_sum__1170_comb = p6_sum__1428_comb + p6_sum__1429_comb;
  assign p6_sum__1171_comb = p6_sum__1430_comb + p6_sum__1431_comb;
  assign p6_sum__1156_comb = p6_sum__1400_comb + p6_sum__1401_comb;
  assign p6_sum__1157_comb = p6_sum__1402_comb + p6_sum__1403_comb;
  assign p6_sum__1142_comb = p6_sum__1372_comb + p6_sum__1373_comb;
  assign p6_sum__1143_comb = p6_sum__1374_comb + p6_sum__1375_comb;
  assign p6_sum__1238_comb = p6_sum__1564_comb + p6_sum__1565_comb;
  assign p6_sum__1239_comb = p6_sum__1566_comb + p6_sum__1567_comb;
  assign p6_sum__1224_comb = p6_sum__1536_comb + p6_sum__1537_comb;
  assign p6_sum__1225_comb = p6_sum__1538_comb + p6_sum__1539_comb;
  assign p6_sum__1210_comb = p6_sum__1508_comb + p6_sum__1509_comb;
  assign p6_sum__1211_comb = p6_sum__1510_comb + p6_sum__1511_comb;
  assign p6_sum__1196_comb = p6_sum__1480_comb + p6_sum__1481_comb;
  assign p6_sum__1197_comb = p6_sum__1482_comb + p6_sum__1483_comb;
  assign p6_sum__1182_comb = p6_sum__1452_comb + p6_sum__1453_comb;
  assign p6_sum__1183_comb = p6_sum__1454_comb + p6_sum__1455_comb;
  assign p6_sum__1168_comb = p6_sum__1424_comb + p6_sum__1425_comb;
  assign p6_sum__1169_comb = p6_sum__1426_comb + p6_sum__1427_comb;
  assign p6_sum__1154_comb = p6_sum__1396_comb + p6_sum__1397_comb;
  assign p6_sum__1155_comb = p6_sum__1398_comb + p6_sum__1399_comb;
  assign p6_sum__1140_comb = p6_sum__1368_comb + p6_sum__1369_comb;
  assign p6_sum__1141_comb = p6_sum__1370_comb + p6_sum__1371_comb;
  assign p6_sum__1234_comb = p6_sum__1556_comb + p6_sum__1557_comb;
  assign p6_sum__1235_comb = p6_sum__1558_comb + p6_sum__1559_comb;
  assign p6_sum__1220_comb = p6_sum__1528_comb + p6_sum__1529_comb;
  assign p6_sum__1221_comb = p6_sum__1530_comb + p6_sum__1531_comb;
  assign p6_sum__1206_comb = p6_sum__1500_comb + p6_sum__1501_comb;
  assign p6_sum__1207_comb = p6_sum__1502_comb + p6_sum__1503_comb;
  assign p6_sum__1192_comb = p6_sum__1472_comb + p6_sum__1473_comb;
  assign p6_sum__1193_comb = p6_sum__1474_comb + p6_sum__1475_comb;
  assign p6_sum__1178_comb = p6_sum__1444_comb + p6_sum__1445_comb;
  assign p6_sum__1179_comb = p6_sum__1446_comb + p6_sum__1447_comb;
  assign p6_sum__1164_comb = p6_sum__1416_comb + p6_sum__1417_comb;
  assign p6_sum__1165_comb = p6_sum__1418_comb + p6_sum__1419_comb;
  assign p6_sum__1150_comb = p6_sum__1388_comb + p6_sum__1389_comb;
  assign p6_sum__1151_comb = p6_sum__1390_comb + p6_sum__1391_comb;
  assign p6_sum__1136_comb = p6_sum__1360_comb + p6_sum__1361_comb;
  assign p6_sum__1137_comb = p6_sum__1362_comb + p6_sum__1363_comb;
  assign p6_sum__1071_comb = p6_sum__1230_comb + p6_sum__1231_comb;
  assign p6_sum__1064_comb = p6_sum__1216_comb + p6_sum__1217_comb;
  assign p6_sum__1057_comb = p6_sum__1202_comb + p6_sum__1203_comb;
  assign p6_sum__1043_comb = p6_sum__1174_comb + p6_sum__1175_comb;
  assign p6_sum__1036_comb = p6_sum__1160_comb + p6_sum__1161_comb;
  assign p6_sum__1029_comb = p6_sum__1146_comb + p6_sum__1147_comb;
  assign p6_sum__1067_comb = p6_sum__1222_comb + p6_sum__1223_comb;
  assign p6_sum__1060_comb = p6_sum__1208_comb + p6_sum__1209_comb;
  assign p6_sum__1053_comb = p6_sum__1194_comb + p6_sum__1195_comb;
  assign p6_sum__1039_comb = p6_sum__1166_comb + p6_sum__1167_comb;
  assign p6_sum__1032_comb = p6_sum__1152_comb + p6_sum__1153_comb;
  assign p6_sum__1025_comb = p6_sum__1138_comb + p6_sum__1139_comb;
  assign p6_add_156701_comb = p6_sum__1078_comb + 25'h000_0001;
  assign p6_add_156702_comb = p6_sum__1050_comb + 25'h000_0001;
  assign p6_add_156703_comb = p6_sum__1074_comb + 25'h000_0001;
  assign p6_add_156704_comb = p6_sum__1046_comb + 25'h000_0001;
  assign p6_sgt_156710_comb = $signed(p6_add_156699_comb[24:1]) > $signed(24'h00_7fff);
  assign p6_bit_slice_156711_comb = p6_add_156699_comb[16:8];
  assign p6_sgt_156713_comb = $signed(p6_add_156700_comb[24:1]) > $signed(24'h00_7fff);
  assign p6_bit_slice_156714_comb = p6_add_156700_comb[16:8];
  assign p6_slt_156715_comb = $signed(p6_add_156699_comb[24:1]) < $signed(24'hff_8000);
  assign p6_slt_156716_comb = $signed(p6_add_156700_comb[24:1]) < $signed(24'hff_8000);

  // Registers for pipe stage 6:
  reg [31:0] p6_umul_156556;
  reg [31:0] p6_umul_156557;
  reg [31:0] p6_umul_156558;
  reg [31:0] p6_umul_156560;
  reg [31:0] p6_umul_156561;
  reg [31:0] p6_umul_156562;
  reg [24:0] p6_sum__1246;
  reg [24:0] p6_sum__1247;
  reg [24:0] p6_sum__1232;
  reg [24:0] p6_sum__1233;
  reg [24:0] p6_sum__1218;
  reg [24:0] p6_sum__1219;
  reg [24:0] p6_sum__1204;
  reg [24:0] p6_sum__1205;
  reg [24:0] p6_sum__1190;
  reg [24:0] p6_sum__1191;
  reg [24:0] p6_sum__1176;
  reg [24:0] p6_sum__1177;
  reg [24:0] p6_sum__1162;
  reg [24:0] p6_sum__1163;
  reg [24:0] p6_sum__1148;
  reg [24:0] p6_sum__1149;
  reg [24:0] p6_sum__1242;
  reg [24:0] p6_sum__1243;
  reg [24:0] p6_sum__1228;
  reg [24:0] p6_sum__1229;
  reg [24:0] p6_sum__1214;
  reg [24:0] p6_sum__1215;
  reg [24:0] p6_sum__1200;
  reg [24:0] p6_sum__1201;
  reg [24:0] p6_sum__1186;
  reg [24:0] p6_sum__1187;
  reg [24:0] p6_sum__1172;
  reg [24:0] p6_sum__1173;
  reg [24:0] p6_sum__1158;
  reg [24:0] p6_sum__1159;
  reg [24:0] p6_sum__1144;
  reg [24:0] p6_sum__1145;
  reg [24:0] p6_sum__1240;
  reg [24:0] p6_sum__1241;
  reg [24:0] p6_sum__1226;
  reg [24:0] p6_sum__1227;
  reg [24:0] p6_sum__1212;
  reg [24:0] p6_sum__1213;
  reg [24:0] p6_sum__1198;
  reg [24:0] p6_sum__1199;
  reg [24:0] p6_sum__1184;
  reg [24:0] p6_sum__1185;
  reg [24:0] p6_sum__1170;
  reg [24:0] p6_sum__1171;
  reg [24:0] p6_sum__1156;
  reg [24:0] p6_sum__1157;
  reg [24:0] p6_sum__1142;
  reg [24:0] p6_sum__1143;
  reg [24:0] p6_sum__1238;
  reg [24:0] p6_sum__1239;
  reg [24:0] p6_sum__1224;
  reg [24:0] p6_sum__1225;
  reg [24:0] p6_sum__1210;
  reg [24:0] p6_sum__1211;
  reg [24:0] p6_sum__1196;
  reg [24:0] p6_sum__1197;
  reg [24:0] p6_sum__1182;
  reg [24:0] p6_sum__1183;
  reg [24:0] p6_sum__1168;
  reg [24:0] p6_sum__1169;
  reg [24:0] p6_sum__1154;
  reg [24:0] p6_sum__1155;
  reg [24:0] p6_sum__1140;
  reg [24:0] p6_sum__1141;
  reg [24:0] p6_sum__1234;
  reg [24:0] p6_sum__1235;
  reg [24:0] p6_sum__1220;
  reg [24:0] p6_sum__1221;
  reg [24:0] p6_sum__1206;
  reg [24:0] p6_sum__1207;
  reg [24:0] p6_sum__1192;
  reg [24:0] p6_sum__1193;
  reg [24:0] p6_sum__1178;
  reg [24:0] p6_sum__1179;
  reg [24:0] p6_sum__1164;
  reg [24:0] p6_sum__1165;
  reg [24:0] p6_sum__1150;
  reg [24:0] p6_sum__1151;
  reg [24:0] p6_sum__1136;
  reg [24:0] p6_sum__1137;
  reg [24:0] p6_sum__1071;
  reg [24:0] p6_sum__1064;
  reg [24:0] p6_sum__1057;
  reg [24:0] p6_sum__1043;
  reg [24:0] p6_sum__1036;
  reg [24:0] p6_sum__1029;
  reg [24:0] p6_sum__1067;
  reg [24:0] p6_sum__1060;
  reg [24:0] p6_sum__1053;
  reg [24:0] p6_sum__1039;
  reg [24:0] p6_sum__1032;
  reg [24:0] p6_sum__1025;
  reg [24:0] p6_add_156701;
  reg [24:0] p6_add_156702;
  reg [24:0] p6_add_156703;
  reg [24:0] p6_add_156704;
  reg p6_sgt_156710;
  reg [8:0] p6_bit_slice_156711;
  reg p6_sgt_156713;
  reg [8:0] p6_bit_slice_156714;
  reg p6_slt_156715;
  reg p6_slt_156716;
  always @ (posedge clk) begin
    p6_umul_156556 <= p6_umul_156556_comb;
    p6_umul_156557 <= p6_umul_156557_comb;
    p6_umul_156558 <= p6_umul_156558_comb;
    p6_umul_156560 <= p6_umul_156560_comb;
    p6_umul_156561 <= p6_umul_156561_comb;
    p6_umul_156562 <= p6_umul_156562_comb;
    p6_sum__1246 <= p6_sum__1246_comb;
    p6_sum__1247 <= p6_sum__1247_comb;
    p6_sum__1232 <= p6_sum__1232_comb;
    p6_sum__1233 <= p6_sum__1233_comb;
    p6_sum__1218 <= p6_sum__1218_comb;
    p6_sum__1219 <= p6_sum__1219_comb;
    p6_sum__1204 <= p6_sum__1204_comb;
    p6_sum__1205 <= p6_sum__1205_comb;
    p6_sum__1190 <= p6_sum__1190_comb;
    p6_sum__1191 <= p6_sum__1191_comb;
    p6_sum__1176 <= p6_sum__1176_comb;
    p6_sum__1177 <= p6_sum__1177_comb;
    p6_sum__1162 <= p6_sum__1162_comb;
    p6_sum__1163 <= p6_sum__1163_comb;
    p6_sum__1148 <= p6_sum__1148_comb;
    p6_sum__1149 <= p6_sum__1149_comb;
    p6_sum__1242 <= p6_sum__1242_comb;
    p6_sum__1243 <= p6_sum__1243_comb;
    p6_sum__1228 <= p6_sum__1228_comb;
    p6_sum__1229 <= p6_sum__1229_comb;
    p6_sum__1214 <= p6_sum__1214_comb;
    p6_sum__1215 <= p6_sum__1215_comb;
    p6_sum__1200 <= p6_sum__1200_comb;
    p6_sum__1201 <= p6_sum__1201_comb;
    p6_sum__1186 <= p6_sum__1186_comb;
    p6_sum__1187 <= p6_sum__1187_comb;
    p6_sum__1172 <= p6_sum__1172_comb;
    p6_sum__1173 <= p6_sum__1173_comb;
    p6_sum__1158 <= p6_sum__1158_comb;
    p6_sum__1159 <= p6_sum__1159_comb;
    p6_sum__1144 <= p6_sum__1144_comb;
    p6_sum__1145 <= p6_sum__1145_comb;
    p6_sum__1240 <= p6_sum__1240_comb;
    p6_sum__1241 <= p6_sum__1241_comb;
    p6_sum__1226 <= p6_sum__1226_comb;
    p6_sum__1227 <= p6_sum__1227_comb;
    p6_sum__1212 <= p6_sum__1212_comb;
    p6_sum__1213 <= p6_sum__1213_comb;
    p6_sum__1198 <= p6_sum__1198_comb;
    p6_sum__1199 <= p6_sum__1199_comb;
    p6_sum__1184 <= p6_sum__1184_comb;
    p6_sum__1185 <= p6_sum__1185_comb;
    p6_sum__1170 <= p6_sum__1170_comb;
    p6_sum__1171 <= p6_sum__1171_comb;
    p6_sum__1156 <= p6_sum__1156_comb;
    p6_sum__1157 <= p6_sum__1157_comb;
    p6_sum__1142 <= p6_sum__1142_comb;
    p6_sum__1143 <= p6_sum__1143_comb;
    p6_sum__1238 <= p6_sum__1238_comb;
    p6_sum__1239 <= p6_sum__1239_comb;
    p6_sum__1224 <= p6_sum__1224_comb;
    p6_sum__1225 <= p6_sum__1225_comb;
    p6_sum__1210 <= p6_sum__1210_comb;
    p6_sum__1211 <= p6_sum__1211_comb;
    p6_sum__1196 <= p6_sum__1196_comb;
    p6_sum__1197 <= p6_sum__1197_comb;
    p6_sum__1182 <= p6_sum__1182_comb;
    p6_sum__1183 <= p6_sum__1183_comb;
    p6_sum__1168 <= p6_sum__1168_comb;
    p6_sum__1169 <= p6_sum__1169_comb;
    p6_sum__1154 <= p6_sum__1154_comb;
    p6_sum__1155 <= p6_sum__1155_comb;
    p6_sum__1140 <= p6_sum__1140_comb;
    p6_sum__1141 <= p6_sum__1141_comb;
    p6_sum__1234 <= p6_sum__1234_comb;
    p6_sum__1235 <= p6_sum__1235_comb;
    p6_sum__1220 <= p6_sum__1220_comb;
    p6_sum__1221 <= p6_sum__1221_comb;
    p6_sum__1206 <= p6_sum__1206_comb;
    p6_sum__1207 <= p6_sum__1207_comb;
    p6_sum__1192 <= p6_sum__1192_comb;
    p6_sum__1193 <= p6_sum__1193_comb;
    p6_sum__1178 <= p6_sum__1178_comb;
    p6_sum__1179 <= p6_sum__1179_comb;
    p6_sum__1164 <= p6_sum__1164_comb;
    p6_sum__1165 <= p6_sum__1165_comb;
    p6_sum__1150 <= p6_sum__1150_comb;
    p6_sum__1151 <= p6_sum__1151_comb;
    p6_sum__1136 <= p6_sum__1136_comb;
    p6_sum__1137 <= p6_sum__1137_comb;
    p6_sum__1071 <= p6_sum__1071_comb;
    p6_sum__1064 <= p6_sum__1064_comb;
    p6_sum__1057 <= p6_sum__1057_comb;
    p6_sum__1043 <= p6_sum__1043_comb;
    p6_sum__1036 <= p6_sum__1036_comb;
    p6_sum__1029 <= p6_sum__1029_comb;
    p6_sum__1067 <= p6_sum__1067_comb;
    p6_sum__1060 <= p6_sum__1060_comb;
    p6_sum__1053 <= p6_sum__1053_comb;
    p6_sum__1039 <= p6_sum__1039_comb;
    p6_sum__1032 <= p6_sum__1032_comb;
    p6_sum__1025 <= p6_sum__1025_comb;
    p6_add_156701 <= p6_add_156701_comb;
    p6_add_156702 <= p6_add_156702_comb;
    p6_add_156703 <= p6_add_156703_comb;
    p6_add_156704 <= p6_add_156704_comb;
    p6_sgt_156710 <= p6_sgt_156710_comb;
    p6_bit_slice_156711 <= p6_bit_slice_156711_comb;
    p6_sgt_156713 <= p6_sgt_156713_comb;
    p6_bit_slice_156714 <= p6_bit_slice_156714_comb;
    p6_slt_156715 <= p6_slt_156715_comb;
    p6_slt_156716 <= p6_slt_156716_comb;
  end

  // ===== Pipe stage 7:
  wire [24:0] p7_sum__1079_comb;
  wire [24:0] p7_sum__1072_comb;
  wire [24:0] p7_sum__1065_comb;
  wire [24:0] p7_sum__1058_comb;
  wire [24:0] p7_sum__1051_comb;
  wire [24:0] p7_sum__1044_comb;
  wire [24:0] p7_sum__1037_comb;
  wire [24:0] p7_sum__1030_comb;
  wire [24:0] p7_sum__1077_comb;
  wire [24:0] p7_sum__1070_comb;
  wire [24:0] p7_sum__1063_comb;
  wire [24:0] p7_sum__1056_comb;
  wire [24:0] p7_sum__1049_comb;
  wire [24:0] p7_sum__1042_comb;
  wire [24:0] p7_sum__1035_comb;
  wire [24:0] p7_sum__1028_comb;
  wire [24:0] p7_sum__1076_comb;
  wire [24:0] p7_sum__1069_comb;
  wire [24:0] p7_sum__1062_comb;
  wire [24:0] p7_sum__1055_comb;
  wire [24:0] p7_sum__1048_comb;
  wire [24:0] p7_sum__1041_comb;
  wire [24:0] p7_sum__1034_comb;
  wire [24:0] p7_sum__1027_comb;
  wire [24:0] p7_sum__1075_comb;
  wire [24:0] p7_sum__1068_comb;
  wire [24:0] p7_sum__1061_comb;
  wire [24:0] p7_sum__1054_comb;
  wire [24:0] p7_sum__1047_comb;
  wire [24:0] p7_sum__1040_comb;
  wire [24:0] p7_sum__1033_comb;
  wire [24:0] p7_sum__1026_comb;
  wire [24:0] p7_sum__1073_comb;
  wire [24:0] p7_sum__1066_comb;
  wire [24:0] p7_sum__1059_comb;
  wire [24:0] p7_sum__1052_comb;
  wire [24:0] p7_sum__1045_comb;
  wire [24:0] p7_sum__1038_comb;
  wire [24:0] p7_sum__1031_comb;
  wire [24:0] p7_sum__1024_comb;
  wire [24:0] p7_add_157051_comb;
  wire [24:0] p7_add_157052_comb;
  wire [24:0] p7_add_157053_comb;
  wire [24:0] p7_add_157054_comb;
  wire [24:0] p7_add_157055_comb;
  wire [24:0] p7_add_157056_comb;
  wire [24:0] p7_add_157081_comb;
  wire [24:0] p7_add_157082_comb;
  wire [24:0] p7_add_157083_comb;
  wire [24:0] p7_add_157084_comb;
  wire [24:0] p7_add_157085_comb;
  wire [24:0] p7_add_157086_comb;
  wire [24:0] p7_add_157037_comb;
  wire [24:0] p7_add_157038_comb;
  wire [24:0] p7_add_157039_comb;
  wire [24:0] p7_add_157040_comb;
  wire [24:0] p7_add_157041_comb;
  wire [24:0] p7_add_157042_comb;
  wire [24:0] p7_add_157043_comb;
  wire [24:0] p7_add_157044_comb;
  wire [24:0] p7_add_157045_comb;
  wire [24:0] p7_add_157046_comb;
  wire [24:0] p7_add_157047_comb;
  wire [24:0] p7_add_157048_comb;
  wire [24:0] p7_add_157049_comb;
  wire [24:0] p7_add_157050_comb;
  wire [24:0] p7_add_157057_comb;
  wire [24:0] p7_add_157058_comb;
  wire [24:0] p7_add_157059_comb;
  wire [24:0] p7_add_157060_comb;
  wire [24:0] p7_add_157061_comb;
  wire [24:0] p7_add_157062_comb;
  wire [24:0] p7_add_157063_comb;
  wire [24:0] p7_add_157064_comb;
  wire [24:0] p7_add_157065_comb;
  wire [24:0] p7_add_157066_comb;
  wire [24:0] p7_add_157067_comb;
  wire [24:0] p7_add_157068_comb;
  wire [24:0] p7_add_157069_comb;
  wire [24:0] p7_add_157070_comb;
  wire [24:0] p7_add_157071_comb;
  wire [24:0] p7_add_157072_comb;
  wire [24:0] p7_add_157073_comb;
  wire [24:0] p7_add_157074_comb;
  wire [24:0] p7_add_157075_comb;
  wire [24:0] p7_add_157076_comb;
  wire [24:0] p7_add_157077_comb;
  wire [24:0] p7_add_157078_comb;
  wire [24:0] p7_add_157079_comb;
  wire [24:0] p7_add_157080_comb;
  wire [24:0] p7_add_157087_comb;
  wire [24:0] p7_add_157088_comb;
  wire [24:0] p7_add_157089_comb;
  wire [24:0] p7_add_157090_comb;
  wire [24:0] p7_add_157091_comb;
  wire [24:0] p7_add_157092_comb;
  wire [24:0] p7_add_157093_comb;
  wire [24:0] p7_add_157094_comb;
  wire [8:0] p7_clipped__320_comb;
  wire [8:0] p7_clipped__324_comb;
  wire [9:0] p7_add_157851_comb;
  wire [9:0] p7_add_157855_comb;
  wire [8:0] p7_clipped__336_comb;
  wire [8:0] p7_clipped__337_comb;
  wire [8:0] p7_clipped__338_comb;
  wire [8:0] p7_clipped__339_comb;
  wire [8:0] p7_clipped__340_comb;
  wire [8:0] p7_clipped__341_comb;
  wire [8:0] p7_clipped__342_comb;
  wire [8:0] p7_clipped__343_comb;
  wire [8:0] p7_clipped__368_comb;
  wire [8:0] p7_clipped__369_comb;
  wire [8:0] p7_clipped__370_comb;
  wire [8:0] p7_clipped__371_comb;
  wire [8:0] p7_clipped__372_comb;
  wire [8:0] p7_clipped__373_comb;
  wire [8:0] p7_clipped__374_comb;
  wire [8:0] p7_clipped__375_comb;
  wire [1:0] p7_bit_slice_157915_comb;
  wire [1:0] p7_bit_slice_157916_comb;
  wire [8:0] p7_clipped__321_comb;
  wire [8:0] p7_clipped__322_comb;
  wire [8:0] p7_clipped__323_comb;
  wire [8:0] p7_clipped__325_comb;
  wire [8:0] p7_clipped__326_comb;
  wire [8:0] p7_clipped__327_comb;
  wire [8:0] p7_clipped__328_comb;
  wire [8:0] p7_clipped__329_comb;
  wire [8:0] p7_clipped__330_comb;
  wire [8:0] p7_clipped__331_comb;
  wire [8:0] p7_clipped__332_comb;
  wire [8:0] p7_clipped__333_comb;
  wire [8:0] p7_clipped__334_comb;
  wire [8:0] p7_clipped__335_comb;
  wire [8:0] p7_clipped__344_comb;
  wire [8:0] p7_clipped__345_comb;
  wire [8:0] p7_clipped__346_comb;
  wire [8:0] p7_clipped__347_comb;
  wire [8:0] p7_clipped__348_comb;
  wire [8:0] p7_clipped__349_comb;
  wire [8:0] p7_clipped__350_comb;
  wire [8:0] p7_clipped__351_comb;
  wire [8:0] p7_clipped__352_comb;
  wire [8:0] p7_clipped__353_comb;
  wire [8:0] p7_clipped__354_comb;
  wire [8:0] p7_clipped__355_comb;
  wire [8:0] p7_clipped__356_comb;
  wire [8:0] p7_clipped__357_comb;
  wire [8:0] p7_clipped__358_comb;
  wire [8:0] p7_clipped__359_comb;
  wire [8:0] p7_clipped__360_comb;
  wire [8:0] p7_clipped__361_comb;
  wire [8:0] p7_clipped__362_comb;
  wire [8:0] p7_clipped__363_comb;
  wire [8:0] p7_clipped__364_comb;
  wire [8:0] p7_clipped__365_comb;
  wire [8:0] p7_clipped__366_comb;
  wire [8:0] p7_clipped__367_comb;
  wire [8:0] p7_clipped__376_comb;
  wire [8:0] p7_clipped__377_comb;
  wire [8:0] p7_clipped__378_comb;
  wire [8:0] p7_clipped__379_comb;
  wire [8:0] p7_clipped__380_comb;
  wire [8:0] p7_clipped__381_comb;
  wire [8:0] p7_clipped__382_comb;
  wire [8:0] p7_clipped__383_comb;
  wire [9:0] p7_add_157867_comb;
  wire [9:0] p7_add_157868_comb;
  wire [9:0] p7_add_157869_comb;
  wire [9:0] p7_add_157870_comb;
  wire [9:0] p7_add_157871_comb;
  wire [9:0] p7_add_157872_comb;
  wire [9:0] p7_add_157873_comb;
  wire [9:0] p7_add_157874_comb;
  wire [9:0] p7_add_157899_comb;
  wire [9:0] p7_add_157900_comb;
  wire [9:0] p7_add_157901_comb;
  wire [9:0] p7_add_157902_comb;
  wire [9:0] p7_add_157903_comb;
  wire [9:0] p7_add_157904_comb;
  wire [9:0] p7_add_157905_comb;
  wire [9:0] p7_add_157906_comb;
  wire [2:0] p7_add_157937_comb;
  wire [2:0] p7_add_157938_comb;
  wire [9:0] p7_add_157852_comb;
  wire [9:0] p7_add_157853_comb;
  wire [9:0] p7_add_157854_comb;
  wire [9:0] p7_add_157856_comb;
  wire [9:0] p7_add_157857_comb;
  wire [9:0] p7_add_157858_comb;
  wire [9:0] p7_add_157859_comb;
  wire [9:0] p7_add_157860_comb;
  wire [9:0] p7_add_157861_comb;
  wire [9:0] p7_add_157862_comb;
  wire [9:0] p7_add_157863_comb;
  wire [9:0] p7_add_157864_comb;
  wire [9:0] p7_add_157865_comb;
  wire [9:0] p7_add_157866_comb;
  wire [9:0] p7_add_157875_comb;
  wire [9:0] p7_add_157876_comb;
  wire [9:0] p7_add_157877_comb;
  wire [9:0] p7_add_157878_comb;
  wire [9:0] p7_add_157879_comb;
  wire [9:0] p7_add_157880_comb;
  wire [9:0] p7_add_157881_comb;
  wire [9:0] p7_add_157882_comb;
  wire [9:0] p7_add_157883_comb;
  wire [9:0] p7_add_157884_comb;
  wire [9:0] p7_add_157885_comb;
  wire [9:0] p7_add_157886_comb;
  wire [9:0] p7_add_157887_comb;
  wire [9:0] p7_add_157888_comb;
  wire [9:0] p7_add_157889_comb;
  wire [9:0] p7_add_157890_comb;
  wire [9:0] p7_add_157891_comb;
  wire [9:0] p7_add_157892_comb;
  wire [9:0] p7_add_157893_comb;
  wire [9:0] p7_add_157894_comb;
  wire [9:0] p7_add_157895_comb;
  wire [9:0] p7_add_157896_comb;
  wire [9:0] p7_add_157897_comb;
  wire [9:0] p7_add_157898_comb;
  wire [9:0] p7_add_157907_comb;
  wire [9:0] p7_add_157908_comb;
  wire [9:0] p7_add_157909_comb;
  wire [9:0] p7_add_157910_comb;
  wire [9:0] p7_add_157911_comb;
  wire [9:0] p7_add_157912_comb;
  wire [9:0] p7_add_157913_comb;
  wire [9:0] p7_add_157914_comb;
  wire [1:0] p7_bit_slice_157917_comb;
  wire [1:0] p7_bit_slice_157918_comb;
  wire [1:0] p7_bit_slice_157919_comb;
  wire [1:0] p7_bit_slice_157920_comb;
  wire [1:0] p7_bit_slice_157921_comb;
  wire [1:0] p7_bit_slice_157922_comb;
  wire [1:0] p7_bit_slice_157923_comb;
  wire [1:0] p7_bit_slice_157924_comb;
  wire [1:0] p7_bit_slice_157925_comb;
  wire [1:0] p7_bit_slice_157926_comb;
  wire [1:0] p7_bit_slice_157927_comb;
  wire [1:0] p7_bit_slice_157928_comb;
  wire [1:0] p7_bit_slice_157929_comb;
  wire [1:0] p7_bit_slice_157930_comb;
  wire [1:0] p7_bit_slice_157931_comb;
  wire [1:0] p7_bit_slice_157932_comb;
  wire p7_bit_slice_157939_comb;
  wire [6:0] p7_bit_slice_157940_comb;
  wire p7_bit_slice_157941_comb;
  wire [6:0] p7_bit_slice_157942_comb;
  wire [6:0] p7_bit_slice_157943_comb;
  wire [6:0] p7_bit_slice_157944_comb;
  wire [6:0] p7_bit_slice_157945_comb;
  wire [6:0] p7_bit_slice_157946_comb;
  wire [6:0] p7_bit_slice_157947_comb;
  wire [6:0] p7_bit_slice_157948_comb;
  wire [6:0] p7_bit_slice_157949_comb;
  wire [6:0] p7_bit_slice_157950_comb;
  wire [6:0] p7_bit_slice_157951_comb;
  wire [6:0] p7_bit_slice_157952_comb;
  wire [6:0] p7_bit_slice_157953_comb;
  wire [6:0] p7_bit_slice_157954_comb;
  wire [6:0] p7_bit_slice_157955_comb;
  wire [6:0] p7_bit_slice_157956_comb;
  wire [6:0] p7_bit_slice_157957_comb;
  wire [6:0] p7_bit_slice_157958_comb;
  wire p7_bit_slice_157959_comb;
  wire p7_bit_slice_157960_comb;
  assign p7_sum__1079_comb = p6_sum__1246 + p6_sum__1247;
  assign p7_sum__1072_comb = p6_sum__1232 + p6_sum__1233;
  assign p7_sum__1065_comb = p6_sum__1218 + p6_sum__1219;
  assign p7_sum__1058_comb = p6_sum__1204 + p6_sum__1205;
  assign p7_sum__1051_comb = p6_sum__1190 + p6_sum__1191;
  assign p7_sum__1044_comb = p6_sum__1176 + p6_sum__1177;
  assign p7_sum__1037_comb = p6_sum__1162 + p6_sum__1163;
  assign p7_sum__1030_comb = p6_sum__1148 + p6_sum__1149;
  assign p7_sum__1077_comb = p6_sum__1242 + p6_sum__1243;
  assign p7_sum__1070_comb = p6_sum__1228 + p6_sum__1229;
  assign p7_sum__1063_comb = p6_sum__1214 + p6_sum__1215;
  assign p7_sum__1056_comb = p6_sum__1200 + p6_sum__1201;
  assign p7_sum__1049_comb = p6_sum__1186 + p6_sum__1187;
  assign p7_sum__1042_comb = p6_sum__1172 + p6_sum__1173;
  assign p7_sum__1035_comb = p6_sum__1158 + p6_sum__1159;
  assign p7_sum__1028_comb = p6_sum__1144 + p6_sum__1145;
  assign p7_sum__1076_comb = p6_sum__1240 + p6_sum__1241;
  assign p7_sum__1069_comb = p6_sum__1226 + p6_sum__1227;
  assign p7_sum__1062_comb = p6_sum__1212 + p6_sum__1213;
  assign p7_sum__1055_comb = p6_sum__1198 + p6_sum__1199;
  assign p7_sum__1048_comb = p6_sum__1184 + p6_sum__1185;
  assign p7_sum__1041_comb = p6_sum__1170 + p6_sum__1171;
  assign p7_sum__1034_comb = p6_sum__1156 + p6_sum__1157;
  assign p7_sum__1027_comb = p6_sum__1142 + p6_sum__1143;
  assign p7_sum__1075_comb = p6_sum__1238 + p6_sum__1239;
  assign p7_sum__1068_comb = p6_sum__1224 + p6_sum__1225;
  assign p7_sum__1061_comb = p6_sum__1210 + p6_sum__1211;
  assign p7_sum__1054_comb = p6_sum__1196 + p6_sum__1197;
  assign p7_sum__1047_comb = p6_sum__1182 + p6_sum__1183;
  assign p7_sum__1040_comb = p6_sum__1168 + p6_sum__1169;
  assign p7_sum__1033_comb = p6_sum__1154 + p6_sum__1155;
  assign p7_sum__1026_comb = p6_sum__1140 + p6_sum__1141;
  assign p7_sum__1073_comb = p6_sum__1234 + p6_sum__1235;
  assign p7_sum__1066_comb = p6_sum__1220 + p6_sum__1221;
  assign p7_sum__1059_comb = p6_sum__1206 + p6_sum__1207;
  assign p7_sum__1052_comb = p6_sum__1192 + p6_sum__1193;
  assign p7_sum__1045_comb = p6_sum__1178 + p6_sum__1179;
  assign p7_sum__1038_comb = p6_sum__1164 + p6_sum__1165;
  assign p7_sum__1031_comb = p6_sum__1150 + p6_sum__1151;
  assign p7_sum__1024_comb = p6_sum__1136 + p6_sum__1137;
  assign p7_add_157051_comb = p6_sum__1071 + 25'h000_0001;
  assign p7_add_157052_comb = p6_sum__1064 + 25'h000_0001;
  assign p7_add_157053_comb = p6_sum__1057 + 25'h000_0001;
  assign p7_add_157054_comb = p6_sum__1043 + 25'h000_0001;
  assign p7_add_157055_comb = p6_sum__1036 + 25'h000_0001;
  assign p7_add_157056_comb = p6_sum__1029 + 25'h000_0001;
  assign p7_add_157081_comb = p6_sum__1067 + 25'h000_0001;
  assign p7_add_157082_comb = p6_sum__1060 + 25'h000_0001;
  assign p7_add_157083_comb = p6_sum__1053 + 25'h000_0001;
  assign p7_add_157084_comb = p6_sum__1039 + 25'h000_0001;
  assign p7_add_157085_comb = p6_sum__1032 + 25'h000_0001;
  assign p7_add_157086_comb = p6_sum__1025 + 25'h000_0001;
  assign p7_add_157037_comb = p6_umul_156556[31:7] + 25'h000_0001;
  assign p7_add_157038_comb = p6_umul_156557[31:7] + 25'h000_0001;
  assign p7_add_157039_comb = p6_umul_156558[31:7] + 25'h000_0001;
  assign p7_add_157040_comb = p6_umul_156560[31:7] + 25'h000_0001;
  assign p7_add_157041_comb = p6_umul_156561[31:7] + 25'h000_0001;
  assign p7_add_157042_comb = p6_umul_156562[31:7] + 25'h000_0001;
  assign p7_add_157043_comb = p7_sum__1079_comb + 25'h000_0001;
  assign p7_add_157044_comb = p7_sum__1072_comb + 25'h000_0001;
  assign p7_add_157045_comb = p7_sum__1065_comb + 25'h000_0001;
  assign p7_add_157046_comb = p7_sum__1058_comb + 25'h000_0001;
  assign p7_add_157047_comb = p7_sum__1051_comb + 25'h000_0001;
  assign p7_add_157048_comb = p7_sum__1044_comb + 25'h000_0001;
  assign p7_add_157049_comb = p7_sum__1037_comb + 25'h000_0001;
  assign p7_add_157050_comb = p7_sum__1030_comb + 25'h000_0001;
  assign p7_add_157057_comb = p7_sum__1077_comb + 25'h000_0001;
  assign p7_add_157058_comb = p7_sum__1070_comb + 25'h000_0001;
  assign p7_add_157059_comb = p7_sum__1063_comb + 25'h000_0001;
  assign p7_add_157060_comb = p7_sum__1056_comb + 25'h000_0001;
  assign p7_add_157061_comb = p7_sum__1049_comb + 25'h000_0001;
  assign p7_add_157062_comb = p7_sum__1042_comb + 25'h000_0001;
  assign p7_add_157063_comb = p7_sum__1035_comb + 25'h000_0001;
  assign p7_add_157064_comb = p7_sum__1028_comb + 25'h000_0001;
  assign p7_add_157065_comb = p7_sum__1076_comb + 25'h000_0001;
  assign p7_add_157066_comb = p7_sum__1069_comb + 25'h000_0001;
  assign p7_add_157067_comb = p7_sum__1062_comb + 25'h000_0001;
  assign p7_add_157068_comb = p7_sum__1055_comb + 25'h000_0001;
  assign p7_add_157069_comb = p7_sum__1048_comb + 25'h000_0001;
  assign p7_add_157070_comb = p7_sum__1041_comb + 25'h000_0001;
  assign p7_add_157071_comb = p7_sum__1034_comb + 25'h000_0001;
  assign p7_add_157072_comb = p7_sum__1027_comb + 25'h000_0001;
  assign p7_add_157073_comb = p7_sum__1075_comb + 25'h000_0001;
  assign p7_add_157074_comb = p7_sum__1068_comb + 25'h000_0001;
  assign p7_add_157075_comb = p7_sum__1061_comb + 25'h000_0001;
  assign p7_add_157076_comb = p7_sum__1054_comb + 25'h000_0001;
  assign p7_add_157077_comb = p7_sum__1047_comb + 25'h000_0001;
  assign p7_add_157078_comb = p7_sum__1040_comb + 25'h000_0001;
  assign p7_add_157079_comb = p7_sum__1033_comb + 25'h000_0001;
  assign p7_add_157080_comb = p7_sum__1026_comb + 25'h000_0001;
  assign p7_add_157087_comb = p7_sum__1073_comb + 25'h000_0001;
  assign p7_add_157088_comb = p7_sum__1066_comb + 25'h000_0001;
  assign p7_add_157089_comb = p7_sum__1059_comb + 25'h000_0001;
  assign p7_add_157090_comb = p7_sum__1052_comb + 25'h000_0001;
  assign p7_add_157091_comb = p7_sum__1045_comb + 25'h000_0001;
  assign p7_add_157092_comb = p7_sum__1038_comb + 25'h000_0001;
  assign p7_add_157093_comb = p7_sum__1031_comb + 25'h000_0001;
  assign p7_add_157094_comb = p7_sum__1024_comb + 25'h000_0001;
  assign p7_clipped__320_comb = p6_slt_156715 ? 9'h100 : (p6_sgt_156710 ? 9'h0ff : p6_bit_slice_156711);
  assign p7_clipped__324_comb = p6_slt_156716 ? 9'h100 : (p6_sgt_156713 ? 9'h0ff : p6_bit_slice_156714);
  assign p7_add_157851_comb = {{1{p7_clipped__320_comb[8]}}, p7_clipped__320_comb} + 10'h001;
  assign p7_add_157855_comb = {{1{p7_clipped__324_comb[8]}}, p7_clipped__324_comb} + 10'h001;
  assign p7_clipped__336_comb = $signed(p6_add_156701[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p6_add_156701[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p6_add_156701[16:8]);
  assign p7_clipped__337_comb = $signed(p7_add_157051_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157051_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157051_comb[16:8]);
  assign p7_clipped__338_comb = $signed(p7_add_157052_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157052_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157052_comb[16:8]);
  assign p7_clipped__339_comb = $signed(p7_add_157053_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157053_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157053_comb[16:8]);
  assign p7_clipped__340_comb = $signed(p6_add_156702[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p6_add_156702[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p6_add_156702[16:8]);
  assign p7_clipped__341_comb = $signed(p7_add_157054_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157054_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157054_comb[16:8]);
  assign p7_clipped__342_comb = $signed(p7_add_157055_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157055_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157055_comb[16:8]);
  assign p7_clipped__343_comb = $signed(p7_add_157056_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157056_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157056_comb[16:8]);
  assign p7_clipped__368_comb = $signed(p6_add_156703[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p6_add_156703[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p6_add_156703[16:8]);
  assign p7_clipped__369_comb = $signed(p7_add_157081_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157081_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157081_comb[16:8]);
  assign p7_clipped__370_comb = $signed(p7_add_157082_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157082_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157082_comb[16:8]);
  assign p7_clipped__371_comb = $signed(p7_add_157083_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157083_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157083_comb[16:8]);
  assign p7_clipped__372_comb = $signed(p6_add_156704[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p6_add_156704[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p6_add_156704[16:8]);
  assign p7_clipped__373_comb = $signed(p7_add_157084_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157084_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157084_comb[16:8]);
  assign p7_clipped__374_comb = $signed(p7_add_157085_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157085_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157085_comb[16:8]);
  assign p7_clipped__375_comb = $signed(p7_add_157086_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157086_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157086_comb[16:8]);
  assign p7_bit_slice_157915_comb = p7_add_157851_comb[9:8];
  assign p7_bit_slice_157916_comb = p7_add_157855_comb[9:8];
  assign p7_clipped__321_comb = $signed(p7_add_157037_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157037_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157037_comb[16:8]);
  assign p7_clipped__322_comb = $signed(p7_add_157038_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157038_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157038_comb[16:8]);
  assign p7_clipped__323_comb = $signed(p7_add_157039_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157039_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157039_comb[16:8]);
  assign p7_clipped__325_comb = $signed(p7_add_157040_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157040_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157040_comb[16:8]);
  assign p7_clipped__326_comb = $signed(p7_add_157041_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157041_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157041_comb[16:8]);
  assign p7_clipped__327_comb = $signed(p7_add_157042_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157042_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157042_comb[16:8]);
  assign p7_clipped__328_comb = $signed(p7_add_157043_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157043_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157043_comb[16:8]);
  assign p7_clipped__329_comb = $signed(p7_add_157044_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157044_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157044_comb[16:8]);
  assign p7_clipped__330_comb = $signed(p7_add_157045_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157045_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157045_comb[16:8]);
  assign p7_clipped__331_comb = $signed(p7_add_157046_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157046_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157046_comb[16:8]);
  assign p7_clipped__332_comb = $signed(p7_add_157047_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157047_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157047_comb[16:8]);
  assign p7_clipped__333_comb = $signed(p7_add_157048_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157048_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157048_comb[16:8]);
  assign p7_clipped__334_comb = $signed(p7_add_157049_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157049_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157049_comb[16:8]);
  assign p7_clipped__335_comb = $signed(p7_add_157050_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157050_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157050_comb[16:8]);
  assign p7_clipped__344_comb = $signed(p7_add_157057_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157057_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157057_comb[16:8]);
  assign p7_clipped__345_comb = $signed(p7_add_157058_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157058_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157058_comb[16:8]);
  assign p7_clipped__346_comb = $signed(p7_add_157059_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157059_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157059_comb[16:8]);
  assign p7_clipped__347_comb = $signed(p7_add_157060_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157060_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157060_comb[16:8]);
  assign p7_clipped__348_comb = $signed(p7_add_157061_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157061_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157061_comb[16:8]);
  assign p7_clipped__349_comb = $signed(p7_add_157062_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157062_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157062_comb[16:8]);
  assign p7_clipped__350_comb = $signed(p7_add_157063_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157063_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157063_comb[16:8]);
  assign p7_clipped__351_comb = $signed(p7_add_157064_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157064_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157064_comb[16:8]);
  assign p7_clipped__352_comb = $signed(p7_add_157065_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157065_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157065_comb[16:8]);
  assign p7_clipped__353_comb = $signed(p7_add_157066_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157066_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157066_comb[16:8]);
  assign p7_clipped__354_comb = $signed(p7_add_157067_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157067_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157067_comb[16:8]);
  assign p7_clipped__355_comb = $signed(p7_add_157068_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157068_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157068_comb[16:8]);
  assign p7_clipped__356_comb = $signed(p7_add_157069_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157069_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157069_comb[16:8]);
  assign p7_clipped__357_comb = $signed(p7_add_157070_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157070_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157070_comb[16:8]);
  assign p7_clipped__358_comb = $signed(p7_add_157071_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157071_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157071_comb[16:8]);
  assign p7_clipped__359_comb = $signed(p7_add_157072_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157072_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157072_comb[16:8]);
  assign p7_clipped__360_comb = $signed(p7_add_157073_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157073_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157073_comb[16:8]);
  assign p7_clipped__361_comb = $signed(p7_add_157074_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157074_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157074_comb[16:8]);
  assign p7_clipped__362_comb = $signed(p7_add_157075_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157075_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157075_comb[16:8]);
  assign p7_clipped__363_comb = $signed(p7_add_157076_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157076_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157076_comb[16:8]);
  assign p7_clipped__364_comb = $signed(p7_add_157077_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157077_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157077_comb[16:8]);
  assign p7_clipped__365_comb = $signed(p7_add_157078_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157078_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157078_comb[16:8]);
  assign p7_clipped__366_comb = $signed(p7_add_157079_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157079_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157079_comb[16:8]);
  assign p7_clipped__367_comb = $signed(p7_add_157080_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157080_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157080_comb[16:8]);
  assign p7_clipped__376_comb = $signed(p7_add_157087_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157087_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157087_comb[16:8]);
  assign p7_clipped__377_comb = $signed(p7_add_157088_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157088_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157088_comb[16:8]);
  assign p7_clipped__378_comb = $signed(p7_add_157089_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157089_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157089_comb[16:8]);
  assign p7_clipped__379_comb = $signed(p7_add_157090_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157090_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157090_comb[16:8]);
  assign p7_clipped__380_comb = $signed(p7_add_157091_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157091_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157091_comb[16:8]);
  assign p7_clipped__381_comb = $signed(p7_add_157092_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157092_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157092_comb[16:8]);
  assign p7_clipped__382_comb = $signed(p7_add_157093_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157093_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157093_comb[16:8]);
  assign p7_clipped__383_comb = $signed(p7_add_157094_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p7_add_157094_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p7_add_157094_comb[16:8]);
  assign p7_add_157867_comb = {{1{p7_clipped__336_comb[8]}}, p7_clipped__336_comb} + 10'h001;
  assign p7_add_157868_comb = {{1{p7_clipped__337_comb[8]}}, p7_clipped__337_comb} + 10'h001;
  assign p7_add_157869_comb = {{1{p7_clipped__338_comb[8]}}, p7_clipped__338_comb} + 10'h001;
  assign p7_add_157870_comb = {{1{p7_clipped__339_comb[8]}}, p7_clipped__339_comb} + 10'h001;
  assign p7_add_157871_comb = {{1{p7_clipped__340_comb[8]}}, p7_clipped__340_comb} + 10'h001;
  assign p7_add_157872_comb = {{1{p7_clipped__341_comb[8]}}, p7_clipped__341_comb} + 10'h001;
  assign p7_add_157873_comb = {{1{p7_clipped__342_comb[8]}}, p7_clipped__342_comb} + 10'h001;
  assign p7_add_157874_comb = {{1{p7_clipped__343_comb[8]}}, p7_clipped__343_comb} + 10'h001;
  assign p7_add_157899_comb = {{1{p7_clipped__368_comb[8]}}, p7_clipped__368_comb} + 10'h001;
  assign p7_add_157900_comb = {{1{p7_clipped__369_comb[8]}}, p7_clipped__369_comb} + 10'h001;
  assign p7_add_157901_comb = {{1{p7_clipped__370_comb[8]}}, p7_clipped__370_comb} + 10'h001;
  assign p7_add_157902_comb = {{1{p7_clipped__371_comb[8]}}, p7_clipped__371_comb} + 10'h001;
  assign p7_add_157903_comb = {{1{p7_clipped__372_comb[8]}}, p7_clipped__372_comb} + 10'h001;
  assign p7_add_157904_comb = {{1{p7_clipped__373_comb[8]}}, p7_clipped__373_comb} + 10'h001;
  assign p7_add_157905_comb = {{1{p7_clipped__374_comb[8]}}, p7_clipped__374_comb} + 10'h001;
  assign p7_add_157906_comb = {{1{p7_clipped__375_comb[8]}}, p7_clipped__375_comb} + 10'h001;
  assign p7_add_157937_comb = {{1{p7_bit_slice_157915_comb[1]}}, p7_bit_slice_157915_comb} + 3'h1;
  assign p7_add_157938_comb = {{1{p7_bit_slice_157916_comb[1]}}, p7_bit_slice_157916_comb} + 3'h1;
  assign p7_add_157852_comb = {{1{p7_clipped__321_comb[8]}}, p7_clipped__321_comb} + 10'h001;
  assign p7_add_157853_comb = {{1{p7_clipped__322_comb[8]}}, p7_clipped__322_comb} + 10'h001;
  assign p7_add_157854_comb = {{1{p7_clipped__323_comb[8]}}, p7_clipped__323_comb} + 10'h001;
  assign p7_add_157856_comb = {{1{p7_clipped__325_comb[8]}}, p7_clipped__325_comb} + 10'h001;
  assign p7_add_157857_comb = {{1{p7_clipped__326_comb[8]}}, p7_clipped__326_comb} + 10'h001;
  assign p7_add_157858_comb = {{1{p7_clipped__327_comb[8]}}, p7_clipped__327_comb} + 10'h001;
  assign p7_add_157859_comb = {{1{p7_clipped__328_comb[8]}}, p7_clipped__328_comb} + 10'h001;
  assign p7_add_157860_comb = {{1{p7_clipped__329_comb[8]}}, p7_clipped__329_comb} + 10'h001;
  assign p7_add_157861_comb = {{1{p7_clipped__330_comb[8]}}, p7_clipped__330_comb} + 10'h001;
  assign p7_add_157862_comb = {{1{p7_clipped__331_comb[8]}}, p7_clipped__331_comb} + 10'h001;
  assign p7_add_157863_comb = {{1{p7_clipped__332_comb[8]}}, p7_clipped__332_comb} + 10'h001;
  assign p7_add_157864_comb = {{1{p7_clipped__333_comb[8]}}, p7_clipped__333_comb} + 10'h001;
  assign p7_add_157865_comb = {{1{p7_clipped__334_comb[8]}}, p7_clipped__334_comb} + 10'h001;
  assign p7_add_157866_comb = {{1{p7_clipped__335_comb[8]}}, p7_clipped__335_comb} + 10'h001;
  assign p7_add_157875_comb = {{1{p7_clipped__344_comb[8]}}, p7_clipped__344_comb} + 10'h001;
  assign p7_add_157876_comb = {{1{p7_clipped__345_comb[8]}}, p7_clipped__345_comb} + 10'h001;
  assign p7_add_157877_comb = {{1{p7_clipped__346_comb[8]}}, p7_clipped__346_comb} + 10'h001;
  assign p7_add_157878_comb = {{1{p7_clipped__347_comb[8]}}, p7_clipped__347_comb} + 10'h001;
  assign p7_add_157879_comb = {{1{p7_clipped__348_comb[8]}}, p7_clipped__348_comb} + 10'h001;
  assign p7_add_157880_comb = {{1{p7_clipped__349_comb[8]}}, p7_clipped__349_comb} + 10'h001;
  assign p7_add_157881_comb = {{1{p7_clipped__350_comb[8]}}, p7_clipped__350_comb} + 10'h001;
  assign p7_add_157882_comb = {{1{p7_clipped__351_comb[8]}}, p7_clipped__351_comb} + 10'h001;
  assign p7_add_157883_comb = {{1{p7_clipped__352_comb[8]}}, p7_clipped__352_comb} + 10'h001;
  assign p7_add_157884_comb = {{1{p7_clipped__353_comb[8]}}, p7_clipped__353_comb} + 10'h001;
  assign p7_add_157885_comb = {{1{p7_clipped__354_comb[8]}}, p7_clipped__354_comb} + 10'h001;
  assign p7_add_157886_comb = {{1{p7_clipped__355_comb[8]}}, p7_clipped__355_comb} + 10'h001;
  assign p7_add_157887_comb = {{1{p7_clipped__356_comb[8]}}, p7_clipped__356_comb} + 10'h001;
  assign p7_add_157888_comb = {{1{p7_clipped__357_comb[8]}}, p7_clipped__357_comb} + 10'h001;
  assign p7_add_157889_comb = {{1{p7_clipped__358_comb[8]}}, p7_clipped__358_comb} + 10'h001;
  assign p7_add_157890_comb = {{1{p7_clipped__359_comb[8]}}, p7_clipped__359_comb} + 10'h001;
  assign p7_add_157891_comb = {{1{p7_clipped__360_comb[8]}}, p7_clipped__360_comb} + 10'h001;
  assign p7_add_157892_comb = {{1{p7_clipped__361_comb[8]}}, p7_clipped__361_comb} + 10'h001;
  assign p7_add_157893_comb = {{1{p7_clipped__362_comb[8]}}, p7_clipped__362_comb} + 10'h001;
  assign p7_add_157894_comb = {{1{p7_clipped__363_comb[8]}}, p7_clipped__363_comb} + 10'h001;
  assign p7_add_157895_comb = {{1{p7_clipped__364_comb[8]}}, p7_clipped__364_comb} + 10'h001;
  assign p7_add_157896_comb = {{1{p7_clipped__365_comb[8]}}, p7_clipped__365_comb} + 10'h001;
  assign p7_add_157897_comb = {{1{p7_clipped__366_comb[8]}}, p7_clipped__366_comb} + 10'h001;
  assign p7_add_157898_comb = {{1{p7_clipped__367_comb[8]}}, p7_clipped__367_comb} + 10'h001;
  assign p7_add_157907_comb = {{1{p7_clipped__376_comb[8]}}, p7_clipped__376_comb} + 10'h001;
  assign p7_add_157908_comb = {{1{p7_clipped__377_comb[8]}}, p7_clipped__377_comb} + 10'h001;
  assign p7_add_157909_comb = {{1{p7_clipped__378_comb[8]}}, p7_clipped__378_comb} + 10'h001;
  assign p7_add_157910_comb = {{1{p7_clipped__379_comb[8]}}, p7_clipped__379_comb} + 10'h001;
  assign p7_add_157911_comb = {{1{p7_clipped__380_comb[8]}}, p7_clipped__380_comb} + 10'h001;
  assign p7_add_157912_comb = {{1{p7_clipped__381_comb[8]}}, p7_clipped__381_comb} + 10'h001;
  assign p7_add_157913_comb = {{1{p7_clipped__382_comb[8]}}, p7_clipped__382_comb} + 10'h001;
  assign p7_add_157914_comb = {{1{p7_clipped__383_comb[8]}}, p7_clipped__383_comb} + 10'h001;
  assign p7_bit_slice_157917_comb = p7_add_157867_comb[9:8];
  assign p7_bit_slice_157918_comb = p7_add_157868_comb[9:8];
  assign p7_bit_slice_157919_comb = p7_add_157869_comb[9:8];
  assign p7_bit_slice_157920_comb = p7_add_157870_comb[9:8];
  assign p7_bit_slice_157921_comb = p7_add_157871_comb[9:8];
  assign p7_bit_slice_157922_comb = p7_add_157872_comb[9:8];
  assign p7_bit_slice_157923_comb = p7_add_157873_comb[9:8];
  assign p7_bit_slice_157924_comb = p7_add_157874_comb[9:8];
  assign p7_bit_slice_157925_comb = p7_add_157899_comb[9:8];
  assign p7_bit_slice_157926_comb = p7_add_157900_comb[9:8];
  assign p7_bit_slice_157927_comb = p7_add_157901_comb[9:8];
  assign p7_bit_slice_157928_comb = p7_add_157902_comb[9:8];
  assign p7_bit_slice_157929_comb = p7_add_157903_comb[9:8];
  assign p7_bit_slice_157930_comb = p7_add_157904_comb[9:8];
  assign p7_bit_slice_157931_comb = p7_add_157905_comb[9:8];
  assign p7_bit_slice_157932_comb = p7_add_157906_comb[9:8];
  assign p7_bit_slice_157939_comb = p7_add_157937_comb[0];
  assign p7_bit_slice_157940_comb = p7_add_157851_comb[7:1];
  assign p7_bit_slice_157941_comb = p7_add_157938_comb[0];
  assign p7_bit_slice_157942_comb = p7_add_157855_comb[7:1];
  assign p7_bit_slice_157943_comb = p7_add_157867_comb[7:1];
  assign p7_bit_slice_157944_comb = p7_add_157868_comb[7:1];
  assign p7_bit_slice_157945_comb = p7_add_157869_comb[7:1];
  assign p7_bit_slice_157946_comb = p7_add_157870_comb[7:1];
  assign p7_bit_slice_157947_comb = p7_add_157871_comb[7:1];
  assign p7_bit_slice_157948_comb = p7_add_157872_comb[7:1];
  assign p7_bit_slice_157949_comb = p7_add_157873_comb[7:1];
  assign p7_bit_slice_157950_comb = p7_add_157874_comb[7:1];
  assign p7_bit_slice_157951_comb = p7_add_157899_comb[7:1];
  assign p7_bit_slice_157952_comb = p7_add_157900_comb[7:1];
  assign p7_bit_slice_157953_comb = p7_add_157901_comb[7:1];
  assign p7_bit_slice_157954_comb = p7_add_157902_comb[7:1];
  assign p7_bit_slice_157955_comb = p7_add_157903_comb[7:1];
  assign p7_bit_slice_157956_comb = p7_add_157904_comb[7:1];
  assign p7_bit_slice_157957_comb = p7_add_157905_comb[7:1];
  assign p7_bit_slice_157958_comb = p7_add_157906_comb[7:1];
  assign p7_bit_slice_157959_comb = p7_add_157937_comb[1];
  assign p7_bit_slice_157960_comb = p7_add_157938_comb[1];

  // Registers for pipe stage 7:
  reg [9:0] p7_add_157852;
  reg [9:0] p7_add_157853;
  reg [9:0] p7_add_157854;
  reg [9:0] p7_add_157856;
  reg [9:0] p7_add_157857;
  reg [9:0] p7_add_157858;
  reg [9:0] p7_add_157859;
  reg [9:0] p7_add_157860;
  reg [9:0] p7_add_157861;
  reg [9:0] p7_add_157862;
  reg [9:0] p7_add_157863;
  reg [9:0] p7_add_157864;
  reg [9:0] p7_add_157865;
  reg [9:0] p7_add_157866;
  reg [9:0] p7_add_157875;
  reg [9:0] p7_add_157876;
  reg [9:0] p7_add_157877;
  reg [9:0] p7_add_157878;
  reg [9:0] p7_add_157879;
  reg [9:0] p7_add_157880;
  reg [9:0] p7_add_157881;
  reg [9:0] p7_add_157882;
  reg [9:0] p7_add_157883;
  reg [9:0] p7_add_157884;
  reg [9:0] p7_add_157885;
  reg [9:0] p7_add_157886;
  reg [9:0] p7_add_157887;
  reg [9:0] p7_add_157888;
  reg [9:0] p7_add_157889;
  reg [9:0] p7_add_157890;
  reg [9:0] p7_add_157891;
  reg [9:0] p7_add_157892;
  reg [9:0] p7_add_157893;
  reg [9:0] p7_add_157894;
  reg [9:0] p7_add_157895;
  reg [9:0] p7_add_157896;
  reg [9:0] p7_add_157897;
  reg [9:0] p7_add_157898;
  reg [9:0] p7_add_157907;
  reg [9:0] p7_add_157908;
  reg [9:0] p7_add_157909;
  reg [9:0] p7_add_157910;
  reg [9:0] p7_add_157911;
  reg [9:0] p7_add_157912;
  reg [9:0] p7_add_157913;
  reg [9:0] p7_add_157914;
  reg [1:0] p7_bit_slice_157917;
  reg [1:0] p7_bit_slice_157918;
  reg [1:0] p7_bit_slice_157919;
  reg [1:0] p7_bit_slice_157920;
  reg [1:0] p7_bit_slice_157921;
  reg [1:0] p7_bit_slice_157922;
  reg [1:0] p7_bit_slice_157923;
  reg [1:0] p7_bit_slice_157924;
  reg [1:0] p7_bit_slice_157925;
  reg [1:0] p7_bit_slice_157926;
  reg [1:0] p7_bit_slice_157927;
  reg [1:0] p7_bit_slice_157928;
  reg [1:0] p7_bit_slice_157929;
  reg [1:0] p7_bit_slice_157930;
  reg [1:0] p7_bit_slice_157931;
  reg [1:0] p7_bit_slice_157932;
  reg p7_bit_slice_157939;
  reg [6:0] p7_bit_slice_157940;
  reg p7_bit_slice_157941;
  reg [6:0] p7_bit_slice_157942;
  reg [6:0] p7_bit_slice_157943;
  reg [6:0] p7_bit_slice_157944;
  reg [6:0] p7_bit_slice_157945;
  reg [6:0] p7_bit_slice_157946;
  reg [6:0] p7_bit_slice_157947;
  reg [6:0] p7_bit_slice_157948;
  reg [6:0] p7_bit_slice_157949;
  reg [6:0] p7_bit_slice_157950;
  reg [6:0] p7_bit_slice_157951;
  reg [6:0] p7_bit_slice_157952;
  reg [6:0] p7_bit_slice_157953;
  reg [6:0] p7_bit_slice_157954;
  reg [6:0] p7_bit_slice_157955;
  reg [6:0] p7_bit_slice_157956;
  reg [6:0] p7_bit_slice_157957;
  reg [6:0] p7_bit_slice_157958;
  reg p7_bit_slice_157959;
  reg p7_bit_slice_157960;
  always @ (posedge clk) begin
    p7_add_157852 <= p7_add_157852_comb;
    p7_add_157853 <= p7_add_157853_comb;
    p7_add_157854 <= p7_add_157854_comb;
    p7_add_157856 <= p7_add_157856_comb;
    p7_add_157857 <= p7_add_157857_comb;
    p7_add_157858 <= p7_add_157858_comb;
    p7_add_157859 <= p7_add_157859_comb;
    p7_add_157860 <= p7_add_157860_comb;
    p7_add_157861 <= p7_add_157861_comb;
    p7_add_157862 <= p7_add_157862_comb;
    p7_add_157863 <= p7_add_157863_comb;
    p7_add_157864 <= p7_add_157864_comb;
    p7_add_157865 <= p7_add_157865_comb;
    p7_add_157866 <= p7_add_157866_comb;
    p7_add_157875 <= p7_add_157875_comb;
    p7_add_157876 <= p7_add_157876_comb;
    p7_add_157877 <= p7_add_157877_comb;
    p7_add_157878 <= p7_add_157878_comb;
    p7_add_157879 <= p7_add_157879_comb;
    p7_add_157880 <= p7_add_157880_comb;
    p7_add_157881 <= p7_add_157881_comb;
    p7_add_157882 <= p7_add_157882_comb;
    p7_add_157883 <= p7_add_157883_comb;
    p7_add_157884 <= p7_add_157884_comb;
    p7_add_157885 <= p7_add_157885_comb;
    p7_add_157886 <= p7_add_157886_comb;
    p7_add_157887 <= p7_add_157887_comb;
    p7_add_157888 <= p7_add_157888_comb;
    p7_add_157889 <= p7_add_157889_comb;
    p7_add_157890 <= p7_add_157890_comb;
    p7_add_157891 <= p7_add_157891_comb;
    p7_add_157892 <= p7_add_157892_comb;
    p7_add_157893 <= p7_add_157893_comb;
    p7_add_157894 <= p7_add_157894_comb;
    p7_add_157895 <= p7_add_157895_comb;
    p7_add_157896 <= p7_add_157896_comb;
    p7_add_157897 <= p7_add_157897_comb;
    p7_add_157898 <= p7_add_157898_comb;
    p7_add_157907 <= p7_add_157907_comb;
    p7_add_157908 <= p7_add_157908_comb;
    p7_add_157909 <= p7_add_157909_comb;
    p7_add_157910 <= p7_add_157910_comb;
    p7_add_157911 <= p7_add_157911_comb;
    p7_add_157912 <= p7_add_157912_comb;
    p7_add_157913 <= p7_add_157913_comb;
    p7_add_157914 <= p7_add_157914_comb;
    p7_bit_slice_157917 <= p7_bit_slice_157917_comb;
    p7_bit_slice_157918 <= p7_bit_slice_157918_comb;
    p7_bit_slice_157919 <= p7_bit_slice_157919_comb;
    p7_bit_slice_157920 <= p7_bit_slice_157920_comb;
    p7_bit_slice_157921 <= p7_bit_slice_157921_comb;
    p7_bit_slice_157922 <= p7_bit_slice_157922_comb;
    p7_bit_slice_157923 <= p7_bit_slice_157923_comb;
    p7_bit_slice_157924 <= p7_bit_slice_157924_comb;
    p7_bit_slice_157925 <= p7_bit_slice_157925_comb;
    p7_bit_slice_157926 <= p7_bit_slice_157926_comb;
    p7_bit_slice_157927 <= p7_bit_slice_157927_comb;
    p7_bit_slice_157928 <= p7_bit_slice_157928_comb;
    p7_bit_slice_157929 <= p7_bit_slice_157929_comb;
    p7_bit_slice_157930 <= p7_bit_slice_157930_comb;
    p7_bit_slice_157931 <= p7_bit_slice_157931_comb;
    p7_bit_slice_157932 <= p7_bit_slice_157932_comb;
    p7_bit_slice_157939 <= p7_bit_slice_157939_comb;
    p7_bit_slice_157940 <= p7_bit_slice_157940_comb;
    p7_bit_slice_157941 <= p7_bit_slice_157941_comb;
    p7_bit_slice_157942 <= p7_bit_slice_157942_comb;
    p7_bit_slice_157943 <= p7_bit_slice_157943_comb;
    p7_bit_slice_157944 <= p7_bit_slice_157944_comb;
    p7_bit_slice_157945 <= p7_bit_slice_157945_comb;
    p7_bit_slice_157946 <= p7_bit_slice_157946_comb;
    p7_bit_slice_157947 <= p7_bit_slice_157947_comb;
    p7_bit_slice_157948 <= p7_bit_slice_157948_comb;
    p7_bit_slice_157949 <= p7_bit_slice_157949_comb;
    p7_bit_slice_157950 <= p7_bit_slice_157950_comb;
    p7_bit_slice_157951 <= p7_bit_slice_157951_comb;
    p7_bit_slice_157952 <= p7_bit_slice_157952_comb;
    p7_bit_slice_157953 <= p7_bit_slice_157953_comb;
    p7_bit_slice_157954 <= p7_bit_slice_157954_comb;
    p7_bit_slice_157955 <= p7_bit_slice_157955_comb;
    p7_bit_slice_157956 <= p7_bit_slice_157956_comb;
    p7_bit_slice_157957 <= p7_bit_slice_157957_comb;
    p7_bit_slice_157958 <= p7_bit_slice_157958_comb;
    p7_bit_slice_157959 <= p7_bit_slice_157959_comb;
    p7_bit_slice_157960 <= p7_bit_slice_157960_comb;
  end

  // ===== Pipe stage 8:
  wire [1:0] p8_bit_slice_158129_comb;
  wire [1:0] p8_bit_slice_158130_comb;
  wire [1:0] p8_bit_slice_158131_comb;
  wire [1:0] p8_bit_slice_158132_comb;
  wire [1:0] p8_bit_slice_158133_comb;
  wire [1:0] p8_bit_slice_158134_comb;
  wire [1:0] p8_bit_slice_158135_comb;
  wire [1:0] p8_bit_slice_158136_comb;
  wire [1:0] p8_bit_slice_158137_comb;
  wire [1:0] p8_bit_slice_158138_comb;
  wire [1:0] p8_bit_slice_158139_comb;
  wire [1:0] p8_bit_slice_158140_comb;
  wire [1:0] p8_bit_slice_158141_comb;
  wire [1:0] p8_bit_slice_158142_comb;
  wire [1:0] p8_bit_slice_158143_comb;
  wire [1:0] p8_bit_slice_158144_comb;
  wire [1:0] p8_bit_slice_158145_comb;
  wire [1:0] p8_bit_slice_158146_comb;
  wire [1:0] p8_bit_slice_158147_comb;
  wire [1:0] p8_bit_slice_158148_comb;
  wire [1:0] p8_bit_slice_158149_comb;
  wire [1:0] p8_bit_slice_158150_comb;
  wire [1:0] p8_bit_slice_158151_comb;
  wire [1:0] p8_bit_slice_158152_comb;
  wire [1:0] p8_bit_slice_158153_comb;
  wire [1:0] p8_bit_slice_158154_comb;
  wire [1:0] p8_bit_slice_158155_comb;
  wire [1:0] p8_bit_slice_158156_comb;
  wire [1:0] p8_bit_slice_158157_comb;
  wire [1:0] p8_bit_slice_158158_comb;
  wire [1:0] p8_bit_slice_158159_comb;
  wire [1:0] p8_bit_slice_158160_comb;
  wire [1:0] p8_bit_slice_158161_comb;
  wire [1:0] p8_bit_slice_158162_comb;
  wire [1:0] p8_bit_slice_158163_comb;
  wire [1:0] p8_bit_slice_158164_comb;
  wire [1:0] p8_bit_slice_158165_comb;
  wire [1:0] p8_bit_slice_158166_comb;
  wire [1:0] p8_bit_slice_158167_comb;
  wire [1:0] p8_bit_slice_158168_comb;
  wire [1:0] p8_bit_slice_158169_comb;
  wire [1:0] p8_bit_slice_158170_comb;
  wire [1:0] p8_bit_slice_158171_comb;
  wire [1:0] p8_bit_slice_158172_comb;
  wire [1:0] p8_bit_slice_158173_comb;
  wire [1:0] p8_bit_slice_158174_comb;
  wire [2:0] p8_add_158299_comb;
  wire [2:0] p8_add_158300_comb;
  wire [2:0] p8_add_158301_comb;
  wire [2:0] p8_add_158302_comb;
  wire [2:0] p8_add_158303_comb;
  wire [2:0] p8_add_158304_comb;
  wire [2:0] p8_add_158305_comb;
  wire [2:0] p8_add_158306_comb;
  wire [2:0] p8_add_158307_comb;
  wire [2:0] p8_add_158308_comb;
  wire [2:0] p8_add_158309_comb;
  wire [2:0] p8_add_158310_comb;
  wire [2:0] p8_add_158311_comb;
  wire [2:0] p8_add_158312_comb;
  wire [2:0] p8_add_158313_comb;
  wire [2:0] p8_add_158314_comb;
  wire [2:0] p8_add_158315_comb;
  wire [2:0] p8_add_158316_comb;
  wire [2:0] p8_add_158317_comb;
  wire [2:0] p8_add_158318_comb;
  wire [2:0] p8_add_158319_comb;
  wire [2:0] p8_add_158320_comb;
  wire [2:0] p8_add_158321_comb;
  wire [2:0] p8_add_158322_comb;
  wire [2:0] p8_add_158323_comb;
  wire [2:0] p8_add_158324_comb;
  wire [2:0] p8_add_158325_comb;
  wire [2:0] p8_add_158326_comb;
  wire [2:0] p8_add_158327_comb;
  wire [2:0] p8_add_158328_comb;
  wire [2:0] p8_add_158329_comb;
  wire [2:0] p8_add_158330_comb;
  wire [2:0] p8_add_158331_comb;
  wire [2:0] p8_add_158332_comb;
  wire [2:0] p8_add_158333_comb;
  wire [2:0] p8_add_158334_comb;
  wire [2:0] p8_add_158335_comb;
  wire [2:0] p8_add_158336_comb;
  wire [2:0] p8_add_158337_comb;
  wire [2:0] p8_add_158338_comb;
  wire [2:0] p8_add_158339_comb;
  wire [2:0] p8_add_158340_comb;
  wire [2:0] p8_add_158341_comb;
  wire [2:0] p8_add_158342_comb;
  wire [2:0] p8_add_158343_comb;
  wire [2:0] p8_add_158344_comb;
  wire [2:0] p8_add_158345_comb;
  wire [2:0] p8_add_158346_comb;
  wire [2:0] p8_add_158347_comb;
  wire [2:0] p8_add_158348_comb;
  wire [2:0] p8_add_158349_comb;
  wire [2:0] p8_add_158350_comb;
  wire [2:0] p8_add_158351_comb;
  wire [2:0] p8_add_158352_comb;
  wire [2:0] p8_add_158353_comb;
  wire [2:0] p8_add_158354_comb;
  wire [2:0] p8_add_158355_comb;
  wire [2:0] p8_add_158356_comb;
  wire [2:0] p8_add_158357_comb;
  wire [2:0] p8_add_158358_comb;
  wire [2:0] p8_add_158359_comb;
  wire [2:0] p8_add_158360_comb;
  wire [7:0] p8_clipped__136_comb;
  wire [7:0] p8_clipped__152_comb;
  wire [7:0] p8_clipped__168_comb;
  wire [7:0] p8_clipped__184_comb;
  wire [7:0] p8_clipped__200_comb;
  wire [7:0] p8_clipped__216_comb;
  wire [7:0] p8_clipped__232_comb;
  wire [7:0] p8_clipped__248_comb;
  wire [7:0] p8_clipped__137_comb;
  wire [7:0] p8_clipped__153_comb;
  wire [7:0] p8_clipped__169_comb;
  wire [7:0] p8_clipped__185_comb;
  wire [7:0] p8_clipped__201_comb;
  wire [7:0] p8_clipped__217_comb;
  wire [7:0] p8_clipped__233_comb;
  wire [7:0] p8_clipped__249_comb;
  wire [7:0] p8_clipped__138_comb;
  wire [7:0] p8_clipped__154_comb;
  wire [7:0] p8_clipped__170_comb;
  wire [7:0] p8_clipped__186_comb;
  wire [7:0] p8_clipped__202_comb;
  wire [7:0] p8_clipped__218_comb;
  wire [7:0] p8_clipped__234_comb;
  wire [7:0] p8_clipped__250_comb;
  wire [7:0] p8_clipped__139_comb;
  wire [7:0] p8_clipped__155_comb;
  wire [7:0] p8_clipped__171_comb;
  wire [7:0] p8_clipped__187_comb;
  wire [7:0] p8_clipped__203_comb;
  wire [7:0] p8_clipped__219_comb;
  wire [7:0] p8_clipped__235_comb;
  wire [7:0] p8_clipped__251_comb;
  wire [7:0] p8_clipped__140_comb;
  wire [7:0] p8_clipped__156_comb;
  wire [7:0] p8_clipped__172_comb;
  wire [7:0] p8_clipped__188_comb;
  wire [7:0] p8_clipped__204_comb;
  wire [7:0] p8_clipped__220_comb;
  wire [7:0] p8_clipped__236_comb;
  wire [7:0] p8_clipped__252_comb;
  wire [7:0] p8_clipped__141_comb;
  wire [7:0] p8_clipped__157_comb;
  wire [7:0] p8_clipped__173_comb;
  wire [7:0] p8_clipped__189_comb;
  wire [7:0] p8_clipped__205_comb;
  wire [7:0] p8_clipped__221_comb;
  wire [7:0] p8_clipped__237_comb;
  wire [7:0] p8_clipped__253_comb;
  wire [7:0] p8_clipped__142_comb;
  wire [7:0] p8_clipped__158_comb;
  wire [7:0] p8_clipped__174_comb;
  wire [7:0] p8_clipped__190_comb;
  wire [7:0] p8_clipped__206_comb;
  wire [7:0] p8_clipped__222_comb;
  wire [7:0] p8_clipped__238_comb;
  wire [7:0] p8_clipped__254_comb;
  wire [7:0] p8_clipped__143_comb;
  wire [7:0] p8_clipped__159_comb;
  wire [7:0] p8_clipped__175_comb;
  wire [7:0] p8_clipped__191_comb;
  wire [7:0] p8_clipped__207_comb;
  wire [7:0] p8_clipped__223_comb;
  wire [7:0] p8_clipped__239_comb;
  wire [7:0] p8_clipped__255_comb;
  wire [7:0] p8_array_158723_comb[0:7];
  wire [7:0] p8_array_158724_comb[0:7];
  wire [7:0] p8_array_158725_comb[0:7];
  wire [7:0] p8_array_158726_comb[0:7];
  wire [7:0] p8_array_158727_comb[0:7];
  wire [7:0] p8_array_158728_comb[0:7];
  wire [7:0] p8_array_158729_comb[0:7];
  wire [7:0] p8_array_158730_comb[0:7];
  wire [7:0] p8_col_transformed_comb[0:7][0:7];
  assign p8_bit_slice_158129_comb = p7_add_157852[9:8];
  assign p8_bit_slice_158130_comb = p7_add_157853[9:8];
  assign p8_bit_slice_158131_comb = p7_add_157854[9:8];
  assign p8_bit_slice_158132_comb = p7_add_157856[9:8];
  assign p8_bit_slice_158133_comb = p7_add_157857[9:8];
  assign p8_bit_slice_158134_comb = p7_add_157858[9:8];
  assign p8_bit_slice_158135_comb = p7_add_157859[9:8];
  assign p8_bit_slice_158136_comb = p7_add_157860[9:8];
  assign p8_bit_slice_158137_comb = p7_add_157861[9:8];
  assign p8_bit_slice_158138_comb = p7_add_157862[9:8];
  assign p8_bit_slice_158139_comb = p7_add_157863[9:8];
  assign p8_bit_slice_158140_comb = p7_add_157864[9:8];
  assign p8_bit_slice_158141_comb = p7_add_157865[9:8];
  assign p8_bit_slice_158142_comb = p7_add_157866[9:8];
  assign p8_bit_slice_158143_comb = p7_add_157875[9:8];
  assign p8_bit_slice_158144_comb = p7_add_157876[9:8];
  assign p8_bit_slice_158145_comb = p7_add_157877[9:8];
  assign p8_bit_slice_158146_comb = p7_add_157878[9:8];
  assign p8_bit_slice_158147_comb = p7_add_157879[9:8];
  assign p8_bit_slice_158148_comb = p7_add_157880[9:8];
  assign p8_bit_slice_158149_comb = p7_add_157881[9:8];
  assign p8_bit_slice_158150_comb = p7_add_157882[9:8];
  assign p8_bit_slice_158151_comb = p7_add_157883[9:8];
  assign p8_bit_slice_158152_comb = p7_add_157884[9:8];
  assign p8_bit_slice_158153_comb = p7_add_157885[9:8];
  assign p8_bit_slice_158154_comb = p7_add_157886[9:8];
  assign p8_bit_slice_158155_comb = p7_add_157887[9:8];
  assign p8_bit_slice_158156_comb = p7_add_157888[9:8];
  assign p8_bit_slice_158157_comb = p7_add_157889[9:8];
  assign p8_bit_slice_158158_comb = p7_add_157890[9:8];
  assign p8_bit_slice_158159_comb = p7_add_157891[9:8];
  assign p8_bit_slice_158160_comb = p7_add_157892[9:8];
  assign p8_bit_slice_158161_comb = p7_add_157893[9:8];
  assign p8_bit_slice_158162_comb = p7_add_157894[9:8];
  assign p8_bit_slice_158163_comb = p7_add_157895[9:8];
  assign p8_bit_slice_158164_comb = p7_add_157896[9:8];
  assign p8_bit_slice_158165_comb = p7_add_157897[9:8];
  assign p8_bit_slice_158166_comb = p7_add_157898[9:8];
  assign p8_bit_slice_158167_comb = p7_add_157907[9:8];
  assign p8_bit_slice_158168_comb = p7_add_157908[9:8];
  assign p8_bit_slice_158169_comb = p7_add_157909[9:8];
  assign p8_bit_slice_158170_comb = p7_add_157910[9:8];
  assign p8_bit_slice_158171_comb = p7_add_157911[9:8];
  assign p8_bit_slice_158172_comb = p7_add_157912[9:8];
  assign p8_bit_slice_158173_comb = p7_add_157913[9:8];
  assign p8_bit_slice_158174_comb = p7_add_157914[9:8];
  assign p8_add_158299_comb = {{1{p8_bit_slice_158129_comb[1]}}, p8_bit_slice_158129_comb} + 3'h1;
  assign p8_add_158300_comb = {{1{p8_bit_slice_158130_comb[1]}}, p8_bit_slice_158130_comb} + 3'h1;
  assign p8_add_158301_comb = {{1{p8_bit_slice_158131_comb[1]}}, p8_bit_slice_158131_comb} + 3'h1;
  assign p8_add_158302_comb = {{1{p8_bit_slice_158132_comb[1]}}, p8_bit_slice_158132_comb} + 3'h1;
  assign p8_add_158303_comb = {{1{p8_bit_slice_158133_comb[1]}}, p8_bit_slice_158133_comb} + 3'h1;
  assign p8_add_158304_comb = {{1{p8_bit_slice_158134_comb[1]}}, p8_bit_slice_158134_comb} + 3'h1;
  assign p8_add_158305_comb = {{1{p8_bit_slice_158135_comb[1]}}, p8_bit_slice_158135_comb} + 3'h1;
  assign p8_add_158306_comb = {{1{p8_bit_slice_158136_comb[1]}}, p8_bit_slice_158136_comb} + 3'h1;
  assign p8_add_158307_comb = {{1{p8_bit_slice_158137_comb[1]}}, p8_bit_slice_158137_comb} + 3'h1;
  assign p8_add_158308_comb = {{1{p8_bit_slice_158138_comb[1]}}, p8_bit_slice_158138_comb} + 3'h1;
  assign p8_add_158309_comb = {{1{p8_bit_slice_158139_comb[1]}}, p8_bit_slice_158139_comb} + 3'h1;
  assign p8_add_158310_comb = {{1{p8_bit_slice_158140_comb[1]}}, p8_bit_slice_158140_comb} + 3'h1;
  assign p8_add_158311_comb = {{1{p8_bit_slice_158141_comb[1]}}, p8_bit_slice_158141_comb} + 3'h1;
  assign p8_add_158312_comb = {{1{p8_bit_slice_158142_comb[1]}}, p8_bit_slice_158142_comb} + 3'h1;
  assign p8_add_158313_comb = {{1{p7_bit_slice_157917[1]}}, p7_bit_slice_157917} + 3'h1;
  assign p8_add_158314_comb = {{1{p7_bit_slice_157918[1]}}, p7_bit_slice_157918} + 3'h1;
  assign p8_add_158315_comb = {{1{p7_bit_slice_157919[1]}}, p7_bit_slice_157919} + 3'h1;
  assign p8_add_158316_comb = {{1{p7_bit_slice_157920[1]}}, p7_bit_slice_157920} + 3'h1;
  assign p8_add_158317_comb = {{1{p7_bit_slice_157921[1]}}, p7_bit_slice_157921} + 3'h1;
  assign p8_add_158318_comb = {{1{p7_bit_slice_157922[1]}}, p7_bit_slice_157922} + 3'h1;
  assign p8_add_158319_comb = {{1{p7_bit_slice_157923[1]}}, p7_bit_slice_157923} + 3'h1;
  assign p8_add_158320_comb = {{1{p7_bit_slice_157924[1]}}, p7_bit_slice_157924} + 3'h1;
  assign p8_add_158321_comb = {{1{p8_bit_slice_158143_comb[1]}}, p8_bit_slice_158143_comb} + 3'h1;
  assign p8_add_158322_comb = {{1{p8_bit_slice_158144_comb[1]}}, p8_bit_slice_158144_comb} + 3'h1;
  assign p8_add_158323_comb = {{1{p8_bit_slice_158145_comb[1]}}, p8_bit_slice_158145_comb} + 3'h1;
  assign p8_add_158324_comb = {{1{p8_bit_slice_158146_comb[1]}}, p8_bit_slice_158146_comb} + 3'h1;
  assign p8_add_158325_comb = {{1{p8_bit_slice_158147_comb[1]}}, p8_bit_slice_158147_comb} + 3'h1;
  assign p8_add_158326_comb = {{1{p8_bit_slice_158148_comb[1]}}, p8_bit_slice_158148_comb} + 3'h1;
  assign p8_add_158327_comb = {{1{p8_bit_slice_158149_comb[1]}}, p8_bit_slice_158149_comb} + 3'h1;
  assign p8_add_158328_comb = {{1{p8_bit_slice_158150_comb[1]}}, p8_bit_slice_158150_comb} + 3'h1;
  assign p8_add_158329_comb = {{1{p8_bit_slice_158151_comb[1]}}, p8_bit_slice_158151_comb} + 3'h1;
  assign p8_add_158330_comb = {{1{p8_bit_slice_158152_comb[1]}}, p8_bit_slice_158152_comb} + 3'h1;
  assign p8_add_158331_comb = {{1{p8_bit_slice_158153_comb[1]}}, p8_bit_slice_158153_comb} + 3'h1;
  assign p8_add_158332_comb = {{1{p8_bit_slice_158154_comb[1]}}, p8_bit_slice_158154_comb} + 3'h1;
  assign p8_add_158333_comb = {{1{p8_bit_slice_158155_comb[1]}}, p8_bit_slice_158155_comb} + 3'h1;
  assign p8_add_158334_comb = {{1{p8_bit_slice_158156_comb[1]}}, p8_bit_slice_158156_comb} + 3'h1;
  assign p8_add_158335_comb = {{1{p8_bit_slice_158157_comb[1]}}, p8_bit_slice_158157_comb} + 3'h1;
  assign p8_add_158336_comb = {{1{p8_bit_slice_158158_comb[1]}}, p8_bit_slice_158158_comb} + 3'h1;
  assign p8_add_158337_comb = {{1{p8_bit_slice_158159_comb[1]}}, p8_bit_slice_158159_comb} + 3'h1;
  assign p8_add_158338_comb = {{1{p8_bit_slice_158160_comb[1]}}, p8_bit_slice_158160_comb} + 3'h1;
  assign p8_add_158339_comb = {{1{p8_bit_slice_158161_comb[1]}}, p8_bit_slice_158161_comb} + 3'h1;
  assign p8_add_158340_comb = {{1{p8_bit_slice_158162_comb[1]}}, p8_bit_slice_158162_comb} + 3'h1;
  assign p8_add_158341_comb = {{1{p8_bit_slice_158163_comb[1]}}, p8_bit_slice_158163_comb} + 3'h1;
  assign p8_add_158342_comb = {{1{p8_bit_slice_158164_comb[1]}}, p8_bit_slice_158164_comb} + 3'h1;
  assign p8_add_158343_comb = {{1{p8_bit_slice_158165_comb[1]}}, p8_bit_slice_158165_comb} + 3'h1;
  assign p8_add_158344_comb = {{1{p8_bit_slice_158166_comb[1]}}, p8_bit_slice_158166_comb} + 3'h1;
  assign p8_add_158345_comb = {{1{p7_bit_slice_157925[1]}}, p7_bit_slice_157925} + 3'h1;
  assign p8_add_158346_comb = {{1{p7_bit_slice_157926[1]}}, p7_bit_slice_157926} + 3'h1;
  assign p8_add_158347_comb = {{1{p7_bit_slice_157927[1]}}, p7_bit_slice_157927} + 3'h1;
  assign p8_add_158348_comb = {{1{p7_bit_slice_157928[1]}}, p7_bit_slice_157928} + 3'h1;
  assign p8_add_158349_comb = {{1{p7_bit_slice_157929[1]}}, p7_bit_slice_157929} + 3'h1;
  assign p8_add_158350_comb = {{1{p7_bit_slice_157930[1]}}, p7_bit_slice_157930} + 3'h1;
  assign p8_add_158351_comb = {{1{p7_bit_slice_157931[1]}}, p7_bit_slice_157931} + 3'h1;
  assign p8_add_158352_comb = {{1{p7_bit_slice_157932[1]}}, p7_bit_slice_157932} + 3'h1;
  assign p8_add_158353_comb = {{1{p8_bit_slice_158167_comb[1]}}, p8_bit_slice_158167_comb} + 3'h1;
  assign p8_add_158354_comb = {{1{p8_bit_slice_158168_comb[1]}}, p8_bit_slice_158168_comb} + 3'h1;
  assign p8_add_158355_comb = {{1{p8_bit_slice_158169_comb[1]}}, p8_bit_slice_158169_comb} + 3'h1;
  assign p8_add_158356_comb = {{1{p8_bit_slice_158170_comb[1]}}, p8_bit_slice_158170_comb} + 3'h1;
  assign p8_add_158357_comb = {{1{p8_bit_slice_158171_comb[1]}}, p8_bit_slice_158171_comb} + 3'h1;
  assign p8_add_158358_comb = {{1{p8_bit_slice_158172_comb[1]}}, p8_bit_slice_158172_comb} + 3'h1;
  assign p8_add_158359_comb = {{1{p8_bit_slice_158173_comb[1]}}, p8_bit_slice_158173_comb} + 3'h1;
  assign p8_add_158360_comb = {{1{p8_bit_slice_158174_comb[1]}}, p8_bit_slice_158174_comb} + 3'h1;
  assign p8_clipped__136_comb = p7_bit_slice_157959 ? 8'hff : {p7_bit_slice_157939, p7_bit_slice_157940};
  assign p8_clipped__152_comb = p8_add_158299_comb[1] ? 8'hff : {p8_add_158299_comb[0], p7_add_157852[7:1]};
  assign p8_clipped__168_comb = p8_add_158300_comb[1] ? 8'hff : {p8_add_158300_comb[0], p7_add_157853[7:1]};
  assign p8_clipped__184_comb = p8_add_158301_comb[1] ? 8'hff : {p8_add_158301_comb[0], p7_add_157854[7:1]};
  assign p8_clipped__200_comb = p7_bit_slice_157960 ? 8'hff : {p7_bit_slice_157941, p7_bit_slice_157942};
  assign p8_clipped__216_comb = p8_add_158302_comb[1] ? 8'hff : {p8_add_158302_comb[0], p7_add_157856[7:1]};
  assign p8_clipped__232_comb = p8_add_158303_comb[1] ? 8'hff : {p8_add_158303_comb[0], p7_add_157857[7:1]};
  assign p8_clipped__248_comb = p8_add_158304_comb[1] ? 8'hff : {p8_add_158304_comb[0], p7_add_157858[7:1]};
  assign p8_clipped__137_comb = p8_add_158305_comb[1] ? 8'hff : {p8_add_158305_comb[0], p7_add_157859[7:1]};
  assign p8_clipped__153_comb = p8_add_158306_comb[1] ? 8'hff : {p8_add_158306_comb[0], p7_add_157860[7:1]};
  assign p8_clipped__169_comb = p8_add_158307_comb[1] ? 8'hff : {p8_add_158307_comb[0], p7_add_157861[7:1]};
  assign p8_clipped__185_comb = p8_add_158308_comb[1] ? 8'hff : {p8_add_158308_comb[0], p7_add_157862[7:1]};
  assign p8_clipped__201_comb = p8_add_158309_comb[1] ? 8'hff : {p8_add_158309_comb[0], p7_add_157863[7:1]};
  assign p8_clipped__217_comb = p8_add_158310_comb[1] ? 8'hff : {p8_add_158310_comb[0], p7_add_157864[7:1]};
  assign p8_clipped__233_comb = p8_add_158311_comb[1] ? 8'hff : {p8_add_158311_comb[0], p7_add_157865[7:1]};
  assign p8_clipped__249_comb = p8_add_158312_comb[1] ? 8'hff : {p8_add_158312_comb[0], p7_add_157866[7:1]};
  assign p8_clipped__138_comb = p8_add_158313_comb[1] ? 8'hff : {p8_add_158313_comb[0], p7_bit_slice_157943};
  assign p8_clipped__154_comb = p8_add_158314_comb[1] ? 8'hff : {p8_add_158314_comb[0], p7_bit_slice_157944};
  assign p8_clipped__170_comb = p8_add_158315_comb[1] ? 8'hff : {p8_add_158315_comb[0], p7_bit_slice_157945};
  assign p8_clipped__186_comb = p8_add_158316_comb[1] ? 8'hff : {p8_add_158316_comb[0], p7_bit_slice_157946};
  assign p8_clipped__202_comb = p8_add_158317_comb[1] ? 8'hff : {p8_add_158317_comb[0], p7_bit_slice_157947};
  assign p8_clipped__218_comb = p8_add_158318_comb[1] ? 8'hff : {p8_add_158318_comb[0], p7_bit_slice_157948};
  assign p8_clipped__234_comb = p8_add_158319_comb[1] ? 8'hff : {p8_add_158319_comb[0], p7_bit_slice_157949};
  assign p8_clipped__250_comb = p8_add_158320_comb[1] ? 8'hff : {p8_add_158320_comb[0], p7_bit_slice_157950};
  assign p8_clipped__139_comb = p8_add_158321_comb[1] ? 8'hff : {p8_add_158321_comb[0], p7_add_157875[7:1]};
  assign p8_clipped__155_comb = p8_add_158322_comb[1] ? 8'hff : {p8_add_158322_comb[0], p7_add_157876[7:1]};
  assign p8_clipped__171_comb = p8_add_158323_comb[1] ? 8'hff : {p8_add_158323_comb[0], p7_add_157877[7:1]};
  assign p8_clipped__187_comb = p8_add_158324_comb[1] ? 8'hff : {p8_add_158324_comb[0], p7_add_157878[7:1]};
  assign p8_clipped__203_comb = p8_add_158325_comb[1] ? 8'hff : {p8_add_158325_comb[0], p7_add_157879[7:1]};
  assign p8_clipped__219_comb = p8_add_158326_comb[1] ? 8'hff : {p8_add_158326_comb[0], p7_add_157880[7:1]};
  assign p8_clipped__235_comb = p8_add_158327_comb[1] ? 8'hff : {p8_add_158327_comb[0], p7_add_157881[7:1]};
  assign p8_clipped__251_comb = p8_add_158328_comb[1] ? 8'hff : {p8_add_158328_comb[0], p7_add_157882[7:1]};
  assign p8_clipped__140_comb = p8_add_158329_comb[1] ? 8'hff : {p8_add_158329_comb[0], p7_add_157883[7:1]};
  assign p8_clipped__156_comb = p8_add_158330_comb[1] ? 8'hff : {p8_add_158330_comb[0], p7_add_157884[7:1]};
  assign p8_clipped__172_comb = p8_add_158331_comb[1] ? 8'hff : {p8_add_158331_comb[0], p7_add_157885[7:1]};
  assign p8_clipped__188_comb = p8_add_158332_comb[1] ? 8'hff : {p8_add_158332_comb[0], p7_add_157886[7:1]};
  assign p8_clipped__204_comb = p8_add_158333_comb[1] ? 8'hff : {p8_add_158333_comb[0], p7_add_157887[7:1]};
  assign p8_clipped__220_comb = p8_add_158334_comb[1] ? 8'hff : {p8_add_158334_comb[0], p7_add_157888[7:1]};
  assign p8_clipped__236_comb = p8_add_158335_comb[1] ? 8'hff : {p8_add_158335_comb[0], p7_add_157889[7:1]};
  assign p8_clipped__252_comb = p8_add_158336_comb[1] ? 8'hff : {p8_add_158336_comb[0], p7_add_157890[7:1]};
  assign p8_clipped__141_comb = p8_add_158337_comb[1] ? 8'hff : {p8_add_158337_comb[0], p7_add_157891[7:1]};
  assign p8_clipped__157_comb = p8_add_158338_comb[1] ? 8'hff : {p8_add_158338_comb[0], p7_add_157892[7:1]};
  assign p8_clipped__173_comb = p8_add_158339_comb[1] ? 8'hff : {p8_add_158339_comb[0], p7_add_157893[7:1]};
  assign p8_clipped__189_comb = p8_add_158340_comb[1] ? 8'hff : {p8_add_158340_comb[0], p7_add_157894[7:1]};
  assign p8_clipped__205_comb = p8_add_158341_comb[1] ? 8'hff : {p8_add_158341_comb[0], p7_add_157895[7:1]};
  assign p8_clipped__221_comb = p8_add_158342_comb[1] ? 8'hff : {p8_add_158342_comb[0], p7_add_157896[7:1]};
  assign p8_clipped__237_comb = p8_add_158343_comb[1] ? 8'hff : {p8_add_158343_comb[0], p7_add_157897[7:1]};
  assign p8_clipped__253_comb = p8_add_158344_comb[1] ? 8'hff : {p8_add_158344_comb[0], p7_add_157898[7:1]};
  assign p8_clipped__142_comb = p8_add_158345_comb[1] ? 8'hff : {p8_add_158345_comb[0], p7_bit_slice_157951};
  assign p8_clipped__158_comb = p8_add_158346_comb[1] ? 8'hff : {p8_add_158346_comb[0], p7_bit_slice_157952};
  assign p8_clipped__174_comb = p8_add_158347_comb[1] ? 8'hff : {p8_add_158347_comb[0], p7_bit_slice_157953};
  assign p8_clipped__190_comb = p8_add_158348_comb[1] ? 8'hff : {p8_add_158348_comb[0], p7_bit_slice_157954};
  assign p8_clipped__206_comb = p8_add_158349_comb[1] ? 8'hff : {p8_add_158349_comb[0], p7_bit_slice_157955};
  assign p8_clipped__222_comb = p8_add_158350_comb[1] ? 8'hff : {p8_add_158350_comb[0], p7_bit_slice_157956};
  assign p8_clipped__238_comb = p8_add_158351_comb[1] ? 8'hff : {p8_add_158351_comb[0], p7_bit_slice_157957};
  assign p8_clipped__254_comb = p8_add_158352_comb[1] ? 8'hff : {p8_add_158352_comb[0], p7_bit_slice_157958};
  assign p8_clipped__143_comb = p8_add_158353_comb[1] ? 8'hff : {p8_add_158353_comb[0], p7_add_157907[7:1]};
  assign p8_clipped__159_comb = p8_add_158354_comb[1] ? 8'hff : {p8_add_158354_comb[0], p7_add_157908[7:1]};
  assign p8_clipped__175_comb = p8_add_158355_comb[1] ? 8'hff : {p8_add_158355_comb[0], p7_add_157909[7:1]};
  assign p8_clipped__191_comb = p8_add_158356_comb[1] ? 8'hff : {p8_add_158356_comb[0], p7_add_157910[7:1]};
  assign p8_clipped__207_comb = p8_add_158357_comb[1] ? 8'hff : {p8_add_158357_comb[0], p7_add_157911[7:1]};
  assign p8_clipped__223_comb = p8_add_158358_comb[1] ? 8'hff : {p8_add_158358_comb[0], p7_add_157912[7:1]};
  assign p8_clipped__239_comb = p8_add_158359_comb[1] ? 8'hff : {p8_add_158359_comb[0], p7_add_157913[7:1]};
  assign p8_clipped__255_comb = p8_add_158360_comb[1] ? 8'hff : {p8_add_158360_comb[0], p7_add_157914[7:1]};
  assign p8_array_158723_comb[0] = p8_clipped__136_comb;
  assign p8_array_158723_comb[1] = p8_clipped__152_comb;
  assign p8_array_158723_comb[2] = p8_clipped__168_comb;
  assign p8_array_158723_comb[3] = p8_clipped__184_comb;
  assign p8_array_158723_comb[4] = p8_clipped__200_comb;
  assign p8_array_158723_comb[5] = p8_clipped__216_comb;
  assign p8_array_158723_comb[6] = p8_clipped__232_comb;
  assign p8_array_158723_comb[7] = p8_clipped__248_comb;
  assign p8_array_158724_comb[0] = p8_clipped__137_comb;
  assign p8_array_158724_comb[1] = p8_clipped__153_comb;
  assign p8_array_158724_comb[2] = p8_clipped__169_comb;
  assign p8_array_158724_comb[3] = p8_clipped__185_comb;
  assign p8_array_158724_comb[4] = p8_clipped__201_comb;
  assign p8_array_158724_comb[5] = p8_clipped__217_comb;
  assign p8_array_158724_comb[6] = p8_clipped__233_comb;
  assign p8_array_158724_comb[7] = p8_clipped__249_comb;
  assign p8_array_158725_comb[0] = p8_clipped__138_comb;
  assign p8_array_158725_comb[1] = p8_clipped__154_comb;
  assign p8_array_158725_comb[2] = p8_clipped__170_comb;
  assign p8_array_158725_comb[3] = p8_clipped__186_comb;
  assign p8_array_158725_comb[4] = p8_clipped__202_comb;
  assign p8_array_158725_comb[5] = p8_clipped__218_comb;
  assign p8_array_158725_comb[6] = p8_clipped__234_comb;
  assign p8_array_158725_comb[7] = p8_clipped__250_comb;
  assign p8_array_158726_comb[0] = p8_clipped__139_comb;
  assign p8_array_158726_comb[1] = p8_clipped__155_comb;
  assign p8_array_158726_comb[2] = p8_clipped__171_comb;
  assign p8_array_158726_comb[3] = p8_clipped__187_comb;
  assign p8_array_158726_comb[4] = p8_clipped__203_comb;
  assign p8_array_158726_comb[5] = p8_clipped__219_comb;
  assign p8_array_158726_comb[6] = p8_clipped__235_comb;
  assign p8_array_158726_comb[7] = p8_clipped__251_comb;
  assign p8_array_158727_comb[0] = p8_clipped__140_comb;
  assign p8_array_158727_comb[1] = p8_clipped__156_comb;
  assign p8_array_158727_comb[2] = p8_clipped__172_comb;
  assign p8_array_158727_comb[3] = p8_clipped__188_comb;
  assign p8_array_158727_comb[4] = p8_clipped__204_comb;
  assign p8_array_158727_comb[5] = p8_clipped__220_comb;
  assign p8_array_158727_comb[6] = p8_clipped__236_comb;
  assign p8_array_158727_comb[7] = p8_clipped__252_comb;
  assign p8_array_158728_comb[0] = p8_clipped__141_comb;
  assign p8_array_158728_comb[1] = p8_clipped__157_comb;
  assign p8_array_158728_comb[2] = p8_clipped__173_comb;
  assign p8_array_158728_comb[3] = p8_clipped__189_comb;
  assign p8_array_158728_comb[4] = p8_clipped__205_comb;
  assign p8_array_158728_comb[5] = p8_clipped__221_comb;
  assign p8_array_158728_comb[6] = p8_clipped__237_comb;
  assign p8_array_158728_comb[7] = p8_clipped__253_comb;
  assign p8_array_158729_comb[0] = p8_clipped__142_comb;
  assign p8_array_158729_comb[1] = p8_clipped__158_comb;
  assign p8_array_158729_comb[2] = p8_clipped__174_comb;
  assign p8_array_158729_comb[3] = p8_clipped__190_comb;
  assign p8_array_158729_comb[4] = p8_clipped__206_comb;
  assign p8_array_158729_comb[5] = p8_clipped__222_comb;
  assign p8_array_158729_comb[6] = p8_clipped__238_comb;
  assign p8_array_158729_comb[7] = p8_clipped__254_comb;
  assign p8_array_158730_comb[0] = p8_clipped__143_comb;
  assign p8_array_158730_comb[1] = p8_clipped__159_comb;
  assign p8_array_158730_comb[2] = p8_clipped__175_comb;
  assign p8_array_158730_comb[3] = p8_clipped__191_comb;
  assign p8_array_158730_comb[4] = p8_clipped__207_comb;
  assign p8_array_158730_comb[5] = p8_clipped__223_comb;
  assign p8_array_158730_comb[6] = p8_clipped__239_comb;
  assign p8_array_158730_comb[7] = p8_clipped__255_comb;
  assign p8_col_transformed_comb[0][0] = p8_array_158723_comb[0];
  assign p8_col_transformed_comb[0][1] = p8_array_158723_comb[1];
  assign p8_col_transformed_comb[0][2] = p8_array_158723_comb[2];
  assign p8_col_transformed_comb[0][3] = p8_array_158723_comb[3];
  assign p8_col_transformed_comb[0][4] = p8_array_158723_comb[4];
  assign p8_col_transformed_comb[0][5] = p8_array_158723_comb[5];
  assign p8_col_transformed_comb[0][6] = p8_array_158723_comb[6];
  assign p8_col_transformed_comb[0][7] = p8_array_158723_comb[7];
  assign p8_col_transformed_comb[1][0] = p8_array_158724_comb[0];
  assign p8_col_transformed_comb[1][1] = p8_array_158724_comb[1];
  assign p8_col_transformed_comb[1][2] = p8_array_158724_comb[2];
  assign p8_col_transformed_comb[1][3] = p8_array_158724_comb[3];
  assign p8_col_transformed_comb[1][4] = p8_array_158724_comb[4];
  assign p8_col_transformed_comb[1][5] = p8_array_158724_comb[5];
  assign p8_col_transformed_comb[1][6] = p8_array_158724_comb[6];
  assign p8_col_transformed_comb[1][7] = p8_array_158724_comb[7];
  assign p8_col_transformed_comb[2][0] = p8_array_158725_comb[0];
  assign p8_col_transformed_comb[2][1] = p8_array_158725_comb[1];
  assign p8_col_transformed_comb[2][2] = p8_array_158725_comb[2];
  assign p8_col_transformed_comb[2][3] = p8_array_158725_comb[3];
  assign p8_col_transformed_comb[2][4] = p8_array_158725_comb[4];
  assign p8_col_transformed_comb[2][5] = p8_array_158725_comb[5];
  assign p8_col_transformed_comb[2][6] = p8_array_158725_comb[6];
  assign p8_col_transformed_comb[2][7] = p8_array_158725_comb[7];
  assign p8_col_transformed_comb[3][0] = p8_array_158726_comb[0];
  assign p8_col_transformed_comb[3][1] = p8_array_158726_comb[1];
  assign p8_col_transformed_comb[3][2] = p8_array_158726_comb[2];
  assign p8_col_transformed_comb[3][3] = p8_array_158726_comb[3];
  assign p8_col_transformed_comb[3][4] = p8_array_158726_comb[4];
  assign p8_col_transformed_comb[3][5] = p8_array_158726_comb[5];
  assign p8_col_transformed_comb[3][6] = p8_array_158726_comb[6];
  assign p8_col_transformed_comb[3][7] = p8_array_158726_comb[7];
  assign p8_col_transformed_comb[4][0] = p8_array_158727_comb[0];
  assign p8_col_transformed_comb[4][1] = p8_array_158727_comb[1];
  assign p8_col_transformed_comb[4][2] = p8_array_158727_comb[2];
  assign p8_col_transformed_comb[4][3] = p8_array_158727_comb[3];
  assign p8_col_transformed_comb[4][4] = p8_array_158727_comb[4];
  assign p8_col_transformed_comb[4][5] = p8_array_158727_comb[5];
  assign p8_col_transformed_comb[4][6] = p8_array_158727_comb[6];
  assign p8_col_transformed_comb[4][7] = p8_array_158727_comb[7];
  assign p8_col_transformed_comb[5][0] = p8_array_158728_comb[0];
  assign p8_col_transformed_comb[5][1] = p8_array_158728_comb[1];
  assign p8_col_transformed_comb[5][2] = p8_array_158728_comb[2];
  assign p8_col_transformed_comb[5][3] = p8_array_158728_comb[3];
  assign p8_col_transformed_comb[5][4] = p8_array_158728_comb[4];
  assign p8_col_transformed_comb[5][5] = p8_array_158728_comb[5];
  assign p8_col_transformed_comb[5][6] = p8_array_158728_comb[6];
  assign p8_col_transformed_comb[5][7] = p8_array_158728_comb[7];
  assign p8_col_transformed_comb[6][0] = p8_array_158729_comb[0];
  assign p8_col_transformed_comb[6][1] = p8_array_158729_comb[1];
  assign p8_col_transformed_comb[6][2] = p8_array_158729_comb[2];
  assign p8_col_transformed_comb[6][3] = p8_array_158729_comb[3];
  assign p8_col_transformed_comb[6][4] = p8_array_158729_comb[4];
  assign p8_col_transformed_comb[6][5] = p8_array_158729_comb[5];
  assign p8_col_transformed_comb[6][6] = p8_array_158729_comb[6];
  assign p8_col_transformed_comb[6][7] = p8_array_158729_comb[7];
  assign p8_col_transformed_comb[7][0] = p8_array_158730_comb[0];
  assign p8_col_transformed_comb[7][1] = p8_array_158730_comb[1];
  assign p8_col_transformed_comb[7][2] = p8_array_158730_comb[2];
  assign p8_col_transformed_comb[7][3] = p8_array_158730_comb[3];
  assign p8_col_transformed_comb[7][4] = p8_array_158730_comb[4];
  assign p8_col_transformed_comb[7][5] = p8_array_158730_comb[5];
  assign p8_col_transformed_comb[7][6] = p8_array_158730_comb[6];
  assign p8_col_transformed_comb[7][7] = p8_array_158730_comb[7];

  // Registers for pipe stage 8:
  reg [7:0] p8_col_transformed[0:7][0:7];
  always @ (posedge clk) begin
    p8_col_transformed[0][0] <= p8_col_transformed_comb[0][0];
    p8_col_transformed[0][1] <= p8_col_transformed_comb[0][1];
    p8_col_transformed[0][2] <= p8_col_transformed_comb[0][2];
    p8_col_transformed[0][3] <= p8_col_transformed_comb[0][3];
    p8_col_transformed[0][4] <= p8_col_transformed_comb[0][4];
    p8_col_transformed[0][5] <= p8_col_transformed_comb[0][5];
    p8_col_transformed[0][6] <= p8_col_transformed_comb[0][6];
    p8_col_transformed[0][7] <= p8_col_transformed_comb[0][7];
    p8_col_transformed[1][0] <= p8_col_transformed_comb[1][0];
    p8_col_transformed[1][1] <= p8_col_transformed_comb[1][1];
    p8_col_transformed[1][2] <= p8_col_transformed_comb[1][2];
    p8_col_transformed[1][3] <= p8_col_transformed_comb[1][3];
    p8_col_transformed[1][4] <= p8_col_transformed_comb[1][4];
    p8_col_transformed[1][5] <= p8_col_transformed_comb[1][5];
    p8_col_transformed[1][6] <= p8_col_transformed_comb[1][6];
    p8_col_transformed[1][7] <= p8_col_transformed_comb[1][7];
    p8_col_transformed[2][0] <= p8_col_transformed_comb[2][0];
    p8_col_transformed[2][1] <= p8_col_transformed_comb[2][1];
    p8_col_transformed[2][2] <= p8_col_transformed_comb[2][2];
    p8_col_transformed[2][3] <= p8_col_transformed_comb[2][3];
    p8_col_transformed[2][4] <= p8_col_transformed_comb[2][4];
    p8_col_transformed[2][5] <= p8_col_transformed_comb[2][5];
    p8_col_transformed[2][6] <= p8_col_transformed_comb[2][6];
    p8_col_transformed[2][7] <= p8_col_transformed_comb[2][7];
    p8_col_transformed[3][0] <= p8_col_transformed_comb[3][0];
    p8_col_transformed[3][1] <= p8_col_transformed_comb[3][1];
    p8_col_transformed[3][2] <= p8_col_transformed_comb[3][2];
    p8_col_transformed[3][3] <= p8_col_transformed_comb[3][3];
    p8_col_transformed[3][4] <= p8_col_transformed_comb[3][4];
    p8_col_transformed[3][5] <= p8_col_transformed_comb[3][5];
    p8_col_transformed[3][6] <= p8_col_transformed_comb[3][6];
    p8_col_transformed[3][7] <= p8_col_transformed_comb[3][7];
    p8_col_transformed[4][0] <= p8_col_transformed_comb[4][0];
    p8_col_transformed[4][1] <= p8_col_transformed_comb[4][1];
    p8_col_transformed[4][2] <= p8_col_transformed_comb[4][2];
    p8_col_transformed[4][3] <= p8_col_transformed_comb[4][3];
    p8_col_transformed[4][4] <= p8_col_transformed_comb[4][4];
    p8_col_transformed[4][5] <= p8_col_transformed_comb[4][5];
    p8_col_transformed[4][6] <= p8_col_transformed_comb[4][6];
    p8_col_transformed[4][7] <= p8_col_transformed_comb[4][7];
    p8_col_transformed[5][0] <= p8_col_transformed_comb[5][0];
    p8_col_transformed[5][1] <= p8_col_transformed_comb[5][1];
    p8_col_transformed[5][2] <= p8_col_transformed_comb[5][2];
    p8_col_transformed[5][3] <= p8_col_transformed_comb[5][3];
    p8_col_transformed[5][4] <= p8_col_transformed_comb[5][4];
    p8_col_transformed[5][5] <= p8_col_transformed_comb[5][5];
    p8_col_transformed[5][6] <= p8_col_transformed_comb[5][6];
    p8_col_transformed[5][7] <= p8_col_transformed_comb[5][7];
    p8_col_transformed[6][0] <= p8_col_transformed_comb[6][0];
    p8_col_transformed[6][1] <= p8_col_transformed_comb[6][1];
    p8_col_transformed[6][2] <= p8_col_transformed_comb[6][2];
    p8_col_transformed[6][3] <= p8_col_transformed_comb[6][3];
    p8_col_transformed[6][4] <= p8_col_transformed_comb[6][4];
    p8_col_transformed[6][5] <= p8_col_transformed_comb[6][5];
    p8_col_transformed[6][6] <= p8_col_transformed_comb[6][6];
    p8_col_transformed[6][7] <= p8_col_transformed_comb[6][7];
    p8_col_transformed[7][0] <= p8_col_transformed_comb[7][0];
    p8_col_transformed[7][1] <= p8_col_transformed_comb[7][1];
    p8_col_transformed[7][2] <= p8_col_transformed_comb[7][2];
    p8_col_transformed[7][3] <= p8_col_transformed_comb[7][3];
    p8_col_transformed[7][4] <= p8_col_transformed_comb[7][4];
    p8_col_transformed[7][5] <= p8_col_transformed_comb[7][5];
    p8_col_transformed[7][6] <= p8_col_transformed_comb[7][6];
    p8_col_transformed[7][7] <= p8_col_transformed_comb[7][7];
  end
  assign out = {{p8_col_transformed[7][7], p8_col_transformed[7][6], p8_col_transformed[7][5], p8_col_transformed[7][4], p8_col_transformed[7][3], p8_col_transformed[7][2], p8_col_transformed[7][1], p8_col_transformed[7][0]}, {p8_col_transformed[6][7], p8_col_transformed[6][6], p8_col_transformed[6][5], p8_col_transformed[6][4], p8_col_transformed[6][3], p8_col_transformed[6][2], p8_col_transformed[6][1], p8_col_transformed[6][0]}, {p8_col_transformed[5][7], p8_col_transformed[5][6], p8_col_transformed[5][5], p8_col_transformed[5][4], p8_col_transformed[5][3], p8_col_transformed[5][2], p8_col_transformed[5][1], p8_col_transformed[5][0]}, {p8_col_transformed[4][7], p8_col_transformed[4][6], p8_col_transformed[4][5], p8_col_transformed[4][4], p8_col_transformed[4][3], p8_col_transformed[4][2], p8_col_transformed[4][1], p8_col_transformed[4][0]}, {p8_col_transformed[3][7], p8_col_transformed[3][6], p8_col_transformed[3][5], p8_col_transformed[3][4], p8_col_transformed[3][3], p8_col_transformed[3][2], p8_col_transformed[3][1], p8_col_transformed[3][0]}, {p8_col_transformed[2][7], p8_col_transformed[2][6], p8_col_transformed[2][5], p8_col_transformed[2][4], p8_col_transformed[2][3], p8_col_transformed[2][2], p8_col_transformed[2][1], p8_col_transformed[2][0]}, {p8_col_transformed[1][7], p8_col_transformed[1][6], p8_col_transformed[1][5], p8_col_transformed[1][4], p8_col_transformed[1][3], p8_col_transformed[1][2], p8_col_transformed[1][1], p8_col_transformed[1][0]}, {p8_col_transformed[0][7], p8_col_transformed[0][6], p8_col_transformed[0][5], p8_col_transformed[0][4], p8_col_transformed[0][3], p8_col_transformed[0][2], p8_col_transformed[0][1], p8_col_transformed[0][0]}};
endmodule
