module dct_2d_u8(
  input wire clk,
  input wire [511:0] x,
  output wire [511:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [15:0] smul16b_8b_x_8b (input reg [7:0] lhs, input reg [7:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [15:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul16b_8b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_6b (input reg [7:0] lhs, input reg [5:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [15:0] smul16b_8b_x_9b (input reg [7:0] lhs, input reg [8:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [15:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul16b_8b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_7b (input reg [31:0] lhs, input reg [6:0] rhs);
    begin
      umul32b_32b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [7:0] x_unflattened[0:7][0:7];
  assign x_unflattened[0][0] = x[7:0];
  assign x_unflattened[0][1] = x[15:8];
  assign x_unflattened[0][2] = x[23:16];
  assign x_unflattened[0][3] = x[31:24];
  assign x_unflattened[0][4] = x[39:32];
  assign x_unflattened[0][5] = x[47:40];
  assign x_unflattened[0][6] = x[55:48];
  assign x_unflattened[0][7] = x[63:56];
  assign x_unflattened[1][0] = x[71:64];
  assign x_unflattened[1][1] = x[79:72];
  assign x_unflattened[1][2] = x[87:80];
  assign x_unflattened[1][3] = x[95:88];
  assign x_unflattened[1][4] = x[103:96];
  assign x_unflattened[1][5] = x[111:104];
  assign x_unflattened[1][6] = x[119:112];
  assign x_unflattened[1][7] = x[127:120];
  assign x_unflattened[2][0] = x[135:128];
  assign x_unflattened[2][1] = x[143:136];
  assign x_unflattened[2][2] = x[151:144];
  assign x_unflattened[2][3] = x[159:152];
  assign x_unflattened[2][4] = x[167:160];
  assign x_unflattened[2][5] = x[175:168];
  assign x_unflattened[2][6] = x[183:176];
  assign x_unflattened[2][7] = x[191:184];
  assign x_unflattened[3][0] = x[199:192];
  assign x_unflattened[3][1] = x[207:200];
  assign x_unflattened[3][2] = x[215:208];
  assign x_unflattened[3][3] = x[223:216];
  assign x_unflattened[3][4] = x[231:224];
  assign x_unflattened[3][5] = x[239:232];
  assign x_unflattened[3][6] = x[247:240];
  assign x_unflattened[3][7] = x[255:248];
  assign x_unflattened[4][0] = x[263:256];
  assign x_unflattened[4][1] = x[271:264];
  assign x_unflattened[4][2] = x[279:272];
  assign x_unflattened[4][3] = x[287:280];
  assign x_unflattened[4][4] = x[295:288];
  assign x_unflattened[4][5] = x[303:296];
  assign x_unflattened[4][6] = x[311:304];
  assign x_unflattened[4][7] = x[319:312];
  assign x_unflattened[5][0] = x[327:320];
  assign x_unflattened[5][1] = x[335:328];
  assign x_unflattened[5][2] = x[343:336];
  assign x_unflattened[5][3] = x[351:344];
  assign x_unflattened[5][4] = x[359:352];
  assign x_unflattened[5][5] = x[367:360];
  assign x_unflattened[5][6] = x[375:368];
  assign x_unflattened[5][7] = x[383:376];
  assign x_unflattened[6][0] = x[391:384];
  assign x_unflattened[6][1] = x[399:392];
  assign x_unflattened[6][2] = x[407:400];
  assign x_unflattened[6][3] = x[415:408];
  assign x_unflattened[6][4] = x[423:416];
  assign x_unflattened[6][5] = x[431:424];
  assign x_unflattened[6][6] = x[439:432];
  assign x_unflattened[6][7] = x[447:440];
  assign x_unflattened[7][0] = x[455:448];
  assign x_unflattened[7][1] = x[463:456];
  assign x_unflattened[7][2] = x[471:464];
  assign x_unflattened[7][3] = x[479:472];
  assign x_unflattened[7][4] = x[487:480];
  assign x_unflattened[7][5] = x[495:488];
  assign x_unflattened[7][6] = x[503:496];
  assign x_unflattened[7][7] = x[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_x[0:7][0:7];
  always @ (posedge clk) begin
    p0_x[0][0] <= x_unflattened[0][0];
    p0_x[0][1] <= x_unflattened[0][1];
    p0_x[0][2] <= x_unflattened[0][2];
    p0_x[0][3] <= x_unflattened[0][3];
    p0_x[0][4] <= x_unflattened[0][4];
    p0_x[0][5] <= x_unflattened[0][5];
    p0_x[0][6] <= x_unflattened[0][6];
    p0_x[0][7] <= x_unflattened[0][7];
    p0_x[1][0] <= x_unflattened[1][0];
    p0_x[1][1] <= x_unflattened[1][1];
    p0_x[1][2] <= x_unflattened[1][2];
    p0_x[1][3] <= x_unflattened[1][3];
    p0_x[1][4] <= x_unflattened[1][4];
    p0_x[1][5] <= x_unflattened[1][5];
    p0_x[1][6] <= x_unflattened[1][6];
    p0_x[1][7] <= x_unflattened[1][7];
    p0_x[2][0] <= x_unflattened[2][0];
    p0_x[2][1] <= x_unflattened[2][1];
    p0_x[2][2] <= x_unflattened[2][2];
    p0_x[2][3] <= x_unflattened[2][3];
    p0_x[2][4] <= x_unflattened[2][4];
    p0_x[2][5] <= x_unflattened[2][5];
    p0_x[2][6] <= x_unflattened[2][6];
    p0_x[2][7] <= x_unflattened[2][7];
    p0_x[3][0] <= x_unflattened[3][0];
    p0_x[3][1] <= x_unflattened[3][1];
    p0_x[3][2] <= x_unflattened[3][2];
    p0_x[3][3] <= x_unflattened[3][3];
    p0_x[3][4] <= x_unflattened[3][4];
    p0_x[3][5] <= x_unflattened[3][5];
    p0_x[3][6] <= x_unflattened[3][6];
    p0_x[3][7] <= x_unflattened[3][7];
    p0_x[4][0] <= x_unflattened[4][0];
    p0_x[4][1] <= x_unflattened[4][1];
    p0_x[4][2] <= x_unflattened[4][2];
    p0_x[4][3] <= x_unflattened[4][3];
    p0_x[4][4] <= x_unflattened[4][4];
    p0_x[4][5] <= x_unflattened[4][5];
    p0_x[4][6] <= x_unflattened[4][6];
    p0_x[4][7] <= x_unflattened[4][7];
    p0_x[5][0] <= x_unflattened[5][0];
    p0_x[5][1] <= x_unflattened[5][1];
    p0_x[5][2] <= x_unflattened[5][2];
    p0_x[5][3] <= x_unflattened[5][3];
    p0_x[5][4] <= x_unflattened[5][4];
    p0_x[5][5] <= x_unflattened[5][5];
    p0_x[5][6] <= x_unflattened[5][6];
    p0_x[5][7] <= x_unflattened[5][7];
    p0_x[6][0] <= x_unflattened[6][0];
    p0_x[6][1] <= x_unflattened[6][1];
    p0_x[6][2] <= x_unflattened[6][2];
    p0_x[6][3] <= x_unflattened[6][3];
    p0_x[6][4] <= x_unflattened[6][4];
    p0_x[6][5] <= x_unflattened[6][5];
    p0_x[6][6] <= x_unflattened[6][6];
    p0_x[6][7] <= x_unflattened[6][7];
    p0_x[7][0] <= x_unflattened[7][0];
    p0_x[7][1] <= x_unflattened[7][1];
    p0_x[7][2] <= x_unflattened[7][2];
    p0_x[7][3] <= x_unflattened[7][3];
    p0_x[7][4] <= x_unflattened[7][4];
    p0_x[7][5] <= x_unflattened[7][5];
    p0_x[7][6] <= x_unflattened[7][6];
    p0_x[7][7] <= x_unflattened[7][7];
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_array_index_130665_comb;
  wire [7:0] p1_array_index_130666_comb;
  wire [7:0] p1_array_index_130667_comb;
  wire [7:0] p1_array_index_130668_comb;
  wire [7:0] p1_array_index_130669_comb;
  wire [7:0] p1_array_index_130670_comb;
  wire [7:0] p1_array_index_130671_comb;
  wire [7:0] p1_array_index_130672_comb;
  wire [7:0] p1_array_index_130673_comb;
  wire [7:0] p1_array_index_130674_comb;
  wire [7:0] p1_array_index_130675_comb;
  wire [7:0] p1_array_index_130676_comb;
  wire [7:0] p1_array_index_130677_comb;
  wire [7:0] p1_array_index_130678_comb;
  wire [7:0] p1_array_index_130679_comb;
  wire [7:0] p1_array_index_130680_comb;
  wire [7:0] p1_array_index_130681_comb;
  wire [7:0] p1_array_index_130682_comb;
  wire [7:0] p1_array_index_130683_comb;
  wire [7:0] p1_array_index_130684_comb;
  wire [7:0] p1_array_index_130685_comb;
  wire [7:0] p1_array_index_130686_comb;
  wire [7:0] p1_array_index_130687_comb;
  wire [7:0] p1_array_index_130688_comb;
  wire [7:0] p1_array_index_130689_comb;
  wire [7:0] p1_array_index_130690_comb;
  wire [7:0] p1_array_index_130691_comb;
  wire [7:0] p1_array_index_130692_comb;
  wire [7:0] p1_array_index_130693_comb;
  wire [7:0] p1_array_index_130694_comb;
  wire [7:0] p1_array_index_130695_comb;
  wire [7:0] p1_array_index_130696_comb;
  wire [7:0] p1_array_index_130697_comb;
  wire [7:0] p1_array_index_130698_comb;
  wire [7:0] p1_array_index_130699_comb;
  wire [7:0] p1_array_index_130700_comb;
  wire [7:0] p1_array_index_130701_comb;
  wire [7:0] p1_array_index_130702_comb;
  wire [7:0] p1_array_index_130703_comb;
  wire [7:0] p1_array_index_130704_comb;
  wire [7:0] p1_array_index_130705_comb;
  wire [7:0] p1_array_index_130706_comb;
  wire [7:0] p1_array_index_130707_comb;
  wire [7:0] p1_array_index_130708_comb;
  wire [7:0] p1_array_index_130709_comb;
  wire [7:0] p1_array_index_130710_comb;
  wire [7:0] p1_array_index_130711_comb;
  wire [7:0] p1_array_index_130712_comb;
  wire [7:0] p1_array_index_130713_comb;
  wire [7:0] p1_array_index_130714_comb;
  wire [7:0] p1_array_index_130715_comb;
  wire [7:0] p1_array_index_130716_comb;
  wire [7:0] p1_array_index_130717_comb;
  wire [7:0] p1_array_index_130718_comb;
  wire [7:0] p1_array_index_130719_comb;
  wire [7:0] p1_array_index_130720_comb;
  wire [7:0] p1_array_index_130721_comb;
  wire [7:0] p1_array_index_130722_comb;
  wire [7:0] p1_array_index_130723_comb;
  wire [7:0] p1_array_index_130724_comb;
  wire [7:0] p1_array_index_130725_comb;
  wire [7:0] p1_array_index_130726_comb;
  wire [7:0] p1_array_index_130727_comb;
  wire [7:0] p1_array_index_130728_comb;
  wire [7:0] p1_shifted__18_squeezed_comb;
  wire [7:0] p1_shifted__19_squeezed_comb;
  wire [7:0] p1_shifted__20_squeezed_comb;
  wire [7:0] p1_shifted__21_squeezed_comb;
  wire [7:0] p1_shifted__26_squeezed_comb;
  wire [7:0] p1_shifted__27_squeezed_comb;
  wire [7:0] p1_shifted__28_squeezed_comb;
  wire [7:0] p1_shifted__29_squeezed_comb;
  wire [7:0] p1_shifted__34_squeezed_comb;
  wire [7:0] p1_shifted__35_squeezed_comb;
  wire [7:0] p1_shifted__36_squeezed_comb;
  wire [7:0] p1_shifted__37_squeezed_comb;
  wire [7:0] p1_shifted__42_squeezed_comb;
  wire [7:0] p1_shifted__43_squeezed_comb;
  wire [7:0] p1_shifted__44_squeezed_comb;
  wire [7:0] p1_shifted__45_squeezed_comb;
  wire [7:0] p1_shifted__16_squeezed_comb;
  wire [7:0] p1_shifted__23_squeezed_comb;
  wire [7:0] p1_shifted__24_squeezed_comb;
  wire [7:0] p1_shifted__31_squeezed_comb;
  wire [7:0] p1_shifted__32_squeezed_comb;
  wire [7:0] p1_shifted__39_squeezed_comb;
  wire [7:0] p1_shifted__40_squeezed_comb;
  wire [7:0] p1_shifted__47_squeezed_comb;
  wire [7:0] p1_shifted__17_squeezed_comb;
  wire [7:0] p1_shifted__22_squeezed_comb;
  wire [7:0] p1_shifted__25_squeezed_comb;
  wire [7:0] p1_shifted__30_squeezed_comb;
  wire [7:0] p1_shifted__33_squeezed_comb;
  wire [7:0] p1_shifted__38_squeezed_comb;
  wire [7:0] p1_shifted__41_squeezed_comb;
  wire [7:0] p1_shifted__46_squeezed_comb;
  wire [7:0] p1_shifted__2_squeezed_comb;
  wire [7:0] p1_shifted__3_squeezed_comb;
  wire [7:0] p1_shifted__4_squeezed_comb;
  wire [7:0] p1_shifted__5_squeezed_comb;
  wire [7:0] p1_shifted__58_squeezed_comb;
  wire [7:0] p1_shifted__59_squeezed_comb;
  wire [7:0] p1_shifted__60_squeezed_comb;
  wire [7:0] p1_shifted__61_squeezed_comb;
  wire [7:0] p1_shifted_squeezed_comb;
  wire [7:0] p1_shifted__7_squeezed_comb;
  wire [7:0] p1_shifted__56_squeezed_comb;
  wire [7:0] p1_shifted__63_squeezed_comb;
  wire [7:0] p1_shifted__1_squeezed_comb;
  wire [7:0] p1_shifted__6_squeezed_comb;
  wire [7:0] p1_shifted__57_squeezed_comb;
  wire [7:0] p1_shifted__62_squeezed_comb;
  wire [7:0] p1_shifted__10_squeezed_comb;
  wire [7:0] p1_shifted__11_squeezed_comb;
  wire [7:0] p1_shifted__12_squeezed_comb;
  wire [7:0] p1_shifted__13_squeezed_comb;
  wire [7:0] p1_shifted__50_squeezed_comb;
  wire [7:0] p1_shifted__51_squeezed_comb;
  wire [7:0] p1_shifted__52_squeezed_comb;
  wire [7:0] p1_shifted__53_squeezed_comb;
  wire [7:0] p1_shifted__8_squeezed_comb;
  wire [7:0] p1_shifted__15_squeezed_comb;
  wire [7:0] p1_shifted__48_squeezed_comb;
  wire [7:0] p1_shifted__55_squeezed_comb;
  wire [7:0] p1_shifted__9_squeezed_comb;
  wire [7:0] p1_shifted__14_squeezed_comb;
  wire [7:0] p1_shifted__49_squeezed_comb;
  wire [7:0] p1_shifted__54_squeezed_comb;
  wire [15:0] p1_smul_57362_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___8_comb;
  wire [13:0] p1_smul_57364_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___9_comb;
  wire [13:0] p1_smul_57366_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___10_comb;
  wire [15:0] p1_smul_57368_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___11_comb;
  wire [15:0] p1_smul_57378_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___12_comb;
  wire [13:0] p1_smul_57380_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___13_comb;
  wire [13:0] p1_smul_57382_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___14_comb;
  wire [15:0] p1_smul_57384_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___15_comb;
  wire [15:0] p1_smul_57394_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___16_comb;
  wire [13:0] p1_smul_57396_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___17_comb;
  wire [13:0] p1_smul_57398_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___18_comb;
  wire [15:0] p1_smul_57400_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___19_comb;
  wire [15:0] p1_smul_57410_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___20_comb;
  wire [13:0] p1_smul_57412_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___21_comb;
  wire [13:0] p1_smul_57414_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___22_comb;
  wire [15:0] p1_smul_57416_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___23_comb;
  wire [14:0] p1_smul_57486_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___8_comb;
  wire [14:0] p1_smul_57492_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___9_comb;
  wire [14:0] p1_smul_57494_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___10_comb;
  wire [14:0] p1_smul_57500_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___11_comb;
  wire [14:0] p1_smul_57502_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___12_comb;
  wire [14:0] p1_smul_57508_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___13_comb;
  wire [14:0] p1_smul_57510_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___14_comb;
  wire [14:0] p1_smul_57516_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___15_comb;
  wire [14:0] p1_smul_57518_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___16_comb;
  wire [14:0] p1_smul_57524_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___17_comb;
  wire [14:0] p1_smul_57526_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___18_comb;
  wire [14:0] p1_smul_57532_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___19_comb;
  wire [14:0] p1_smul_57534_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___20_comb;
  wire [14:0] p1_smul_57540_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___21_comb;
  wire [14:0] p1_smul_57542_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___22_comb;
  wire [14:0] p1_smul_57548_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___23_comb;
  wire [13:0] p1_smul_57616_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___40_comb;
  wire [15:0] p1_smul_57620_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___41_comb;
  wire [15:0] p1_smul_57622_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___42_comb;
  wire [13:0] p1_smul_57626_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___43_comb;
  wire [13:0] p1_smul_57632_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___44_comb;
  wire [15:0] p1_smul_57636_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___45_comb;
  wire [15:0] p1_smul_57638_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___46_comb;
  wire [13:0] p1_smul_57642_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___47_comb;
  wire [13:0] p1_smul_57648_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___48_comb;
  wire [15:0] p1_smul_57652_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___49_comb;
  wire [15:0] p1_smul_57654_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___50_comb;
  wire [13:0] p1_smul_57658_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___51_comb;
  wire [13:0] p1_smul_57664_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___52_comb;
  wire [15:0] p1_smul_57668_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___53_comb;
  wire [15:0] p1_smul_57670_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___54_comb;
  wire [13:0] p1_smul_57674_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___55_comb;
  wire [15:0] p1_smul_57870_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___72_comb;
  wire [13:0] p1_smul_57874_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___73_comb;
  wire [13:0] p1_smul_57880_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___74_comb;
  wire [15:0] p1_smul_57884_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___75_comb;
  wire [15:0] p1_smul_57886_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___76_comb;
  wire [13:0] p1_smul_57890_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___77_comb;
  wire [13:0] p1_smul_57896_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___78_comb;
  wire [15:0] p1_smul_57900_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___79_comb;
  wire [15:0] p1_smul_57902_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___80_comb;
  wire [13:0] p1_smul_57906_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___81_comb;
  wire [13:0] p1_smul_57912_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___82_comb;
  wire [15:0] p1_smul_57916_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___83_comb;
  wire [15:0] p1_smul_57918_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___84_comb;
  wire [13:0] p1_smul_57922_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___85_comb;
  wire [13:0] p1_smul_57928_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___86_comb;
  wire [15:0] p1_smul_57932_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___87_comb;
  wire [14:0] p1_smul_58000_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___40_comb;
  wire [14:0] p1_smul_58004_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___41_comb;
  wire [14:0] p1_smul_58006_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___42_comb;
  wire [14:0] p1_smul_58010_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___43_comb;
  wire [14:0] p1_smul_58016_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___44_comb;
  wire [14:0] p1_smul_58020_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___45_comb;
  wire [14:0] p1_smul_58022_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___46_comb;
  wire [14:0] p1_smul_58026_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___47_comb;
  wire [14:0] p1_smul_58032_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___48_comb;
  wire [14:0] p1_smul_58036_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___49_comb;
  wire [14:0] p1_smul_58038_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___50_comb;
  wire [14:0] p1_smul_58042_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___51_comb;
  wire [14:0] p1_smul_58048_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___52_comb;
  wire [14:0] p1_smul_58052_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___53_comb;
  wire [14:0] p1_smul_58054_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___54_comb;
  wire [14:0] p1_smul_58058_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___55_comb;
  wire [13:0] p1_smul_58126_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___104_comb;
  wire [15:0] p1_smul_58128_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___105_comb;
  wire [15:0] p1_smul_58138_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___106_comb;
  wire [13:0] p1_smul_58140_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___107_comb;
  wire [13:0] p1_smul_58142_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___108_comb;
  wire [15:0] p1_smul_58144_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___109_comb;
  wire [15:0] p1_smul_58154_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___110_comb;
  wire [13:0] p1_smul_58156_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___111_comb;
  wire [13:0] p1_smul_58158_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___112_comb;
  wire [15:0] p1_smul_58160_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___113_comb;
  wire [15:0] p1_smul_58170_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___114_comb;
  wire [13:0] p1_smul_58172_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___115_comb;
  wire [13:0] p1_smul_58174_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___116_comb;
  wire [15:0] p1_smul_58176_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___117_comb;
  wire [15:0] p1_smul_58186_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___118_comb;
  wire [13:0] p1_smul_58188_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___119_comb;
  wire [15:0] p1_smul_57330_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits__comb;
  wire [13:0] p1_smul_57332_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___1_comb;
  wire [13:0] p1_smul_57334_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___2_comb;
  wire [15:0] p1_smul_57336_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___3_comb;
  wire [15:0] p1_smul_57442_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___28_comb;
  wire [13:0] p1_smul_57444_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___29_comb;
  wire [13:0] p1_smul_57446_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___30_comb;
  wire [15:0] p1_smul_57448_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___31_comb;
  wire [14:0] p1_smul_57454_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits__comb;
  wire [14:0] p1_smul_57460_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___1_comb;
  wire [14:0] p1_smul_57462_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___2_comb;
  wire [14:0] p1_smul_57468_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___3_comb;
  wire [14:0] p1_smul_57566_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___28_comb;
  wire [14:0] p1_smul_57572_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___29_comb;
  wire [14:0] p1_smul_57574_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___30_comb;
  wire [14:0] p1_smul_57580_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___31_comb;
  wire [13:0] p1_smul_57584_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___32_comb;
  wire [15:0] p1_smul_57588_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___33_comb;
  wire [15:0] p1_smul_57590_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___34_comb;
  wire [13:0] p1_smul_57594_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___35_comb;
  wire [13:0] p1_smul_57696_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___60_comb;
  wire [15:0] p1_smul_57700_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___61_comb;
  wire [15:0] p1_smul_57702_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___62_comb;
  wire [13:0] p1_smul_57706_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___63_comb;
  wire [15:0] p1_smul_57838_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___64_comb;
  wire [13:0] p1_smul_57842_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___65_comb;
  wire [13:0] p1_smul_57848_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___66_comb;
  wire [15:0] p1_smul_57852_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___67_comb;
  wire [15:0] p1_smul_57950_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___92_comb;
  wire [13:0] p1_smul_57954_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___93_comb;
  wire [13:0] p1_smul_57960_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___94_comb;
  wire [15:0] p1_smul_57964_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___95_comb;
  wire [14:0] p1_smul_57968_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___32_comb;
  wire [14:0] p1_smul_57972_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___33_comb;
  wire [14:0] p1_smul_57974_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___34_comb;
  wire [14:0] p1_smul_57978_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___35_comb;
  wire [14:0] p1_smul_58080_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___60_comb;
  wire [14:0] p1_smul_58084_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___61_comb;
  wire [14:0] p1_smul_58086_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___62_comb;
  wire [14:0] p1_smul_58090_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___63_comb;
  wire [13:0] p1_smul_58094_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___96_comb;
  wire [15:0] p1_smul_58096_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___97_comb;
  wire [15:0] p1_smul_58106_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___98_comb;
  wire [13:0] p1_smul_58108_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___99_comb;
  wire [13:0] p1_smul_58206_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___124_comb;
  wire [15:0] p1_smul_58208_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___125_comb;
  wire [15:0] p1_smul_58218_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___126_comb;
  wire [13:0] p1_smul_58220_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___127_comb;
  wire [15:0] p1_smul_57346_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___4_comb;
  wire [13:0] p1_smul_57348_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___5_comb;
  wire [13:0] p1_smul_57350_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___6_comb;
  wire [15:0] p1_smul_57352_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___7_comb;
  wire [15:0] p1_smul_57426_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___24_comb;
  wire [13:0] p1_smul_57428_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___25_comb;
  wire [13:0] p1_smul_57430_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___26_comb;
  wire [15:0] p1_smul_57432_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___27_comb;
  wire [14:0] p1_smul_57470_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___4_comb;
  wire [14:0] p1_smul_57476_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___5_comb;
  wire [14:0] p1_smul_57478_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___6_comb;
  wire [14:0] p1_smul_57484_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___7_comb;
  wire [14:0] p1_smul_57550_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___24_comb;
  wire [14:0] p1_smul_57556_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___25_comb;
  wire [14:0] p1_smul_57558_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___26_comb;
  wire [14:0] p1_smul_57564_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___27_comb;
  wire [13:0] p1_smul_57600_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___36_comb;
  wire [15:0] p1_smul_57604_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___37_comb;
  wire [15:0] p1_smul_57606_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___38_comb;
  wire [13:0] p1_smul_57610_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___39_comb;
  wire [13:0] p1_smul_57680_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___56_comb;
  wire [15:0] p1_smul_57684_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___57_comb;
  wire [15:0] p1_smul_57686_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___58_comb;
  wire [13:0] p1_smul_57690_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___59_comb;
  wire [15:0] p1_smul_57854_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___68_comb;
  wire [13:0] p1_smul_57858_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___69_comb;
  wire [13:0] p1_smul_57864_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___70_comb;
  wire [15:0] p1_smul_57868_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___71_comb;
  wire [15:0] p1_smul_57934_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___88_comb;
  wire [13:0] p1_smul_57938_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___89_comb;
  wire [13:0] p1_smul_57944_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___90_comb;
  wire [15:0] p1_smul_57948_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___91_comb;
  wire [14:0] p1_smul_57984_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___36_comb;
  wire [14:0] p1_smul_57988_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___37_comb;
  wire [14:0] p1_smul_57990_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___38_comb;
  wire [14:0] p1_smul_57994_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___39_comb;
  wire [14:0] p1_smul_58064_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___56_comb;
  wire [14:0] p1_smul_58068_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___57_comb;
  wire [14:0] p1_smul_58070_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___58_comb;
  wire [14:0] p1_smul_58074_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___59_comb;
  wire [13:0] p1_smul_58110_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___100_comb;
  wire [15:0] p1_smul_58112_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___101_comb;
  wire [15:0] p1_smul_58122_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___102_comb;
  wire [13:0] p1_smul_58124_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___103_comb;
  wire [13:0] p1_smul_58190_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___120_comb;
  wire [15:0] p1_smul_58192_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___121_comb;
  wire [15:0] p1_smul_58202_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___122_comb;
  wire [13:0] p1_smul_58204_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___123_comb;
  wire [7:0] p1_smul_57326_TrailingBits___144_comb;
  wire [7:0] p1_smul_57326_TrailingBits___145_comb;
  wire [7:0] p1_smul_57326_TrailingBits___146_comb;
  wire [7:0] p1_smul_57326_TrailingBits___147_comb;
  wire [7:0] p1_smul_57326_TrailingBits___148_comb;
  wire [7:0] p1_smul_57326_TrailingBits___149_comb;
  wire [7:0] p1_smul_57326_TrailingBits___150_comb;
  wire [7:0] p1_smul_57326_TrailingBits___151_comb;
  wire [7:0] p1_smul_57326_TrailingBits___152_comb;
  wire [7:0] p1_smul_57326_TrailingBits___153_comb;
  wire [7:0] p1_smul_57326_TrailingBits___154_comb;
  wire [7:0] p1_smul_57326_TrailingBits___155_comb;
  wire [7:0] p1_smul_57326_TrailingBits___156_comb;
  wire [7:0] p1_smul_57326_TrailingBits___157_comb;
  wire [7:0] p1_smul_57326_TrailingBits___158_comb;
  wire [7:0] p1_smul_57326_TrailingBits___159_comb;
  wire [7:0] p1_smul_57326_TrailingBits___160_comb;
  wire [7:0] p1_smul_57326_TrailingBits___161_comb;
  wire [7:0] p1_smul_57326_TrailingBits___162_comb;
  wire [7:0] p1_smul_57326_TrailingBits___163_comb;
  wire [7:0] p1_smul_57326_TrailingBits___164_comb;
  wire [7:0] p1_smul_57326_TrailingBits___165_comb;
  wire [7:0] p1_smul_57326_TrailingBits___166_comb;
  wire [7:0] p1_smul_57326_TrailingBits___167_comb;
  wire [7:0] p1_smul_57326_TrailingBits___168_comb;
  wire [7:0] p1_smul_57326_TrailingBits___169_comb;
  wire [7:0] p1_smul_57326_TrailingBits___170_comb;
  wire [7:0] p1_smul_57326_TrailingBits___171_comb;
  wire [7:0] p1_smul_57326_TrailingBits___172_comb;
  wire [7:0] p1_smul_57326_TrailingBits___173_comb;
  wire [7:0] p1_smul_57326_TrailingBits___174_comb;
  wire [7:0] p1_smul_57326_TrailingBits___175_comb;
  wire [24:0] p1_concat_131721_comb;
  wire [22:0] p1_concat_131722_comb;
  wire [22:0] p1_concat_131723_comb;
  wire [24:0] p1_concat_131724_comb;
  wire [24:0] p1_concat_131725_comb;
  wire [22:0] p1_concat_131726_comb;
  wire [22:0] p1_concat_131727_comb;
  wire [24:0] p1_concat_131728_comb;
  wire [24:0] p1_concat_131729_comb;
  wire [22:0] p1_concat_131730_comb;
  wire [22:0] p1_concat_131731_comb;
  wire [24:0] p1_concat_131732_comb;
  wire [24:0] p1_concat_131733_comb;
  wire [22:0] p1_concat_131734_comb;
  wire [22:0] p1_concat_131735_comb;
  wire [24:0] p1_concat_131736_comb;
  wire [24:0] p1_concat_131737_comb;
  wire [24:0] p1_concat_131738_comb;
  wire [24:0] p1_concat_131739_comb;
  wire [24:0] p1_concat_131740_comb;
  wire [24:0] p1_concat_131741_comb;
  wire [24:0] p1_concat_131742_comb;
  wire [24:0] p1_concat_131743_comb;
  wire [24:0] p1_concat_131744_comb;
  wire [24:0] p1_concat_131745_comb;
  wire [24:0] p1_concat_131746_comb;
  wire [24:0] p1_concat_131747_comb;
  wire [24:0] p1_concat_131748_comb;
  wire [24:0] p1_concat_131749_comb;
  wire [24:0] p1_concat_131750_comb;
  wire [24:0] p1_concat_131751_comb;
  wire [24:0] p1_concat_131752_comb;
  wire [22:0] p1_concat_131753_comb;
  wire [24:0] p1_concat_131754_comb;
  wire [24:0] p1_concat_131755_comb;
  wire [22:0] p1_concat_131756_comb;
  wire [22:0] p1_concat_131757_comb;
  wire [24:0] p1_concat_131758_comb;
  wire [24:0] p1_concat_131759_comb;
  wire [22:0] p1_concat_131760_comb;
  wire [22:0] p1_concat_131761_comb;
  wire [24:0] p1_concat_131762_comb;
  wire [24:0] p1_concat_131763_comb;
  wire [22:0] p1_concat_131764_comb;
  wire [22:0] p1_concat_131765_comb;
  wire [24:0] p1_concat_131766_comb;
  wire [24:0] p1_concat_131767_comb;
  wire [22:0] p1_concat_131768_comb;
  wire [24:0] p1_concat_131769_comb;
  wire [22:0] p1_concat_131770_comb;
  wire [22:0] p1_concat_131771_comb;
  wire [24:0] p1_concat_131772_comb;
  wire [24:0] p1_concat_131773_comb;
  wire [22:0] p1_concat_131774_comb;
  wire [22:0] p1_concat_131775_comb;
  wire [24:0] p1_concat_131776_comb;
  wire [24:0] p1_concat_131777_comb;
  wire [22:0] p1_concat_131778_comb;
  wire [22:0] p1_concat_131779_comb;
  wire [24:0] p1_concat_131780_comb;
  wire [24:0] p1_concat_131781_comb;
  wire [22:0] p1_concat_131782_comb;
  wire [22:0] p1_concat_131783_comb;
  wire [24:0] p1_concat_131784_comb;
  wire [24:0] p1_concat_131785_comb;
  wire [24:0] p1_concat_131786_comb;
  wire [24:0] p1_concat_131787_comb;
  wire [24:0] p1_concat_131788_comb;
  wire [24:0] p1_concat_131789_comb;
  wire [24:0] p1_concat_131790_comb;
  wire [24:0] p1_concat_131791_comb;
  wire [24:0] p1_concat_131792_comb;
  wire [24:0] p1_concat_131793_comb;
  wire [24:0] p1_concat_131794_comb;
  wire [24:0] p1_concat_131795_comb;
  wire [24:0] p1_concat_131796_comb;
  wire [24:0] p1_concat_131797_comb;
  wire [24:0] p1_concat_131798_comb;
  wire [24:0] p1_concat_131799_comb;
  wire [24:0] p1_concat_131800_comb;
  wire [22:0] p1_concat_131801_comb;
  wire [24:0] p1_concat_131802_comb;
  wire [24:0] p1_concat_131803_comb;
  wire [22:0] p1_concat_131804_comb;
  wire [22:0] p1_concat_131805_comb;
  wire [24:0] p1_concat_131806_comb;
  wire [24:0] p1_concat_131807_comb;
  wire [22:0] p1_concat_131808_comb;
  wire [22:0] p1_concat_131809_comb;
  wire [24:0] p1_concat_131810_comb;
  wire [24:0] p1_concat_131811_comb;
  wire [22:0] p1_concat_131812_comb;
  wire [22:0] p1_concat_131813_comb;
  wire [24:0] p1_concat_131814_comb;
  wire [24:0] p1_concat_131815_comb;
  wire [22:0] p1_concat_131816_comb;
  wire [7:0] p1_smul_57326_TrailingBits___128_comb;
  wire [7:0] p1_smul_57326_TrailingBits___129_comb;
  wire [7:0] p1_smul_57326_TrailingBits___130_comb;
  wire [7:0] p1_smul_57326_TrailingBits___131_comb;
  wire [7:0] p1_smul_57326_TrailingBits___132_comb;
  wire [7:0] p1_smul_57326_TrailingBits___133_comb;
  wire [7:0] p1_smul_57326_TrailingBits___134_comb;
  wire [7:0] p1_smul_57326_TrailingBits___135_comb;
  wire [7:0] p1_smul_57326_TrailingBits___184_comb;
  wire [7:0] p1_smul_57326_TrailingBits___185_comb;
  wire [7:0] p1_smul_57326_TrailingBits___186_comb;
  wire [7:0] p1_smul_57326_TrailingBits___187_comb;
  wire [7:0] p1_smul_57326_TrailingBits___188_comb;
  wire [7:0] p1_smul_57326_TrailingBits___189_comb;
  wire [7:0] p1_smul_57326_TrailingBits___190_comb;
  wire [7:0] p1_smul_57326_TrailingBits___191_comb;
  wire [24:0] p1_concat_131865_comb;
  wire [22:0] p1_concat_131866_comb;
  wire [22:0] p1_concat_131867_comb;
  wire [24:0] p1_concat_131868_comb;
  wire [24:0] p1_concat_131869_comb;
  wire [22:0] p1_concat_131870_comb;
  wire [22:0] p1_concat_131871_comb;
  wire [24:0] p1_concat_131872_comb;
  wire [24:0] p1_concat_131873_comb;
  wire [24:0] p1_concat_131874_comb;
  wire [24:0] p1_concat_131875_comb;
  wire [24:0] p1_concat_131876_comb;
  wire [24:0] p1_concat_131877_comb;
  wire [24:0] p1_concat_131878_comb;
  wire [24:0] p1_concat_131879_comb;
  wire [24:0] p1_concat_131880_comb;
  wire [22:0] p1_concat_131881_comb;
  wire [24:0] p1_concat_131882_comb;
  wire [24:0] p1_concat_131883_comb;
  wire [22:0] p1_concat_131884_comb;
  wire [22:0] p1_concat_131885_comb;
  wire [24:0] p1_concat_131886_comb;
  wire [24:0] p1_concat_131887_comb;
  wire [22:0] p1_concat_131888_comb;
  wire [24:0] p1_concat_131889_comb;
  wire [22:0] p1_concat_131890_comb;
  wire [22:0] p1_concat_131891_comb;
  wire [24:0] p1_concat_131892_comb;
  wire [24:0] p1_concat_131893_comb;
  wire [22:0] p1_concat_131894_comb;
  wire [22:0] p1_concat_131895_comb;
  wire [24:0] p1_concat_131896_comb;
  wire [24:0] p1_concat_131897_comb;
  wire [24:0] p1_concat_131898_comb;
  wire [24:0] p1_concat_131899_comb;
  wire [24:0] p1_concat_131900_comb;
  wire [24:0] p1_concat_131901_comb;
  wire [24:0] p1_concat_131902_comb;
  wire [24:0] p1_concat_131903_comb;
  wire [24:0] p1_concat_131904_comb;
  wire [22:0] p1_concat_131905_comb;
  wire [24:0] p1_concat_131906_comb;
  wire [24:0] p1_concat_131907_comb;
  wire [22:0] p1_concat_131908_comb;
  wire [22:0] p1_concat_131909_comb;
  wire [24:0] p1_concat_131910_comb;
  wire [24:0] p1_concat_131911_comb;
  wire [22:0] p1_concat_131912_comb;
  wire [7:0] p1_smul_57326_TrailingBits___136_comb;
  wire [7:0] p1_smul_57326_TrailingBits___137_comb;
  wire [7:0] p1_smul_57326_TrailingBits___138_comb;
  wire [7:0] p1_smul_57326_TrailingBits___139_comb;
  wire [7:0] p1_smul_57326_TrailingBits___140_comb;
  wire [7:0] p1_smul_57326_TrailingBits___141_comb;
  wire [7:0] p1_smul_57326_TrailingBits___142_comb;
  wire [7:0] p1_smul_57326_TrailingBits___143_comb;
  wire [7:0] p1_smul_57326_TrailingBits___176_comb;
  wire [7:0] p1_smul_57326_TrailingBits___177_comb;
  wire [7:0] p1_smul_57326_TrailingBits___178_comb;
  wire [7:0] p1_smul_57326_TrailingBits___179_comb;
  wire [7:0] p1_smul_57326_TrailingBits___180_comb;
  wire [7:0] p1_smul_57326_TrailingBits___181_comb;
  wire [7:0] p1_smul_57326_TrailingBits___182_comb;
  wire [7:0] p1_smul_57326_TrailingBits___183_comb;
  wire [24:0] p1_concat_131961_comb;
  wire [22:0] p1_concat_131962_comb;
  wire [22:0] p1_concat_131963_comb;
  wire [24:0] p1_concat_131964_comb;
  wire [24:0] p1_concat_131965_comb;
  wire [22:0] p1_concat_131966_comb;
  wire [22:0] p1_concat_131967_comb;
  wire [24:0] p1_concat_131968_comb;
  wire [24:0] p1_concat_131969_comb;
  wire [24:0] p1_concat_131970_comb;
  wire [24:0] p1_concat_131971_comb;
  wire [24:0] p1_concat_131972_comb;
  wire [24:0] p1_concat_131973_comb;
  wire [24:0] p1_concat_131974_comb;
  wire [24:0] p1_concat_131975_comb;
  wire [24:0] p1_concat_131976_comb;
  wire [22:0] p1_concat_131977_comb;
  wire [24:0] p1_concat_131978_comb;
  wire [24:0] p1_concat_131979_comb;
  wire [22:0] p1_concat_131980_comb;
  wire [22:0] p1_concat_131981_comb;
  wire [24:0] p1_concat_131982_comb;
  wire [24:0] p1_concat_131983_comb;
  wire [22:0] p1_concat_131984_comb;
  wire [24:0] p1_concat_131985_comb;
  wire [22:0] p1_concat_131986_comb;
  wire [22:0] p1_concat_131987_comb;
  wire [24:0] p1_concat_131988_comb;
  wire [24:0] p1_concat_131989_comb;
  wire [22:0] p1_concat_131990_comb;
  wire [22:0] p1_concat_131991_comb;
  wire [24:0] p1_concat_131992_comb;
  wire [24:0] p1_concat_131993_comb;
  wire [24:0] p1_concat_131994_comb;
  wire [24:0] p1_concat_131995_comb;
  wire [24:0] p1_concat_131996_comb;
  wire [24:0] p1_concat_131997_comb;
  wire [24:0] p1_concat_131998_comb;
  wire [24:0] p1_concat_131999_comb;
  wire [24:0] p1_concat_132000_comb;
  wire [22:0] p1_concat_132001_comb;
  wire [24:0] p1_concat_132002_comb;
  wire [24:0] p1_concat_132003_comb;
  wire [22:0] p1_concat_132004_comb;
  wire [22:0] p1_concat_132005_comb;
  wire [24:0] p1_concat_132006_comb;
  wire [24:0] p1_concat_132007_comb;
  wire [22:0] p1_concat_132008_comb;
  wire [15:0] p1_shifted__16_comb;
  wire [7:0] p1_smul_57326_TrailingBits___16_comb;
  wire [15:0] p1_shifted__17_comb;
  wire [7:0] p1_smul_57326_TrailingBits___17_comb;
  wire [15:0] p1_shifted__18_comb;
  wire [7:0] p1_smul_57326_TrailingBits___18_comb;
  wire [15:0] p1_shifted__19_comb;
  wire [7:0] p1_smul_57326_TrailingBits___19_comb;
  wire [15:0] p1_shifted__20_comb;
  wire [7:0] p1_smul_57326_TrailingBits___20_comb;
  wire [15:0] p1_shifted__21_comb;
  wire [7:0] p1_smul_57326_TrailingBits___21_comb;
  wire [15:0] p1_shifted__22_comb;
  wire [7:0] p1_smul_57326_TrailingBits___22_comb;
  wire [15:0] p1_shifted__23_comb;
  wire [7:0] p1_smul_57326_TrailingBits___23_comb;
  wire [15:0] p1_shifted__24_comb;
  wire [7:0] p1_smul_57326_TrailingBits___24_comb;
  wire [15:0] p1_shifted__25_comb;
  wire [7:0] p1_smul_57326_TrailingBits___25_comb;
  wire [15:0] p1_shifted__26_comb;
  wire [7:0] p1_smul_57326_TrailingBits___26_comb;
  wire [15:0] p1_shifted__27_comb;
  wire [7:0] p1_smul_57326_TrailingBits___27_comb;
  wire [15:0] p1_shifted__28_comb;
  wire [7:0] p1_smul_57326_TrailingBits___28_comb;
  wire [15:0] p1_shifted__29_comb;
  wire [7:0] p1_smul_57326_TrailingBits___29_comb;
  wire [15:0] p1_shifted__30_comb;
  wire [7:0] p1_smul_57326_TrailingBits___30_comb;
  wire [15:0] p1_shifted__31_comb;
  wire [7:0] p1_smul_57326_TrailingBits___31_comb;
  wire [15:0] p1_shifted__32_comb;
  wire [7:0] p1_smul_57326_TrailingBits___32_comb;
  wire [15:0] p1_shifted__33_comb;
  wire [7:0] p1_smul_57326_TrailingBits___33_comb;
  wire [15:0] p1_shifted__34_comb;
  wire [7:0] p1_smul_57326_TrailingBits___34_comb;
  wire [15:0] p1_shifted__35_comb;
  wire [7:0] p1_smul_57326_TrailingBits___35_comb;
  wire [15:0] p1_shifted__36_comb;
  wire [7:0] p1_smul_57326_TrailingBits___36_comb;
  wire [15:0] p1_shifted__37_comb;
  wire [7:0] p1_smul_57326_TrailingBits___37_comb;
  wire [15:0] p1_shifted__38_comb;
  wire [7:0] p1_smul_57326_TrailingBits___38_comb;
  wire [15:0] p1_shifted__39_comb;
  wire [7:0] p1_smul_57326_TrailingBits___39_comb;
  wire [15:0] p1_shifted__40_comb;
  wire [7:0] p1_smul_57326_TrailingBits___40_comb;
  wire [15:0] p1_shifted__41_comb;
  wire [7:0] p1_smul_57326_TrailingBits___41_comb;
  wire [15:0] p1_shifted__42_comb;
  wire [7:0] p1_smul_57326_TrailingBits___42_comb;
  wire [15:0] p1_shifted__43_comb;
  wire [7:0] p1_smul_57326_TrailingBits___43_comb;
  wire [15:0] p1_shifted__44_comb;
  wire [7:0] p1_smul_57326_TrailingBits___44_comb;
  wire [15:0] p1_shifted__45_comb;
  wire [7:0] p1_smul_57326_TrailingBits___45_comb;
  wire [15:0] p1_shifted__46_comb;
  wire [7:0] p1_smul_57326_TrailingBits___46_comb;
  wire [15:0] p1_shifted__47_comb;
  wire [7:0] p1_smul_57326_TrailingBits___47_comb;
  wire [31:0] p1_prod__135_comb;
  wire [31:0] p1_prod__139_comb;
  wire [31:0] p1_prod__144_comb;
  wire [31:0] p1_prod__150_comb;
  wire [31:0] p1_prod__199_comb;
  wire [31:0] p1_prod__203_comb;
  wire [31:0] p1_prod__208_comb;
  wire [31:0] p1_prod__214_comb;
  wire [31:0] p1_prod__263_comb;
  wire [31:0] p1_prod__267_comb;
  wire [31:0] p1_prod__272_comb;
  wire [31:0] p1_prod__278_comb;
  wire [31:0] p1_prod__327_comb;
  wire [31:0] p1_prod__331_comb;
  wire [31:0] p1_prod__336_comb;
  wire [31:0] p1_prod__342_comb;
  wire [31:0] p1_prod__133_comb;
  wire [31:0] p1_prod__145_comb;
  wire [31:0] p1_prod__151_comb;
  wire [31:0] p1_prod__171_comb;
  wire [31:0] p1_prod__197_comb;
  wire [31:0] p1_prod__209_comb;
  wire [31:0] p1_prod__215_comb;
  wire [31:0] p1_prod__235_comb;
  wire [31:0] p1_prod__261_comb;
  wire [31:0] p1_prod__273_comb;
  wire [31:0] p1_prod__279_comb;
  wire [31:0] p1_prod__299_comb;
  wire [31:0] p1_prod__325_comb;
  wire [31:0] p1_prod__337_comb;
  wire [31:0] p1_prod__343_comb;
  wire [31:0] p1_prod__363_comb;
  wire [31:0] p1_prod__141_comb;
  wire [31:0] p1_prod__152_comb;
  wire [31:0] p1_prod__159_comb;
  wire [31:0] p1_prod__172_comb;
  wire [31:0] p1_prod__205_comb;
  wire [31:0] p1_prod__216_comb;
  wire [31:0] p1_prod__223_comb;
  wire [31:0] p1_prod__236_comb;
  wire [31:0] p1_prod__269_comb;
  wire [31:0] p1_prod__280_comb;
  wire [31:0] p1_prod__287_comb;
  wire [31:0] p1_prod__300_comb;
  wire [31:0] p1_prod__333_comb;
  wire [31:0] p1_prod__344_comb;
  wire [31:0] p1_prod__351_comb;
  wire [31:0] p1_prod__364_comb;
  wire [31:0] p1_prod__148_comb;
  wire [31:0] p1_prod__161_comb;
  wire [31:0] p1_prod__179_comb;
  wire [31:0] p1_prod__186_comb;
  wire [31:0] p1_prod__212_comb;
  wire [31:0] p1_prod__225_comb;
  wire [31:0] p1_prod__243_comb;
  wire [31:0] p1_prod__250_comb;
  wire [31:0] p1_prod__276_comb;
  wire [31:0] p1_prod__289_comb;
  wire [31:0] p1_prod__307_comb;
  wire [31:0] p1_prod__314_comb;
  wire [31:0] p1_prod__340_comb;
  wire [31:0] p1_prod__353_comb;
  wire [31:0] p1_prod__371_comb;
  wire [31:0] p1_prod__378_comb;
  wire [31:0] p1_prod__162_comb;
  wire [31:0] p1_prod__175_comb;
  wire [31:0] p1_prod__180_comb;
  wire [31:0] p1_prod__187_comb;
  wire [31:0] p1_prod__226_comb;
  wire [31:0] p1_prod__239_comb;
  wire [31:0] p1_prod__244_comb;
  wire [31:0] p1_prod__251_comb;
  wire [31:0] p1_prod__290_comb;
  wire [31:0] p1_prod__303_comb;
  wire [31:0] p1_prod__308_comb;
  wire [31:0] p1_prod__315_comb;
  wire [31:0] p1_prod__354_comb;
  wire [31:0] p1_prod__367_comb;
  wire [31:0] p1_prod__372_comb;
  wire [31:0] p1_prod__379_comb;
  wire [31:0] p1_prod__163_comb;
  wire [31:0] p1_prod__170_comb;
  wire [31:0] p1_prod__190_comb;
  wire [31:0] p1_prod__191_comb;
  wire [31:0] p1_prod__227_comb;
  wire [31:0] p1_prod__234_comb;
  wire [31:0] p1_prod__254_comb;
  wire [31:0] p1_prod__255_comb;
  wire [31:0] p1_prod__291_comb;
  wire [31:0] p1_prod__298_comb;
  wire [31:0] p1_prod__318_comb;
  wire [31:0] p1_prod__319_comb;
  wire [31:0] p1_prod__355_comb;
  wire [31:0] p1_prod__362_comb;
  wire [31:0] p1_prod__382_comb;
  wire [31:0] p1_prod__383_comb;
  wire [15:0] p1_shifted_comb;
  wire [7:0] p1_smul_57326_TrailingBits__comb;
  wire [15:0] p1_shifted__1_comb;
  wire [7:0] p1_smul_57326_TrailingBits___1_comb;
  wire [15:0] p1_shifted__2_comb;
  wire [7:0] p1_smul_57326_TrailingBits___2_comb;
  wire [15:0] p1_shifted__3_comb;
  wire [7:0] p1_smul_57326_TrailingBits___3_comb;
  wire [15:0] p1_shifted__4_comb;
  wire [7:0] p1_smul_57326_TrailingBits___4_comb;
  wire [15:0] p1_shifted__5_comb;
  wire [7:0] p1_smul_57326_TrailingBits___5_comb;
  wire [15:0] p1_shifted__6_comb;
  wire [7:0] p1_smul_57326_TrailingBits___6_comb;
  wire [15:0] p1_shifted__7_comb;
  wire [7:0] p1_smul_57326_TrailingBits___7_comb;
  wire [15:0] p1_shifted__56_comb;
  wire [7:0] p1_smul_57326_TrailingBits___56_comb;
  wire [15:0] p1_shifted__57_comb;
  wire [7:0] p1_smul_57326_TrailingBits___57_comb;
  wire [15:0] p1_shifted__58_comb;
  wire [7:0] p1_smul_57326_TrailingBits___58_comb;
  wire [15:0] p1_shifted__59_comb;
  wire [7:0] p1_smul_57326_TrailingBits___59_comb;
  wire [15:0] p1_shifted__60_comb;
  wire [7:0] p1_smul_57326_TrailingBits___60_comb;
  wire [15:0] p1_shifted__61_comb;
  wire [7:0] p1_smul_57326_TrailingBits___61_comb;
  wire [15:0] p1_shifted__62_comb;
  wire [7:0] p1_smul_57326_TrailingBits___62_comb;
  wire [15:0] p1_shifted__63_comb;
  wire [7:0] p1_smul_57326_TrailingBits___63_comb;
  wire [31:0] p1_prod__10_comb;
  wire [31:0] p1_prod__11_comb;
  wire [31:0] p1_prod__12_comb;
  wire [31:0] p1_prod__13_comb;
  wire [31:0] p1_prod__455_comb;
  wire [31:0] p1_prod__459_comb;
  wire [31:0] p1_prod__464_comb;
  wire [31:0] p1_prod__470_comb;
  wire [31:0] p1_prod__16_comb;
  wire [31:0] p1_prod__19_comb;
  wire [31:0] p1_prod__20_comb;
  wire [31:0] p1_prod__23_comb;
  wire [31:0] p1_prod__453_comb;
  wire [31:0] p1_prod__465_comb;
  wire [31:0] p1_prod__471_comb;
  wire [31:0] p1_prod__491_comb;
  wire [31:0] p1_prod__25_comb;
  wire [31:0] p1_prod__27_comb;
  wire [31:0] p1_prod__28_comb;
  wire [31:0] p1_prod__30_comb;
  wire [31:0] p1_prod__461_comb;
  wire [31:0] p1_prod__472_comb;
  wire [31:0] p1_prod__479_comb;
  wire [31:0] p1_prod__492_comb;
  wire [31:0] p1_prod__40_comb;
  wire [31:0] p1_prod__42_comb;
  wire [31:0] p1_prod__45_comb;
  wire [31:0] p1_prod__47_comb;
  wire [31:0] p1_prod__468_comb;
  wire [31:0] p1_prod__481_comb;
  wire [31:0] p1_prod__499_comb;
  wire [31:0] p1_prod__506_comb;
  wire [31:0] p1_prod__49_comb;
  wire [31:0] p1_prod__51_comb;
  wire [31:0] p1_prod__52_comb;
  wire [31:0] p1_prod__54_comb;
  wire [31:0] p1_prod__482_comb;
  wire [31:0] p1_prod__495_comb;
  wire [31:0] p1_prod__500_comb;
  wire [31:0] p1_prod__507_comb;
  wire [31:0] p1_prod__56_comb;
  wire [31:0] p1_prod__57_comb;
  wire [31:0] p1_prod__62_comb;
  wire [31:0] p1_prod__63_comb;
  wire [31:0] p1_prod__483_comb;
  wire [31:0] p1_prod__490_comb;
  wire [31:0] p1_prod__510_comb;
  wire [31:0] p1_prod__511_comb;
  wire [15:0] p1_shifted__8_comb;
  wire [7:0] p1_smul_57326_TrailingBits___8_comb;
  wire [15:0] p1_shifted__9_comb;
  wire [7:0] p1_smul_57326_TrailingBits___9_comb;
  wire [15:0] p1_shifted__10_comb;
  wire [7:0] p1_smul_57326_TrailingBits___10_comb;
  wire [15:0] p1_shifted__11_comb;
  wire [7:0] p1_smul_57326_TrailingBits___11_comb;
  wire [15:0] p1_shifted__12_comb;
  wire [7:0] p1_smul_57326_TrailingBits___12_comb;
  wire [15:0] p1_shifted__13_comb;
  wire [7:0] p1_smul_57326_TrailingBits___13_comb;
  wire [15:0] p1_shifted__14_comb;
  wire [7:0] p1_smul_57326_TrailingBits___14_comb;
  wire [15:0] p1_shifted__15_comb;
  wire [7:0] p1_smul_57326_TrailingBits___15_comb;
  wire [15:0] p1_shifted__48_comb;
  wire [7:0] p1_smul_57326_TrailingBits___48_comb;
  wire [15:0] p1_shifted__49_comb;
  wire [7:0] p1_smul_57326_TrailingBits___49_comb;
  wire [15:0] p1_shifted__50_comb;
  wire [7:0] p1_smul_57326_TrailingBits___50_comb;
  wire [15:0] p1_shifted__51_comb;
  wire [7:0] p1_smul_57326_TrailingBits___51_comb;
  wire [15:0] p1_shifted__52_comb;
  wire [7:0] p1_smul_57326_TrailingBits___52_comb;
  wire [15:0] p1_shifted__53_comb;
  wire [7:0] p1_smul_57326_TrailingBits___53_comb;
  wire [15:0] p1_shifted__54_comb;
  wire [7:0] p1_smul_57326_TrailingBits___54_comb;
  wire [15:0] p1_shifted__55_comb;
  wire [7:0] p1_smul_57326_TrailingBits___55_comb;
  wire [31:0] p1_prod__71_comb;
  wire [31:0] p1_prod__75_comb;
  wire [31:0] p1_prod__80_comb;
  wire [31:0] p1_prod__86_comb;
  wire [31:0] p1_prod__391_comb;
  wire [31:0] p1_prod__395_comb;
  wire [31:0] p1_prod__400_comb;
  wire [31:0] p1_prod__406_comb;
  wire [31:0] p1_prod__69_comb;
  wire [31:0] p1_prod__81_comb;
  wire [31:0] p1_prod__87_comb;
  wire [31:0] p1_prod__107_comb;
  wire [31:0] p1_prod__389_comb;
  wire [31:0] p1_prod__401_comb;
  wire [31:0] p1_prod__407_comb;
  wire [31:0] p1_prod__427_comb;
  wire [31:0] p1_prod__77_comb;
  wire [31:0] p1_prod__88_comb;
  wire [31:0] p1_prod__95_comb;
  wire [31:0] p1_prod__108_comb;
  wire [31:0] p1_prod__397_comb;
  wire [31:0] p1_prod__408_comb;
  wire [31:0] p1_prod__415_comb;
  wire [31:0] p1_prod__428_comb;
  wire [31:0] p1_prod__84_comb;
  wire [31:0] p1_prod__97_comb;
  wire [31:0] p1_prod__115_comb;
  wire [31:0] p1_prod__122_comb;
  wire [31:0] p1_prod__404_comb;
  wire [31:0] p1_prod__417_comb;
  wire [31:0] p1_prod__435_comb;
  wire [31:0] p1_prod__442_comb;
  wire [31:0] p1_prod__98_comb;
  wire [31:0] p1_prod__111_comb;
  wire [31:0] p1_prod__116_comb;
  wire [31:0] p1_prod__123_comb;
  wire [31:0] p1_prod__418_comb;
  wire [31:0] p1_prod__431_comb;
  wire [31:0] p1_prod__436_comb;
  wire [31:0] p1_prod__443_comb;
  wire [31:0] p1_prod__99_comb;
  wire [31:0] p1_prod__106_comb;
  wire [31:0] p1_prod__126_comb;
  wire [31:0] p1_prod__127_comb;
  wire [31:0] p1_prod__419_comb;
  wire [31:0] p1_prod__426_comb;
  wire [31:0] p1_prod__446_comb;
  wire [31:0] p1_prod__447_comb;
  wire [31:0] p1_or_132809_comb;
  wire [31:0] p1_or_132810_comb;
  wire [31:0] p1_or_132811_comb;
  wire [31:0] p1_or_132812_comb;
  wire [31:0] p1_or_132813_comb;
  wire [31:0] p1_or_132814_comb;
  wire [31:0] p1_or_132815_comb;
  wire [31:0] p1_or_132816_comb;
  wire [31:0] p1_or_132817_comb;
  wire [31:0] p1_or_132818_comb;
  wire [31:0] p1_or_132819_comb;
  wire [31:0] p1_or_132820_comb;
  wire [31:0] p1_or_132821_comb;
  wire [31:0] p1_or_132822_comb;
  wire [31:0] p1_or_132823_comb;
  wire [31:0] p1_or_132824_comb;
  wire [31:0] p1_or_132825_comb;
  wire [14:0] p1_smul_57488_NarrowedMult__comb;
  wire [14:0] p1_smul_57490_NarrowedMult__comb;
  wire [31:0] p1_or_132830_comb;
  wire [31:0] p1_or_132831_comb;
  wire [14:0] p1_smul_57496_NarrowedMult__comb;
  wire [14:0] p1_smul_57498_NarrowedMult__comb;
  wire [31:0] p1_or_132836_comb;
  wire [31:0] p1_or_132837_comb;
  wire [14:0] p1_smul_57504_NarrowedMult__comb;
  wire [14:0] p1_smul_57506_NarrowedMult__comb;
  wire [31:0] p1_or_132842_comb;
  wire [31:0] p1_or_132843_comb;
  wire [14:0] p1_smul_57512_NarrowedMult__comb;
  wire [14:0] p1_smul_57514_NarrowedMult__comb;
  wire [31:0] p1_or_132848_comb;
  wire [31:0] p1_or_132849_comb;
  wire [14:0] p1_smul_57520_NarrowedMult__comb;
  wire [14:0] p1_smul_57522_NarrowedMult__comb;
  wire [31:0] p1_or_132854_comb;
  wire [31:0] p1_or_132855_comb;
  wire [14:0] p1_smul_57528_NarrowedMult__comb;
  wire [14:0] p1_smul_57530_NarrowedMult__comb;
  wire [31:0] p1_or_132860_comb;
  wire [31:0] p1_or_132861_comb;
  wire [14:0] p1_smul_57536_NarrowedMult__comb;
  wire [14:0] p1_smul_57538_NarrowedMult__comb;
  wire [31:0] p1_or_132866_comb;
  wire [31:0] p1_or_132867_comb;
  wire [14:0] p1_smul_57544_NarrowedMult__comb;
  wire [14:0] p1_smul_57546_NarrowedMult__comb;
  wire [31:0] p1_or_132872_comb;
  wire [31:0] p1_or_132873_comb;
  wire [31:0] p1_or_132874_comb;
  wire [31:0] p1_or_132875_comb;
  wire [31:0] p1_or_132876_comb;
  wire [31:0] p1_or_132877_comb;
  wire [31:0] p1_or_132878_comb;
  wire [31:0] p1_or_132879_comb;
  wire [31:0] p1_or_132880_comb;
  wire [31:0] p1_or_132881_comb;
  wire [31:0] p1_or_132882_comb;
  wire [31:0] p1_or_132883_comb;
  wire [31:0] p1_or_132884_comb;
  wire [31:0] p1_or_132885_comb;
  wire [31:0] p1_or_132886_comb;
  wire [31:0] p1_or_132887_comb;
  wire [31:0] p1_or_132888_comb;
  wire [31:0] p1_or_132889_comb;
  wire [31:0] p1_or_132890_comb;
  wire [31:0] p1_or_132891_comb;
  wire [31:0] p1_or_132892_comb;
  wire [31:0] p1_or_132893_comb;
  wire [31:0] p1_or_132894_comb;
  wire [31:0] p1_or_132895_comb;
  wire [31:0] p1_or_132896_comb;
  wire [31:0] p1_or_132897_comb;
  wire [31:0] p1_or_132898_comb;
  wire [31:0] p1_or_132899_comb;
  wire [31:0] p1_or_132900_comb;
  wire [31:0] p1_or_132901_comb;
  wire [31:0] p1_or_132902_comb;
  wire [31:0] p1_or_132903_comb;
  wire [31:0] p1_or_132904_comb;
  wire [14:0] p1_smul_57998_NarrowedMult__comb;
  wire [31:0] p1_or_132907_comb;
  wire [14:0] p1_smul_58002_NarrowedMult__comb;
  wire [31:0] p1_or_132910_comb;
  wire [31:0] p1_or_132911_comb;
  wire [14:0] p1_smul_58008_NarrowedMult__comb;
  wire [31:0] p1_or_132914_comb;
  wire [14:0] p1_smul_58012_NarrowedMult__comb;
  wire [14:0] p1_smul_58014_NarrowedMult__comb;
  wire [31:0] p1_or_132919_comb;
  wire [14:0] p1_smul_58018_NarrowedMult__comb;
  wire [31:0] p1_or_132922_comb;
  wire [31:0] p1_or_132923_comb;
  wire [14:0] p1_smul_58024_NarrowedMult__comb;
  wire [31:0] p1_or_132926_comb;
  wire [14:0] p1_smul_58028_NarrowedMult__comb;
  wire [14:0] p1_smul_58030_NarrowedMult__comb;
  wire [31:0] p1_or_132931_comb;
  wire [14:0] p1_smul_58034_NarrowedMult__comb;
  wire [31:0] p1_or_132934_comb;
  wire [31:0] p1_or_132935_comb;
  wire [14:0] p1_smul_58040_NarrowedMult__comb;
  wire [31:0] p1_or_132938_comb;
  wire [14:0] p1_smul_58044_NarrowedMult__comb;
  wire [14:0] p1_smul_58046_NarrowedMult__comb;
  wire [31:0] p1_or_132943_comb;
  wire [14:0] p1_smul_58050_NarrowedMult__comb;
  wire [31:0] p1_or_132946_comb;
  wire [31:0] p1_or_132947_comb;
  wire [14:0] p1_smul_58056_NarrowedMult__comb;
  wire [31:0] p1_or_132950_comb;
  wire [14:0] p1_smul_58060_NarrowedMult__comb;
  wire [31:0] p1_or_132953_comb;
  wire [31:0] p1_or_132954_comb;
  wire [31:0] p1_or_132955_comb;
  wire [31:0] p1_or_132956_comb;
  wire [31:0] p1_or_132957_comb;
  wire [31:0] p1_or_132958_comb;
  wire [31:0] p1_or_132959_comb;
  wire [31:0] p1_or_132960_comb;
  wire [31:0] p1_or_132961_comb;
  wire [31:0] p1_or_132962_comb;
  wire [31:0] p1_or_132963_comb;
  wire [31:0] p1_or_132964_comb;
  wire [31:0] p1_or_132965_comb;
  wire [31:0] p1_or_132966_comb;
  wire [31:0] p1_or_132967_comb;
  wire [31:0] p1_or_132968_comb;
  wire [31:0] p1_or_133017_comb;
  wire [31:0] p1_or_133018_comb;
  wire [31:0] p1_or_133019_comb;
  wire [31:0] p1_or_133020_comb;
  wire [31:0] p1_or_133021_comb;
  wire [31:0] p1_or_133022_comb;
  wire [31:0] p1_or_133023_comb;
  wire [31:0] p1_or_133024_comb;
  wire [31:0] p1_or_133025_comb;
  wire [14:0] p1_smul_57456_NarrowedMult__comb;
  wire [14:0] p1_smul_57458_NarrowedMult__comb;
  wire [31:0] p1_or_133030_comb;
  wire [31:0] p1_or_133031_comb;
  wire [14:0] p1_smul_57464_NarrowedMult__comb;
  wire [14:0] p1_smul_57466_NarrowedMult__comb;
  wire [31:0] p1_or_133036_comb;
  wire [31:0] p1_or_133037_comb;
  wire [14:0] p1_smul_57568_NarrowedMult__comb;
  wire [14:0] p1_smul_57570_NarrowedMult__comb;
  wire [31:0] p1_or_133042_comb;
  wire [31:0] p1_or_133043_comb;
  wire [14:0] p1_smul_57576_NarrowedMult__comb;
  wire [14:0] p1_smul_57578_NarrowedMult__comb;
  wire [31:0] p1_or_133048_comb;
  wire [31:0] p1_or_133049_comb;
  wire [31:0] p1_or_133050_comb;
  wire [31:0] p1_or_133051_comb;
  wire [31:0] p1_or_133052_comb;
  wire [31:0] p1_or_133053_comb;
  wire [31:0] p1_or_133054_comb;
  wire [31:0] p1_or_133055_comb;
  wire [31:0] p1_or_133056_comb;
  wire [31:0] p1_or_133057_comb;
  wire [31:0] p1_or_133058_comb;
  wire [31:0] p1_or_133059_comb;
  wire [31:0] p1_or_133060_comb;
  wire [31:0] p1_or_133061_comb;
  wire [31:0] p1_or_133062_comb;
  wire [31:0] p1_or_133063_comb;
  wire [31:0] p1_or_133064_comb;
  wire [14:0] p1_smul_57966_NarrowedMult__comb;
  wire [31:0] p1_or_133067_comb;
  wire [14:0] p1_smul_57970_NarrowedMult__comb;
  wire [31:0] p1_or_133070_comb;
  wire [31:0] p1_or_133071_comb;
  wire [14:0] p1_smul_57976_NarrowedMult__comb;
  wire [31:0] p1_or_133074_comb;
  wire [14:0] p1_smul_57980_NarrowedMult__comb;
  wire [14:0] p1_smul_58078_NarrowedMult__comb;
  wire [31:0] p1_or_133079_comb;
  wire [14:0] p1_smul_58082_NarrowedMult__comb;
  wire [31:0] p1_or_133082_comb;
  wire [31:0] p1_or_133083_comb;
  wire [14:0] p1_smul_58088_NarrowedMult__comb;
  wire [31:0] p1_or_133086_comb;
  wire [14:0] p1_smul_58092_NarrowedMult__comb;
  wire [31:0] p1_or_133089_comb;
  wire [31:0] p1_or_133090_comb;
  wire [31:0] p1_or_133091_comb;
  wire [31:0] p1_or_133092_comb;
  wire [31:0] p1_or_133093_comb;
  wire [31:0] p1_or_133094_comb;
  wire [31:0] p1_or_133095_comb;
  wire [31:0] p1_or_133096_comb;
  wire [31:0] p1_or_133145_comb;
  wire [31:0] p1_or_133146_comb;
  wire [31:0] p1_or_133147_comb;
  wire [31:0] p1_or_133148_comb;
  wire [31:0] p1_or_133149_comb;
  wire [31:0] p1_or_133150_comb;
  wire [31:0] p1_or_133151_comb;
  wire [31:0] p1_or_133152_comb;
  wire [31:0] p1_or_133153_comb;
  wire [14:0] p1_smul_57472_NarrowedMult__comb;
  wire [14:0] p1_smul_57474_NarrowedMult__comb;
  wire [31:0] p1_or_133158_comb;
  wire [31:0] p1_or_133159_comb;
  wire [14:0] p1_smul_57480_NarrowedMult__comb;
  wire [14:0] p1_smul_57482_NarrowedMult__comb;
  wire [31:0] p1_or_133164_comb;
  wire [31:0] p1_or_133165_comb;
  wire [14:0] p1_smul_57552_NarrowedMult__comb;
  wire [14:0] p1_smul_57554_NarrowedMult__comb;
  wire [31:0] p1_or_133170_comb;
  wire [31:0] p1_or_133171_comb;
  wire [14:0] p1_smul_57560_NarrowedMult__comb;
  wire [14:0] p1_smul_57562_NarrowedMult__comb;
  wire [31:0] p1_or_133176_comb;
  wire [31:0] p1_or_133177_comb;
  wire [31:0] p1_or_133178_comb;
  wire [31:0] p1_or_133179_comb;
  wire [31:0] p1_or_133180_comb;
  wire [31:0] p1_or_133181_comb;
  wire [31:0] p1_or_133182_comb;
  wire [31:0] p1_or_133183_comb;
  wire [31:0] p1_or_133184_comb;
  wire [31:0] p1_or_133185_comb;
  wire [31:0] p1_or_133186_comb;
  wire [31:0] p1_or_133187_comb;
  wire [31:0] p1_or_133188_comb;
  wire [31:0] p1_or_133189_comb;
  wire [31:0] p1_or_133190_comb;
  wire [31:0] p1_or_133191_comb;
  wire [31:0] p1_or_133192_comb;
  wire [14:0] p1_smul_57982_NarrowedMult__comb;
  wire [31:0] p1_or_133195_comb;
  wire [14:0] p1_smul_57986_NarrowedMult__comb;
  wire [31:0] p1_or_133198_comb;
  wire [31:0] p1_or_133199_comb;
  wire [14:0] p1_smul_57992_NarrowedMult__comb;
  wire [31:0] p1_or_133202_comb;
  wire [14:0] p1_smul_57996_NarrowedMult__comb;
  wire [14:0] p1_smul_58062_NarrowedMult__comb;
  wire [31:0] p1_or_133207_comb;
  wire [14:0] p1_smul_58066_NarrowedMult__comb;
  wire [31:0] p1_or_133210_comb;
  wire [31:0] p1_or_133211_comb;
  wire [14:0] p1_smul_58072_NarrowedMult__comb;
  wire [31:0] p1_or_133214_comb;
  wire [14:0] p1_smul_58076_NarrowedMult__comb;
  wire [31:0] p1_or_133217_comb;
  wire [31:0] p1_or_133218_comb;
  wire [31:0] p1_or_133219_comb;
  wire [31:0] p1_or_133220_comb;
  wire [31:0] p1_or_133221_comb;
  wire [31:0] p1_or_133222_comb;
  wire [31:0] p1_or_133223_comb;
  wire [31:0] p1_or_133224_comb;
  wire [15:0] p1_sel_133225_comb;
  wire [15:0] p1_sel_133226_comb;
  wire [15:0] p1_sel_133227_comb;
  wire [15:0] p1_sel_133228_comb;
  wire [15:0] p1_sel_133229_comb;
  wire [15:0] p1_sel_133230_comb;
  wire [15:0] p1_sel_133231_comb;
  wire [15:0] p1_sel_133232_comb;
  wire [15:0] p1_sel_133233_comb;
  wire [15:0] p1_sel_133234_comb;
  wire [15:0] p1_sel_133235_comb;
  wire [15:0] p1_sel_133236_comb;
  wire [15:0] p1_sel_133237_comb;
  wire [15:0] p1_sel_133238_comb;
  wire [15:0] p1_sel_133239_comb;
  wire [15:0] p1_sel_133240_comb;
  wire [15:0] p1_sel_133241_comb;
  wire [15:0] p1_sel_133242_comb;
  wire [15:0] p1_sel_133243_comb;
  wire [15:0] p1_sel_133244_comb;
  wire [15:0] p1_sel_133245_comb;
  wire [15:0] p1_sel_133246_comb;
  wire [15:0] p1_sel_133247_comb;
  wire [15:0] p1_sel_133248_comb;
  wire [15:0] p1_sel_133249_comb;
  wire [15:0] p1_sel_133250_comb;
  wire [15:0] p1_sel_133251_comb;
  wire [15:0] p1_sel_133252_comb;
  wire [15:0] p1_sel_133253_comb;
  wire [15:0] p1_sel_133254_comb;
  wire [15:0] p1_sel_133255_comb;
  wire [15:0] p1_sel_133256_comb;
  wire [15:0] p1_concat_133325_comb;
  wire [15:0] p1_concat_133327_comb;
  wire [15:0] p1_concat_133337_comb;
  wire [15:0] p1_concat_133339_comb;
  wire [15:0] p1_concat_133349_comb;
  wire [15:0] p1_concat_133351_comb;
  wire [15:0] p1_concat_133361_comb;
  wire [15:0] p1_concat_133363_comb;
  wire [15:0] p1_concat_133373_comb;
  wire [15:0] p1_concat_133375_comb;
  wire [15:0] p1_concat_133385_comb;
  wire [15:0] p1_concat_133387_comb;
  wire [15:0] p1_concat_133397_comb;
  wire [15:0] p1_concat_133399_comb;
  wire [15:0] p1_concat_133409_comb;
  wire [15:0] p1_concat_133411_comb;
  wire [15:0] p1_concat_133545_comb;
  wire [15:0] p1_concat_133551_comb;
  wire [15:0] p1_concat_133561_comb;
  wire [15:0] p1_concat_133567_comb;
  wire [15:0] p1_concat_133569_comb;
  wire [15:0] p1_concat_133575_comb;
  wire [15:0] p1_concat_133585_comb;
  wire [15:0] p1_concat_133591_comb;
  wire [15:0] p1_concat_133593_comb;
  wire [15:0] p1_concat_133599_comb;
  wire [15:0] p1_concat_133609_comb;
  wire [15:0] p1_concat_133615_comb;
  wire [15:0] p1_concat_133617_comb;
  wire [15:0] p1_concat_133623_comb;
  wire [15:0] p1_concat_133633_comb;
  wire [15:0] p1_concat_133639_comb;
  wire [15:0] p1_sel_133705_comb;
  wire [15:0] p1_sel_133706_comb;
  wire [15:0] p1_sel_133707_comb;
  wire [15:0] p1_sel_133708_comb;
  wire [15:0] p1_sel_133709_comb;
  wire [15:0] p1_sel_133710_comb;
  wire [15:0] p1_sel_133711_comb;
  wire [15:0] p1_sel_133712_comb;
  wire [15:0] p1_sel_133713_comb;
  wire [15:0] p1_sel_133714_comb;
  wire [15:0] p1_sel_133715_comb;
  wire [15:0] p1_sel_133716_comb;
  wire [15:0] p1_sel_133717_comb;
  wire [15:0] p1_sel_133718_comb;
  wire [15:0] p1_sel_133719_comb;
  wire [15:0] p1_sel_133720_comb;
  wire [15:0] p1_concat_133757_comb;
  wire [15:0] p1_concat_133759_comb;
  wire [15:0] p1_concat_133769_comb;
  wire [15:0] p1_concat_133771_comb;
  wire [15:0] p1_concat_133781_comb;
  wire [15:0] p1_concat_133783_comb;
  wire [15:0] p1_concat_133793_comb;
  wire [15:0] p1_concat_133795_comb;
  wire [15:0] p1_concat_133865_comb;
  wire [15:0] p1_concat_133871_comb;
  wire [15:0] p1_concat_133881_comb;
  wire [15:0] p1_concat_133887_comb;
  wire [15:0] p1_concat_133889_comb;
  wire [15:0] p1_concat_133895_comb;
  wire [15:0] p1_concat_133905_comb;
  wire [15:0] p1_concat_133911_comb;
  wire [15:0] p1_sel_133945_comb;
  wire [15:0] p1_sel_133946_comb;
  wire [15:0] p1_sel_133947_comb;
  wire [15:0] p1_sel_133948_comb;
  wire [15:0] p1_sel_133949_comb;
  wire [15:0] p1_sel_133950_comb;
  wire [15:0] p1_sel_133951_comb;
  wire [15:0] p1_sel_133952_comb;
  wire [15:0] p1_sel_133953_comb;
  wire [15:0] p1_sel_133954_comb;
  wire [15:0] p1_sel_133955_comb;
  wire [15:0] p1_sel_133956_comb;
  wire [15:0] p1_sel_133957_comb;
  wire [15:0] p1_sel_133958_comb;
  wire [15:0] p1_sel_133959_comb;
  wire [15:0] p1_sel_133960_comb;
  wire [15:0] p1_concat_133997_comb;
  wire [15:0] p1_concat_133999_comb;
  wire [15:0] p1_concat_134009_comb;
  wire [15:0] p1_concat_134011_comb;
  wire [15:0] p1_concat_134021_comb;
  wire [15:0] p1_concat_134023_comb;
  wire [15:0] p1_concat_134033_comb;
  wire [15:0] p1_concat_134035_comb;
  wire [15:0] p1_concat_134105_comb;
  wire [15:0] p1_concat_134111_comb;
  wire [15:0] p1_concat_134121_comb;
  wire [15:0] p1_concat_134127_comb;
  wire [15:0] p1_concat_134129_comb;
  wire [15:0] p1_concat_134135_comb;
  wire [15:0] p1_concat_134145_comb;
  wire [15:0] p1_concat_134151_comb;
  wire [16:0] p1_add_135145_comb;
  wire [16:0] p1_add_135146_comb;
  wire [16:0] p1_add_135147_comb;
  wire [16:0] p1_add_135148_comb;
  wire [16:0] p1_add_135149_comb;
  wire [16:0] p1_add_135150_comb;
  wire [16:0] p1_add_135151_comb;
  wire [16:0] p1_add_135152_comb;
  wire [16:0] p1_add_135153_comb;
  wire [16:0] p1_add_135154_comb;
  wire [16:0] p1_add_135155_comb;
  wire [16:0] p1_add_135156_comb;
  wire [16:0] p1_add_135157_comb;
  wire [16:0] p1_add_135158_comb;
  wire [16:0] p1_add_135159_comb;
  wire [16:0] p1_add_135160_comb;
  wire [15:0] p1_smul_135161_comb;
  wire [15:0] p1_smul_135162_comb;
  wire [15:0] p1_sel_135163_comb;
  wire [15:0] p1_sel_135164_comb;
  wire [15:0] p1_sel_135165_comb;
  wire [15:0] p1_sel_135166_comb;
  wire [15:0] p1_smul_135167_comb;
  wire [15:0] p1_smul_135168_comb;
  wire [15:0] p1_smul_135169_comb;
  wire [15:0] p1_smul_135170_comb;
  wire [15:0] p1_sel_135171_comb;
  wire [15:0] p1_sel_135172_comb;
  wire [15:0] p1_sel_135173_comb;
  wire [15:0] p1_sel_135174_comb;
  wire [15:0] p1_smul_135175_comb;
  wire [15:0] p1_smul_135176_comb;
  wire [15:0] p1_smul_135177_comb;
  wire [15:0] p1_smul_135178_comb;
  wire [15:0] p1_sel_135179_comb;
  wire [15:0] p1_sel_135180_comb;
  wire [15:0] p1_sel_135181_comb;
  wire [15:0] p1_sel_135182_comb;
  wire [15:0] p1_smul_135183_comb;
  wire [15:0] p1_smul_135184_comb;
  wire [15:0] p1_smul_135185_comb;
  wire [15:0] p1_smul_135186_comb;
  wire [15:0] p1_sel_135187_comb;
  wire [15:0] p1_sel_135188_comb;
  wire [15:0] p1_sel_135189_comb;
  wire [15:0] p1_sel_135190_comb;
  wire [15:0] p1_smul_135191_comb;
  wire [15:0] p1_smul_135192_comb;
  wire [15:0] p1_sel_135193_comb;
  wire [15:0] p1_sel_135194_comb;
  wire [15:0] p1_sel_135195_comb;
  wire [15:0] p1_sel_135196_comb;
  wire [15:0] p1_sel_135197_comb;
  wire [15:0] p1_sel_135198_comb;
  wire [15:0] p1_sel_135199_comb;
  wire [15:0] p1_sel_135200_comb;
  wire [15:0] p1_sel_135201_comb;
  wire [15:0] p1_sel_135202_comb;
  wire [15:0] p1_sel_135203_comb;
  wire [15:0] p1_sel_135204_comb;
  wire [15:0] p1_sel_135205_comb;
  wire [15:0] p1_sel_135206_comb;
  wire [15:0] p1_sel_135207_comb;
  wire [15:0] p1_sel_135208_comb;
  wire [15:0] p1_sel_135209_comb;
  wire [15:0] p1_sel_135210_comb;
  wire [15:0] p1_sel_135211_comb;
  wire [15:0] p1_sel_135212_comb;
  wire [15:0] p1_sel_135213_comb;
  wire [15:0] p1_sel_135214_comb;
  wire [15:0] p1_sel_135215_comb;
  wire [15:0] p1_sel_135216_comb;
  wire [15:0] p1_sel_135217_comb;
  wire [15:0] p1_sel_135218_comb;
  wire [15:0] p1_sel_135219_comb;
  wire [15:0] p1_sel_135220_comb;
  wire [15:0] p1_sel_135221_comb;
  wire [15:0] p1_sel_135222_comb;
  wire [15:0] p1_sel_135223_comb;
  wire [15:0] p1_sel_135224_comb;
  wire [15:0] p1_smul_135225_comb;
  wire [15:0] p1_sel_135226_comb;
  wire [15:0] p1_smul_135227_comb;
  wire [15:0] p1_sel_135228_comb;
  wire [15:0] p1_sel_135229_comb;
  wire [15:0] p1_smul_135230_comb;
  wire [15:0] p1_sel_135231_comb;
  wire [15:0] p1_smul_135232_comb;
  wire [15:0] p1_smul_135233_comb;
  wire [15:0] p1_sel_135234_comb;
  wire [15:0] p1_smul_135235_comb;
  wire [15:0] p1_sel_135236_comb;
  wire [15:0] p1_sel_135237_comb;
  wire [15:0] p1_smul_135238_comb;
  wire [15:0] p1_sel_135239_comb;
  wire [15:0] p1_smul_135240_comb;
  wire [15:0] p1_smul_135241_comb;
  wire [15:0] p1_sel_135242_comb;
  wire [15:0] p1_smul_135243_comb;
  wire [15:0] p1_sel_135244_comb;
  wire [15:0] p1_sel_135245_comb;
  wire [15:0] p1_smul_135246_comb;
  wire [15:0] p1_sel_135247_comb;
  wire [15:0] p1_smul_135248_comb;
  wire [15:0] p1_smul_135249_comb;
  wire [15:0] p1_sel_135250_comb;
  wire [15:0] p1_smul_135251_comb;
  wire [15:0] p1_sel_135252_comb;
  wire [15:0] p1_sel_135253_comb;
  wire [15:0] p1_smul_135254_comb;
  wire [15:0] p1_sel_135255_comb;
  wire [15:0] p1_smul_135256_comb;
  wire [15:0] p1_smul_135257_comb;
  wire [15:0] p1_smul_135258_comb;
  wire [15:0] p1_smul_135259_comb;
  wire [15:0] p1_smul_135260_comb;
  wire [15:0] p1_smul_135261_comb;
  wire [15:0] p1_smul_135262_comb;
  wire [15:0] p1_smul_135263_comb;
  wire [15:0] p1_smul_135264_comb;
  wire [15:0] p1_smul_135265_comb;
  wire [15:0] p1_smul_135266_comb;
  wire [15:0] p1_smul_135267_comb;
  wire [15:0] p1_smul_135268_comb;
  wire [15:0] p1_smul_135269_comb;
  wire [15:0] p1_smul_135270_comb;
  wire [15:0] p1_smul_135271_comb;
  wire [15:0] p1_smul_135272_comb;
  wire [15:0] p1_smul_135273_comb;
  wire [15:0] p1_smul_135274_comb;
  wire [15:0] p1_smul_135275_comb;
  wire [15:0] p1_smul_135276_comb;
  wire [15:0] p1_smul_135277_comb;
  wire [15:0] p1_smul_135278_comb;
  wire [15:0] p1_smul_135279_comb;
  wire [15:0] p1_smul_135280_comb;
  wire [15:0] p1_smul_135281_comb;
  wire [15:0] p1_smul_135282_comb;
  wire [15:0] p1_smul_135283_comb;
  wire [15:0] p1_smul_135284_comb;
  wire [15:0] p1_smul_135285_comb;
  wire [15:0] p1_smul_135286_comb;
  wire [15:0] p1_smul_135287_comb;
  wire [15:0] p1_smul_135288_comb;
  wire [15:0] p1_sel_135289_comb;
  wire [15:0] p1_smul_135290_comb;
  wire [15:0] p1_sel_135291_comb;
  wire [15:0] p1_smul_135292_comb;
  wire [15:0] p1_smul_135293_comb;
  wire [15:0] p1_sel_135294_comb;
  wire [15:0] p1_smul_135295_comb;
  wire [15:0] p1_sel_135296_comb;
  wire [15:0] p1_sel_135297_comb;
  wire [15:0] p1_smul_135298_comb;
  wire [15:0] p1_sel_135299_comb;
  wire [15:0] p1_smul_135300_comb;
  wire [15:0] p1_smul_135301_comb;
  wire [15:0] p1_sel_135302_comb;
  wire [15:0] p1_smul_135303_comb;
  wire [15:0] p1_sel_135304_comb;
  wire [15:0] p1_sel_135305_comb;
  wire [15:0] p1_smul_135306_comb;
  wire [15:0] p1_sel_135307_comb;
  wire [15:0] p1_smul_135308_comb;
  wire [15:0] p1_smul_135309_comb;
  wire [15:0] p1_sel_135310_comb;
  wire [15:0] p1_smul_135311_comb;
  wire [15:0] p1_sel_135312_comb;
  wire [15:0] p1_sel_135313_comb;
  wire [15:0] p1_smul_135314_comb;
  wire [15:0] p1_sel_135315_comb;
  wire [15:0] p1_smul_135316_comb;
  wire [15:0] p1_smul_135317_comb;
  wire [15:0] p1_sel_135318_comb;
  wire [15:0] p1_smul_135319_comb;
  wire [15:0] p1_sel_135320_comb;
  wire [15:0] p1_sel_135321_comb;
  wire [15:0] p1_sel_135322_comb;
  wire [15:0] p1_sel_135323_comb;
  wire [15:0] p1_sel_135324_comb;
  wire [15:0] p1_sel_135325_comb;
  wire [15:0] p1_sel_135326_comb;
  wire [15:0] p1_sel_135327_comb;
  wire [15:0] p1_sel_135328_comb;
  wire [15:0] p1_sel_135329_comb;
  wire [15:0] p1_sel_135330_comb;
  wire [15:0] p1_sel_135331_comb;
  wire [15:0] p1_sel_135332_comb;
  wire [15:0] p1_sel_135333_comb;
  wire [15:0] p1_sel_135334_comb;
  wire [15:0] p1_sel_135335_comb;
  wire [15:0] p1_sel_135336_comb;
  wire [15:0] p1_sel_135337_comb;
  wire [15:0] p1_sel_135338_comb;
  wire [15:0] p1_sel_135339_comb;
  wire [15:0] p1_sel_135340_comb;
  wire [15:0] p1_sel_135341_comb;
  wire [15:0] p1_sel_135342_comb;
  wire [15:0] p1_sel_135343_comb;
  wire [15:0] p1_sel_135344_comb;
  wire [15:0] p1_sel_135345_comb;
  wire [15:0] p1_sel_135346_comb;
  wire [15:0] p1_sel_135347_comb;
  wire [15:0] p1_sel_135348_comb;
  wire [15:0] p1_sel_135349_comb;
  wire [15:0] p1_sel_135350_comb;
  wire [15:0] p1_sel_135351_comb;
  wire [15:0] p1_sel_135352_comb;
  wire [15:0] p1_sel_135353_comb;
  wire [15:0] p1_sel_135354_comb;
  wire [15:0] p1_smul_135355_comb;
  wire [15:0] p1_smul_135356_comb;
  wire [15:0] p1_smul_135357_comb;
  wire [15:0] p1_smul_135358_comb;
  wire [15:0] p1_sel_135359_comb;
  wire [15:0] p1_sel_135360_comb;
  wire [15:0] p1_sel_135361_comb;
  wire [15:0] p1_sel_135362_comb;
  wire [15:0] p1_smul_135363_comb;
  wire [15:0] p1_smul_135364_comb;
  wire [15:0] p1_smul_135365_comb;
  wire [15:0] p1_smul_135366_comb;
  wire [15:0] p1_sel_135367_comb;
  wire [15:0] p1_sel_135368_comb;
  wire [15:0] p1_sel_135369_comb;
  wire [15:0] p1_sel_135370_comb;
  wire [15:0] p1_smul_135371_comb;
  wire [15:0] p1_smul_135372_comb;
  wire [15:0] p1_smul_135373_comb;
  wire [15:0] p1_smul_135374_comb;
  wire [15:0] p1_sel_135375_comb;
  wire [15:0] p1_sel_135376_comb;
  wire [15:0] p1_sel_135377_comb;
  wire [15:0] p1_sel_135378_comb;
  wire [15:0] p1_smul_135379_comb;
  wire [15:0] p1_smul_135380_comb;
  wire [15:0] p1_smul_135381_comb;
  wire [15:0] p1_smul_135382_comb;
  wire [15:0] p1_sel_135383_comb;
  wire [15:0] p1_sel_135384_comb;
  wire [16:0] p1_add_135385_comb;
  wire [16:0] p1_add_135386_comb;
  wire [16:0] p1_add_135387_comb;
  wire [16:0] p1_add_135388_comb;
  wire [16:0] p1_add_135389_comb;
  wire [16:0] p1_add_135390_comb;
  wire [16:0] p1_add_135391_comb;
  wire [16:0] p1_add_135392_comb;
  wire [15:0] p1_smul_135393_comb;
  wire [15:0] p1_smul_135394_comb;
  wire [15:0] p1_sel_135395_comb;
  wire [15:0] p1_sel_135396_comb;
  wire [15:0] p1_sel_135397_comb;
  wire [15:0] p1_sel_135398_comb;
  wire [15:0] p1_smul_135399_comb;
  wire [15:0] p1_smul_135400_comb;
  wire [15:0] p1_smul_135401_comb;
  wire [15:0] p1_smul_135402_comb;
  wire [15:0] p1_sel_135403_comb;
  wire [15:0] p1_sel_135404_comb;
  wire [15:0] p1_sel_135405_comb;
  wire [15:0] p1_sel_135406_comb;
  wire [15:0] p1_smul_135407_comb;
  wire [15:0] p1_smul_135408_comb;
  wire [15:0] p1_sel_135409_comb;
  wire [15:0] p1_sel_135410_comb;
  wire [15:0] p1_sel_135411_comb;
  wire [15:0] p1_sel_135412_comb;
  wire [15:0] p1_sel_135413_comb;
  wire [15:0] p1_sel_135414_comb;
  wire [15:0] p1_sel_135415_comb;
  wire [15:0] p1_sel_135416_comb;
  wire [15:0] p1_sel_135417_comb;
  wire [15:0] p1_sel_135418_comb;
  wire [15:0] p1_sel_135419_comb;
  wire [15:0] p1_sel_135420_comb;
  wire [15:0] p1_sel_135421_comb;
  wire [15:0] p1_sel_135422_comb;
  wire [15:0] p1_sel_135423_comb;
  wire [15:0] p1_sel_135424_comb;
  wire [15:0] p1_smul_135425_comb;
  wire [15:0] p1_sel_135426_comb;
  wire [15:0] p1_smul_135427_comb;
  wire [15:0] p1_sel_135428_comb;
  wire [15:0] p1_sel_135429_comb;
  wire [15:0] p1_smul_135430_comb;
  wire [15:0] p1_sel_135431_comb;
  wire [15:0] p1_smul_135432_comb;
  wire [15:0] p1_smul_135433_comb;
  wire [15:0] p1_sel_135434_comb;
  wire [15:0] p1_smul_135435_comb;
  wire [15:0] p1_sel_135436_comb;
  wire [15:0] p1_sel_135437_comb;
  wire [15:0] p1_smul_135438_comb;
  wire [15:0] p1_sel_135439_comb;
  wire [15:0] p1_smul_135440_comb;
  wire [15:0] p1_smul_135441_comb;
  wire [15:0] p1_smul_135442_comb;
  wire [15:0] p1_smul_135443_comb;
  wire [15:0] p1_smul_135444_comb;
  wire [15:0] p1_smul_135445_comb;
  wire [15:0] p1_smul_135446_comb;
  wire [15:0] p1_smul_135447_comb;
  wire [15:0] p1_smul_135448_comb;
  wire [15:0] p1_smul_135449_comb;
  wire [15:0] p1_smul_135450_comb;
  wire [15:0] p1_smul_135451_comb;
  wire [15:0] p1_smul_135452_comb;
  wire [15:0] p1_smul_135453_comb;
  wire [15:0] p1_smul_135454_comb;
  wire [15:0] p1_smul_135455_comb;
  wire [15:0] p1_smul_135456_comb;
  wire [15:0] p1_sel_135457_comb;
  wire [15:0] p1_smul_135458_comb;
  wire [15:0] p1_sel_135459_comb;
  wire [15:0] p1_smul_135460_comb;
  wire [15:0] p1_smul_135461_comb;
  wire [15:0] p1_sel_135462_comb;
  wire [15:0] p1_smul_135463_comb;
  wire [15:0] p1_sel_135464_comb;
  wire [15:0] p1_sel_135465_comb;
  wire [15:0] p1_smul_135466_comb;
  wire [15:0] p1_sel_135467_comb;
  wire [15:0] p1_smul_135468_comb;
  wire [15:0] p1_smul_135469_comb;
  wire [15:0] p1_sel_135470_comb;
  wire [15:0] p1_smul_135471_comb;
  wire [15:0] p1_sel_135472_comb;
  wire [15:0] p1_sel_135473_comb;
  wire [15:0] p1_sel_135474_comb;
  wire [15:0] p1_sel_135475_comb;
  wire [15:0] p1_sel_135476_comb;
  wire [15:0] p1_sel_135477_comb;
  wire [15:0] p1_sel_135478_comb;
  wire [15:0] p1_sel_135479_comb;
  wire [15:0] p1_sel_135480_comb;
  wire [15:0] p1_sel_135481_comb;
  wire [15:0] p1_sel_135482_comb;
  wire [15:0] p1_sel_135483_comb;
  wire [15:0] p1_sel_135484_comb;
  wire [15:0] p1_sel_135485_comb;
  wire [15:0] p1_sel_135486_comb;
  wire [15:0] p1_sel_135487_comb;
  wire [15:0] p1_sel_135488_comb;
  wire [15:0] p1_sel_135489_comb;
  wire [15:0] p1_sel_135490_comb;
  wire [15:0] p1_smul_135491_comb;
  wire [15:0] p1_smul_135492_comb;
  wire [15:0] p1_smul_135493_comb;
  wire [15:0] p1_smul_135494_comb;
  wire [15:0] p1_sel_135495_comb;
  wire [15:0] p1_sel_135496_comb;
  wire [15:0] p1_sel_135497_comb;
  wire [15:0] p1_sel_135498_comb;
  wire [15:0] p1_smul_135499_comb;
  wire [15:0] p1_smul_135500_comb;
  wire [15:0] p1_smul_135501_comb;
  wire [15:0] p1_smul_135502_comb;
  wire [15:0] p1_sel_135503_comb;
  wire [15:0] p1_sel_135504_comb;
  wire [16:0] p1_add_135505_comb;
  wire [16:0] p1_add_135506_comb;
  wire [16:0] p1_add_135507_comb;
  wire [16:0] p1_add_135508_comb;
  wire [16:0] p1_add_135509_comb;
  wire [16:0] p1_add_135510_comb;
  wire [16:0] p1_add_135511_comb;
  wire [16:0] p1_add_135512_comb;
  wire [15:0] p1_smul_135513_comb;
  wire [15:0] p1_smul_135514_comb;
  wire [15:0] p1_sel_135515_comb;
  wire [15:0] p1_sel_135516_comb;
  wire [15:0] p1_sel_135517_comb;
  wire [15:0] p1_sel_135518_comb;
  wire [15:0] p1_smul_135519_comb;
  wire [15:0] p1_smul_135520_comb;
  wire [15:0] p1_smul_135521_comb;
  wire [15:0] p1_smul_135522_comb;
  wire [15:0] p1_sel_135523_comb;
  wire [15:0] p1_sel_135524_comb;
  wire [15:0] p1_sel_135525_comb;
  wire [15:0] p1_sel_135526_comb;
  wire [15:0] p1_smul_135527_comb;
  wire [15:0] p1_smul_135528_comb;
  wire [15:0] p1_sel_135529_comb;
  wire [15:0] p1_sel_135530_comb;
  wire [15:0] p1_sel_135531_comb;
  wire [15:0] p1_sel_135532_comb;
  wire [15:0] p1_sel_135533_comb;
  wire [15:0] p1_sel_135534_comb;
  wire [15:0] p1_sel_135535_comb;
  wire [15:0] p1_sel_135536_comb;
  wire [15:0] p1_sel_135537_comb;
  wire [15:0] p1_sel_135538_comb;
  wire [15:0] p1_sel_135539_comb;
  wire [15:0] p1_sel_135540_comb;
  wire [15:0] p1_sel_135541_comb;
  wire [15:0] p1_sel_135542_comb;
  wire [15:0] p1_sel_135543_comb;
  wire [15:0] p1_sel_135544_comb;
  wire [15:0] p1_smul_135545_comb;
  wire [15:0] p1_sel_135546_comb;
  wire [15:0] p1_smul_135547_comb;
  wire [15:0] p1_sel_135548_comb;
  wire [15:0] p1_sel_135549_comb;
  wire [15:0] p1_smul_135550_comb;
  wire [15:0] p1_sel_135551_comb;
  wire [15:0] p1_smul_135552_comb;
  wire [15:0] p1_smul_135553_comb;
  wire [15:0] p1_sel_135554_comb;
  wire [15:0] p1_smul_135555_comb;
  wire [15:0] p1_sel_135556_comb;
  wire [15:0] p1_sel_135557_comb;
  wire [15:0] p1_smul_135558_comb;
  wire [15:0] p1_sel_135559_comb;
  wire [15:0] p1_smul_135560_comb;
  wire [15:0] p1_smul_135561_comb;
  wire [15:0] p1_smul_135562_comb;
  wire [15:0] p1_smul_135563_comb;
  wire [15:0] p1_smul_135564_comb;
  wire [15:0] p1_smul_135565_comb;
  wire [15:0] p1_smul_135566_comb;
  wire [15:0] p1_smul_135567_comb;
  wire [15:0] p1_smul_135568_comb;
  wire [15:0] p1_smul_135569_comb;
  wire [15:0] p1_smul_135570_comb;
  wire [15:0] p1_smul_135571_comb;
  wire [15:0] p1_smul_135572_comb;
  wire [15:0] p1_smul_135573_comb;
  wire [15:0] p1_smul_135574_comb;
  wire [15:0] p1_smul_135575_comb;
  wire [15:0] p1_smul_135576_comb;
  wire [15:0] p1_sel_135577_comb;
  wire [15:0] p1_smul_135578_comb;
  wire [15:0] p1_sel_135579_comb;
  wire [15:0] p1_smul_135580_comb;
  wire [15:0] p1_smul_135581_comb;
  wire [15:0] p1_sel_135582_comb;
  wire [15:0] p1_smul_135583_comb;
  wire [15:0] p1_sel_135584_comb;
  wire [15:0] p1_sel_135585_comb;
  wire [15:0] p1_smul_135586_comb;
  wire [15:0] p1_sel_135587_comb;
  wire [15:0] p1_smul_135588_comb;
  wire [15:0] p1_smul_135589_comb;
  wire [15:0] p1_sel_135590_comb;
  wire [15:0] p1_smul_135591_comb;
  wire [15:0] p1_sel_135592_comb;
  wire [15:0] p1_sel_135593_comb;
  wire [15:0] p1_sel_135594_comb;
  wire [15:0] p1_sel_135595_comb;
  wire [15:0] p1_sel_135596_comb;
  wire [15:0] p1_sel_135597_comb;
  wire [15:0] p1_sel_135598_comb;
  wire [15:0] p1_sel_135599_comb;
  wire [15:0] p1_sel_135600_comb;
  wire [15:0] p1_sel_135601_comb;
  wire [15:0] p1_sel_135602_comb;
  wire [15:0] p1_sel_135603_comb;
  wire [15:0] p1_sel_135604_comb;
  wire [15:0] p1_sel_135605_comb;
  wire [15:0] p1_sel_135606_comb;
  wire [15:0] p1_sel_135607_comb;
  wire [15:0] p1_sel_135608_comb;
  wire [15:0] p1_sel_135609_comb;
  wire [15:0] p1_sel_135610_comb;
  wire [15:0] p1_smul_135611_comb;
  wire [15:0] p1_smul_135612_comb;
  wire [15:0] p1_smul_135613_comb;
  wire [15:0] p1_smul_135614_comb;
  wire [15:0] p1_sel_135615_comb;
  wire [15:0] p1_sel_135616_comb;
  wire [15:0] p1_sel_135617_comb;
  wire [15:0] p1_sel_135618_comb;
  wire [15:0] p1_smul_135619_comb;
  wire [15:0] p1_smul_135620_comb;
  wire [15:0] p1_smul_135621_comb;
  wire [15:0] p1_smul_135622_comb;
  wire [15:0] p1_sel_135623_comb;
  wire [15:0] p1_sel_135624_comb;
  wire [31:0] p1_sum__989_comb;
  wire [31:0] p1_sum__990_comb;
  wire [31:0] p1_sum__991_comb;
  wire [31:0] p1_sum__992_comb;
  wire [31:0] p1_sum__961_comb;
  wire [31:0] p1_sum__962_comb;
  wire [31:0] p1_sum__963_comb;
  wire [31:0] p1_sum__964_comb;
  wire [31:0] p1_sum__926_comb;
  wire [31:0] p1_sum__927_comb;
  wire [31:0] p1_sum__928_comb;
  wire [31:0] p1_sum__929_comb;
  wire [31:0] p1_sum__884_comb;
  wire [31:0] p1_sum__885_comb;
  wire [31:0] p1_sum__886_comb;
  wire [31:0] p1_sum__887_comb;
  wire [31:0] p1_sum__1017_comb;
  wire [31:0] p1_sum__1018_comb;
  wire [31:0] p1_sum__1019_comb;
  wire [31:0] p1_sum__1020_comb;
  wire [31:0] p1_sum__779_comb;
  wire [31:0] p1_sum__780_comb;
  wire [31:0] p1_sum__781_comb;
  wire [31:0] p1_sum__782_comb;
  wire [31:0] p1_sum__1010_comb;
  wire [31:0] p1_sum__1011_comb;
  wire [31:0] p1_sum__1012_comb;
  wire [31:0] p1_sum__1013_comb;
  wire [31:0] p1_sum__835_comb;
  wire [31:0] p1_sum__836_comb;
  wire [31:0] p1_sum__837_comb;
  wire [31:0] p1_sum__838_comb;
  wire [31:0] p1_sum__993_comb;
  wire [31:0] p1_sum__994_comb;
  wire [31:0] p1_sum__965_comb;
  wire [31:0] p1_sum__966_comb;
  wire [31:0] p1_sum__930_comb;
  wire [31:0] p1_sum__931_comb;
  wire [31:0] p1_sum__888_comb;
  wire [31:0] p1_sum__889_comb;
  wire [16:0] p1_add_136113_comb;
  wire [16:0] p1_add_136114_comb;
  wire [16:0] p1_add_136115_comb;
  wire [16:0] p1_add_136116_comb;
  wire [16:0] p1_add_136117_comb;
  wire [16:0] p1_add_136118_comb;
  wire [16:0] p1_add_136119_comb;
  wire [16:0] p1_add_136120_comb;
  wire [16:0] p1_add_136121_comb;
  wire [16:0] p1_add_136122_comb;
  wire [16:0] p1_add_136123_comb;
  wire [16:0] p1_add_136124_comb;
  wire [16:0] p1_add_136125_comb;
  wire [16:0] p1_add_136126_comb;
  wire [16:0] p1_add_136127_comb;
  wire [16:0] p1_add_136128_comb;
  wire [16:0] p1_add_136129_comb;
  wire [16:0] p1_add_136130_comb;
  wire [16:0] p1_add_136131_comb;
  wire [16:0] p1_add_136132_comb;
  wire [16:0] p1_add_136133_comb;
  wire [16:0] p1_add_136134_comb;
  wire [16:0] p1_add_136135_comb;
  wire [16:0] p1_add_136136_comb;
  wire [16:0] p1_add_136137_comb;
  wire [16:0] p1_add_136138_comb;
  wire [16:0] p1_add_136139_comb;
  wire [16:0] p1_add_136140_comb;
  wire [16:0] p1_add_136141_comb;
  wire [16:0] p1_add_136142_comb;
  wire [16:0] p1_add_136143_comb;
  wire [16:0] p1_add_136144_comb;
  wire [16:0] p1_add_136145_comb;
  wire [16:0] p1_add_136146_comb;
  wire [16:0] p1_add_136147_comb;
  wire [16:0] p1_add_136148_comb;
  wire [16:0] p1_add_136149_comb;
  wire [16:0] p1_add_136150_comb;
  wire [16:0] p1_add_136151_comb;
  wire [16:0] p1_add_136152_comb;
  wire [16:0] p1_add_136153_comb;
  wire [16:0] p1_add_136154_comb;
  wire [16:0] p1_add_136155_comb;
  wire [16:0] p1_add_136156_comb;
  wire [16:0] p1_add_136157_comb;
  wire [16:0] p1_add_136158_comb;
  wire [16:0] p1_add_136159_comb;
  wire [16:0] p1_add_136160_comb;
  wire [16:0] p1_add_136161_comb;
  wire [16:0] p1_add_136162_comb;
  wire [16:0] p1_add_136163_comb;
  wire [16:0] p1_add_136164_comb;
  wire [16:0] p1_add_136165_comb;
  wire [16:0] p1_add_136166_comb;
  wire [16:0] p1_add_136167_comb;
  wire [16:0] p1_add_136168_comb;
  wire [16:0] p1_add_136169_comb;
  wire [16:0] p1_add_136170_comb;
  wire [16:0] p1_add_136171_comb;
  wire [16:0] p1_add_136172_comb;
  wire [16:0] p1_add_136173_comb;
  wire [16:0] p1_add_136174_comb;
  wire [16:0] p1_add_136175_comb;
  wire [16:0] p1_add_136176_comb;
  wire [16:0] p1_add_136177_comb;
  wire [16:0] p1_add_136178_comb;
  wire [16:0] p1_add_136179_comb;
  wire [16:0] p1_add_136180_comb;
  wire [16:0] p1_add_136181_comb;
  wire [16:0] p1_add_136182_comb;
  wire [16:0] p1_add_136183_comb;
  wire [16:0] p1_add_136184_comb;
  wire [16:0] p1_add_136185_comb;
  wire [16:0] p1_add_136186_comb;
  wire [16:0] p1_add_136187_comb;
  wire [16:0] p1_add_136188_comb;
  wire [16:0] p1_add_136189_comb;
  wire [16:0] p1_add_136190_comb;
  wire [16:0] p1_add_136191_comb;
  wire [16:0] p1_add_136192_comb;
  wire [16:0] p1_add_136193_comb;
  wire [16:0] p1_add_136194_comb;
  wire [16:0] p1_add_136195_comb;
  wire [16:0] p1_add_136196_comb;
  wire [16:0] p1_add_136197_comb;
  wire [16:0] p1_add_136198_comb;
  wire [16:0] p1_add_136199_comb;
  wire [16:0] p1_add_136200_comb;
  wire [16:0] p1_add_136201_comb;
  wire [16:0] p1_add_136202_comb;
  wire [16:0] p1_add_136203_comb;
  wire [16:0] p1_add_136204_comb;
  wire [16:0] p1_add_136205_comb;
  wire [16:0] p1_add_136206_comb;
  wire [16:0] p1_add_136207_comb;
  wire [16:0] p1_add_136208_comb;
  wire [16:0] p1_add_136209_comb;
  wire [16:0] p1_add_136210_comb;
  wire [16:0] p1_add_136211_comb;
  wire [16:0] p1_add_136212_comb;
  wire [16:0] p1_add_136213_comb;
  wire [16:0] p1_add_136214_comb;
  wire [16:0] p1_add_136215_comb;
  wire [16:0] p1_add_136216_comb;
  wire [16:0] p1_add_136217_comb;
  wire [16:0] p1_add_136218_comb;
  wire [16:0] p1_add_136219_comb;
  wire [16:0] p1_add_136220_comb;
  wire [16:0] p1_add_136221_comb;
  wire [16:0] p1_add_136222_comb;
  wire [16:0] p1_add_136223_comb;
  wire [16:0] p1_add_136224_comb;
  wire [31:0] p1_sum__1021_comb;
  wire [31:0] p1_sum__1022_comb;
  wire [31:0] p1_sum__783_comb;
  wire [31:0] p1_sum__784_comb;
  wire [16:0] p1_add_136229_comb;
  wire [16:0] p1_add_136230_comb;
  wire [16:0] p1_add_136231_comb;
  wire [16:0] p1_add_136232_comb;
  wire [16:0] p1_add_136233_comb;
  wire [16:0] p1_add_136234_comb;
  wire [16:0] p1_add_136235_comb;
  wire [16:0] p1_add_136236_comb;
  wire [16:0] p1_add_136237_comb;
  wire [16:0] p1_add_136238_comb;
  wire [16:0] p1_add_136239_comb;
  wire [16:0] p1_add_136240_comb;
  wire [16:0] p1_add_136241_comb;
  wire [16:0] p1_add_136242_comb;
  wire [16:0] p1_add_136243_comb;
  wire [16:0] p1_add_136244_comb;
  wire [16:0] p1_add_136245_comb;
  wire [16:0] p1_add_136246_comb;
  wire [16:0] p1_add_136247_comb;
  wire [16:0] p1_add_136248_comb;
  wire [16:0] p1_add_136249_comb;
  wire [16:0] p1_add_136250_comb;
  wire [16:0] p1_add_136251_comb;
  wire [16:0] p1_add_136252_comb;
  wire [16:0] p1_add_136253_comb;
  wire [16:0] p1_add_136254_comb;
  wire [16:0] p1_add_136255_comb;
  wire [16:0] p1_add_136256_comb;
  wire [16:0] p1_add_136257_comb;
  wire [16:0] p1_add_136258_comb;
  wire [16:0] p1_add_136259_comb;
  wire [16:0] p1_add_136260_comb;
  wire [16:0] p1_add_136261_comb;
  wire [16:0] p1_add_136262_comb;
  wire [16:0] p1_add_136263_comb;
  wire [16:0] p1_add_136264_comb;
  wire [16:0] p1_add_136265_comb;
  wire [16:0] p1_add_136266_comb;
  wire [16:0] p1_add_136267_comb;
  wire [16:0] p1_add_136268_comb;
  wire [16:0] p1_add_136269_comb;
  wire [16:0] p1_add_136270_comb;
  wire [16:0] p1_add_136271_comb;
  wire [16:0] p1_add_136272_comb;
  wire [16:0] p1_add_136273_comb;
  wire [16:0] p1_add_136274_comb;
  wire [16:0] p1_add_136275_comb;
  wire [16:0] p1_add_136276_comb;
  wire [16:0] p1_add_136277_comb;
  wire [16:0] p1_add_136278_comb;
  wire [16:0] p1_add_136279_comb;
  wire [16:0] p1_add_136280_comb;
  wire [16:0] p1_add_136281_comb;
  wire [16:0] p1_add_136282_comb;
  wire [16:0] p1_add_136283_comb;
  wire [16:0] p1_add_136284_comb;
  wire [31:0] p1_sum__1014_comb;
  wire [31:0] p1_sum__1015_comb;
  wire [31:0] p1_sum__839_comb;
  wire [31:0] p1_sum__840_comb;
  wire [16:0] p1_add_136289_comb;
  wire [16:0] p1_add_136290_comb;
  wire [16:0] p1_add_136291_comb;
  wire [16:0] p1_add_136292_comb;
  wire [16:0] p1_add_136293_comb;
  wire [16:0] p1_add_136294_comb;
  wire [16:0] p1_add_136295_comb;
  wire [16:0] p1_add_136296_comb;
  wire [16:0] p1_add_136297_comb;
  wire [16:0] p1_add_136298_comb;
  wire [16:0] p1_add_136299_comb;
  wire [16:0] p1_add_136300_comb;
  wire [16:0] p1_add_136301_comb;
  wire [16:0] p1_add_136302_comb;
  wire [16:0] p1_add_136303_comb;
  wire [16:0] p1_add_136304_comb;
  wire [16:0] p1_add_136305_comb;
  wire [16:0] p1_add_136306_comb;
  wire [16:0] p1_add_136307_comb;
  wire [16:0] p1_add_136308_comb;
  wire [16:0] p1_add_136309_comb;
  wire [16:0] p1_add_136310_comb;
  wire [16:0] p1_add_136311_comb;
  wire [16:0] p1_add_136312_comb;
  wire [16:0] p1_add_136313_comb;
  wire [16:0] p1_add_136314_comb;
  wire [16:0] p1_add_136315_comb;
  wire [16:0] p1_add_136316_comb;
  wire [16:0] p1_add_136317_comb;
  wire [16:0] p1_add_136318_comb;
  wire [16:0] p1_add_136319_comb;
  wire [16:0] p1_add_136320_comb;
  wire [16:0] p1_add_136321_comb;
  wire [16:0] p1_add_136322_comb;
  wire [16:0] p1_add_136323_comb;
  wire [16:0] p1_add_136324_comb;
  wire [16:0] p1_add_136325_comb;
  wire [16:0] p1_add_136326_comb;
  wire [16:0] p1_add_136327_comb;
  wire [16:0] p1_add_136328_comb;
  wire [16:0] p1_add_136329_comb;
  wire [16:0] p1_add_136330_comb;
  wire [16:0] p1_add_136331_comb;
  wire [16:0] p1_add_136332_comb;
  wire [16:0] p1_add_136333_comb;
  wire [16:0] p1_add_136334_comb;
  wire [16:0] p1_add_136335_comb;
  wire [16:0] p1_add_136336_comb;
  wire [16:0] p1_add_136337_comb;
  wire [16:0] p1_add_136338_comb;
  wire [16:0] p1_add_136339_comb;
  wire [16:0] p1_add_136340_comb;
  wire [16:0] p1_add_136341_comb;
  wire [16:0] p1_add_136342_comb;
  wire [16:0] p1_add_136343_comb;
  wire [16:0] p1_add_136344_comb;
  wire [31:0] p1_sum__995_comb;
  wire [31:0] p1_sum__967_comb;
  wire [31:0] p1_sum__932_comb;
  wire [31:0] p1_sum__890_comb;
  wire [24:0] p1_sum__1784_comb;
  wire [24:0] p1_sum__1785_comb;
  wire [24:0] p1_sum__1786_comb;
  wire [24:0] p1_sum__1787_comb;
  wire [24:0] p1_sum__1768_comb;
  wire [24:0] p1_sum__1769_comb;
  wire [24:0] p1_sum__1770_comb;
  wire [24:0] p1_sum__1771_comb;
  wire [24:0] p1_sum__1748_comb;
  wire [24:0] p1_sum__1749_comb;
  wire [24:0] p1_sum__1750_comb;
  wire [24:0] p1_sum__1751_comb;
  wire [24:0] p1_sum__1724_comb;
  wire [24:0] p1_sum__1725_comb;
  wire [24:0] p1_sum__1726_comb;
  wire [24:0] p1_sum__1727_comb;
  wire [24:0] p1_sum__1772_comb;
  wire [24:0] p1_sum__1773_comb;
  wire [24:0] p1_sum__1774_comb;
  wire [24:0] p1_sum__1775_comb;
  wire [24:0] p1_sum__1752_comb;
  wire [24:0] p1_sum__1753_comb;
  wire [24:0] p1_sum__1754_comb;
  wire [24:0] p1_sum__1755_comb;
  wire [24:0] p1_sum__1728_comb;
  wire [24:0] p1_sum__1729_comb;
  wire [24:0] p1_sum__1730_comb;
  wire [24:0] p1_sum__1731_comb;
  wire [24:0] p1_sum__1700_comb;
  wire [24:0] p1_sum__1701_comb;
  wire [24:0] p1_sum__1702_comb;
  wire [24:0] p1_sum__1703_comb;
  wire [24:0] p1_sum__1756_comb;
  wire [24:0] p1_sum__1757_comb;
  wire [24:0] p1_sum__1758_comb;
  wire [24:0] p1_sum__1759_comb;
  wire [24:0] p1_sum__1732_comb;
  wire [24:0] p1_sum__1733_comb;
  wire [24:0] p1_sum__1734_comb;
  wire [24:0] p1_sum__1735_comb;
  wire [24:0] p1_sum__1704_comb;
  wire [24:0] p1_sum__1705_comb;
  wire [24:0] p1_sum__1706_comb;
  wire [24:0] p1_sum__1707_comb;
  wire [24:0] p1_sum__1676_comb;
  wire [24:0] p1_sum__1677_comb;
  wire [24:0] p1_sum__1678_comb;
  wire [24:0] p1_sum__1679_comb;
  wire [24:0] p1_sum__1736_comb;
  wire [24:0] p1_sum__1737_comb;
  wire [24:0] p1_sum__1738_comb;
  wire [24:0] p1_sum__1739_comb;
  wire [24:0] p1_sum__1708_comb;
  wire [24:0] p1_sum__1709_comb;
  wire [24:0] p1_sum__1710_comb;
  wire [24:0] p1_sum__1711_comb;
  wire [24:0] p1_sum__1680_comb;
  wire [24:0] p1_sum__1681_comb;
  wire [24:0] p1_sum__1682_comb;
  wire [24:0] p1_sum__1683_comb;
  wire [24:0] p1_sum__1652_comb;
  wire [24:0] p1_sum__1653_comb;
  wire [24:0] p1_sum__1654_comb;
  wire [24:0] p1_sum__1655_comb;
  wire [24:0] p1_sum__1712_comb;
  wire [24:0] p1_sum__1713_comb;
  wire [24:0] p1_sum__1714_comb;
  wire [24:0] p1_sum__1715_comb;
  wire [24:0] p1_sum__1684_comb;
  wire [24:0] p1_sum__1685_comb;
  wire [24:0] p1_sum__1686_comb;
  wire [24:0] p1_sum__1687_comb;
  wire [24:0] p1_sum__1656_comb;
  wire [24:0] p1_sum__1657_comb;
  wire [24:0] p1_sum__1658_comb;
  wire [24:0] p1_sum__1659_comb;
  wire [24:0] p1_sum__1632_comb;
  wire [24:0] p1_sum__1633_comb;
  wire [24:0] p1_sum__1634_comb;
  wire [24:0] p1_sum__1635_comb;
  wire [24:0] p1_sum__1688_comb;
  wire [24:0] p1_sum__1689_comb;
  wire [24:0] p1_sum__1690_comb;
  wire [24:0] p1_sum__1691_comb;
  wire [24:0] p1_sum__1660_comb;
  wire [24:0] p1_sum__1661_comb;
  wire [24:0] p1_sum__1662_comb;
  wire [24:0] p1_sum__1663_comb;
  wire [24:0] p1_sum__1636_comb;
  wire [24:0] p1_sum__1637_comb;
  wire [24:0] p1_sum__1638_comb;
  wire [24:0] p1_sum__1639_comb;
  wire [24:0] p1_sum__1616_comb;
  wire [24:0] p1_sum__1617_comb;
  wire [24:0] p1_sum__1618_comb;
  wire [24:0] p1_sum__1619_comb;
  wire [24:0] p1_sum__1664_comb;
  wire [24:0] p1_sum__1665_comb;
  wire [24:0] p1_sum__1666_comb;
  wire [24:0] p1_sum__1667_comb;
  wire [24:0] p1_sum__1640_comb;
  wire [24:0] p1_sum__1641_comb;
  wire [24:0] p1_sum__1642_comb;
  wire [24:0] p1_sum__1643_comb;
  wire [24:0] p1_sum__1620_comb;
  wire [24:0] p1_sum__1621_comb;
  wire [24:0] p1_sum__1622_comb;
  wire [24:0] p1_sum__1623_comb;
  wire [24:0] p1_sum__1604_comb;
  wire [24:0] p1_sum__1605_comb;
  wire [24:0] p1_sum__1606_comb;
  wire [24:0] p1_sum__1607_comb;
  wire [31:0] p1_sum__1023_comb;
  wire [31:0] p1_sum__785_comb;
  wire [24:0] p1_sum__1804_comb;
  wire [24:0] p1_sum__1805_comb;
  wire [24:0] p1_sum__1806_comb;
  wire [24:0] p1_sum__1807_comb;
  wire [24:0] p1_sum__1668_comb;
  wire [24:0] p1_sum__1669_comb;
  wire [24:0] p1_sum__1670_comb;
  wire [24:0] p1_sum__1671_comb;
  wire [24:0] p1_sum__1800_comb;
  wire [24:0] p1_sum__1801_comb;
  wire [24:0] p1_sum__1802_comb;
  wire [24:0] p1_sum__1803_comb;
  wire [24:0] p1_sum__1644_comb;
  wire [24:0] p1_sum__1645_comb;
  wire [24:0] p1_sum__1646_comb;
  wire [24:0] p1_sum__1647_comb;
  wire [24:0] p1_sum__1792_comb;
  wire [24:0] p1_sum__1793_comb;
  wire [24:0] p1_sum__1794_comb;
  wire [24:0] p1_sum__1795_comb;
  wire [24:0] p1_sum__1624_comb;
  wire [24:0] p1_sum__1625_comb;
  wire [24:0] p1_sum__1626_comb;
  wire [24:0] p1_sum__1627_comb;
  wire [24:0] p1_sum__1780_comb;
  wire [24:0] p1_sum__1781_comb;
  wire [24:0] p1_sum__1782_comb;
  wire [24:0] p1_sum__1783_comb;
  wire [24:0] p1_sum__1608_comb;
  wire [24:0] p1_sum__1609_comb;
  wire [24:0] p1_sum__1610_comb;
  wire [24:0] p1_sum__1611_comb;
  wire [24:0] p1_sum__1764_comb;
  wire [24:0] p1_sum__1765_comb;
  wire [24:0] p1_sum__1766_comb;
  wire [24:0] p1_sum__1767_comb;
  wire [24:0] p1_sum__1596_comb;
  wire [24:0] p1_sum__1597_comb;
  wire [24:0] p1_sum__1598_comb;
  wire [24:0] p1_sum__1599_comb;
  wire [24:0] p1_sum__1744_comb;
  wire [24:0] p1_sum__1745_comb;
  wire [24:0] p1_sum__1746_comb;
  wire [24:0] p1_sum__1747_comb;
  wire [24:0] p1_sum__1588_comb;
  wire [24:0] p1_sum__1589_comb;
  wire [24:0] p1_sum__1590_comb;
  wire [24:0] p1_sum__1591_comb;
  wire [24:0] p1_sum__1720_comb;
  wire [24:0] p1_sum__1721_comb;
  wire [24:0] p1_sum__1722_comb;
  wire [24:0] p1_sum__1723_comb;
  wire [24:0] p1_sum__1584_comb;
  wire [24:0] p1_sum__1585_comb;
  wire [24:0] p1_sum__1586_comb;
  wire [24:0] p1_sum__1587_comb;
  wire [31:0] p1_sum__1016_comb;
  wire [31:0] p1_sum__841_comb;
  wire [24:0] p1_sum__1796_comb;
  wire [24:0] p1_sum__1797_comb;
  wire [24:0] p1_sum__1798_comb;
  wire [24:0] p1_sum__1799_comb;
  wire [24:0] p1_sum__1696_comb;
  wire [24:0] p1_sum__1697_comb;
  wire [24:0] p1_sum__1698_comb;
  wire [24:0] p1_sum__1699_comb;
  wire [24:0] p1_sum__1788_comb;
  wire [24:0] p1_sum__1789_comb;
  wire [24:0] p1_sum__1790_comb;
  wire [24:0] p1_sum__1791_comb;
  wire [24:0] p1_sum__1672_comb;
  wire [24:0] p1_sum__1673_comb;
  wire [24:0] p1_sum__1674_comb;
  wire [24:0] p1_sum__1675_comb;
  wire [24:0] p1_sum__1776_comb;
  wire [24:0] p1_sum__1777_comb;
  wire [24:0] p1_sum__1778_comb;
  wire [24:0] p1_sum__1779_comb;
  wire [24:0] p1_sum__1648_comb;
  wire [24:0] p1_sum__1649_comb;
  wire [24:0] p1_sum__1650_comb;
  wire [24:0] p1_sum__1651_comb;
  wire [24:0] p1_sum__1760_comb;
  wire [24:0] p1_sum__1761_comb;
  wire [24:0] p1_sum__1762_comb;
  wire [24:0] p1_sum__1763_comb;
  wire [24:0] p1_sum__1628_comb;
  wire [24:0] p1_sum__1629_comb;
  wire [24:0] p1_sum__1630_comb;
  wire [24:0] p1_sum__1631_comb;
  wire [24:0] p1_sum__1740_comb;
  wire [24:0] p1_sum__1741_comb;
  wire [24:0] p1_sum__1742_comb;
  wire [24:0] p1_sum__1743_comb;
  wire [24:0] p1_sum__1612_comb;
  wire [24:0] p1_sum__1613_comb;
  wire [24:0] p1_sum__1614_comb;
  wire [24:0] p1_sum__1615_comb;
  wire [24:0] p1_sum__1716_comb;
  wire [24:0] p1_sum__1717_comb;
  wire [24:0] p1_sum__1718_comb;
  wire [24:0] p1_sum__1719_comb;
  wire [24:0] p1_sum__1600_comb;
  wire [24:0] p1_sum__1601_comb;
  wire [24:0] p1_sum__1602_comb;
  wire [24:0] p1_sum__1603_comb;
  wire [24:0] p1_sum__1692_comb;
  wire [24:0] p1_sum__1693_comb;
  wire [24:0] p1_sum__1694_comb;
  wire [24:0] p1_sum__1695_comb;
  wire [24:0] p1_sum__1592_comb;
  wire [24:0] p1_sum__1593_comb;
  wire [24:0] p1_sum__1594_comb;
  wire [24:0] p1_sum__1595_comb;
  wire [31:0] p1_umul_136585_comb;
  wire [31:0] p1_umul_136586_comb;
  wire [31:0] p1_umul_136587_comb;
  wire [31:0] p1_umul_136588_comb;
  wire [24:0] p1_sum__1348_comb;
  wire [24:0] p1_sum__1349_comb;
  wire [24:0] p1_sum__1340_comb;
  wire [24:0] p1_sum__1341_comb;
  wire [24:0] p1_sum__1330_comb;
  wire [24:0] p1_sum__1331_comb;
  wire [24:0] p1_sum__1318_comb;
  wire [24:0] p1_sum__1319_comb;
  wire [24:0] p1_sum__1342_comb;
  wire [24:0] p1_sum__1343_comb;
  wire [24:0] p1_sum__1332_comb;
  wire [24:0] p1_sum__1333_comb;
  wire [24:0] p1_sum__1320_comb;
  wire [24:0] p1_sum__1321_comb;
  wire [24:0] p1_sum__1306_comb;
  wire [24:0] p1_sum__1307_comb;
  wire [24:0] p1_sum__1334_comb;
  wire [24:0] p1_sum__1335_comb;
  wire [24:0] p1_sum__1322_comb;
  wire [24:0] p1_sum__1323_comb;
  wire [24:0] p1_sum__1308_comb;
  wire [24:0] p1_sum__1309_comb;
  wire [24:0] p1_sum__1294_comb;
  wire [24:0] p1_sum__1295_comb;
  wire [24:0] p1_sum__1324_comb;
  wire [24:0] p1_sum__1325_comb;
  wire [24:0] p1_sum__1310_comb;
  wire [24:0] p1_sum__1311_comb;
  wire [24:0] p1_sum__1296_comb;
  wire [24:0] p1_sum__1297_comb;
  wire [24:0] p1_sum__1282_comb;
  wire [24:0] p1_sum__1283_comb;
  wire [24:0] p1_sum__1312_comb;
  wire [24:0] p1_sum__1313_comb;
  wire [24:0] p1_sum__1298_comb;
  wire [24:0] p1_sum__1299_comb;
  wire [24:0] p1_sum__1284_comb;
  wire [24:0] p1_sum__1285_comb;
  wire [24:0] p1_sum__1272_comb;
  wire [24:0] p1_sum__1273_comb;
  wire [24:0] p1_sum__1300_comb;
  wire [24:0] p1_sum__1301_comb;
  wire [24:0] p1_sum__1286_comb;
  wire [24:0] p1_sum__1287_comb;
  wire [24:0] p1_sum__1274_comb;
  wire [24:0] p1_sum__1275_comb;
  wire [24:0] p1_sum__1264_comb;
  wire [24:0] p1_sum__1265_comb;
  wire [24:0] p1_sum__1288_comb;
  wire [24:0] p1_sum__1289_comb;
  wire [24:0] p1_sum__1276_comb;
  wire [24:0] p1_sum__1277_comb;
  wire [24:0] p1_sum__1266_comb;
  wire [24:0] p1_sum__1267_comb;
  wire [24:0] p1_sum__1258_comb;
  wire [24:0] p1_sum__1259_comb;
  wire [31:0] p1_umul_136645_comb;
  wire [31:0] p1_umul_136646_comb;
  wire [24:0] p1_sum__1358_comb;
  wire [24:0] p1_sum__1359_comb;
  wire [24:0] p1_sum__1290_comb;
  wire [24:0] p1_sum__1291_comb;
  wire [24:0] p1_sum__1356_comb;
  wire [24:0] p1_sum__1357_comb;
  wire [24:0] p1_sum__1278_comb;
  wire [24:0] p1_sum__1279_comb;
  wire [24:0] p1_sum__1352_comb;
  wire [24:0] p1_sum__1353_comb;
  wire [24:0] p1_sum__1268_comb;
  wire [24:0] p1_sum__1269_comb;
  wire [24:0] p1_sum__1346_comb;
  wire [24:0] p1_sum__1347_comb;
  wire [24:0] p1_sum__1260_comb;
  wire [24:0] p1_sum__1261_comb;
  wire [24:0] p1_sum__1338_comb;
  wire [24:0] p1_sum__1339_comb;
  wire [24:0] p1_sum__1254_comb;
  wire [24:0] p1_sum__1255_comb;
  wire [24:0] p1_sum__1328_comb;
  wire [24:0] p1_sum__1329_comb;
  wire [24:0] p1_sum__1250_comb;
  wire [24:0] p1_sum__1251_comb;
  wire [24:0] p1_sum__1316_comb;
  wire [24:0] p1_sum__1317_comb;
  wire [24:0] p1_sum__1248_comb;
  wire [24:0] p1_sum__1249_comb;
  wire [31:0] p1_umul_136675_comb;
  wire [31:0] p1_umul_136676_comb;
  wire [24:0] p1_sum__1354_comb;
  wire [24:0] p1_sum__1355_comb;
  wire [24:0] p1_sum__1304_comb;
  wire [24:0] p1_sum__1305_comb;
  wire [24:0] p1_sum__1350_comb;
  wire [24:0] p1_sum__1351_comb;
  wire [24:0] p1_sum__1292_comb;
  wire [24:0] p1_sum__1293_comb;
  wire [24:0] p1_sum__1344_comb;
  wire [24:0] p1_sum__1345_comb;
  wire [24:0] p1_sum__1280_comb;
  wire [24:0] p1_sum__1281_comb;
  wire [24:0] p1_sum__1336_comb;
  wire [24:0] p1_sum__1337_comb;
  wire [24:0] p1_sum__1270_comb;
  wire [24:0] p1_sum__1271_comb;
  wire [24:0] p1_sum__1326_comb;
  wire [24:0] p1_sum__1327_comb;
  wire [24:0] p1_sum__1262_comb;
  wire [24:0] p1_sum__1263_comb;
  wire [24:0] p1_sum__1314_comb;
  wire [24:0] p1_sum__1315_comb;
  wire [24:0] p1_sum__1256_comb;
  wire [24:0] p1_sum__1257_comb;
  wire [24:0] p1_sum__1302_comb;
  wire [24:0] p1_sum__1303_comb;
  wire [24:0] p1_sum__1252_comb;
  wire [24:0] p1_sum__1253_comb;
  wire [24:0] p1_sum__1130_comb;
  wire [24:0] p1_sum__1126_comb;
  wire [24:0] p1_sum__1121_comb;
  wire [24:0] p1_sum__1115_comb;
  wire [24:0] p1_sum__1127_comb;
  wire [24:0] p1_sum__1122_comb;
  wire [24:0] p1_sum__1116_comb;
  wire [24:0] p1_sum__1109_comb;
  wire [24:0] p1_sum__1123_comb;
  wire [24:0] p1_sum__1117_comb;
  wire [24:0] p1_sum__1110_comb;
  wire [24:0] p1_sum__1103_comb;
  wire [24:0] p1_sum__1118_comb;
  wire [24:0] p1_sum__1111_comb;
  wire [24:0] p1_sum__1104_comb;
  wire [24:0] p1_sum__1097_comb;
  wire [24:0] p1_sum__1112_comb;
  wire [24:0] p1_sum__1105_comb;
  wire [24:0] p1_sum__1098_comb;
  wire [24:0] p1_sum__1092_comb;
  wire [24:0] p1_sum__1106_comb;
  wire [24:0] p1_sum__1099_comb;
  wire [24:0] p1_sum__1093_comb;
  wire [24:0] p1_sum__1088_comb;
  wire [24:0] p1_sum__1100_comb;
  wire [24:0] p1_sum__1094_comb;
  wire [24:0] p1_sum__1089_comb;
  wire [24:0] p1_sum__1085_comb;
  wire [24:0] p1_sum__1135_comb;
  wire [24:0] p1_sum__1101_comb;
  wire [24:0] p1_sum__1134_comb;
  wire [24:0] p1_sum__1095_comb;
  wire [24:0] p1_sum__1132_comb;
  wire [24:0] p1_sum__1090_comb;
  wire [24:0] p1_sum__1129_comb;
  wire [24:0] p1_sum__1086_comb;
  wire [24:0] p1_sum__1125_comb;
  wire [24:0] p1_sum__1083_comb;
  wire [24:0] p1_sum__1120_comb;
  wire [24:0] p1_sum__1081_comb;
  wire [24:0] p1_sum__1114_comb;
  wire [24:0] p1_sum__1080_comb;
  wire [24:0] p1_sum__1133_comb;
  wire [24:0] p1_sum__1108_comb;
  wire [24:0] p1_sum__1131_comb;
  wire [24:0] p1_sum__1102_comb;
  wire [24:0] p1_sum__1128_comb;
  wire [24:0] p1_sum__1096_comb;
  wire [24:0] p1_sum__1124_comb;
  wire [24:0] p1_sum__1091_comb;
  wire [24:0] p1_sum__1119_comb;
  wire [24:0] p1_sum__1087_comb;
  wire [24:0] p1_sum__1113_comb;
  wire [24:0] p1_sum__1084_comb;
  wire [24:0] p1_sum__1107_comb;
  wire [24:0] p1_sum__1082_comb;
  wire [24:0] p1_add_136833_comb;
  wire [24:0] p1_add_136834_comb;
  wire [24:0] p1_add_136835_comb;
  wire [24:0] p1_add_136836_comb;
  wire [24:0] p1_add_136837_comb;
  wire [24:0] p1_add_136838_comb;
  wire [24:0] p1_add_136839_comb;
  wire [24:0] p1_add_136840_comb;
  wire [24:0] p1_add_136841_comb;
  wire [24:0] p1_add_136842_comb;
  wire [24:0] p1_add_136843_comb;
  wire [24:0] p1_add_136844_comb;
  wire [24:0] p1_add_136845_comb;
  wire [24:0] p1_add_136846_comb;
  wire [24:0] p1_add_136847_comb;
  wire [24:0] p1_add_136848_comb;
  wire [24:0] p1_add_136849_comb;
  wire [24:0] p1_add_136850_comb;
  wire [24:0] p1_add_136851_comb;
  wire [24:0] p1_add_136852_comb;
  wire [24:0] p1_add_136853_comb;
  wire [24:0] p1_add_136854_comb;
  wire [24:0] p1_add_136855_comb;
  wire [24:0] p1_add_136856_comb;
  wire [24:0] p1_add_136857_comb;
  wire [24:0] p1_add_136858_comb;
  wire [24:0] p1_add_136859_comb;
  wire [24:0] p1_add_136860_comb;
  wire [24:0] p1_add_136861_comb;
  wire [24:0] p1_add_136862_comb;
  wire [24:0] p1_add_136863_comb;
  wire [24:0] p1_add_136864_comb;
  wire [24:0] p1_add_136865_comb;
  wire [24:0] p1_add_136866_comb;
  wire [24:0] p1_add_136867_comb;
  wire [24:0] p1_add_136868_comb;
  wire [24:0] p1_add_136869_comb;
  wire [24:0] p1_add_136870_comb;
  wire [24:0] p1_add_136871_comb;
  wire [24:0] p1_add_136872_comb;
  wire [24:0] p1_add_136873_comb;
  wire [24:0] p1_add_136874_comb;
  wire [24:0] p1_add_136875_comb;
  wire [24:0] p1_add_136876_comb;
  wire [24:0] p1_add_136877_comb;
  wire [24:0] p1_add_136878_comb;
  wire [24:0] p1_add_136879_comb;
  wire [24:0] p1_add_136880_comb;
  wire [24:0] p1_add_136881_comb;
  wire [24:0] p1_add_136882_comb;
  wire [24:0] p1_add_136883_comb;
  wire [24:0] p1_add_136884_comb;
  wire [24:0] p1_add_136885_comb;
  wire [24:0] p1_add_136886_comb;
  wire [24:0] p1_add_136887_comb;
  wire [24:0] p1_add_136888_comb;
  wire [24:0] p1_add_136889_comb;
  wire [24:0] p1_add_136890_comb;
  wire [24:0] p1_add_136891_comb;
  wire [24:0] p1_add_136892_comb;
  wire [24:0] p1_add_136893_comb;
  wire [24:0] p1_add_136894_comb;
  wire [24:0] p1_add_136895_comb;
  wire [24:0] p1_add_136896_comb;
  wire [8:0] p1_clipped__256_comb;
  wire [8:0] p1_clipped__257_comb;
  wire [8:0] p1_clipped__258_comb;
  wire [8:0] p1_clipped__259_comb;
  wire [8:0] p1_clipped__260_comb;
  wire [8:0] p1_clipped__261_comb;
  wire [8:0] p1_clipped__262_comb;
  wire [8:0] p1_clipped__263_comb;
  wire [8:0] p1_clipped__264_comb;
  wire [8:0] p1_clipped__265_comb;
  wire [8:0] p1_clipped__266_comb;
  wire [8:0] p1_clipped__267_comb;
  wire [8:0] p1_clipped__268_comb;
  wire [8:0] p1_clipped__269_comb;
  wire [8:0] p1_clipped__270_comb;
  wire [8:0] p1_clipped__271_comb;
  wire [8:0] p1_clipped__272_comb;
  wire [8:0] p1_clipped__273_comb;
  wire [8:0] p1_clipped__274_comb;
  wire [8:0] p1_clipped__275_comb;
  wire [8:0] p1_clipped__276_comb;
  wire [8:0] p1_clipped__277_comb;
  wire [8:0] p1_clipped__278_comb;
  wire [8:0] p1_clipped__279_comb;
  wire [8:0] p1_clipped__280_comb;
  wire [8:0] p1_clipped__281_comb;
  wire [8:0] p1_clipped__282_comb;
  wire [8:0] p1_clipped__283_comb;
  wire [8:0] p1_clipped__284_comb;
  wire [8:0] p1_clipped__285_comb;
  wire [8:0] p1_clipped__286_comb;
  wire [8:0] p1_clipped__287_comb;
  wire [8:0] p1_clipped__288_comb;
  wire [8:0] p1_clipped__291_comb;
  wire [8:0] p1_clipped__292_comb;
  wire [8:0] p1_clipped__295_comb;
  wire [8:0] p1_clipped__296_comb;
  wire [8:0] p1_clipped__299_comb;
  wire [8:0] p1_clipped__300_comb;
  wire [8:0] p1_clipped__303_comb;
  wire [8:0] p1_clipped__304_comb;
  wire [8:0] p1_clipped__307_comb;
  wire [8:0] p1_clipped__308_comb;
  wire [8:0] p1_clipped__311_comb;
  wire [8:0] p1_clipped__312_comb;
  wire [8:0] p1_clipped__315_comb;
  wire [8:0] p1_clipped__316_comb;
  wire [8:0] p1_clipped__319_comb;
  wire [8:0] p1_clipped__289_comb;
  wire [8:0] p1_clipped__290_comb;
  wire [8:0] p1_clipped__293_comb;
  wire [8:0] p1_clipped__294_comb;
  wire [8:0] p1_clipped__297_comb;
  wire [8:0] p1_clipped__298_comb;
  wire [8:0] p1_clipped__301_comb;
  wire [8:0] p1_clipped__302_comb;
  wire [8:0] p1_clipped__305_comb;
  wire [8:0] p1_clipped__306_comb;
  wire [8:0] p1_clipped__309_comb;
  wire [8:0] p1_clipped__310_comb;
  wire [8:0] p1_clipped__313_comb;
  wire [8:0] p1_clipped__314_comb;
  wire [8:0] p1_clipped__317_comb;
  wire [8:0] p1_clipped__318_comb;
  wire [9:0] p1_add_137665_comb;
  wire [9:0] p1_add_137666_comb;
  wire [9:0] p1_add_137667_comb;
  wire [9:0] p1_add_137668_comb;
  wire [9:0] p1_add_137669_comb;
  wire [9:0] p1_add_137670_comb;
  wire [9:0] p1_add_137671_comb;
  wire [9:0] p1_add_137672_comb;
  wire [9:0] p1_add_137673_comb;
  wire [9:0] p1_add_137674_comb;
  wire [9:0] p1_add_137675_comb;
  wire [9:0] p1_add_137676_comb;
  wire [9:0] p1_add_137677_comb;
  wire [9:0] p1_add_137678_comb;
  wire [9:0] p1_add_137679_comb;
  wire [9:0] p1_add_137680_comb;
  wire [9:0] p1_add_137681_comb;
  wire [9:0] p1_add_137682_comb;
  wire [9:0] p1_add_137683_comb;
  wire [9:0] p1_add_137684_comb;
  wire [9:0] p1_add_137685_comb;
  wire [9:0] p1_add_137686_comb;
  wire [9:0] p1_add_137687_comb;
  wire [9:0] p1_add_137688_comb;
  wire [9:0] p1_add_137689_comb;
  wire [9:0] p1_add_137690_comb;
  wire [9:0] p1_add_137691_comb;
  wire [9:0] p1_add_137692_comb;
  wire [9:0] p1_add_137693_comb;
  wire [9:0] p1_add_137694_comb;
  wire [9:0] p1_add_137695_comb;
  wire [9:0] p1_add_137696_comb;
  wire [9:0] p1_add_137697_comb;
  wire [9:0] p1_add_137698_comb;
  wire [9:0] p1_add_137699_comb;
  wire [9:0] p1_add_137700_comb;
  wire [9:0] p1_add_137701_comb;
  wire [9:0] p1_add_137702_comb;
  wire [9:0] p1_add_137703_comb;
  wire [9:0] p1_add_137704_comb;
  wire [9:0] p1_add_137705_comb;
  wire [9:0] p1_add_137706_comb;
  wire [9:0] p1_add_137707_comb;
  wire [9:0] p1_add_137708_comb;
  wire [9:0] p1_add_137709_comb;
  wire [9:0] p1_add_137710_comb;
  wire [9:0] p1_add_137711_comb;
  wire [9:0] p1_add_137712_comb;
  wire [9:0] p1_add_137713_comb;
  wire [9:0] p1_add_137714_comb;
  wire [9:0] p1_add_137715_comb;
  wire [9:0] p1_add_137716_comb;
  wire [9:0] p1_add_137717_comb;
  wire [9:0] p1_add_137718_comb;
  wire [9:0] p1_add_137719_comb;
  wire [9:0] p1_add_137720_comb;
  wire [9:0] p1_add_137721_comb;
  wire [9:0] p1_add_137722_comb;
  wire [9:0] p1_add_137723_comb;
  wire [9:0] p1_add_137724_comb;
  wire [9:0] p1_add_137725_comb;
  wire [9:0] p1_add_137726_comb;
  wire [9:0] p1_add_137727_comb;
  wire [9:0] p1_add_137728_comb;
  wire [1:0] p1_bit_slice_137729_comb;
  wire [1:0] p1_bit_slice_137730_comb;
  wire [1:0] p1_bit_slice_137731_comb;
  wire [1:0] p1_bit_slice_137732_comb;
  wire [1:0] p1_bit_slice_137733_comb;
  wire [1:0] p1_bit_slice_137734_comb;
  wire [1:0] p1_bit_slice_137735_comb;
  wire [1:0] p1_bit_slice_137736_comb;
  wire [1:0] p1_bit_slice_137737_comb;
  wire [1:0] p1_bit_slice_137738_comb;
  wire [1:0] p1_bit_slice_137739_comb;
  wire [1:0] p1_bit_slice_137740_comb;
  wire [1:0] p1_bit_slice_137741_comb;
  wire [1:0] p1_bit_slice_137742_comb;
  wire [1:0] p1_bit_slice_137743_comb;
  wire [1:0] p1_bit_slice_137744_comb;
  wire [1:0] p1_bit_slice_137745_comb;
  wire [1:0] p1_bit_slice_137746_comb;
  wire [1:0] p1_bit_slice_137747_comb;
  wire [1:0] p1_bit_slice_137748_comb;
  wire [1:0] p1_bit_slice_137749_comb;
  wire [1:0] p1_bit_slice_137750_comb;
  wire [1:0] p1_bit_slice_137751_comb;
  wire [1:0] p1_bit_slice_137752_comb;
  wire [1:0] p1_bit_slice_137753_comb;
  wire [1:0] p1_bit_slice_137754_comb;
  wire [1:0] p1_bit_slice_137755_comb;
  wire [1:0] p1_bit_slice_137756_comb;
  wire [1:0] p1_bit_slice_137757_comb;
  wire [1:0] p1_bit_slice_137758_comb;
  wire [1:0] p1_bit_slice_137759_comb;
  wire [1:0] p1_bit_slice_137760_comb;
  wire [1:0] p1_bit_slice_137761_comb;
  wire [1:0] p1_bit_slice_137762_comb;
  wire [1:0] p1_bit_slice_137763_comb;
  wire [1:0] p1_bit_slice_137764_comb;
  wire [1:0] p1_bit_slice_137765_comb;
  wire [1:0] p1_bit_slice_137766_comb;
  wire [1:0] p1_bit_slice_137767_comb;
  wire [1:0] p1_bit_slice_137768_comb;
  wire [1:0] p1_bit_slice_137769_comb;
  wire [1:0] p1_bit_slice_137770_comb;
  wire [1:0] p1_bit_slice_137771_comb;
  wire [1:0] p1_bit_slice_137772_comb;
  wire [1:0] p1_bit_slice_137773_comb;
  wire [1:0] p1_bit_slice_137774_comb;
  wire [1:0] p1_bit_slice_137775_comb;
  wire [1:0] p1_bit_slice_137776_comb;
  wire [1:0] p1_bit_slice_137777_comb;
  wire [1:0] p1_bit_slice_137778_comb;
  wire [1:0] p1_bit_slice_137779_comb;
  wire [1:0] p1_bit_slice_137780_comb;
  wire [1:0] p1_bit_slice_137781_comb;
  wire [1:0] p1_bit_slice_137782_comb;
  wire [1:0] p1_bit_slice_137783_comb;
  wire [1:0] p1_bit_slice_137784_comb;
  wire [1:0] p1_bit_slice_137785_comb;
  wire [1:0] p1_bit_slice_137786_comb;
  wire [1:0] p1_bit_slice_137787_comb;
  wire [1:0] p1_bit_slice_137788_comb;
  wire [1:0] p1_bit_slice_137789_comb;
  wire [1:0] p1_bit_slice_137790_comb;
  wire [1:0] p1_bit_slice_137791_comb;
  wire [1:0] p1_bit_slice_137792_comb;
  wire [2:0] p1_add_137921_comb;
  wire [2:0] p1_add_137922_comb;
  wire [2:0] p1_add_137923_comb;
  wire [2:0] p1_add_137924_comb;
  wire [2:0] p1_add_137925_comb;
  wire [2:0] p1_add_137926_comb;
  wire [2:0] p1_add_137927_comb;
  wire [2:0] p1_add_137928_comb;
  wire [2:0] p1_add_137929_comb;
  wire [2:0] p1_add_137930_comb;
  wire [2:0] p1_add_137931_comb;
  wire [2:0] p1_add_137932_comb;
  wire [2:0] p1_add_137933_comb;
  wire [2:0] p1_add_137934_comb;
  wire [2:0] p1_add_137935_comb;
  wire [2:0] p1_add_137936_comb;
  wire [2:0] p1_add_137937_comb;
  wire [2:0] p1_add_137938_comb;
  wire [2:0] p1_add_137939_comb;
  wire [2:0] p1_add_137940_comb;
  wire [2:0] p1_add_137941_comb;
  wire [2:0] p1_add_137942_comb;
  wire [2:0] p1_add_137943_comb;
  wire [2:0] p1_add_137944_comb;
  wire [2:0] p1_add_137945_comb;
  wire [2:0] p1_add_137946_comb;
  wire [2:0] p1_add_137947_comb;
  wire [2:0] p1_add_137948_comb;
  wire [2:0] p1_add_137949_comb;
  wire [2:0] p1_add_137950_comb;
  wire [2:0] p1_add_137951_comb;
  wire [2:0] p1_add_137952_comb;
  wire [2:0] p1_add_137953_comb;
  wire [2:0] p1_add_137954_comb;
  wire [2:0] p1_add_137955_comb;
  wire [2:0] p1_add_137956_comb;
  wire [2:0] p1_add_137957_comb;
  wire [2:0] p1_add_137958_comb;
  wire [2:0] p1_add_137959_comb;
  wire [2:0] p1_add_137960_comb;
  wire [2:0] p1_add_137961_comb;
  wire [2:0] p1_add_137962_comb;
  wire [2:0] p1_add_137963_comb;
  wire [2:0] p1_add_137964_comb;
  wire [2:0] p1_add_137965_comb;
  wire [2:0] p1_add_137966_comb;
  wire [2:0] p1_add_137967_comb;
  wire [2:0] p1_add_137968_comb;
  wire [2:0] p1_add_137969_comb;
  wire [2:0] p1_add_137970_comb;
  wire [2:0] p1_add_137971_comb;
  wire [2:0] p1_add_137972_comb;
  wire [2:0] p1_add_137973_comb;
  wire [2:0] p1_add_137974_comb;
  wire [2:0] p1_add_137975_comb;
  wire [2:0] p1_add_137976_comb;
  wire [2:0] p1_add_137977_comb;
  wire [2:0] p1_add_137978_comb;
  wire [2:0] p1_add_137979_comb;
  wire [2:0] p1_add_137980_comb;
  wire [2:0] p1_add_137981_comb;
  wire [2:0] p1_add_137982_comb;
  wire [2:0] p1_add_137983_comb;
  wire [2:0] p1_add_137984_comb;
  wire [7:0] p1_clipped__40_comb;
  wire [7:0] p1_clipped__56_comb;
  wire [7:0] p1_clipped__72_comb;
  wire [7:0] p1_clipped__88_comb;
  wire [7:0] p1_clipped__41_comb;
  wire [7:0] p1_clipped__57_comb;
  wire [7:0] p1_clipped__73_comb;
  wire [7:0] p1_clipped__89_comb;
  wire [7:0] p1_clipped__42_comb;
  wire [7:0] p1_clipped__58_comb;
  wire [7:0] p1_clipped__74_comb;
  wire [7:0] p1_clipped__90_comb;
  wire [7:0] p1_clipped__43_comb;
  wire [7:0] p1_clipped__59_comb;
  wire [7:0] p1_clipped__75_comb;
  wire [7:0] p1_clipped__91_comb;
  wire [7:0] p1_clipped__44_comb;
  wire [7:0] p1_clipped__60_comb;
  wire [7:0] p1_clipped__76_comb;
  wire [7:0] p1_clipped__92_comb;
  wire [7:0] p1_clipped__45_comb;
  wire [7:0] p1_clipped__61_comb;
  wire [7:0] p1_clipped__77_comb;
  wire [7:0] p1_clipped__93_comb;
  wire [7:0] p1_clipped__46_comb;
  wire [7:0] p1_clipped__62_comb;
  wire [7:0] p1_clipped__78_comb;
  wire [7:0] p1_clipped__94_comb;
  wire [7:0] p1_clipped__47_comb;
  wire [7:0] p1_clipped__63_comb;
  wire [7:0] p1_clipped__79_comb;
  wire [7:0] p1_clipped__95_comb;
  wire [7:0] p1_clipped__8_comb;
  wire [7:0] p1_clipped__120_comb;
  wire [7:0] p1_clipped__9_comb;
  wire [7:0] p1_clipped__121_comb;
  wire [7:0] p1_clipped__10_comb;
  wire [7:0] p1_clipped__122_comb;
  wire [7:0] p1_clipped__11_comb;
  wire [7:0] p1_clipped__123_comb;
  wire [7:0] p1_clipped__12_comb;
  wire [7:0] p1_clipped__124_comb;
  wire [7:0] p1_clipped__13_comb;
  wire [7:0] p1_clipped__125_comb;
  wire [7:0] p1_clipped__14_comb;
  wire [7:0] p1_clipped__126_comb;
  wire [7:0] p1_clipped__15_comb;
  wire [7:0] p1_clipped__127_comb;
  wire [7:0] p1_clipped__24_comb;
  wire [7:0] p1_clipped__104_comb;
  wire [7:0] p1_clipped__25_comb;
  wire [7:0] p1_clipped__105_comb;
  wire [7:0] p1_clipped__26_comb;
  wire [7:0] p1_clipped__106_comb;
  wire [7:0] p1_clipped__27_comb;
  wire [7:0] p1_clipped__107_comb;
  wire [7:0] p1_clipped__28_comb;
  wire [7:0] p1_clipped__108_comb;
  wire [7:0] p1_clipped__29_comb;
  wire [7:0] p1_clipped__109_comb;
  wire [7:0] p1_clipped__30_comb;
  wire [7:0] p1_clipped__110_comb;
  wire [7:0] p1_clipped__31_comb;
  wire [7:0] p1_clipped__111_comb;
  wire [7:0] p1_shifted__66_squeezed_comb;
  wire [7:0] p1_shifted__67_squeezed_comb;
  wire [7:0] p1_shifted__68_squeezed_comb;
  wire [7:0] p1_shifted__69_squeezed_comb;
  wire [7:0] p1_shifted__74_squeezed_comb;
  wire [7:0] p1_shifted__75_squeezed_comb;
  wire [7:0] p1_shifted__76_squeezed_comb;
  wire [7:0] p1_shifted__77_squeezed_comb;
  wire [7:0] p1_shifted__82_squeezed_comb;
  wire [7:0] p1_shifted__83_squeezed_comb;
  wire [7:0] p1_shifted__84_squeezed_comb;
  wire [7:0] p1_shifted__85_squeezed_comb;
  wire [7:0] p1_shifted__90_squeezed_comb;
  wire [7:0] p1_shifted__91_squeezed_comb;
  wire [7:0] p1_shifted__92_squeezed_comb;
  wire [7:0] p1_shifted__93_squeezed_comb;
  wire [7:0] p1_shifted__98_squeezed_comb;
  wire [7:0] p1_shifted__99_squeezed_comb;
  wire [7:0] p1_shifted__100_squeezed_comb;
  wire [7:0] p1_shifted__101_squeezed_comb;
  wire [7:0] p1_shifted__106_squeezed_comb;
  wire [7:0] p1_shifted__107_squeezed_comb;
  wire [7:0] p1_shifted__108_squeezed_comb;
  wire [7:0] p1_shifted__109_squeezed_comb;
  wire [7:0] p1_shifted__114_squeezed_comb;
  wire [7:0] p1_shifted__115_squeezed_comb;
  wire [7:0] p1_shifted__116_squeezed_comb;
  wire [7:0] p1_shifted__117_squeezed_comb;
  wire [7:0] p1_shifted__122_squeezed_comb;
  wire [7:0] p1_shifted__123_squeezed_comb;
  wire [7:0] p1_shifted__124_squeezed_comb;
  wire [7:0] p1_shifted__125_squeezed_comb;
  wire [7:0] p1_shifted__64_squeezed_comb;
  wire [7:0] p1_shifted__71_squeezed_comb;
  wire [7:0] p1_shifted__72_squeezed_comb;
  wire [7:0] p1_shifted__79_squeezed_comb;
  wire [7:0] p1_shifted__80_squeezed_comb;
  wire [7:0] p1_shifted__87_squeezed_comb;
  wire [7:0] p1_shifted__88_squeezed_comb;
  wire [7:0] p1_shifted__95_squeezed_comb;
  wire [7:0] p1_shifted__96_squeezed_comb;
  wire [7:0] p1_shifted__103_squeezed_comb;
  wire [7:0] p1_shifted__104_squeezed_comb;
  wire [7:0] p1_shifted__111_squeezed_comb;
  wire [7:0] p1_shifted__112_squeezed_comb;
  wire [7:0] p1_shifted__119_squeezed_comb;
  wire [7:0] p1_shifted__120_squeezed_comb;
  wire [7:0] p1_shifted__127_squeezed_comb;
  wire [7:0] p1_shifted__65_squeezed_comb;
  wire [7:0] p1_shifted__70_squeezed_comb;
  wire [7:0] p1_shifted__73_squeezed_comb;
  wire [7:0] p1_shifted__78_squeezed_comb;
  wire [7:0] p1_shifted__81_squeezed_comb;
  wire [7:0] p1_shifted__86_squeezed_comb;
  wire [7:0] p1_shifted__89_squeezed_comb;
  wire [7:0] p1_shifted__94_squeezed_comb;
  wire [7:0] p1_shifted__97_squeezed_comb;
  wire [7:0] p1_shifted__102_squeezed_comb;
  wire [7:0] p1_shifted__105_squeezed_comb;
  wire [7:0] p1_shifted__110_squeezed_comb;
  wire [7:0] p1_shifted__113_squeezed_comb;
  wire [7:0] p1_shifted__118_squeezed_comb;
  wire [7:0] p1_shifted__121_squeezed_comb;
  wire [7:0] p1_shifted__126_squeezed_comb;
  wire [15:0] p1_smul_58226_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___128_comb;
  wire [13:0] p1_smul_58228_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___129_comb;
  wire [13:0] p1_smul_58230_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___130_comb;
  wire [15:0] p1_smul_58232_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___131_comb;
  wire [15:0] p1_smul_58242_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___132_comb;
  wire [13:0] p1_smul_58244_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___133_comb;
  wire [13:0] p1_smul_58246_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___134_comb;
  wire [15:0] p1_smul_58248_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___135_comb;
  wire [15:0] p1_smul_58258_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___136_comb;
  wire [13:0] p1_smul_58260_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___137_comb;
  wire [13:0] p1_smul_58262_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___138_comb;
  wire [15:0] p1_smul_58264_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___139_comb;
  wire [15:0] p1_smul_58274_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___140_comb;
  wire [13:0] p1_smul_58276_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___141_comb;
  wire [13:0] p1_smul_58278_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___142_comb;
  wire [15:0] p1_smul_58280_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___143_comb;
  wire [15:0] p1_smul_58290_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___144_comb;
  wire [13:0] p1_smul_58292_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___145_comb;
  wire [13:0] p1_smul_58294_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___146_comb;
  wire [15:0] p1_smul_58296_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___147_comb;
  wire [15:0] p1_smul_58306_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___148_comb;
  wire [13:0] p1_smul_58308_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___149_comb;
  wire [13:0] p1_smul_58310_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___150_comb;
  wire [15:0] p1_smul_58312_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___151_comb;
  wire [15:0] p1_smul_58322_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___152_comb;
  wire [13:0] p1_smul_58324_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___153_comb;
  wire [13:0] p1_smul_58326_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___154_comb;
  wire [15:0] p1_smul_58328_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___155_comb;
  wire [15:0] p1_smul_58338_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___156_comb;
  wire [13:0] p1_smul_58340_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___157_comb;
  wire [13:0] p1_smul_58342_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___158_comb;
  wire [15:0] p1_smul_58344_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___159_comb;
  wire [14:0] p1_smul_58350_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___64_comb;
  wire [14:0] p1_smul_58356_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___65_comb;
  wire [14:0] p1_smul_58358_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___66_comb;
  wire [14:0] p1_smul_58364_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___67_comb;
  wire [14:0] p1_smul_58366_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___68_comb;
  wire [14:0] p1_smul_58372_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___69_comb;
  wire [14:0] p1_smul_58374_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___70_comb;
  wire [14:0] p1_smul_58380_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___71_comb;
  wire [14:0] p1_smul_58382_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___72_comb;
  wire [14:0] p1_smul_58388_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___73_comb;
  wire [14:0] p1_smul_58390_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___74_comb;
  wire [14:0] p1_smul_58396_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___75_comb;
  wire [14:0] p1_smul_58398_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___76_comb;
  wire [14:0] p1_smul_58404_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___77_comb;
  wire [14:0] p1_smul_58406_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___78_comb;
  wire [14:0] p1_smul_58412_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___79_comb;
  wire [14:0] p1_smul_58414_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___80_comb;
  wire [14:0] p1_smul_58420_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___81_comb;
  wire [14:0] p1_smul_58422_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___82_comb;
  wire [14:0] p1_smul_58428_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___83_comb;
  wire [14:0] p1_smul_58430_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___84_comb;
  wire [14:0] p1_smul_58436_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___85_comb;
  wire [14:0] p1_smul_58438_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___86_comb;
  wire [14:0] p1_smul_58444_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___87_comb;
  wire [14:0] p1_smul_58446_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___88_comb;
  wire [14:0] p1_smul_58452_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___89_comb;
  wire [14:0] p1_smul_58454_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___90_comb;
  wire [14:0] p1_smul_58460_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___91_comb;
  wire [14:0] p1_smul_58462_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___92_comb;
  wire [14:0] p1_smul_58468_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___93_comb;
  wire [14:0] p1_smul_58470_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___94_comb;
  wire [14:0] p1_smul_58476_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___95_comb;
  wire [13:0] p1_smul_58480_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___160_comb;
  wire [15:0] p1_smul_58484_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___161_comb;
  wire [15:0] p1_smul_58486_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___162_comb;
  wire [13:0] p1_smul_58490_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___163_comb;
  wire [13:0] p1_smul_58496_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___164_comb;
  wire [15:0] p1_smul_58500_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___165_comb;
  wire [15:0] p1_smul_58502_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___166_comb;
  wire [13:0] p1_smul_58506_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___167_comb;
  wire [13:0] p1_smul_58512_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___168_comb;
  wire [15:0] p1_smul_58516_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___169_comb;
  wire [15:0] p1_smul_58518_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___170_comb;
  wire [13:0] p1_smul_58522_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___171_comb;
  wire [13:0] p1_smul_58528_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___172_comb;
  wire [15:0] p1_smul_58532_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___173_comb;
  wire [15:0] p1_smul_58534_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___174_comb;
  wire [13:0] p1_smul_58538_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___175_comb;
  wire [13:0] p1_smul_58544_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___176_comb;
  wire [15:0] p1_smul_58548_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___177_comb;
  wire [15:0] p1_smul_58550_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___178_comb;
  wire [13:0] p1_smul_58554_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___179_comb;
  wire [13:0] p1_smul_58560_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___180_comb;
  wire [15:0] p1_smul_58564_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___181_comb;
  wire [15:0] p1_smul_58566_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___182_comb;
  wire [13:0] p1_smul_58570_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___183_comb;
  wire [13:0] p1_smul_58576_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___184_comb;
  wire [15:0] p1_smul_58580_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___185_comb;
  wire [15:0] p1_smul_58582_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___186_comb;
  wire [13:0] p1_smul_58586_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___187_comb;
  wire [13:0] p1_smul_58592_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___188_comb;
  wire [15:0] p1_smul_58596_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___189_comb;
  wire [15:0] p1_smul_58598_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___190_comb;
  wire [13:0] p1_smul_58602_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___191_comb;
  wire [15:0] p1_smul_58734_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___192_comb;
  wire [13:0] p1_smul_58738_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___193_comb;
  wire [13:0] p1_smul_58744_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___194_comb;
  wire [15:0] p1_smul_58748_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___195_comb;
  wire [15:0] p1_smul_58750_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___196_comb;
  wire [13:0] p1_smul_58754_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___197_comb;
  wire [13:0] p1_smul_58760_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___198_comb;
  wire [15:0] p1_smul_58764_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___199_comb;
  wire [15:0] p1_smul_58766_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___200_comb;
  wire [13:0] p1_smul_58770_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___201_comb;
  wire [13:0] p1_smul_58776_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___202_comb;
  wire [15:0] p1_smul_58780_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___203_comb;
  wire [15:0] p1_smul_58782_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___204_comb;
  wire [13:0] p1_smul_58786_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___205_comb;
  wire [13:0] p1_smul_58792_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___206_comb;
  wire [15:0] p1_smul_58796_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___207_comb;
  wire [15:0] p1_smul_58798_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___208_comb;
  wire [13:0] p1_smul_58802_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___209_comb;
  wire [13:0] p1_smul_58808_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___210_comb;
  wire [15:0] p1_smul_58812_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___211_comb;
  wire [15:0] p1_smul_58814_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___212_comb;
  wire [13:0] p1_smul_58818_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___213_comb;
  wire [13:0] p1_smul_58824_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___214_comb;
  wire [15:0] p1_smul_58828_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___215_comb;
  wire [15:0] p1_smul_58830_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___216_comb;
  wire [13:0] p1_smul_58834_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___217_comb;
  wire [13:0] p1_smul_58840_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___218_comb;
  wire [15:0] p1_smul_58844_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___219_comb;
  wire [15:0] p1_smul_58846_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___220_comb;
  wire [13:0] p1_smul_58850_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___221_comb;
  wire [13:0] p1_smul_58856_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___222_comb;
  wire [15:0] p1_smul_58860_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___223_comb;
  wire [14:0] p1_smul_58864_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___96_comb;
  wire [14:0] p1_smul_58868_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___97_comb;
  wire [14:0] p1_smul_58870_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___98_comb;
  wire [14:0] p1_smul_58874_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___99_comb;
  wire [14:0] p1_smul_58880_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___100_comb;
  wire [14:0] p1_smul_58884_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___101_comb;
  wire [14:0] p1_smul_58886_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___102_comb;
  wire [14:0] p1_smul_58890_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___103_comb;
  wire [14:0] p1_smul_58896_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___104_comb;
  wire [14:0] p1_smul_58900_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___105_comb;
  wire [14:0] p1_smul_58902_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___106_comb;
  wire [14:0] p1_smul_58906_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___107_comb;
  wire [14:0] p1_smul_58912_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___108_comb;
  wire [14:0] p1_smul_58916_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___109_comb;
  wire [14:0] p1_smul_58918_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___110_comb;
  wire [14:0] p1_smul_58922_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___111_comb;
  wire [14:0] p1_smul_58928_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___112_comb;
  wire [14:0] p1_smul_58932_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___113_comb;
  wire [14:0] p1_smul_58934_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___114_comb;
  wire [14:0] p1_smul_58938_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___115_comb;
  wire [14:0] p1_smul_58944_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___116_comb;
  wire [14:0] p1_smul_58948_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___117_comb;
  wire [14:0] p1_smul_58950_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___118_comb;
  wire [14:0] p1_smul_58954_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___119_comb;
  wire [14:0] p1_smul_58960_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___120_comb;
  wire [14:0] p1_smul_58964_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___121_comb;
  wire [14:0] p1_smul_58966_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___122_comb;
  wire [14:0] p1_smul_58970_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___123_comb;
  wire [14:0] p1_smul_58976_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___124_comb;
  wire [14:0] p1_smul_58980_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___125_comb;
  wire [14:0] p1_smul_58982_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___126_comb;
  wire [14:0] p1_smul_58986_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___127_comb;
  wire [13:0] p1_smul_58990_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___224_comb;
  wire [15:0] p1_smul_58992_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___225_comb;
  wire [15:0] p1_smul_59002_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___226_comb;
  wire [13:0] p1_smul_59004_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___227_comb;
  wire [13:0] p1_smul_59006_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___228_comb;
  wire [15:0] p1_smul_59008_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___229_comb;
  wire [15:0] p1_smul_59018_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___230_comb;
  wire [13:0] p1_smul_59020_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___231_comb;
  wire [13:0] p1_smul_59022_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___232_comb;
  wire [15:0] p1_smul_59024_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___233_comb;
  wire [15:0] p1_smul_59034_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___234_comb;
  wire [13:0] p1_smul_59036_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___235_comb;
  wire [13:0] p1_smul_59038_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___236_comb;
  wire [15:0] p1_smul_59040_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___237_comb;
  wire [15:0] p1_smul_59050_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___238_comb;
  wire [13:0] p1_smul_59052_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___239_comb;
  wire [13:0] p1_smul_59054_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___240_comb;
  wire [15:0] p1_smul_59056_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___241_comb;
  wire [15:0] p1_smul_59066_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___242_comb;
  wire [13:0] p1_smul_59068_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___243_comb;
  wire [13:0] p1_smul_59070_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___244_comb;
  wire [15:0] p1_smul_59072_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___245_comb;
  wire [15:0] p1_smul_59082_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___246_comb;
  wire [13:0] p1_smul_59084_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___247_comb;
  wire [13:0] p1_smul_59086_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___248_comb;
  wire [15:0] p1_smul_59088_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___249_comb;
  wire [15:0] p1_smul_59098_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___250_comb;
  wire [13:0] p1_smul_59100_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___251_comb;
  wire [13:0] p1_smul_59102_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___252_comb;
  wire [15:0] p1_smul_59104_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___253_comb;
  wire [15:0] p1_smul_59114_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___254_comb;
  wire [13:0] p1_smul_59116_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___255_comb;
  wire [7:0] p1_smul_57326_TrailingBits___192_comb;
  wire [7:0] p1_smul_57326_TrailingBits___193_comb;
  wire [7:0] p1_smul_57326_TrailingBits___194_comb;
  wire [7:0] p1_smul_57326_TrailingBits___195_comb;
  wire [7:0] p1_smul_57326_TrailingBits___196_comb;
  wire [7:0] p1_smul_57326_TrailingBits___197_comb;
  wire [7:0] p1_smul_57326_TrailingBits___198_comb;
  wire [7:0] p1_smul_57326_TrailingBits___199_comb;
  wire [7:0] p1_smul_57326_TrailingBits___200_comb;
  wire [7:0] p1_smul_57326_TrailingBits___201_comb;
  wire [7:0] p1_smul_57326_TrailingBits___202_comb;
  wire [7:0] p1_smul_57326_TrailingBits___203_comb;
  wire [7:0] p1_smul_57326_TrailingBits___204_comb;
  wire [7:0] p1_smul_57326_TrailingBits___205_comb;
  wire [7:0] p1_smul_57326_TrailingBits___206_comb;
  wire [7:0] p1_smul_57326_TrailingBits___207_comb;
  wire [7:0] p1_smul_57326_TrailingBits___208_comb;
  wire [7:0] p1_smul_57326_TrailingBits___209_comb;
  wire [7:0] p1_smul_57326_TrailingBits___210_comb;
  wire [7:0] p1_smul_57326_TrailingBits___211_comb;
  wire [7:0] p1_smul_57326_TrailingBits___212_comb;
  wire [7:0] p1_smul_57326_TrailingBits___213_comb;
  wire [7:0] p1_smul_57326_TrailingBits___214_comb;
  wire [7:0] p1_smul_57326_TrailingBits___215_comb;
  wire [7:0] p1_smul_57326_TrailingBits___216_comb;
  wire [7:0] p1_smul_57326_TrailingBits___217_comb;
  wire [7:0] p1_smul_57326_TrailingBits___218_comb;
  wire [7:0] p1_smul_57326_TrailingBits___219_comb;
  wire [7:0] p1_smul_57326_TrailingBits___220_comb;
  wire [7:0] p1_smul_57326_TrailingBits___221_comb;
  wire [7:0] p1_smul_57326_TrailingBits___222_comb;
  wire [7:0] p1_smul_57326_TrailingBits___223_comb;
  wire [7:0] p1_smul_57326_TrailingBits___224_comb;
  wire [7:0] p1_smul_57326_TrailingBits___225_comb;
  wire [7:0] p1_smul_57326_TrailingBits___226_comb;
  wire [7:0] p1_smul_57326_TrailingBits___227_comb;
  wire [7:0] p1_smul_57326_TrailingBits___228_comb;
  wire [7:0] p1_smul_57326_TrailingBits___229_comb;
  wire [7:0] p1_smul_57326_TrailingBits___230_comb;
  wire [7:0] p1_smul_57326_TrailingBits___231_comb;
  wire [7:0] p1_smul_57326_TrailingBits___232_comb;
  wire [7:0] p1_smul_57326_TrailingBits___233_comb;
  wire [7:0] p1_smul_57326_TrailingBits___234_comb;
  wire [7:0] p1_smul_57326_TrailingBits___235_comb;
  wire [7:0] p1_smul_57326_TrailingBits___236_comb;
  wire [7:0] p1_smul_57326_TrailingBits___237_comb;
  wire [7:0] p1_smul_57326_TrailingBits___238_comb;
  wire [7:0] p1_smul_57326_TrailingBits___239_comb;
  wire [7:0] p1_smul_57326_TrailingBits___240_comb;
  wire [7:0] p1_smul_57326_TrailingBits___241_comb;
  wire [7:0] p1_smul_57326_TrailingBits___242_comb;
  wire [7:0] p1_smul_57326_TrailingBits___243_comb;
  wire [7:0] p1_smul_57326_TrailingBits___244_comb;
  wire [7:0] p1_smul_57326_TrailingBits___245_comb;
  wire [7:0] p1_smul_57326_TrailingBits___246_comb;
  wire [7:0] p1_smul_57326_TrailingBits___247_comb;
  wire [7:0] p1_smul_57326_TrailingBits___248_comb;
  wire [7:0] p1_smul_57326_TrailingBits___249_comb;
  wire [7:0] p1_smul_57326_TrailingBits___250_comb;
  wire [7:0] p1_smul_57326_TrailingBits___251_comb;
  wire [7:0] p1_smul_57326_TrailingBits___252_comb;
  wire [7:0] p1_smul_57326_TrailingBits___253_comb;
  wire [7:0] p1_smul_57326_TrailingBits___254_comb;
  wire [7:0] p1_smul_57326_TrailingBits___255_comb;
  wire [24:0] p1_concat_139457_comb;
  wire [22:0] p1_concat_139458_comb;
  wire [22:0] p1_concat_139459_comb;
  wire [24:0] p1_concat_139460_comb;
  wire [24:0] p1_concat_139461_comb;
  wire [22:0] p1_concat_139462_comb;
  wire [22:0] p1_concat_139463_comb;
  wire [24:0] p1_concat_139464_comb;
  wire [24:0] p1_concat_139465_comb;
  wire [22:0] p1_concat_139466_comb;
  wire [22:0] p1_concat_139467_comb;
  wire [24:0] p1_concat_139468_comb;
  wire [24:0] p1_concat_139469_comb;
  wire [22:0] p1_concat_139470_comb;
  wire [22:0] p1_concat_139471_comb;
  wire [24:0] p1_concat_139472_comb;
  wire [24:0] p1_concat_139473_comb;
  wire [22:0] p1_concat_139474_comb;
  wire [22:0] p1_concat_139475_comb;
  wire [24:0] p1_concat_139476_comb;
  wire [24:0] p1_concat_139477_comb;
  wire [22:0] p1_concat_139478_comb;
  wire [22:0] p1_concat_139479_comb;
  wire [24:0] p1_concat_139480_comb;
  wire [24:0] p1_concat_139481_comb;
  wire [22:0] p1_concat_139482_comb;
  wire [22:0] p1_concat_139483_comb;
  wire [24:0] p1_concat_139484_comb;
  wire [24:0] p1_concat_139485_comb;
  wire [22:0] p1_concat_139486_comb;
  wire [22:0] p1_concat_139487_comb;
  wire [24:0] p1_concat_139488_comb;
  wire [24:0] p1_concat_139489_comb;
  wire [24:0] p1_concat_139490_comb;
  wire [24:0] p1_concat_139491_comb;
  wire [24:0] p1_concat_139492_comb;
  wire [24:0] p1_concat_139493_comb;
  wire [24:0] p1_concat_139494_comb;
  wire [24:0] p1_concat_139495_comb;
  wire [24:0] p1_concat_139496_comb;
  wire [24:0] p1_concat_139497_comb;
  wire [24:0] p1_concat_139498_comb;
  wire [24:0] p1_concat_139499_comb;
  wire [24:0] p1_concat_139500_comb;
  wire [24:0] p1_concat_139501_comb;
  wire [24:0] p1_concat_139502_comb;
  wire [24:0] p1_concat_139503_comb;
  wire [24:0] p1_concat_139504_comb;
  wire [24:0] p1_concat_139505_comb;
  wire [24:0] p1_concat_139506_comb;
  wire [24:0] p1_concat_139507_comb;
  wire [24:0] p1_concat_139508_comb;
  wire [24:0] p1_concat_139509_comb;
  wire [24:0] p1_concat_139510_comb;
  wire [24:0] p1_concat_139511_comb;
  wire [24:0] p1_concat_139512_comb;
  wire [24:0] p1_concat_139513_comb;
  wire [24:0] p1_concat_139514_comb;
  wire [24:0] p1_concat_139515_comb;
  wire [24:0] p1_concat_139516_comb;
  wire [24:0] p1_concat_139517_comb;
  wire [24:0] p1_concat_139518_comb;
  wire [24:0] p1_concat_139519_comb;
  wire [24:0] p1_concat_139520_comb;
  wire [22:0] p1_concat_139521_comb;
  wire [24:0] p1_concat_139522_comb;
  wire [24:0] p1_concat_139523_comb;
  wire [22:0] p1_concat_139524_comb;
  wire [22:0] p1_concat_139525_comb;
  wire [24:0] p1_concat_139526_comb;
  wire [24:0] p1_concat_139527_comb;
  wire [22:0] p1_concat_139528_comb;
  wire [22:0] p1_concat_139529_comb;
  wire [24:0] p1_concat_139530_comb;
  wire [24:0] p1_concat_139531_comb;
  wire [22:0] p1_concat_139532_comb;
  wire [22:0] p1_concat_139533_comb;
  wire [24:0] p1_concat_139534_comb;
  wire [24:0] p1_concat_139535_comb;
  wire [22:0] p1_concat_139536_comb;
  wire [22:0] p1_concat_139537_comb;
  wire [24:0] p1_concat_139538_comb;
  wire [24:0] p1_concat_139539_comb;
  wire [22:0] p1_concat_139540_comb;
  wire [22:0] p1_concat_139541_comb;
  wire [24:0] p1_concat_139542_comb;
  wire [24:0] p1_concat_139543_comb;
  wire [22:0] p1_concat_139544_comb;
  wire [22:0] p1_concat_139545_comb;
  wire [24:0] p1_concat_139546_comb;
  wire [24:0] p1_concat_139547_comb;
  wire [22:0] p1_concat_139548_comb;
  wire [22:0] p1_concat_139549_comb;
  wire [24:0] p1_concat_139550_comb;
  wire [24:0] p1_concat_139551_comb;
  wire [22:0] p1_concat_139552_comb;
  wire [24:0] p1_concat_139553_comb;
  wire [22:0] p1_concat_139554_comb;
  wire [22:0] p1_concat_139555_comb;
  wire [24:0] p1_concat_139556_comb;
  wire [24:0] p1_concat_139557_comb;
  wire [22:0] p1_concat_139558_comb;
  wire [22:0] p1_concat_139559_comb;
  wire [24:0] p1_concat_139560_comb;
  wire [24:0] p1_concat_139561_comb;
  wire [22:0] p1_concat_139562_comb;
  wire [22:0] p1_concat_139563_comb;
  wire [24:0] p1_concat_139564_comb;
  wire [24:0] p1_concat_139565_comb;
  wire [22:0] p1_concat_139566_comb;
  wire [22:0] p1_concat_139567_comb;
  wire [24:0] p1_concat_139568_comb;
  wire [24:0] p1_concat_139569_comb;
  wire [22:0] p1_concat_139570_comb;
  wire [22:0] p1_concat_139571_comb;
  wire [24:0] p1_concat_139572_comb;
  wire [24:0] p1_concat_139573_comb;
  wire [22:0] p1_concat_139574_comb;
  wire [22:0] p1_concat_139575_comb;
  wire [24:0] p1_concat_139576_comb;
  wire [24:0] p1_concat_139577_comb;
  wire [22:0] p1_concat_139578_comb;
  wire [22:0] p1_concat_139579_comb;
  wire [24:0] p1_concat_139580_comb;
  wire [24:0] p1_concat_139581_comb;
  wire [22:0] p1_concat_139582_comb;
  wire [22:0] p1_concat_139583_comb;
  wire [24:0] p1_concat_139584_comb;
  wire [24:0] p1_concat_139585_comb;
  wire [24:0] p1_concat_139586_comb;
  wire [24:0] p1_concat_139587_comb;
  wire [24:0] p1_concat_139588_comb;
  wire [24:0] p1_concat_139589_comb;
  wire [24:0] p1_concat_139590_comb;
  wire [24:0] p1_concat_139591_comb;
  wire [24:0] p1_concat_139592_comb;
  wire [24:0] p1_concat_139593_comb;
  wire [24:0] p1_concat_139594_comb;
  wire [24:0] p1_concat_139595_comb;
  wire [24:0] p1_concat_139596_comb;
  wire [24:0] p1_concat_139597_comb;
  wire [24:0] p1_concat_139598_comb;
  wire [24:0] p1_concat_139599_comb;
  wire [24:0] p1_concat_139600_comb;
  wire [24:0] p1_concat_139601_comb;
  wire [24:0] p1_concat_139602_comb;
  wire [24:0] p1_concat_139603_comb;
  wire [24:0] p1_concat_139604_comb;
  wire [24:0] p1_concat_139605_comb;
  wire [24:0] p1_concat_139606_comb;
  wire [24:0] p1_concat_139607_comb;
  wire [24:0] p1_concat_139608_comb;
  wire [24:0] p1_concat_139609_comb;
  wire [24:0] p1_concat_139610_comb;
  wire [24:0] p1_concat_139611_comb;
  wire [24:0] p1_concat_139612_comb;
  wire [24:0] p1_concat_139613_comb;
  wire [24:0] p1_concat_139614_comb;
  wire [24:0] p1_concat_139615_comb;
  wire [24:0] p1_concat_139616_comb;
  wire [22:0] p1_concat_139617_comb;
  wire [24:0] p1_concat_139618_comb;
  wire [24:0] p1_concat_139619_comb;
  wire [22:0] p1_concat_139620_comb;
  wire [22:0] p1_concat_139621_comb;
  wire [24:0] p1_concat_139622_comb;
  wire [24:0] p1_concat_139623_comb;
  wire [22:0] p1_concat_139624_comb;
  wire [22:0] p1_concat_139625_comb;
  wire [24:0] p1_concat_139626_comb;
  wire [24:0] p1_concat_139627_comb;
  wire [22:0] p1_concat_139628_comb;
  wire [22:0] p1_concat_139629_comb;
  wire [24:0] p1_concat_139630_comb;
  wire [24:0] p1_concat_139631_comb;
  wire [22:0] p1_concat_139632_comb;
  wire [22:0] p1_concat_139633_comb;
  wire [24:0] p1_concat_139634_comb;
  wire [24:0] p1_concat_139635_comb;
  wire [22:0] p1_concat_139636_comb;
  wire [22:0] p1_concat_139637_comb;
  wire [24:0] p1_concat_139638_comb;
  wire [24:0] p1_concat_139639_comb;
  wire [22:0] p1_concat_139640_comb;
  wire [22:0] p1_concat_139641_comb;
  wire [24:0] p1_concat_139642_comb;
  wire [24:0] p1_concat_139643_comb;
  wire [22:0] p1_concat_139644_comb;
  wire [22:0] p1_concat_139645_comb;
  wire [24:0] p1_concat_139646_comb;
  wire [24:0] p1_concat_139647_comb;
  wire [22:0] p1_concat_139648_comb;
  wire [15:0] p1_shifted__64_comb;
  wire [7:0] p1_smul_57326_TrailingBits___64_comb;
  wire [15:0] p1_shifted__65_comb;
  wire [7:0] p1_smul_57326_TrailingBits___65_comb;
  wire [15:0] p1_shifted__66_comb;
  wire [7:0] p1_smul_57326_TrailingBits___66_comb;
  wire [15:0] p1_shifted__67_comb;
  wire [7:0] p1_smul_57326_TrailingBits___67_comb;
  wire [15:0] p1_shifted__68_comb;
  wire [7:0] p1_smul_57326_TrailingBits___68_comb;
  wire [15:0] p1_shifted__69_comb;
  wire [7:0] p1_smul_57326_TrailingBits___69_comb;
  wire [15:0] p1_shifted__70_comb;
  wire [7:0] p1_smul_57326_TrailingBits___70_comb;
  wire [15:0] p1_shifted__71_comb;
  wire [7:0] p1_smul_57326_TrailingBits___71_comb;
  wire [15:0] p1_shifted__72_comb;
  wire [7:0] p1_smul_57326_TrailingBits___72_comb;
  wire [15:0] p1_shifted__73_comb;
  wire [7:0] p1_smul_57326_TrailingBits___73_comb;
  wire [15:0] p1_shifted__74_comb;
  wire [7:0] p1_smul_57326_TrailingBits___74_comb;
  wire [15:0] p1_shifted__75_comb;
  wire [7:0] p1_smul_57326_TrailingBits___75_comb;
  wire [15:0] p1_shifted__76_comb;
  wire [7:0] p1_smul_57326_TrailingBits___76_comb;
  wire [15:0] p1_shifted__77_comb;
  wire [7:0] p1_smul_57326_TrailingBits___77_comb;
  wire [15:0] p1_shifted__78_comb;
  wire [7:0] p1_smul_57326_TrailingBits___78_comb;
  wire [15:0] p1_shifted__79_comb;
  wire [7:0] p1_smul_57326_TrailingBits___79_comb;
  wire [15:0] p1_shifted__80_comb;
  wire [7:0] p1_smul_57326_TrailingBits___80_comb;
  wire [15:0] p1_shifted__81_comb;
  wire [7:0] p1_smul_57326_TrailingBits___81_comb;
  wire [15:0] p1_shifted__82_comb;
  wire [7:0] p1_smul_57326_TrailingBits___82_comb;
  wire [15:0] p1_shifted__83_comb;
  wire [7:0] p1_smul_57326_TrailingBits___83_comb;
  wire [15:0] p1_shifted__84_comb;
  wire [7:0] p1_smul_57326_TrailingBits___84_comb;
  wire [15:0] p1_shifted__85_comb;
  wire [7:0] p1_smul_57326_TrailingBits___85_comb;
  wire [15:0] p1_shifted__86_comb;
  wire [7:0] p1_smul_57326_TrailingBits___86_comb;
  wire [15:0] p1_shifted__87_comb;
  wire [7:0] p1_smul_57326_TrailingBits___87_comb;
  wire [15:0] p1_shifted__88_comb;
  wire [7:0] p1_smul_57326_TrailingBits___88_comb;
  wire [15:0] p1_shifted__89_comb;
  wire [7:0] p1_smul_57326_TrailingBits___89_comb;
  wire [15:0] p1_shifted__90_comb;
  wire [7:0] p1_smul_57326_TrailingBits___90_comb;
  wire [15:0] p1_shifted__91_comb;
  wire [7:0] p1_smul_57326_TrailingBits___91_comb;
  wire [15:0] p1_shifted__92_comb;
  wire [7:0] p1_smul_57326_TrailingBits___92_comb;
  wire [15:0] p1_shifted__93_comb;
  wire [7:0] p1_smul_57326_TrailingBits___93_comb;
  wire [15:0] p1_shifted__94_comb;
  wire [7:0] p1_smul_57326_TrailingBits___94_comb;
  wire [15:0] p1_shifted__95_comb;
  wire [7:0] p1_smul_57326_TrailingBits___95_comb;
  wire [15:0] p1_shifted__96_comb;
  wire [7:0] p1_smul_57326_TrailingBits___96_comb;
  wire [15:0] p1_shifted__97_comb;
  wire [7:0] p1_smul_57326_TrailingBits___97_comb;
  wire [15:0] p1_shifted__98_comb;
  wire [7:0] p1_smul_57326_TrailingBits___98_comb;
  wire [15:0] p1_shifted__99_comb;
  wire [7:0] p1_smul_57326_TrailingBits___99_comb;
  wire [15:0] p1_shifted__100_comb;
  wire [7:0] p1_smul_57326_TrailingBits___100_comb;
  wire [15:0] p1_shifted__101_comb;
  wire [7:0] p1_smul_57326_TrailingBits___101_comb;
  wire [15:0] p1_shifted__102_comb;
  wire [7:0] p1_smul_57326_TrailingBits___102_comb;
  wire [15:0] p1_shifted__103_comb;
  wire [7:0] p1_smul_57326_TrailingBits___103_comb;
  wire [15:0] p1_shifted__104_comb;
  wire [7:0] p1_smul_57326_TrailingBits___104_comb;
  wire [15:0] p1_shifted__105_comb;
  wire [7:0] p1_smul_57326_TrailingBits___105_comb;
  wire [15:0] p1_shifted__106_comb;
  wire [7:0] p1_smul_57326_TrailingBits___106_comb;
  wire [15:0] p1_shifted__107_comb;
  wire [7:0] p1_smul_57326_TrailingBits___107_comb;
  wire [15:0] p1_shifted__108_comb;
  wire [7:0] p1_smul_57326_TrailingBits___108_comb;
  wire [15:0] p1_shifted__109_comb;
  wire [7:0] p1_smul_57326_TrailingBits___109_comb;
  wire [15:0] p1_shifted__110_comb;
  wire [7:0] p1_smul_57326_TrailingBits___110_comb;
  wire [15:0] p1_shifted__111_comb;
  wire [7:0] p1_smul_57326_TrailingBits___111_comb;
  wire [15:0] p1_shifted__112_comb;
  wire [7:0] p1_smul_57326_TrailingBits___112_comb;
  wire [15:0] p1_shifted__113_comb;
  wire [7:0] p1_smul_57326_TrailingBits___113_comb;
  wire [15:0] p1_shifted__114_comb;
  wire [7:0] p1_smul_57326_TrailingBits___114_comb;
  wire [15:0] p1_shifted__115_comb;
  wire [7:0] p1_smul_57326_TrailingBits___115_comb;
  wire [15:0] p1_shifted__116_comb;
  wire [7:0] p1_smul_57326_TrailingBits___116_comb;
  wire [15:0] p1_shifted__117_comb;
  wire [7:0] p1_smul_57326_TrailingBits___117_comb;
  wire [15:0] p1_shifted__118_comb;
  wire [7:0] p1_smul_57326_TrailingBits___118_comb;
  wire [15:0] p1_shifted__119_comb;
  wire [7:0] p1_smul_57326_TrailingBits___119_comb;
  wire [15:0] p1_shifted__120_comb;
  wire [7:0] p1_smul_57326_TrailingBits___120_comb;
  wire [15:0] p1_shifted__121_comb;
  wire [7:0] p1_smul_57326_TrailingBits___121_comb;
  wire [15:0] p1_shifted__122_comb;
  wire [7:0] p1_smul_57326_TrailingBits___122_comb;
  wire [15:0] p1_shifted__123_comb;
  wire [7:0] p1_smul_57326_TrailingBits___123_comb;
  wire [15:0] p1_shifted__124_comb;
  wire [7:0] p1_smul_57326_TrailingBits___124_comb;
  wire [15:0] p1_shifted__125_comb;
  wire [7:0] p1_smul_57326_TrailingBits___125_comb;
  wire [15:0] p1_shifted__126_comb;
  wire [7:0] p1_smul_57326_TrailingBits___126_comb;
  wire [15:0] p1_shifted__127_comb;
  wire [7:0] p1_smul_57326_TrailingBits___127_comb;
  wire [31:0] p1_prod__519_comb;
  wire [31:0] p1_prod__523_comb;
  wire [31:0] p1_prod__528_comb;
  wire [31:0] p1_prod__534_comb;
  wire [31:0] p1_prod__583_comb;
  wire [31:0] p1_prod__587_comb;
  wire [31:0] p1_prod__592_comb;
  wire [31:0] p1_prod__598_comb;
  wire [31:0] p1_prod__647_comb;
  wire [31:0] p1_prod__651_comb;
  wire [31:0] p1_prod__656_comb;
  wire [31:0] p1_prod__662_comb;
  wire [31:0] p1_prod__711_comb;
  wire [31:0] p1_prod__715_comb;
  wire [31:0] p1_prod__720_comb;
  wire [31:0] p1_prod__726_comb;
  wire [31:0] p1_prod__775_comb;
  wire [31:0] p1_prod__779_comb;
  wire [31:0] p1_prod__784_comb;
  wire [31:0] p1_prod__790_comb;
  wire [31:0] p1_prod__839_comb;
  wire [31:0] p1_prod__843_comb;
  wire [31:0] p1_prod__848_comb;
  wire [31:0] p1_prod__854_comb;
  wire [31:0] p1_prod__903_comb;
  wire [31:0] p1_prod__907_comb;
  wire [31:0] p1_prod__912_comb;
  wire [31:0] p1_prod__918_comb;
  wire [31:0] p1_prod__967_comb;
  wire [31:0] p1_prod__971_comb;
  wire [31:0] p1_prod__976_comb;
  wire [31:0] p1_prod__982_comb;
  wire [31:0] p1_prod__517_comb;
  wire [31:0] p1_prod__529_comb;
  wire [31:0] p1_prod__535_comb;
  wire [31:0] p1_prod__555_comb;
  wire [31:0] p1_prod__581_comb;
  wire [31:0] p1_prod__593_comb;
  wire [31:0] p1_prod__599_comb;
  wire [31:0] p1_prod__619_comb;
  wire [31:0] p1_prod__645_comb;
  wire [31:0] p1_prod__657_comb;
  wire [31:0] p1_prod__663_comb;
  wire [31:0] p1_prod__683_comb;
  wire [31:0] p1_prod__709_comb;
  wire [31:0] p1_prod__721_comb;
  wire [31:0] p1_prod__727_comb;
  wire [31:0] p1_prod__747_comb;
  wire [31:0] p1_prod__773_comb;
  wire [31:0] p1_prod__785_comb;
  wire [31:0] p1_prod__791_comb;
  wire [31:0] p1_prod__811_comb;
  wire [31:0] p1_prod__837_comb;
  wire [31:0] p1_prod__849_comb;
  wire [31:0] p1_prod__855_comb;
  wire [31:0] p1_prod__875_comb;
  wire [31:0] p1_prod__901_comb;
  wire [31:0] p1_prod__913_comb;
  wire [31:0] p1_prod__919_comb;
  wire [31:0] p1_prod__939_comb;
  wire [31:0] p1_prod__965_comb;
  wire [31:0] p1_prod__977_comb;
  wire [31:0] p1_prod__983_comb;
  wire [31:0] p1_prod__1003_comb;
  wire [31:0] p1_prod__525_comb;
  wire [31:0] p1_prod__536_comb;
  wire [31:0] p1_prod__543_comb;
  wire [31:0] p1_prod__556_comb;
  wire [31:0] p1_prod__589_comb;
  wire [31:0] p1_prod__600_comb;
  wire [31:0] p1_prod__607_comb;
  wire [31:0] p1_prod__620_comb;
  wire [31:0] p1_prod__653_comb;
  wire [31:0] p1_prod__664_comb;
  wire [31:0] p1_prod__671_comb;
  wire [31:0] p1_prod__684_comb;
  wire [31:0] p1_prod__717_comb;
  wire [31:0] p1_prod__728_comb;
  wire [31:0] p1_prod__735_comb;
  wire [31:0] p1_prod__748_comb;
  wire [31:0] p1_prod__781_comb;
  wire [31:0] p1_prod__792_comb;
  wire [31:0] p1_prod__799_comb;
  wire [31:0] p1_prod__812_comb;
  wire [31:0] p1_prod__845_comb;
  wire [31:0] p1_prod__856_comb;
  wire [31:0] p1_prod__863_comb;
  wire [31:0] p1_prod__876_comb;
  wire [31:0] p1_prod__909_comb;
  wire [31:0] p1_prod__920_comb;
  wire [31:0] p1_prod__927_comb;
  wire [31:0] p1_prod__940_comb;
  wire [31:0] p1_prod__973_comb;
  wire [31:0] p1_prod__984_comb;
  wire [31:0] p1_prod__991_comb;
  wire [31:0] p1_prod__1004_comb;
  wire [31:0] p1_prod__532_comb;
  wire [31:0] p1_prod__545_comb;
  wire [31:0] p1_prod__563_comb;
  wire [31:0] p1_prod__570_comb;
  wire [31:0] p1_prod__596_comb;
  wire [31:0] p1_prod__609_comb;
  wire [31:0] p1_prod__627_comb;
  wire [31:0] p1_prod__634_comb;
  wire [31:0] p1_prod__660_comb;
  wire [31:0] p1_prod__673_comb;
  wire [31:0] p1_prod__691_comb;
  wire [31:0] p1_prod__698_comb;
  wire [31:0] p1_prod__724_comb;
  wire [31:0] p1_prod__737_comb;
  wire [31:0] p1_prod__755_comb;
  wire [31:0] p1_prod__762_comb;
  wire [31:0] p1_prod__788_comb;
  wire [31:0] p1_prod__801_comb;
  wire [31:0] p1_prod__819_comb;
  wire [31:0] p1_prod__826_comb;
  wire [31:0] p1_prod__852_comb;
  wire [31:0] p1_prod__865_comb;
  wire [31:0] p1_prod__883_comb;
  wire [31:0] p1_prod__890_comb;
  wire [31:0] p1_prod__916_comb;
  wire [31:0] p1_prod__929_comb;
  wire [31:0] p1_prod__947_comb;
  wire [31:0] p1_prod__954_comb;
  wire [31:0] p1_prod__980_comb;
  wire [31:0] p1_prod__993_comb;
  wire [31:0] p1_prod__1011_comb;
  wire [31:0] p1_prod__1018_comb;
  wire [31:0] p1_prod__546_comb;
  wire [31:0] p1_prod__559_comb;
  wire [31:0] p1_prod__564_comb;
  wire [31:0] p1_prod__571_comb;
  wire [31:0] p1_prod__610_comb;
  wire [31:0] p1_prod__623_comb;
  wire [31:0] p1_prod__628_comb;
  wire [31:0] p1_prod__635_comb;
  wire [31:0] p1_prod__674_comb;
  wire [31:0] p1_prod__687_comb;
  wire [31:0] p1_prod__692_comb;
  wire [31:0] p1_prod__699_comb;
  wire [31:0] p1_prod__738_comb;
  wire [31:0] p1_prod__751_comb;
  wire [31:0] p1_prod__756_comb;
  wire [31:0] p1_prod__763_comb;
  wire [31:0] p1_prod__802_comb;
  wire [31:0] p1_prod__815_comb;
  wire [31:0] p1_prod__820_comb;
  wire [31:0] p1_prod__827_comb;
  wire [31:0] p1_prod__866_comb;
  wire [31:0] p1_prod__879_comb;
  wire [31:0] p1_prod__884_comb;
  wire [31:0] p1_prod__891_comb;
  wire [31:0] p1_prod__930_comb;
  wire [31:0] p1_prod__943_comb;
  wire [31:0] p1_prod__948_comb;
  wire [31:0] p1_prod__955_comb;
  wire [31:0] p1_prod__994_comb;
  wire [31:0] p1_prod__1007_comb;
  wire [31:0] p1_prod__1012_comb;
  wire [31:0] p1_prod__1019_comb;
  wire [31:0] p1_prod__547_comb;
  wire [31:0] p1_prod__554_comb;
  wire [31:0] p1_prod__574_comb;
  wire [31:0] p1_prod__575_comb;
  wire [31:0] p1_prod__611_comb;
  wire [31:0] p1_prod__618_comb;
  wire [31:0] p1_prod__638_comb;
  wire [31:0] p1_prod__639_comb;
  wire [31:0] p1_prod__675_comb;
  wire [31:0] p1_prod__682_comb;
  wire [31:0] p1_prod__702_comb;
  wire [31:0] p1_prod__703_comb;
  wire [31:0] p1_prod__739_comb;
  wire [31:0] p1_prod__746_comb;
  wire [31:0] p1_prod__766_comb;
  wire [31:0] p1_prod__767_comb;
  wire [31:0] p1_prod__803_comb;
  wire [31:0] p1_prod__810_comb;
  wire [31:0] p1_prod__830_comb;
  wire [31:0] p1_prod__831_comb;
  wire [31:0] p1_prod__867_comb;
  wire [31:0] p1_prod__874_comb;
  wire [31:0] p1_prod__894_comb;
  wire [31:0] p1_prod__895_comb;
  wire [31:0] p1_prod__931_comb;
  wire [31:0] p1_prod__938_comb;
  wire [31:0] p1_prod__958_comb;
  wire [31:0] p1_prod__959_comb;
  wire [31:0] p1_prod__995_comb;
  wire [31:0] p1_prod__1002_comb;
  wire [31:0] p1_prod__1022_comb;
  wire [31:0] p1_prod__1023_comb;
  wire [31:0] p1_or_140545_comb;
  wire [31:0] p1_or_140546_comb;
  wire [31:0] p1_or_140547_comb;
  wire [31:0] p1_or_140548_comb;
  wire [31:0] p1_or_140549_comb;
  wire [31:0] p1_or_140550_comb;
  wire [31:0] p1_or_140551_comb;
  wire [31:0] p1_or_140552_comb;
  wire [31:0] p1_or_140553_comb;
  wire [31:0] p1_or_140554_comb;
  wire [31:0] p1_or_140555_comb;
  wire [31:0] p1_or_140556_comb;
  wire [31:0] p1_or_140557_comb;
  wire [31:0] p1_or_140558_comb;
  wire [31:0] p1_or_140559_comb;
  wire [31:0] p1_or_140560_comb;
  wire [31:0] p1_or_140561_comb;
  wire [31:0] p1_or_140562_comb;
  wire [31:0] p1_or_140563_comb;
  wire [31:0] p1_or_140564_comb;
  wire [31:0] p1_or_140565_comb;
  wire [31:0] p1_or_140566_comb;
  wire [31:0] p1_or_140567_comb;
  wire [31:0] p1_or_140568_comb;
  wire [31:0] p1_or_140569_comb;
  wire [31:0] p1_or_140570_comb;
  wire [31:0] p1_or_140571_comb;
  wire [31:0] p1_or_140572_comb;
  wire [31:0] p1_or_140573_comb;
  wire [31:0] p1_or_140574_comb;
  wire [31:0] p1_or_140575_comb;
  wire [31:0] p1_or_140576_comb;
  wire [31:0] p1_or_140577_comb;
  wire [14:0] p1_smul_58352_NarrowedMult__comb;
  wire [14:0] p1_smul_58354_NarrowedMult__comb;
  wire [31:0] p1_or_140582_comb;
  wire [31:0] p1_or_140583_comb;
  wire [14:0] p1_smul_58360_NarrowedMult__comb;
  wire [14:0] p1_smul_58362_NarrowedMult__comb;
  wire [31:0] p1_or_140588_comb;
  wire [31:0] p1_or_140589_comb;
  wire [14:0] p1_smul_58368_NarrowedMult__comb;
  wire [14:0] p1_smul_58370_NarrowedMult__comb;
  wire [31:0] p1_or_140594_comb;
  wire [31:0] p1_or_140595_comb;
  wire [14:0] p1_smul_58376_NarrowedMult__comb;
  wire [14:0] p1_smul_58378_NarrowedMult__comb;
  wire [31:0] p1_or_140600_comb;
  wire [31:0] p1_or_140601_comb;
  wire [14:0] p1_smul_58384_NarrowedMult__comb;
  wire [14:0] p1_smul_58386_NarrowedMult__comb;
  wire [31:0] p1_or_140606_comb;
  wire [31:0] p1_or_140607_comb;
  wire [14:0] p1_smul_58392_NarrowedMult__comb;
  wire [14:0] p1_smul_58394_NarrowedMult__comb;
  wire [31:0] p1_or_140612_comb;
  wire [31:0] p1_or_140613_comb;
  wire [14:0] p1_smul_58400_NarrowedMult__comb;
  wire [14:0] p1_smul_58402_NarrowedMult__comb;
  wire [31:0] p1_or_140618_comb;
  wire [31:0] p1_or_140619_comb;
  wire [14:0] p1_smul_58408_NarrowedMult__comb;
  wire [14:0] p1_smul_58410_NarrowedMult__comb;
  wire [31:0] p1_or_140624_comb;
  wire [31:0] p1_or_140625_comb;
  wire [14:0] p1_smul_58416_NarrowedMult__comb;
  wire [14:0] p1_smul_58418_NarrowedMult__comb;
  wire [31:0] p1_or_140630_comb;
  wire [31:0] p1_or_140631_comb;
  wire [14:0] p1_smul_58424_NarrowedMult__comb;
  wire [14:0] p1_smul_58426_NarrowedMult__comb;
  wire [31:0] p1_or_140636_comb;
  wire [31:0] p1_or_140637_comb;
  wire [14:0] p1_smul_58432_NarrowedMult__comb;
  wire [14:0] p1_smul_58434_NarrowedMult__comb;
  wire [31:0] p1_or_140642_comb;
  wire [31:0] p1_or_140643_comb;
  wire [14:0] p1_smul_58440_NarrowedMult__comb;
  wire [14:0] p1_smul_58442_NarrowedMult__comb;
  wire [31:0] p1_or_140648_comb;
  wire [31:0] p1_or_140649_comb;
  wire [14:0] p1_smul_58448_NarrowedMult__comb;
  wire [14:0] p1_smul_58450_NarrowedMult__comb;
  wire [31:0] p1_or_140654_comb;
  wire [31:0] p1_or_140655_comb;
  wire [14:0] p1_smul_58456_NarrowedMult__comb;
  wire [14:0] p1_smul_58458_NarrowedMult__comb;
  wire [31:0] p1_or_140660_comb;
  wire [31:0] p1_or_140661_comb;
  wire [14:0] p1_smul_58464_NarrowedMult__comb;
  wire [14:0] p1_smul_58466_NarrowedMult__comb;
  wire [31:0] p1_or_140666_comb;
  wire [31:0] p1_or_140667_comb;
  wire [14:0] p1_smul_58472_NarrowedMult__comb;
  wire [14:0] p1_smul_58474_NarrowedMult__comb;
  wire [31:0] p1_or_140672_comb;
  wire [31:0] p1_or_140673_comb;
  wire [31:0] p1_or_140674_comb;
  wire [31:0] p1_or_140675_comb;
  wire [31:0] p1_or_140676_comb;
  wire [31:0] p1_or_140677_comb;
  wire [31:0] p1_or_140678_comb;
  wire [31:0] p1_or_140679_comb;
  wire [31:0] p1_or_140680_comb;
  wire [31:0] p1_or_140681_comb;
  wire [31:0] p1_or_140682_comb;
  wire [31:0] p1_or_140683_comb;
  wire [31:0] p1_or_140684_comb;
  wire [31:0] p1_or_140685_comb;
  wire [31:0] p1_or_140686_comb;
  wire [31:0] p1_or_140687_comb;
  wire [31:0] p1_or_140688_comb;
  wire [31:0] p1_or_140689_comb;
  wire [31:0] p1_or_140690_comb;
  wire [31:0] p1_or_140691_comb;
  wire [31:0] p1_or_140692_comb;
  wire [31:0] p1_or_140693_comb;
  wire [31:0] p1_or_140694_comb;
  wire [31:0] p1_or_140695_comb;
  wire [31:0] p1_or_140696_comb;
  wire [31:0] p1_or_140697_comb;
  wire [31:0] p1_or_140698_comb;
  wire [31:0] p1_or_140699_comb;
  wire [31:0] p1_or_140700_comb;
  wire [31:0] p1_or_140701_comb;
  wire [31:0] p1_or_140702_comb;
  wire [31:0] p1_or_140703_comb;
  wire [31:0] p1_or_140704_comb;
  wire [31:0] p1_or_140705_comb;
  wire [31:0] p1_or_140706_comb;
  wire [31:0] p1_or_140707_comb;
  wire [31:0] p1_or_140708_comb;
  wire [31:0] p1_or_140709_comb;
  wire [31:0] p1_or_140710_comb;
  wire [31:0] p1_or_140711_comb;
  wire [31:0] p1_or_140712_comb;
  wire [31:0] p1_or_140713_comb;
  wire [31:0] p1_or_140714_comb;
  wire [31:0] p1_or_140715_comb;
  wire [31:0] p1_or_140716_comb;
  wire [31:0] p1_or_140717_comb;
  wire [31:0] p1_or_140718_comb;
  wire [31:0] p1_or_140719_comb;
  wire [31:0] p1_or_140720_comb;
  wire [31:0] p1_or_140721_comb;
  wire [31:0] p1_or_140722_comb;
  wire [31:0] p1_or_140723_comb;
  wire [31:0] p1_or_140724_comb;
  wire [31:0] p1_or_140725_comb;
  wire [31:0] p1_or_140726_comb;
  wire [31:0] p1_or_140727_comb;
  wire [31:0] p1_or_140728_comb;
  wire [31:0] p1_or_140729_comb;
  wire [31:0] p1_or_140730_comb;
  wire [31:0] p1_or_140731_comb;
  wire [31:0] p1_or_140732_comb;
  wire [31:0] p1_or_140733_comb;
  wire [31:0] p1_or_140734_comb;
  wire [31:0] p1_or_140735_comb;
  wire [31:0] p1_or_140736_comb;
  wire [14:0] p1_smul_58862_NarrowedMult__comb;
  wire [31:0] p1_or_140739_comb;
  wire [14:0] p1_smul_58866_NarrowedMult__comb;
  wire [31:0] p1_or_140742_comb;
  wire [31:0] p1_or_140743_comb;
  wire [14:0] p1_smul_58872_NarrowedMult__comb;
  wire [31:0] p1_or_140746_comb;
  wire [14:0] p1_smul_58876_NarrowedMult__comb;
  wire [14:0] p1_smul_58878_NarrowedMult__comb;
  wire [31:0] p1_or_140751_comb;
  wire [14:0] p1_smul_58882_NarrowedMult__comb;
  wire [31:0] p1_or_140754_comb;
  wire [31:0] p1_or_140755_comb;
  wire [14:0] p1_smul_58888_NarrowedMult__comb;
  wire [31:0] p1_or_140758_comb;
  wire [14:0] p1_smul_58892_NarrowedMult__comb;
  wire [14:0] p1_smul_58894_NarrowedMult__comb;
  wire [31:0] p1_or_140763_comb;
  wire [14:0] p1_smul_58898_NarrowedMult__comb;
  wire [31:0] p1_or_140766_comb;
  wire [31:0] p1_or_140767_comb;
  wire [14:0] p1_smul_58904_NarrowedMult__comb;
  wire [31:0] p1_or_140770_comb;
  wire [14:0] p1_smul_58908_NarrowedMult__comb;
  wire [14:0] p1_smul_58910_NarrowedMult__comb;
  wire [31:0] p1_or_140775_comb;
  wire [14:0] p1_smul_58914_NarrowedMult__comb;
  wire [31:0] p1_or_140778_comb;
  wire [31:0] p1_or_140779_comb;
  wire [14:0] p1_smul_58920_NarrowedMult__comb;
  wire [31:0] p1_or_140782_comb;
  wire [14:0] p1_smul_58924_NarrowedMult__comb;
  wire [14:0] p1_smul_58926_NarrowedMult__comb;
  wire [31:0] p1_or_140787_comb;
  wire [14:0] p1_smul_58930_NarrowedMult__comb;
  wire [31:0] p1_or_140790_comb;
  wire [31:0] p1_or_140791_comb;
  wire [14:0] p1_smul_58936_NarrowedMult__comb;
  wire [31:0] p1_or_140794_comb;
  wire [14:0] p1_smul_58940_NarrowedMult__comb;
  wire [14:0] p1_smul_58942_NarrowedMult__comb;
  wire [31:0] p1_or_140799_comb;
  wire [14:0] p1_smul_58946_NarrowedMult__comb;
  wire [31:0] p1_or_140802_comb;
  wire [31:0] p1_or_140803_comb;
  wire [14:0] p1_smul_58952_NarrowedMult__comb;
  wire [31:0] p1_or_140806_comb;
  wire [14:0] p1_smul_58956_NarrowedMult__comb;
  wire [14:0] p1_smul_58958_NarrowedMult__comb;
  wire [31:0] p1_or_140811_comb;
  wire [14:0] p1_smul_58962_NarrowedMult__comb;
  wire [31:0] p1_or_140814_comb;
  wire [31:0] p1_or_140815_comb;
  wire [14:0] p1_smul_58968_NarrowedMult__comb;
  wire [31:0] p1_or_140818_comb;
  wire [14:0] p1_smul_58972_NarrowedMult__comb;
  wire [14:0] p1_smul_58974_NarrowedMult__comb;
  wire [31:0] p1_or_140823_comb;
  wire [14:0] p1_smul_58978_NarrowedMult__comb;
  wire [31:0] p1_or_140826_comb;
  wire [31:0] p1_or_140827_comb;
  wire [14:0] p1_smul_58984_NarrowedMult__comb;
  wire [31:0] p1_or_140830_comb;
  wire [14:0] p1_smul_58988_NarrowedMult__comb;
  wire [31:0] p1_or_140833_comb;
  wire [31:0] p1_or_140834_comb;
  wire [31:0] p1_or_140835_comb;
  wire [31:0] p1_or_140836_comb;
  wire [31:0] p1_or_140837_comb;
  wire [31:0] p1_or_140838_comb;
  wire [31:0] p1_or_140839_comb;
  wire [31:0] p1_or_140840_comb;
  wire [31:0] p1_or_140841_comb;
  wire [31:0] p1_or_140842_comb;
  wire [31:0] p1_or_140843_comb;
  wire [31:0] p1_or_140844_comb;
  wire [31:0] p1_or_140845_comb;
  wire [31:0] p1_or_140846_comb;
  wire [31:0] p1_or_140847_comb;
  wire [31:0] p1_or_140848_comb;
  wire [31:0] p1_or_140849_comb;
  wire [31:0] p1_or_140850_comb;
  wire [31:0] p1_or_140851_comb;
  wire [31:0] p1_or_140852_comb;
  wire [31:0] p1_or_140853_comb;
  wire [31:0] p1_or_140854_comb;
  wire [31:0] p1_or_140855_comb;
  wire [31:0] p1_or_140856_comb;
  wire [31:0] p1_or_140857_comb;
  wire [31:0] p1_or_140858_comb;
  wire [31:0] p1_or_140859_comb;
  wire [31:0] p1_or_140860_comb;
  wire [31:0] p1_or_140861_comb;
  wire [31:0] p1_or_140862_comb;
  wire [31:0] p1_or_140863_comb;
  wire [31:0] p1_or_140864_comb;
  wire [15:0] p1_sel_140865_comb;
  wire [15:0] p1_sel_140866_comb;
  wire [15:0] p1_sel_140867_comb;
  wire [15:0] p1_sel_140868_comb;
  wire [15:0] p1_sel_140869_comb;
  wire [15:0] p1_sel_140870_comb;
  wire [15:0] p1_sel_140871_comb;
  wire [15:0] p1_sel_140872_comb;
  wire [15:0] p1_sel_140873_comb;
  wire [15:0] p1_sel_140874_comb;
  wire [15:0] p1_sel_140875_comb;
  wire [15:0] p1_sel_140876_comb;
  wire [15:0] p1_sel_140877_comb;
  wire [15:0] p1_sel_140878_comb;
  wire [15:0] p1_sel_140879_comb;
  wire [15:0] p1_sel_140880_comb;
  wire [15:0] p1_sel_140881_comb;
  wire [15:0] p1_sel_140882_comb;
  wire [15:0] p1_sel_140883_comb;
  wire [15:0] p1_sel_140884_comb;
  wire [15:0] p1_sel_140885_comb;
  wire [15:0] p1_sel_140886_comb;
  wire [15:0] p1_sel_140887_comb;
  wire [15:0] p1_sel_140888_comb;
  wire [15:0] p1_sel_140889_comb;
  wire [15:0] p1_sel_140890_comb;
  wire [15:0] p1_sel_140891_comb;
  wire [15:0] p1_sel_140892_comb;
  wire [15:0] p1_sel_140893_comb;
  wire [15:0] p1_sel_140894_comb;
  wire [15:0] p1_sel_140895_comb;
  wire [15:0] p1_sel_140896_comb;
  wire [15:0] p1_sel_140897_comb;
  wire [15:0] p1_sel_140898_comb;
  wire [15:0] p1_sel_140899_comb;
  wire [15:0] p1_sel_140900_comb;
  wire [15:0] p1_sel_140901_comb;
  wire [15:0] p1_sel_140902_comb;
  wire [15:0] p1_sel_140903_comb;
  wire [15:0] p1_sel_140904_comb;
  wire [15:0] p1_sel_140905_comb;
  wire [15:0] p1_sel_140906_comb;
  wire [15:0] p1_sel_140907_comb;
  wire [15:0] p1_sel_140908_comb;
  wire [15:0] p1_sel_140909_comb;
  wire [15:0] p1_sel_140910_comb;
  wire [15:0] p1_sel_140911_comb;
  wire [15:0] p1_sel_140912_comb;
  wire [15:0] p1_sel_140913_comb;
  wire [15:0] p1_sel_140914_comb;
  wire [15:0] p1_sel_140915_comb;
  wire [15:0] p1_sel_140916_comb;
  wire [15:0] p1_sel_140917_comb;
  wire [15:0] p1_sel_140918_comb;
  wire [15:0] p1_sel_140919_comb;
  wire [15:0] p1_sel_140920_comb;
  wire [15:0] p1_sel_140921_comb;
  wire [15:0] p1_sel_140922_comb;
  wire [15:0] p1_sel_140923_comb;
  wire [15:0] p1_sel_140924_comb;
  wire [15:0] p1_sel_140925_comb;
  wire [15:0] p1_sel_140926_comb;
  wire [15:0] p1_sel_140927_comb;
  wire [15:0] p1_sel_140928_comb;
  wire [15:0] p1_concat_141061_comb;
  wire [15:0] p1_concat_141063_comb;
  wire [15:0] p1_concat_141073_comb;
  wire [15:0] p1_concat_141075_comb;
  wire [15:0] p1_concat_141085_comb;
  wire [15:0] p1_concat_141087_comb;
  wire [15:0] p1_concat_141097_comb;
  wire [15:0] p1_concat_141099_comb;
  wire [15:0] p1_concat_141109_comb;
  wire [15:0] p1_concat_141111_comb;
  wire [15:0] p1_concat_141121_comb;
  wire [15:0] p1_concat_141123_comb;
  wire [15:0] p1_concat_141133_comb;
  wire [15:0] p1_concat_141135_comb;
  wire [15:0] p1_concat_141145_comb;
  wire [15:0] p1_concat_141147_comb;
  wire [15:0] p1_concat_141157_comb;
  wire [15:0] p1_concat_141159_comb;
  wire [15:0] p1_concat_141169_comb;
  wire [15:0] p1_concat_141171_comb;
  wire [15:0] p1_concat_141181_comb;
  wire [15:0] p1_concat_141183_comb;
  wire [15:0] p1_concat_141193_comb;
  wire [15:0] p1_concat_141195_comb;
  wire [15:0] p1_concat_141205_comb;
  wire [15:0] p1_concat_141207_comb;
  wire [15:0] p1_concat_141217_comb;
  wire [15:0] p1_concat_141219_comb;
  wire [15:0] p1_concat_141229_comb;
  wire [15:0] p1_concat_141231_comb;
  wire [15:0] p1_concat_141241_comb;
  wire [15:0] p1_concat_141243_comb;
  wire [15:0] p1_concat_141505_comb;
  wire [15:0] p1_concat_141511_comb;
  wire [15:0] p1_concat_141521_comb;
  wire [15:0] p1_concat_141527_comb;
  wire [15:0] p1_concat_141529_comb;
  wire [15:0] p1_concat_141535_comb;
  wire [15:0] p1_concat_141545_comb;
  wire [15:0] p1_concat_141551_comb;
  wire [15:0] p1_concat_141553_comb;
  wire [15:0] p1_concat_141559_comb;
  wire [15:0] p1_concat_141569_comb;
  wire [15:0] p1_concat_141575_comb;
  wire [15:0] p1_concat_141577_comb;
  wire [15:0] p1_concat_141583_comb;
  wire [15:0] p1_concat_141593_comb;
  wire [15:0] p1_concat_141599_comb;
  wire [15:0] p1_concat_141601_comb;
  wire [15:0] p1_concat_141607_comb;
  wire [15:0] p1_concat_141617_comb;
  wire [15:0] p1_concat_141623_comb;
  wire [15:0] p1_concat_141625_comb;
  wire [15:0] p1_concat_141631_comb;
  wire [15:0] p1_concat_141641_comb;
  wire [15:0] p1_concat_141647_comb;
  wire [15:0] p1_concat_141649_comb;
  wire [15:0] p1_concat_141655_comb;
  wire [15:0] p1_concat_141665_comb;
  wire [15:0] p1_concat_141671_comb;
  wire [15:0] p1_concat_141673_comb;
  wire [15:0] p1_concat_141679_comb;
  wire [15:0] p1_concat_141689_comb;
  wire [15:0] p1_concat_141695_comb;
  wire [16:0] p1_add_142785_comb;
  wire [16:0] p1_add_142786_comb;
  wire [16:0] p1_add_142787_comb;
  wire [16:0] p1_add_142788_comb;
  wire [16:0] p1_add_142789_comb;
  wire [16:0] p1_add_142790_comb;
  wire [16:0] p1_add_142791_comb;
  wire [16:0] p1_add_142792_comb;
  wire [16:0] p1_add_142793_comb;
  wire [16:0] p1_add_142794_comb;
  wire [16:0] p1_add_142795_comb;
  wire [16:0] p1_add_142796_comb;
  wire [16:0] p1_add_142797_comb;
  wire [16:0] p1_add_142798_comb;
  wire [16:0] p1_add_142799_comb;
  wire [16:0] p1_add_142800_comb;
  wire [16:0] p1_add_142801_comb;
  wire [16:0] p1_add_142802_comb;
  wire [16:0] p1_add_142803_comb;
  wire [16:0] p1_add_142804_comb;
  wire [16:0] p1_add_142805_comb;
  wire [16:0] p1_add_142806_comb;
  wire [16:0] p1_add_142807_comb;
  wire [16:0] p1_add_142808_comb;
  wire [16:0] p1_add_142809_comb;
  wire [16:0] p1_add_142810_comb;
  wire [16:0] p1_add_142811_comb;
  wire [16:0] p1_add_142812_comb;
  wire [16:0] p1_add_142813_comb;
  wire [16:0] p1_add_142814_comb;
  wire [16:0] p1_add_142815_comb;
  wire [16:0] p1_add_142816_comb;
  wire [15:0] p1_smul_142817_comb;
  wire [15:0] p1_smul_142818_comb;
  wire [15:0] p1_sel_142819_comb;
  wire [15:0] p1_sel_142820_comb;
  wire [15:0] p1_sel_142821_comb;
  wire [15:0] p1_sel_142822_comb;
  wire [15:0] p1_smul_142823_comb;
  wire [15:0] p1_smul_142824_comb;
  wire [15:0] p1_smul_142825_comb;
  wire [15:0] p1_smul_142826_comb;
  wire [15:0] p1_sel_142827_comb;
  wire [15:0] p1_sel_142828_comb;
  wire [15:0] p1_sel_142829_comb;
  wire [15:0] p1_sel_142830_comb;
  wire [15:0] p1_smul_142831_comb;
  wire [15:0] p1_smul_142832_comb;
  wire [15:0] p1_smul_142833_comb;
  wire [15:0] p1_smul_142834_comb;
  wire [15:0] p1_sel_142835_comb;
  wire [15:0] p1_sel_142836_comb;
  wire [15:0] p1_sel_142837_comb;
  wire [15:0] p1_sel_142838_comb;
  wire [15:0] p1_smul_142839_comb;
  wire [15:0] p1_smul_142840_comb;
  wire [15:0] p1_smul_142841_comb;
  wire [15:0] p1_smul_142842_comb;
  wire [15:0] p1_sel_142843_comb;
  wire [15:0] p1_sel_142844_comb;
  wire [15:0] p1_sel_142845_comb;
  wire [15:0] p1_sel_142846_comb;
  wire [15:0] p1_smul_142847_comb;
  wire [15:0] p1_smul_142848_comb;
  wire [15:0] p1_smul_142849_comb;
  wire [15:0] p1_smul_142850_comb;
  wire [15:0] p1_sel_142851_comb;
  wire [15:0] p1_sel_142852_comb;
  wire [15:0] p1_sel_142853_comb;
  wire [15:0] p1_sel_142854_comb;
  wire [15:0] p1_smul_142855_comb;
  wire [15:0] p1_smul_142856_comb;
  wire [15:0] p1_smul_142857_comb;
  wire [15:0] p1_smul_142858_comb;
  wire [15:0] p1_sel_142859_comb;
  wire [15:0] p1_sel_142860_comb;
  wire [15:0] p1_sel_142861_comb;
  wire [15:0] p1_sel_142862_comb;
  wire [15:0] p1_smul_142863_comb;
  wire [15:0] p1_smul_142864_comb;
  wire [15:0] p1_smul_142865_comb;
  wire [15:0] p1_smul_142866_comb;
  wire [15:0] p1_sel_142867_comb;
  wire [15:0] p1_sel_142868_comb;
  wire [15:0] p1_sel_142869_comb;
  wire [15:0] p1_sel_142870_comb;
  wire [15:0] p1_smul_142871_comb;
  wire [15:0] p1_smul_142872_comb;
  wire [15:0] p1_smul_142873_comb;
  wire [15:0] p1_smul_142874_comb;
  wire [15:0] p1_sel_142875_comb;
  wire [15:0] p1_sel_142876_comb;
  wire [15:0] p1_sel_142877_comb;
  wire [15:0] p1_sel_142878_comb;
  wire [15:0] p1_smul_142879_comb;
  wire [15:0] p1_smul_142880_comb;
  wire [15:0] p1_sel_142881_comb;
  wire [15:0] p1_sel_142882_comb;
  wire [15:0] p1_sel_142883_comb;
  wire [15:0] p1_sel_142884_comb;
  wire [15:0] p1_sel_142885_comb;
  wire [15:0] p1_sel_142886_comb;
  wire [15:0] p1_sel_142887_comb;
  wire [15:0] p1_sel_142888_comb;
  wire [15:0] p1_sel_142889_comb;
  wire [15:0] p1_sel_142890_comb;
  wire [15:0] p1_sel_142891_comb;
  wire [15:0] p1_sel_142892_comb;
  wire [15:0] p1_sel_142893_comb;
  wire [15:0] p1_sel_142894_comb;
  wire [15:0] p1_sel_142895_comb;
  wire [15:0] p1_sel_142896_comb;
  wire [15:0] p1_sel_142897_comb;
  wire [15:0] p1_sel_142898_comb;
  wire [15:0] p1_sel_142899_comb;
  wire [15:0] p1_sel_142900_comb;
  wire [15:0] p1_sel_142901_comb;
  wire [15:0] p1_sel_142902_comb;
  wire [15:0] p1_sel_142903_comb;
  wire [15:0] p1_sel_142904_comb;
  wire [15:0] p1_sel_142905_comb;
  wire [15:0] p1_sel_142906_comb;
  wire [15:0] p1_sel_142907_comb;
  wire [15:0] p1_sel_142908_comb;
  wire [15:0] p1_sel_142909_comb;
  wire [15:0] p1_sel_142910_comb;
  wire [15:0] p1_sel_142911_comb;
  wire [15:0] p1_sel_142912_comb;
  wire [15:0] p1_sel_142913_comb;
  wire [15:0] p1_sel_142914_comb;
  wire [15:0] p1_sel_142915_comb;
  wire [15:0] p1_sel_142916_comb;
  wire [15:0] p1_sel_142917_comb;
  wire [15:0] p1_sel_142918_comb;
  wire [15:0] p1_sel_142919_comb;
  wire [15:0] p1_sel_142920_comb;
  wire [15:0] p1_sel_142921_comb;
  wire [15:0] p1_sel_142922_comb;
  wire [15:0] p1_sel_142923_comb;
  wire [15:0] p1_sel_142924_comb;
  wire [15:0] p1_sel_142925_comb;
  wire [15:0] p1_sel_142926_comb;
  wire [15:0] p1_sel_142927_comb;
  wire [15:0] p1_sel_142928_comb;
  wire [15:0] p1_sel_142929_comb;
  wire [15:0] p1_sel_142930_comb;
  wire [15:0] p1_sel_142931_comb;
  wire [15:0] p1_sel_142932_comb;
  wire [15:0] p1_sel_142933_comb;
  wire [15:0] p1_sel_142934_comb;
  wire [15:0] p1_sel_142935_comb;
  wire [15:0] p1_sel_142936_comb;
  wire [15:0] p1_sel_142937_comb;
  wire [15:0] p1_sel_142938_comb;
  wire [15:0] p1_sel_142939_comb;
  wire [15:0] p1_sel_142940_comb;
  wire [15:0] p1_sel_142941_comb;
  wire [15:0] p1_sel_142942_comb;
  wire [15:0] p1_sel_142943_comb;
  wire [15:0] p1_sel_142944_comb;
  wire [15:0] p1_smul_142945_comb;
  wire [15:0] p1_sel_142946_comb;
  wire [15:0] p1_smul_142947_comb;
  wire [15:0] p1_sel_142948_comb;
  wire [15:0] p1_sel_142949_comb;
  wire [15:0] p1_smul_142950_comb;
  wire [15:0] p1_sel_142951_comb;
  wire [15:0] p1_smul_142952_comb;
  wire [15:0] p1_smul_142953_comb;
  wire [15:0] p1_sel_142954_comb;
  wire [15:0] p1_smul_142955_comb;
  wire [15:0] p1_sel_142956_comb;
  wire [15:0] p1_sel_142957_comb;
  wire [15:0] p1_smul_142958_comb;
  wire [15:0] p1_sel_142959_comb;
  wire [15:0] p1_smul_142960_comb;
  wire [15:0] p1_smul_142961_comb;
  wire [15:0] p1_sel_142962_comb;
  wire [15:0] p1_smul_142963_comb;
  wire [15:0] p1_sel_142964_comb;
  wire [15:0] p1_sel_142965_comb;
  wire [15:0] p1_smul_142966_comb;
  wire [15:0] p1_sel_142967_comb;
  wire [15:0] p1_smul_142968_comb;
  wire [15:0] p1_smul_142969_comb;
  wire [15:0] p1_sel_142970_comb;
  wire [15:0] p1_smul_142971_comb;
  wire [15:0] p1_sel_142972_comb;
  wire [15:0] p1_sel_142973_comb;
  wire [15:0] p1_smul_142974_comb;
  wire [15:0] p1_sel_142975_comb;
  wire [15:0] p1_smul_142976_comb;
  wire [15:0] p1_smul_142977_comb;
  wire [15:0] p1_sel_142978_comb;
  wire [15:0] p1_smul_142979_comb;
  wire [15:0] p1_sel_142980_comb;
  wire [15:0] p1_sel_142981_comb;
  wire [15:0] p1_smul_142982_comb;
  wire [15:0] p1_sel_142983_comb;
  wire [15:0] p1_smul_142984_comb;
  wire [15:0] p1_smul_142985_comb;
  wire [15:0] p1_sel_142986_comb;
  wire [15:0] p1_smul_142987_comb;
  wire [15:0] p1_sel_142988_comb;
  wire [15:0] p1_sel_142989_comb;
  wire [15:0] p1_smul_142990_comb;
  wire [15:0] p1_sel_142991_comb;
  wire [15:0] p1_smul_142992_comb;
  wire [15:0] p1_smul_142993_comb;
  wire [15:0] p1_sel_142994_comb;
  wire [15:0] p1_smul_142995_comb;
  wire [15:0] p1_sel_142996_comb;
  wire [15:0] p1_sel_142997_comb;
  wire [15:0] p1_smul_142998_comb;
  wire [15:0] p1_sel_142999_comb;
  wire [15:0] p1_smul_143000_comb;
  wire [15:0] p1_smul_143001_comb;
  wire [15:0] p1_sel_143002_comb;
  wire [15:0] p1_smul_143003_comb;
  wire [15:0] p1_sel_143004_comb;
  wire [15:0] p1_sel_143005_comb;
  wire [15:0] p1_smul_143006_comb;
  wire [15:0] p1_sel_143007_comb;
  wire [15:0] p1_smul_143008_comb;
  wire [15:0] p1_smul_143009_comb;
  wire [15:0] p1_smul_143010_comb;
  wire [15:0] p1_smul_143011_comb;
  wire [15:0] p1_smul_143012_comb;
  wire [15:0] p1_smul_143013_comb;
  wire [15:0] p1_smul_143014_comb;
  wire [15:0] p1_smul_143015_comb;
  wire [15:0] p1_smul_143016_comb;
  wire [15:0] p1_smul_143017_comb;
  wire [15:0] p1_smul_143018_comb;
  wire [15:0] p1_smul_143019_comb;
  wire [15:0] p1_smul_143020_comb;
  wire [15:0] p1_smul_143021_comb;
  wire [15:0] p1_smul_143022_comb;
  wire [15:0] p1_smul_143023_comb;
  wire [15:0] p1_smul_143024_comb;
  wire [15:0] p1_smul_143025_comb;
  wire [15:0] p1_smul_143026_comb;
  wire [15:0] p1_smul_143027_comb;
  wire [15:0] p1_smul_143028_comb;
  wire [15:0] p1_smul_143029_comb;
  wire [15:0] p1_smul_143030_comb;
  wire [15:0] p1_smul_143031_comb;
  wire [15:0] p1_smul_143032_comb;
  wire [15:0] p1_smul_143033_comb;
  wire [15:0] p1_smul_143034_comb;
  wire [15:0] p1_smul_143035_comb;
  wire [15:0] p1_smul_143036_comb;
  wire [15:0] p1_smul_143037_comb;
  wire [15:0] p1_smul_143038_comb;
  wire [15:0] p1_smul_143039_comb;
  wire [15:0] p1_smul_143040_comb;
  wire [15:0] p1_smul_143041_comb;
  wire [15:0] p1_smul_143042_comb;
  wire [15:0] p1_smul_143043_comb;
  wire [15:0] p1_smul_143044_comb;
  wire [15:0] p1_smul_143045_comb;
  wire [15:0] p1_smul_143046_comb;
  wire [15:0] p1_smul_143047_comb;
  wire [15:0] p1_smul_143048_comb;
  wire [15:0] p1_smul_143049_comb;
  wire [15:0] p1_smul_143050_comb;
  wire [15:0] p1_smul_143051_comb;
  wire [15:0] p1_smul_143052_comb;
  wire [15:0] p1_smul_143053_comb;
  wire [15:0] p1_smul_143054_comb;
  wire [15:0] p1_smul_143055_comb;
  wire [15:0] p1_smul_143056_comb;
  wire [15:0] p1_smul_143057_comb;
  wire [15:0] p1_smul_143058_comb;
  wire [15:0] p1_smul_143059_comb;
  wire [15:0] p1_smul_143060_comb;
  wire [15:0] p1_smul_143061_comb;
  wire [15:0] p1_smul_143062_comb;
  wire [15:0] p1_smul_143063_comb;
  wire [15:0] p1_smul_143064_comb;
  wire [15:0] p1_smul_143065_comb;
  wire [15:0] p1_smul_143066_comb;
  wire [15:0] p1_smul_143067_comb;
  wire [15:0] p1_smul_143068_comb;
  wire [15:0] p1_smul_143069_comb;
  wire [15:0] p1_smul_143070_comb;
  wire [15:0] p1_smul_143071_comb;
  wire [15:0] p1_smul_143072_comb;
  wire [15:0] p1_sel_143073_comb;
  wire [15:0] p1_smul_143074_comb;
  wire [15:0] p1_sel_143075_comb;
  wire [15:0] p1_smul_143076_comb;
  wire [15:0] p1_smul_143077_comb;
  wire [15:0] p1_sel_143078_comb;
  wire [15:0] p1_smul_143079_comb;
  wire [15:0] p1_sel_143080_comb;
  wire [15:0] p1_sel_143081_comb;
  wire [15:0] p1_smul_143082_comb;
  wire [15:0] p1_sel_143083_comb;
  wire [15:0] p1_smul_143084_comb;
  wire [15:0] p1_smul_143085_comb;
  wire [15:0] p1_sel_143086_comb;
  wire [15:0] p1_smul_143087_comb;
  wire [15:0] p1_sel_143088_comb;
  wire [15:0] p1_sel_143089_comb;
  wire [15:0] p1_smul_143090_comb;
  wire [15:0] p1_sel_143091_comb;
  wire [15:0] p1_smul_143092_comb;
  wire [15:0] p1_smul_143093_comb;
  wire [15:0] p1_sel_143094_comb;
  wire [15:0] p1_smul_143095_comb;
  wire [15:0] p1_sel_143096_comb;
  wire [15:0] p1_sel_143097_comb;
  wire [15:0] p1_smul_143098_comb;
  wire [15:0] p1_sel_143099_comb;
  wire [15:0] p1_smul_143100_comb;
  wire [15:0] p1_smul_143101_comb;
  wire [15:0] p1_sel_143102_comb;
  wire [15:0] p1_smul_143103_comb;
  wire [15:0] p1_sel_143104_comb;
  wire [15:0] p1_sel_143105_comb;
  wire [15:0] p1_smul_143106_comb;
  wire [15:0] p1_sel_143107_comb;
  wire [15:0] p1_smul_143108_comb;
  wire [15:0] p1_smul_143109_comb;
  wire [15:0] p1_sel_143110_comb;
  wire [15:0] p1_smul_143111_comb;
  wire [15:0] p1_sel_143112_comb;
  wire [15:0] p1_sel_143113_comb;
  wire [15:0] p1_smul_143114_comb;
  wire [15:0] p1_sel_143115_comb;
  wire [15:0] p1_smul_143116_comb;
  wire [15:0] p1_smul_143117_comb;
  wire [15:0] p1_sel_143118_comb;
  wire [15:0] p1_smul_143119_comb;
  wire [15:0] p1_sel_143120_comb;
  wire [15:0] p1_sel_143121_comb;
  wire [15:0] p1_smul_143122_comb;
  wire [15:0] p1_sel_143123_comb;
  wire [15:0] p1_smul_143124_comb;
  wire [15:0] p1_smul_143125_comb;
  wire [15:0] p1_sel_143126_comb;
  wire [15:0] p1_smul_143127_comb;
  wire [15:0] p1_sel_143128_comb;
  wire [15:0] p1_sel_143129_comb;
  wire [15:0] p1_smul_143130_comb;
  wire [15:0] p1_sel_143131_comb;
  wire [15:0] p1_smul_143132_comb;
  wire [15:0] p1_smul_143133_comb;
  wire [15:0] p1_sel_143134_comb;
  wire [15:0] p1_smul_143135_comb;
  wire [15:0] p1_sel_143136_comb;
  wire [15:0] p1_sel_143137_comb;
  wire [15:0] p1_sel_143138_comb;
  wire [15:0] p1_sel_143139_comb;
  wire [15:0] p1_sel_143140_comb;
  wire [15:0] p1_sel_143141_comb;
  wire [15:0] p1_sel_143142_comb;
  wire [15:0] p1_sel_143143_comb;
  wire [15:0] p1_sel_143144_comb;
  wire [15:0] p1_sel_143145_comb;
  wire [15:0] p1_sel_143146_comb;
  wire [15:0] p1_sel_143147_comb;
  wire [15:0] p1_sel_143148_comb;
  wire [15:0] p1_sel_143149_comb;
  wire [15:0] p1_sel_143150_comb;
  wire [15:0] p1_sel_143151_comb;
  wire [15:0] p1_sel_143152_comb;
  wire [15:0] p1_sel_143153_comb;
  wire [15:0] p1_sel_143154_comb;
  wire [15:0] p1_sel_143155_comb;
  wire [15:0] p1_sel_143156_comb;
  wire [15:0] p1_sel_143157_comb;
  wire [15:0] p1_sel_143158_comb;
  wire [15:0] p1_sel_143159_comb;
  wire [15:0] p1_sel_143160_comb;
  wire [15:0] p1_sel_143161_comb;
  wire [15:0] p1_sel_143162_comb;
  wire [15:0] p1_sel_143163_comb;
  wire [15:0] p1_sel_143164_comb;
  wire [15:0] p1_sel_143165_comb;
  wire [15:0] p1_sel_143166_comb;
  wire [15:0] p1_sel_143167_comb;
  wire [15:0] p1_sel_143168_comb;
  wire [15:0] p1_sel_143169_comb;
  wire [15:0] p1_sel_143170_comb;
  wire [15:0] p1_sel_143171_comb;
  wire [15:0] p1_sel_143172_comb;
  wire [15:0] p1_sel_143173_comb;
  wire [15:0] p1_sel_143174_comb;
  wire [15:0] p1_sel_143175_comb;
  wire [15:0] p1_sel_143176_comb;
  wire [15:0] p1_sel_143177_comb;
  wire [15:0] p1_sel_143178_comb;
  wire [15:0] p1_sel_143179_comb;
  wire [15:0] p1_sel_143180_comb;
  wire [15:0] p1_sel_143181_comb;
  wire [15:0] p1_sel_143182_comb;
  wire [15:0] p1_sel_143183_comb;
  wire [15:0] p1_sel_143184_comb;
  wire [15:0] p1_sel_143185_comb;
  wire [15:0] p1_sel_143186_comb;
  wire [15:0] p1_sel_143187_comb;
  wire [15:0] p1_sel_143188_comb;
  wire [15:0] p1_sel_143189_comb;
  wire [15:0] p1_sel_143190_comb;
  wire [15:0] p1_sel_143191_comb;
  wire [15:0] p1_sel_143192_comb;
  wire [15:0] p1_sel_143193_comb;
  wire [15:0] p1_sel_143194_comb;
  wire [15:0] p1_sel_143195_comb;
  wire [15:0] p1_sel_143196_comb;
  wire [15:0] p1_sel_143197_comb;
  wire [15:0] p1_sel_143198_comb;
  wire [15:0] p1_sel_143199_comb;
  wire [15:0] p1_sel_143200_comb;
  wire [15:0] p1_sel_143201_comb;
  wire [15:0] p1_sel_143202_comb;
  wire [15:0] p1_smul_143203_comb;
  wire [15:0] p1_smul_143204_comb;
  wire [15:0] p1_smul_143205_comb;
  wire [15:0] p1_smul_143206_comb;
  wire [15:0] p1_sel_143207_comb;
  wire [15:0] p1_sel_143208_comb;
  wire [15:0] p1_sel_143209_comb;
  wire [15:0] p1_sel_143210_comb;
  wire [15:0] p1_smul_143211_comb;
  wire [15:0] p1_smul_143212_comb;
  wire [15:0] p1_smul_143213_comb;
  wire [15:0] p1_smul_143214_comb;
  wire [15:0] p1_sel_143215_comb;
  wire [15:0] p1_sel_143216_comb;
  wire [15:0] p1_sel_143217_comb;
  wire [15:0] p1_sel_143218_comb;
  wire [15:0] p1_smul_143219_comb;
  wire [15:0] p1_smul_143220_comb;
  wire [15:0] p1_smul_143221_comb;
  wire [15:0] p1_smul_143222_comb;
  wire [15:0] p1_sel_143223_comb;
  wire [15:0] p1_sel_143224_comb;
  wire [15:0] p1_sel_143225_comb;
  wire [15:0] p1_sel_143226_comb;
  wire [15:0] p1_smul_143227_comb;
  wire [15:0] p1_smul_143228_comb;
  wire [15:0] p1_smul_143229_comb;
  wire [15:0] p1_smul_143230_comb;
  wire [15:0] p1_sel_143231_comb;
  wire [15:0] p1_sel_143232_comb;
  wire [15:0] p1_sel_143233_comb;
  wire [15:0] p1_sel_143234_comb;
  wire [15:0] p1_smul_143235_comb;
  wire [15:0] p1_smul_143236_comb;
  wire [15:0] p1_smul_143237_comb;
  wire [15:0] p1_smul_143238_comb;
  wire [15:0] p1_sel_143239_comb;
  wire [15:0] p1_sel_143240_comb;
  wire [15:0] p1_sel_143241_comb;
  wire [15:0] p1_sel_143242_comb;
  wire [15:0] p1_smul_143243_comb;
  wire [15:0] p1_smul_143244_comb;
  wire [15:0] p1_smul_143245_comb;
  wire [15:0] p1_smul_143246_comb;
  wire [15:0] p1_sel_143247_comb;
  wire [15:0] p1_sel_143248_comb;
  wire [15:0] p1_sel_143249_comb;
  wire [15:0] p1_sel_143250_comb;
  wire [15:0] p1_smul_143251_comb;
  wire [15:0] p1_smul_143252_comb;
  wire [15:0] p1_smul_143253_comb;
  wire [15:0] p1_smul_143254_comb;
  wire [15:0] p1_sel_143255_comb;
  wire [15:0] p1_sel_143256_comb;
  wire [15:0] p1_sel_143257_comb;
  wire [15:0] p1_sel_143258_comb;
  wire [15:0] p1_smul_143259_comb;
  wire [15:0] p1_smul_143260_comb;
  wire [15:0] p1_smul_143261_comb;
  wire [15:0] p1_smul_143262_comb;
  wire [15:0] p1_sel_143263_comb;
  wire [15:0] p1_sel_143264_comb;
  wire [31:0] p1_sum__520_comb;
  wire [31:0] p1_sum__521_comb;
  wire [31:0] p1_sum__522_comb;
  wire [31:0] p1_sum__523_comb;
  wire [31:0] p1_sum__464_comb;
  wire [31:0] p1_sum__465_comb;
  wire [31:0] p1_sum__466_comb;
  wire [31:0] p1_sum__467_comb;
  wire [31:0] p1_sum__408_comb;
  wire [31:0] p1_sum__409_comb;
  wire [31:0] p1_sum__410_comb;
  wire [31:0] p1_sum__411_comb;
  wire [31:0] p1_sum__352_comb;
  wire [31:0] p1_sum__353_comb;
  wire [31:0] p1_sum__354_comb;
  wire [31:0] p1_sum__355_comb;
  wire [31:0] p1_sum__296_comb;
  wire [31:0] p1_sum__297_comb;
  wire [31:0] p1_sum__298_comb;
  wire [31:0] p1_sum__299_comb;
  wire [31:0] p1_sum__240_comb;
  wire [31:0] p1_sum__241_comb;
  wire [31:0] p1_sum__242_comb;
  wire [31:0] p1_sum__243_comb;
  wire [31:0] p1_sum__184_comb;
  wire [31:0] p1_sum__185_comb;
  wire [31:0] p1_sum__186_comb;
  wire [31:0] p1_sum__187_comb;
  wire [31:0] p1_sum__128_comb;
  wire [31:0] p1_sum__129_comb;
  wire [31:0] p1_sum__130_comb;
  wire [31:0] p1_sum__131_comb;
  wire [31:0] p1_sum__524_comb;
  wire [31:0] p1_sum__525_comb;
  wire [31:0] p1_sum__468_comb;
  wire [31:0] p1_sum__469_comb;
  wire [31:0] p1_sum__412_comb;
  wire [31:0] p1_sum__413_comb;
  wire [31:0] p1_sum__356_comb;
  wire [31:0] p1_sum__357_comb;
  wire [31:0] p1_sum__300_comb;
  wire [31:0] p1_sum__301_comb;
  wire [31:0] p1_sum__244_comb;
  wire [31:0] p1_sum__245_comb;
  wire [31:0] p1_sum__188_comb;
  wire [31:0] p1_sum__189_comb;
  wire [31:0] p1_sum__132_comb;
  wire [31:0] p1_sum__133_comb;
  wire [16:0] p1_add_143761_comb;
  wire [16:0] p1_add_143762_comb;
  wire [16:0] p1_add_143763_comb;
  wire [16:0] p1_add_143764_comb;
  wire [16:0] p1_add_143765_comb;
  wire [16:0] p1_add_143766_comb;
  wire [16:0] p1_add_143767_comb;
  wire [16:0] p1_add_143768_comb;
  wire [16:0] p1_add_143769_comb;
  wire [16:0] p1_add_143770_comb;
  wire [16:0] p1_add_143771_comb;
  wire [16:0] p1_add_143772_comb;
  wire [16:0] p1_add_143773_comb;
  wire [16:0] p1_add_143774_comb;
  wire [16:0] p1_add_143775_comb;
  wire [16:0] p1_add_143776_comb;
  wire [16:0] p1_add_143777_comb;
  wire [16:0] p1_add_143778_comb;
  wire [16:0] p1_add_143779_comb;
  wire [16:0] p1_add_143780_comb;
  wire [16:0] p1_add_143781_comb;
  wire [16:0] p1_add_143782_comb;
  wire [16:0] p1_add_143783_comb;
  wire [16:0] p1_add_143784_comb;
  wire [16:0] p1_add_143785_comb;
  wire [16:0] p1_add_143786_comb;
  wire [16:0] p1_add_143787_comb;
  wire [16:0] p1_add_143788_comb;
  wire [16:0] p1_add_143789_comb;
  wire [16:0] p1_add_143790_comb;
  wire [16:0] p1_add_143791_comb;
  wire [16:0] p1_add_143792_comb;
  wire [16:0] p1_add_143793_comb;
  wire [16:0] p1_add_143794_comb;
  wire [16:0] p1_add_143795_comb;
  wire [16:0] p1_add_143796_comb;
  wire [16:0] p1_add_143797_comb;
  wire [16:0] p1_add_143798_comb;
  wire [16:0] p1_add_143799_comb;
  wire [16:0] p1_add_143800_comb;
  wire [16:0] p1_add_143801_comb;
  wire [16:0] p1_add_143802_comb;
  wire [16:0] p1_add_143803_comb;
  wire [16:0] p1_add_143804_comb;
  wire [16:0] p1_add_143805_comb;
  wire [16:0] p1_add_143806_comb;
  wire [16:0] p1_add_143807_comb;
  wire [16:0] p1_add_143808_comb;
  wire [16:0] p1_add_143809_comb;
  wire [16:0] p1_add_143810_comb;
  wire [16:0] p1_add_143811_comb;
  wire [16:0] p1_add_143812_comb;
  wire [16:0] p1_add_143813_comb;
  wire [16:0] p1_add_143814_comb;
  wire [16:0] p1_add_143815_comb;
  wire [16:0] p1_add_143816_comb;
  wire [16:0] p1_add_143817_comb;
  wire [16:0] p1_add_143818_comb;
  wire [16:0] p1_add_143819_comb;
  wire [16:0] p1_add_143820_comb;
  wire [16:0] p1_add_143821_comb;
  wire [16:0] p1_add_143822_comb;
  wire [16:0] p1_add_143823_comb;
  wire [16:0] p1_add_143824_comb;
  wire [16:0] p1_add_143825_comb;
  wire [16:0] p1_add_143826_comb;
  wire [16:0] p1_add_143827_comb;
  wire [16:0] p1_add_143828_comb;
  wire [16:0] p1_add_143829_comb;
  wire [16:0] p1_add_143830_comb;
  wire [16:0] p1_add_143831_comb;
  wire [16:0] p1_add_143832_comb;
  wire [16:0] p1_add_143833_comb;
  wire [16:0] p1_add_143834_comb;
  wire [16:0] p1_add_143835_comb;
  wire [16:0] p1_add_143836_comb;
  wire [16:0] p1_add_143837_comb;
  wire [16:0] p1_add_143838_comb;
  wire [16:0] p1_add_143839_comb;
  wire [16:0] p1_add_143840_comb;
  wire [16:0] p1_add_143841_comb;
  wire [16:0] p1_add_143842_comb;
  wire [16:0] p1_add_143843_comb;
  wire [16:0] p1_add_143844_comb;
  wire [16:0] p1_add_143845_comb;
  wire [16:0] p1_add_143846_comb;
  wire [16:0] p1_add_143847_comb;
  wire [16:0] p1_add_143848_comb;
  wire [16:0] p1_add_143849_comb;
  wire [16:0] p1_add_143850_comb;
  wire [16:0] p1_add_143851_comb;
  wire [16:0] p1_add_143852_comb;
  wire [16:0] p1_add_143853_comb;
  wire [16:0] p1_add_143854_comb;
  wire [16:0] p1_add_143855_comb;
  wire [16:0] p1_add_143856_comb;
  wire [16:0] p1_add_143857_comb;
  wire [16:0] p1_add_143858_comb;
  wire [16:0] p1_add_143859_comb;
  wire [16:0] p1_add_143860_comb;
  wire [16:0] p1_add_143861_comb;
  wire [16:0] p1_add_143862_comb;
  wire [16:0] p1_add_143863_comb;
  wire [16:0] p1_add_143864_comb;
  wire [16:0] p1_add_143865_comb;
  wire [16:0] p1_add_143866_comb;
  wire [16:0] p1_add_143867_comb;
  wire [16:0] p1_add_143868_comb;
  wire [16:0] p1_add_143869_comb;
  wire [16:0] p1_add_143870_comb;
  wire [16:0] p1_add_143871_comb;
  wire [16:0] p1_add_143872_comb;
  wire [16:0] p1_add_143873_comb;
  wire [16:0] p1_add_143874_comb;
  wire [16:0] p1_add_143875_comb;
  wire [16:0] p1_add_143876_comb;
  wire [16:0] p1_add_143877_comb;
  wire [16:0] p1_add_143878_comb;
  wire [16:0] p1_add_143879_comb;
  wire [16:0] p1_add_143880_comb;
  wire [16:0] p1_add_143881_comb;
  wire [16:0] p1_add_143882_comb;
  wire [16:0] p1_add_143883_comb;
  wire [16:0] p1_add_143884_comb;
  wire [16:0] p1_add_143885_comb;
  wire [16:0] p1_add_143886_comb;
  wire [16:0] p1_add_143887_comb;
  wire [16:0] p1_add_143888_comb;
  wire [16:0] p1_add_143889_comb;
  wire [16:0] p1_add_143890_comb;
  wire [16:0] p1_add_143891_comb;
  wire [16:0] p1_add_143892_comb;
  wire [16:0] p1_add_143893_comb;
  wire [16:0] p1_add_143894_comb;
  wire [16:0] p1_add_143895_comb;
  wire [16:0] p1_add_143896_comb;
  wire [16:0] p1_add_143897_comb;
  wire [16:0] p1_add_143898_comb;
  wire [16:0] p1_add_143899_comb;
  wire [16:0] p1_add_143900_comb;
  wire [16:0] p1_add_143901_comb;
  wire [16:0] p1_add_143902_comb;
  wire [16:0] p1_add_143903_comb;
  wire [16:0] p1_add_143904_comb;
  wire [16:0] p1_add_143905_comb;
  wire [16:0] p1_add_143906_comb;
  wire [16:0] p1_add_143907_comb;
  wire [16:0] p1_add_143908_comb;
  wire [16:0] p1_add_143909_comb;
  wire [16:0] p1_add_143910_comb;
  wire [16:0] p1_add_143911_comb;
  wire [16:0] p1_add_143912_comb;
  wire [16:0] p1_add_143913_comb;
  wire [16:0] p1_add_143914_comb;
  wire [16:0] p1_add_143915_comb;
  wire [16:0] p1_add_143916_comb;
  wire [16:0] p1_add_143917_comb;
  wire [16:0] p1_add_143918_comb;
  wire [16:0] p1_add_143919_comb;
  wire [16:0] p1_add_143920_comb;
  wire [16:0] p1_add_143921_comb;
  wire [16:0] p1_add_143922_comb;
  wire [16:0] p1_add_143923_comb;
  wire [16:0] p1_add_143924_comb;
  wire [16:0] p1_add_143925_comb;
  wire [16:0] p1_add_143926_comb;
  wire [16:0] p1_add_143927_comb;
  wire [16:0] p1_add_143928_comb;
  wire [16:0] p1_add_143929_comb;
  wire [16:0] p1_add_143930_comb;
  wire [16:0] p1_add_143931_comb;
  wire [16:0] p1_add_143932_comb;
  wire [16:0] p1_add_143933_comb;
  wire [16:0] p1_add_143934_comb;
  wire [16:0] p1_add_143935_comb;
  wire [16:0] p1_add_143936_comb;
  wire [16:0] p1_add_143937_comb;
  wire [16:0] p1_add_143938_comb;
  wire [16:0] p1_add_143939_comb;
  wire [16:0] p1_add_143940_comb;
  wire [16:0] p1_add_143941_comb;
  wire [16:0] p1_add_143942_comb;
  wire [16:0] p1_add_143943_comb;
  wire [16:0] p1_add_143944_comb;
  wire [16:0] p1_add_143945_comb;
  wire [16:0] p1_add_143946_comb;
  wire [16:0] p1_add_143947_comb;
  wire [16:0] p1_add_143948_comb;
  wire [16:0] p1_add_143949_comb;
  wire [16:0] p1_add_143950_comb;
  wire [16:0] p1_add_143951_comb;
  wire [16:0] p1_add_143952_comb;
  wire [16:0] p1_add_143953_comb;
  wire [16:0] p1_add_143954_comb;
  wire [16:0] p1_add_143955_comb;
  wire [16:0] p1_add_143956_comb;
  wire [16:0] p1_add_143957_comb;
  wire [16:0] p1_add_143958_comb;
  wire [16:0] p1_add_143959_comb;
  wire [16:0] p1_add_143960_comb;
  wire [16:0] p1_add_143961_comb;
  wire [16:0] p1_add_143962_comb;
  wire [16:0] p1_add_143963_comb;
  wire [16:0] p1_add_143964_comb;
  wire [16:0] p1_add_143965_comb;
  wire [16:0] p1_add_143966_comb;
  wire [16:0] p1_add_143967_comb;
  wire [16:0] p1_add_143968_comb;
  wire [16:0] p1_add_143969_comb;
  wire [16:0] p1_add_143970_comb;
  wire [16:0] p1_add_143971_comb;
  wire [16:0] p1_add_143972_comb;
  wire [16:0] p1_add_143973_comb;
  wire [16:0] p1_add_143974_comb;
  wire [16:0] p1_add_143975_comb;
  wire [16:0] p1_add_143976_comb;
  wire [16:0] p1_add_143977_comb;
  wire [16:0] p1_add_143978_comb;
  wire [16:0] p1_add_143979_comb;
  wire [16:0] p1_add_143980_comb;
  wire [16:0] p1_add_143981_comb;
  wire [16:0] p1_add_143982_comb;
  wire [16:0] p1_add_143983_comb;
  wire [16:0] p1_add_143984_comb;
  wire [31:0] p1_sum__526_comb;
  wire [31:0] p1_sum__470_comb;
  wire [31:0] p1_sum__414_comb;
  wire [31:0] p1_sum__358_comb;
  wire [31:0] p1_sum__302_comb;
  wire [31:0] p1_sum__246_comb;
  wire [31:0] p1_sum__190_comb;
  wire [31:0] p1_sum__134_comb;
  wire [24:0] p1_sum__1580_comb;
  wire [24:0] p1_sum__1581_comb;
  wire [24:0] p1_sum__1582_comb;
  wire [24:0] p1_sum__1583_comb;
  wire [24:0] p1_sum__1552_comb;
  wire [24:0] p1_sum__1553_comb;
  wire [24:0] p1_sum__1554_comb;
  wire [24:0] p1_sum__1555_comb;
  wire [24:0] p1_sum__1524_comb;
  wire [24:0] p1_sum__1525_comb;
  wire [24:0] p1_sum__1526_comb;
  wire [24:0] p1_sum__1527_comb;
  wire [24:0] p1_sum__1496_comb;
  wire [24:0] p1_sum__1497_comb;
  wire [24:0] p1_sum__1498_comb;
  wire [24:0] p1_sum__1499_comb;
  wire [24:0] p1_sum__1468_comb;
  wire [24:0] p1_sum__1469_comb;
  wire [24:0] p1_sum__1470_comb;
  wire [24:0] p1_sum__1471_comb;
  wire [24:0] p1_sum__1440_comb;
  wire [24:0] p1_sum__1441_comb;
  wire [24:0] p1_sum__1442_comb;
  wire [24:0] p1_sum__1443_comb;
  wire [24:0] p1_sum__1412_comb;
  wire [24:0] p1_sum__1413_comb;
  wire [24:0] p1_sum__1414_comb;
  wire [24:0] p1_sum__1415_comb;
  wire [24:0] p1_sum__1384_comb;
  wire [24:0] p1_sum__1385_comb;
  wire [24:0] p1_sum__1386_comb;
  wire [24:0] p1_sum__1387_comb;
  wire [24:0] p1_sum__1576_comb;
  wire [24:0] p1_sum__1577_comb;
  wire [24:0] p1_sum__1578_comb;
  wire [24:0] p1_sum__1579_comb;
  wire [24:0] p1_sum__1548_comb;
  wire [24:0] p1_sum__1549_comb;
  wire [24:0] p1_sum__1550_comb;
  wire [24:0] p1_sum__1551_comb;
  wire [24:0] p1_sum__1520_comb;
  wire [24:0] p1_sum__1521_comb;
  wire [24:0] p1_sum__1522_comb;
  wire [24:0] p1_sum__1523_comb;
  wire [24:0] p1_sum__1492_comb;
  wire [24:0] p1_sum__1493_comb;
  wire [24:0] p1_sum__1494_comb;
  wire [24:0] p1_sum__1495_comb;
  wire [24:0] p1_sum__1464_comb;
  wire [24:0] p1_sum__1465_comb;
  wire [24:0] p1_sum__1466_comb;
  wire [24:0] p1_sum__1467_comb;
  wire [24:0] p1_sum__1436_comb;
  wire [24:0] p1_sum__1437_comb;
  wire [24:0] p1_sum__1438_comb;
  wire [24:0] p1_sum__1439_comb;
  wire [24:0] p1_sum__1408_comb;
  wire [24:0] p1_sum__1409_comb;
  wire [24:0] p1_sum__1410_comb;
  wire [24:0] p1_sum__1411_comb;
  wire [24:0] p1_sum__1380_comb;
  wire [24:0] p1_sum__1381_comb;
  wire [24:0] p1_sum__1382_comb;
  wire [24:0] p1_sum__1383_comb;
  wire [24:0] p1_sum__1572_comb;
  wire [24:0] p1_sum__1573_comb;
  wire [24:0] p1_sum__1574_comb;
  wire [24:0] p1_sum__1575_comb;
  wire [24:0] p1_sum__1544_comb;
  wire [24:0] p1_sum__1545_comb;
  wire [24:0] p1_sum__1546_comb;
  wire [24:0] p1_sum__1547_comb;
  wire [24:0] p1_sum__1516_comb;
  wire [24:0] p1_sum__1517_comb;
  wire [24:0] p1_sum__1518_comb;
  wire [24:0] p1_sum__1519_comb;
  wire [24:0] p1_sum__1488_comb;
  wire [24:0] p1_sum__1489_comb;
  wire [24:0] p1_sum__1490_comb;
  wire [24:0] p1_sum__1491_comb;
  wire [24:0] p1_sum__1460_comb;
  wire [24:0] p1_sum__1461_comb;
  wire [24:0] p1_sum__1462_comb;
  wire [24:0] p1_sum__1463_comb;
  wire [24:0] p1_sum__1432_comb;
  wire [24:0] p1_sum__1433_comb;
  wire [24:0] p1_sum__1434_comb;
  wire [24:0] p1_sum__1435_comb;
  wire [24:0] p1_sum__1404_comb;
  wire [24:0] p1_sum__1405_comb;
  wire [24:0] p1_sum__1406_comb;
  wire [24:0] p1_sum__1407_comb;
  wire [24:0] p1_sum__1376_comb;
  wire [24:0] p1_sum__1377_comb;
  wire [24:0] p1_sum__1378_comb;
  wire [24:0] p1_sum__1379_comb;
  wire [24:0] p1_sum__1568_comb;
  wire [24:0] p1_sum__1569_comb;
  wire [24:0] p1_sum__1570_comb;
  wire [24:0] p1_sum__1571_comb;
  wire [24:0] p1_sum__1540_comb;
  wire [24:0] p1_sum__1541_comb;
  wire [24:0] p1_sum__1542_comb;
  wire [24:0] p1_sum__1543_comb;
  wire [24:0] p1_sum__1512_comb;
  wire [24:0] p1_sum__1513_comb;
  wire [24:0] p1_sum__1514_comb;
  wire [24:0] p1_sum__1515_comb;
  wire [24:0] p1_sum__1484_comb;
  wire [24:0] p1_sum__1485_comb;
  wire [24:0] p1_sum__1486_comb;
  wire [24:0] p1_sum__1487_comb;
  wire [24:0] p1_sum__1456_comb;
  wire [24:0] p1_sum__1457_comb;
  wire [24:0] p1_sum__1458_comb;
  wire [24:0] p1_sum__1459_comb;
  wire [24:0] p1_sum__1428_comb;
  wire [24:0] p1_sum__1429_comb;
  wire [24:0] p1_sum__1430_comb;
  wire [24:0] p1_sum__1431_comb;
  wire [24:0] p1_sum__1400_comb;
  wire [24:0] p1_sum__1401_comb;
  wire [24:0] p1_sum__1402_comb;
  wire [24:0] p1_sum__1403_comb;
  wire [24:0] p1_sum__1372_comb;
  wire [24:0] p1_sum__1373_comb;
  wire [24:0] p1_sum__1374_comb;
  wire [24:0] p1_sum__1375_comb;
  wire [24:0] p1_sum__1564_comb;
  wire [24:0] p1_sum__1565_comb;
  wire [24:0] p1_sum__1566_comb;
  wire [24:0] p1_sum__1567_comb;
  wire [24:0] p1_sum__1536_comb;
  wire [24:0] p1_sum__1537_comb;
  wire [24:0] p1_sum__1538_comb;
  wire [24:0] p1_sum__1539_comb;
  wire [24:0] p1_sum__1508_comb;
  wire [24:0] p1_sum__1509_comb;
  wire [24:0] p1_sum__1510_comb;
  wire [24:0] p1_sum__1511_comb;
  wire [24:0] p1_sum__1480_comb;
  wire [24:0] p1_sum__1481_comb;
  wire [24:0] p1_sum__1482_comb;
  wire [24:0] p1_sum__1483_comb;
  wire [24:0] p1_sum__1452_comb;
  wire [24:0] p1_sum__1453_comb;
  wire [24:0] p1_sum__1454_comb;
  wire [24:0] p1_sum__1455_comb;
  wire [24:0] p1_sum__1424_comb;
  wire [24:0] p1_sum__1425_comb;
  wire [24:0] p1_sum__1426_comb;
  wire [24:0] p1_sum__1427_comb;
  wire [24:0] p1_sum__1396_comb;
  wire [24:0] p1_sum__1397_comb;
  wire [24:0] p1_sum__1398_comb;
  wire [24:0] p1_sum__1399_comb;
  wire [24:0] p1_sum__1368_comb;
  wire [24:0] p1_sum__1369_comb;
  wire [24:0] p1_sum__1370_comb;
  wire [24:0] p1_sum__1371_comb;
  wire [24:0] p1_sum__1560_comb;
  wire [24:0] p1_sum__1561_comb;
  wire [24:0] p1_sum__1562_comb;
  wire [24:0] p1_sum__1563_comb;
  wire [24:0] p1_sum__1532_comb;
  wire [24:0] p1_sum__1533_comb;
  wire [24:0] p1_sum__1534_comb;
  wire [24:0] p1_sum__1535_comb;
  wire [24:0] p1_sum__1504_comb;
  wire [24:0] p1_sum__1505_comb;
  wire [24:0] p1_sum__1506_comb;
  wire [24:0] p1_sum__1507_comb;
  wire [24:0] p1_sum__1476_comb;
  wire [24:0] p1_sum__1477_comb;
  wire [24:0] p1_sum__1478_comb;
  wire [24:0] p1_sum__1479_comb;
  wire [24:0] p1_sum__1448_comb;
  wire [24:0] p1_sum__1449_comb;
  wire [24:0] p1_sum__1450_comb;
  wire [24:0] p1_sum__1451_comb;
  wire [24:0] p1_sum__1420_comb;
  wire [24:0] p1_sum__1421_comb;
  wire [24:0] p1_sum__1422_comb;
  wire [24:0] p1_sum__1423_comb;
  wire [24:0] p1_sum__1392_comb;
  wire [24:0] p1_sum__1393_comb;
  wire [24:0] p1_sum__1394_comb;
  wire [24:0] p1_sum__1395_comb;
  wire [24:0] p1_sum__1364_comb;
  wire [24:0] p1_sum__1365_comb;
  wire [24:0] p1_sum__1366_comb;
  wire [24:0] p1_sum__1367_comb;
  wire [24:0] p1_sum__1556_comb;
  wire [24:0] p1_sum__1557_comb;
  wire [24:0] p1_sum__1558_comb;
  wire [24:0] p1_sum__1559_comb;
  wire [24:0] p1_sum__1528_comb;
  wire [24:0] p1_sum__1529_comb;
  wire [24:0] p1_sum__1530_comb;
  wire [24:0] p1_sum__1531_comb;
  wire [24:0] p1_sum__1500_comb;
  wire [24:0] p1_sum__1501_comb;
  wire [24:0] p1_sum__1502_comb;
  wire [24:0] p1_sum__1503_comb;
  wire [24:0] p1_sum__1472_comb;
  wire [24:0] p1_sum__1473_comb;
  wire [24:0] p1_sum__1474_comb;
  wire [24:0] p1_sum__1475_comb;
  wire [24:0] p1_sum__1444_comb;
  wire [24:0] p1_sum__1445_comb;
  wire [24:0] p1_sum__1446_comb;
  wire [24:0] p1_sum__1447_comb;
  wire [24:0] p1_sum__1416_comb;
  wire [24:0] p1_sum__1417_comb;
  wire [24:0] p1_sum__1418_comb;
  wire [24:0] p1_sum__1419_comb;
  wire [24:0] p1_sum__1388_comb;
  wire [24:0] p1_sum__1389_comb;
  wire [24:0] p1_sum__1390_comb;
  wire [24:0] p1_sum__1391_comb;
  wire [24:0] p1_sum__1360_comb;
  wire [24:0] p1_sum__1361_comb;
  wire [24:0] p1_sum__1362_comb;
  wire [24:0] p1_sum__1363_comb;
  wire [31:0] p1_umul_144225_comb;
  wire [31:0] p1_umul_144226_comb;
  wire [31:0] p1_umul_144227_comb;
  wire [31:0] p1_umul_144228_comb;
  wire [31:0] p1_umul_144229_comb;
  wire [31:0] p1_umul_144230_comb;
  wire [31:0] p1_umul_144231_comb;
  wire [31:0] p1_umul_144232_comb;
  wire [24:0] p1_sum__1246_comb;
  wire [24:0] p1_sum__1247_comb;
  wire [24:0] p1_sum__1232_comb;
  wire [24:0] p1_sum__1233_comb;
  wire [24:0] p1_sum__1218_comb;
  wire [24:0] p1_sum__1219_comb;
  wire [24:0] p1_sum__1204_comb;
  wire [24:0] p1_sum__1205_comb;
  wire [24:0] p1_sum__1190_comb;
  wire [24:0] p1_sum__1191_comb;
  wire [24:0] p1_sum__1176_comb;
  wire [24:0] p1_sum__1177_comb;
  wire [24:0] p1_sum__1162_comb;
  wire [24:0] p1_sum__1163_comb;
  wire [24:0] p1_sum__1148_comb;
  wire [24:0] p1_sum__1149_comb;
  wire [24:0] p1_sum__1244_comb;
  wire [24:0] p1_sum__1245_comb;
  wire [24:0] p1_sum__1230_comb;
  wire [24:0] p1_sum__1231_comb;
  wire [24:0] p1_sum__1216_comb;
  wire [24:0] p1_sum__1217_comb;
  wire [24:0] p1_sum__1202_comb;
  wire [24:0] p1_sum__1203_comb;
  wire [24:0] p1_sum__1188_comb;
  wire [24:0] p1_sum__1189_comb;
  wire [24:0] p1_sum__1174_comb;
  wire [24:0] p1_sum__1175_comb;
  wire [24:0] p1_sum__1160_comb;
  wire [24:0] p1_sum__1161_comb;
  wire [24:0] p1_sum__1146_comb;
  wire [24:0] p1_sum__1147_comb;
  wire [24:0] p1_sum__1242_comb;
  wire [24:0] p1_sum__1243_comb;
  wire [24:0] p1_sum__1228_comb;
  wire [24:0] p1_sum__1229_comb;
  wire [24:0] p1_sum__1214_comb;
  wire [24:0] p1_sum__1215_comb;
  wire [24:0] p1_sum__1200_comb;
  wire [24:0] p1_sum__1201_comb;
  wire [24:0] p1_sum__1186_comb;
  wire [24:0] p1_sum__1187_comb;
  wire [24:0] p1_sum__1172_comb;
  wire [24:0] p1_sum__1173_comb;
  wire [24:0] p1_sum__1158_comb;
  wire [24:0] p1_sum__1159_comb;
  wire [24:0] p1_sum__1144_comb;
  wire [24:0] p1_sum__1145_comb;
  wire [24:0] p1_sum__1240_comb;
  wire [24:0] p1_sum__1241_comb;
  wire [24:0] p1_sum__1226_comb;
  wire [24:0] p1_sum__1227_comb;
  wire [24:0] p1_sum__1212_comb;
  wire [24:0] p1_sum__1213_comb;
  wire [24:0] p1_sum__1198_comb;
  wire [24:0] p1_sum__1199_comb;
  wire [24:0] p1_sum__1184_comb;
  wire [24:0] p1_sum__1185_comb;
  wire [24:0] p1_sum__1170_comb;
  wire [24:0] p1_sum__1171_comb;
  wire [24:0] p1_sum__1156_comb;
  wire [24:0] p1_sum__1157_comb;
  wire [24:0] p1_sum__1142_comb;
  wire [24:0] p1_sum__1143_comb;
  wire [24:0] p1_sum__1238_comb;
  wire [24:0] p1_sum__1239_comb;
  wire [24:0] p1_sum__1224_comb;
  wire [24:0] p1_sum__1225_comb;
  wire [24:0] p1_sum__1210_comb;
  wire [24:0] p1_sum__1211_comb;
  wire [24:0] p1_sum__1196_comb;
  wire [24:0] p1_sum__1197_comb;
  wire [24:0] p1_sum__1182_comb;
  wire [24:0] p1_sum__1183_comb;
  wire [24:0] p1_sum__1168_comb;
  wire [24:0] p1_sum__1169_comb;
  wire [24:0] p1_sum__1154_comb;
  wire [24:0] p1_sum__1155_comb;
  wire [24:0] p1_sum__1140_comb;
  wire [24:0] p1_sum__1141_comb;
  wire [24:0] p1_sum__1236_comb;
  wire [24:0] p1_sum__1237_comb;
  wire [24:0] p1_sum__1222_comb;
  wire [24:0] p1_sum__1223_comb;
  wire [24:0] p1_sum__1208_comb;
  wire [24:0] p1_sum__1209_comb;
  wire [24:0] p1_sum__1194_comb;
  wire [24:0] p1_sum__1195_comb;
  wire [24:0] p1_sum__1180_comb;
  wire [24:0] p1_sum__1181_comb;
  wire [24:0] p1_sum__1166_comb;
  wire [24:0] p1_sum__1167_comb;
  wire [24:0] p1_sum__1152_comb;
  wire [24:0] p1_sum__1153_comb;
  wire [24:0] p1_sum__1138_comb;
  wire [24:0] p1_sum__1139_comb;
  wire [24:0] p1_sum__1234_comb;
  wire [24:0] p1_sum__1235_comb;
  wire [24:0] p1_sum__1220_comb;
  wire [24:0] p1_sum__1221_comb;
  wire [24:0] p1_sum__1206_comb;
  wire [24:0] p1_sum__1207_comb;
  wire [24:0] p1_sum__1192_comb;
  wire [24:0] p1_sum__1193_comb;
  wire [24:0] p1_sum__1178_comb;
  wire [24:0] p1_sum__1179_comb;
  wire [24:0] p1_sum__1164_comb;
  wire [24:0] p1_sum__1165_comb;
  wire [24:0] p1_sum__1150_comb;
  wire [24:0] p1_sum__1151_comb;
  wire [24:0] p1_sum__1136_comb;
  wire [24:0] p1_sum__1137_comb;
  wire [24:0] p1_sum__1079_comb;
  wire [24:0] p1_sum__1072_comb;
  wire [24:0] p1_sum__1065_comb;
  wire [24:0] p1_sum__1058_comb;
  wire [24:0] p1_sum__1051_comb;
  wire [24:0] p1_sum__1044_comb;
  wire [24:0] p1_sum__1037_comb;
  wire [24:0] p1_sum__1030_comb;
  wire [24:0] p1_sum__1078_comb;
  wire [24:0] p1_sum__1071_comb;
  wire [24:0] p1_sum__1064_comb;
  wire [24:0] p1_sum__1057_comb;
  wire [24:0] p1_sum__1050_comb;
  wire [24:0] p1_sum__1043_comb;
  wire [24:0] p1_sum__1036_comb;
  wire [24:0] p1_sum__1029_comb;
  wire [24:0] p1_sum__1077_comb;
  wire [24:0] p1_sum__1070_comb;
  wire [24:0] p1_sum__1063_comb;
  wire [24:0] p1_sum__1056_comb;
  wire [24:0] p1_sum__1049_comb;
  wire [24:0] p1_sum__1042_comb;
  wire [24:0] p1_sum__1035_comb;
  wire [24:0] p1_sum__1028_comb;
  wire [24:0] p1_sum__1076_comb;
  wire [24:0] p1_sum__1069_comb;
  wire [24:0] p1_sum__1062_comb;
  wire [24:0] p1_sum__1055_comb;
  wire [24:0] p1_sum__1048_comb;
  wire [24:0] p1_sum__1041_comb;
  wire [24:0] p1_sum__1034_comb;
  wire [24:0] p1_sum__1027_comb;
  wire [24:0] p1_sum__1075_comb;
  wire [24:0] p1_sum__1068_comb;
  wire [24:0] p1_sum__1061_comb;
  wire [24:0] p1_sum__1054_comb;
  wire [24:0] p1_sum__1047_comb;
  wire [24:0] p1_sum__1040_comb;
  wire [24:0] p1_sum__1033_comb;
  wire [24:0] p1_sum__1026_comb;
  wire [24:0] p1_sum__1074_comb;
  wire [24:0] p1_sum__1067_comb;
  wire [24:0] p1_sum__1060_comb;
  wire [24:0] p1_sum__1053_comb;
  wire [24:0] p1_sum__1046_comb;
  wire [24:0] p1_sum__1039_comb;
  wire [24:0] p1_sum__1032_comb;
  wire [24:0] p1_sum__1025_comb;
  wire [24:0] p1_sum__1073_comb;
  wire [24:0] p1_sum__1066_comb;
  wire [24:0] p1_sum__1059_comb;
  wire [24:0] p1_sum__1052_comb;
  wire [24:0] p1_sum__1045_comb;
  wire [24:0] p1_sum__1038_comb;
  wire [24:0] p1_sum__1031_comb;
  wire [24:0] p1_sum__1024_comb;
  wire [24:0] p1_add_144473_comb;
  wire [24:0] p1_add_144474_comb;
  wire [24:0] p1_add_144475_comb;
  wire [24:0] p1_add_144476_comb;
  wire [24:0] p1_add_144477_comb;
  wire [24:0] p1_add_144478_comb;
  wire [24:0] p1_add_144479_comb;
  wire [24:0] p1_add_144480_comb;
  wire [24:0] p1_add_144481_comb;
  wire [24:0] p1_add_144482_comb;
  wire [24:0] p1_add_144483_comb;
  wire [24:0] p1_add_144484_comb;
  wire [24:0] p1_add_144485_comb;
  wire [24:0] p1_add_144486_comb;
  wire [24:0] p1_add_144487_comb;
  wire [24:0] p1_add_144488_comb;
  wire [24:0] p1_add_144489_comb;
  wire [24:0] p1_add_144490_comb;
  wire [24:0] p1_add_144491_comb;
  wire [24:0] p1_add_144492_comb;
  wire [24:0] p1_add_144493_comb;
  wire [24:0] p1_add_144494_comb;
  wire [24:0] p1_add_144495_comb;
  wire [24:0] p1_add_144496_comb;
  wire [24:0] p1_add_144497_comb;
  wire [24:0] p1_add_144498_comb;
  wire [24:0] p1_add_144499_comb;
  wire [24:0] p1_add_144500_comb;
  wire [24:0] p1_add_144501_comb;
  wire [24:0] p1_add_144502_comb;
  wire [24:0] p1_add_144503_comb;
  wire [24:0] p1_add_144504_comb;
  wire [24:0] p1_add_144505_comb;
  wire [24:0] p1_add_144506_comb;
  wire [24:0] p1_add_144507_comb;
  wire [24:0] p1_add_144508_comb;
  wire [24:0] p1_add_144509_comb;
  wire [24:0] p1_add_144510_comb;
  wire [24:0] p1_add_144511_comb;
  wire [24:0] p1_add_144512_comb;
  wire [24:0] p1_add_144513_comb;
  wire [24:0] p1_add_144514_comb;
  wire [24:0] p1_add_144515_comb;
  wire [24:0] p1_add_144516_comb;
  wire [24:0] p1_add_144517_comb;
  wire [24:0] p1_add_144518_comb;
  wire [24:0] p1_add_144519_comb;
  wire [24:0] p1_add_144520_comb;
  wire [24:0] p1_add_144521_comb;
  wire [24:0] p1_add_144522_comb;
  wire [24:0] p1_add_144523_comb;
  wire [24:0] p1_add_144524_comb;
  wire [24:0] p1_add_144525_comb;
  wire [24:0] p1_add_144526_comb;
  wire [24:0] p1_add_144527_comb;
  wire [24:0] p1_add_144528_comb;
  wire [24:0] p1_add_144529_comb;
  wire [24:0] p1_add_144530_comb;
  wire [24:0] p1_add_144531_comb;
  wire [24:0] p1_add_144532_comb;
  wire [24:0] p1_add_144533_comb;
  wire [24:0] p1_add_144534_comb;
  wire [24:0] p1_add_144535_comb;
  wire [24:0] p1_add_144536_comb;
  wire [8:0] p1_clipped__320_comb;
  wire [8:0] p1_clipped__321_comb;
  wire [8:0] p1_clipped__322_comb;
  wire [8:0] p1_clipped__323_comb;
  wire [8:0] p1_clipped__324_comb;
  wire [8:0] p1_clipped__325_comb;
  wire [8:0] p1_clipped__326_comb;
  wire [8:0] p1_clipped__327_comb;
  wire [8:0] p1_clipped__328_comb;
  wire [8:0] p1_clipped__329_comb;
  wire [8:0] p1_clipped__330_comb;
  wire [8:0] p1_clipped__331_comb;
  wire [8:0] p1_clipped__332_comb;
  wire [8:0] p1_clipped__333_comb;
  wire [8:0] p1_clipped__334_comb;
  wire [8:0] p1_clipped__335_comb;
  wire [8:0] p1_clipped__336_comb;
  wire [8:0] p1_clipped__337_comb;
  wire [8:0] p1_clipped__338_comb;
  wire [8:0] p1_clipped__339_comb;
  wire [8:0] p1_clipped__340_comb;
  wire [8:0] p1_clipped__341_comb;
  wire [8:0] p1_clipped__342_comb;
  wire [8:0] p1_clipped__343_comb;
  wire [8:0] p1_clipped__344_comb;
  wire [8:0] p1_clipped__345_comb;
  wire [8:0] p1_clipped__346_comb;
  wire [8:0] p1_clipped__347_comb;
  wire [8:0] p1_clipped__348_comb;
  wire [8:0] p1_clipped__349_comb;
  wire [8:0] p1_clipped__350_comb;
  wire [8:0] p1_clipped__351_comb;
  wire [8:0] p1_clipped__352_comb;
  wire [8:0] p1_clipped__353_comb;
  wire [8:0] p1_clipped__354_comb;
  wire [8:0] p1_clipped__355_comb;
  wire [8:0] p1_clipped__356_comb;
  wire [8:0] p1_clipped__357_comb;
  wire [8:0] p1_clipped__358_comb;
  wire [8:0] p1_clipped__359_comb;
  wire [8:0] p1_clipped__360_comb;
  wire [8:0] p1_clipped__361_comb;
  wire [8:0] p1_clipped__362_comb;
  wire [8:0] p1_clipped__363_comb;
  wire [8:0] p1_clipped__364_comb;
  wire [8:0] p1_clipped__365_comb;
  wire [8:0] p1_clipped__366_comb;
  wire [8:0] p1_clipped__367_comb;
  wire [8:0] p1_clipped__368_comb;
  wire [8:0] p1_clipped__369_comb;
  wire [8:0] p1_clipped__370_comb;
  wire [8:0] p1_clipped__371_comb;
  wire [8:0] p1_clipped__372_comb;
  wire [8:0] p1_clipped__373_comb;
  wire [8:0] p1_clipped__374_comb;
  wire [8:0] p1_clipped__375_comb;
  wire [8:0] p1_clipped__376_comb;
  wire [8:0] p1_clipped__377_comb;
  wire [8:0] p1_clipped__378_comb;
  wire [8:0] p1_clipped__379_comb;
  wire [8:0] p1_clipped__380_comb;
  wire [8:0] p1_clipped__381_comb;
  wire [8:0] p1_clipped__382_comb;
  wire [8:0] p1_clipped__383_comb;
  wire [9:0] p1_add_145305_comb;
  wire [9:0] p1_add_145306_comb;
  wire [9:0] p1_add_145307_comb;
  wire [9:0] p1_add_145308_comb;
  wire [9:0] p1_add_145309_comb;
  wire [9:0] p1_add_145310_comb;
  wire [9:0] p1_add_145311_comb;
  wire [9:0] p1_add_145312_comb;
  wire [9:0] p1_add_145313_comb;
  wire [9:0] p1_add_145314_comb;
  wire [9:0] p1_add_145315_comb;
  wire [9:0] p1_add_145316_comb;
  wire [9:0] p1_add_145317_comb;
  wire [9:0] p1_add_145318_comb;
  wire [9:0] p1_add_145319_comb;
  wire [9:0] p1_add_145320_comb;
  wire [9:0] p1_add_145321_comb;
  wire [9:0] p1_add_145322_comb;
  wire [9:0] p1_add_145323_comb;
  wire [9:0] p1_add_145324_comb;
  wire [9:0] p1_add_145325_comb;
  wire [9:0] p1_add_145326_comb;
  wire [9:0] p1_add_145327_comb;
  wire [9:0] p1_add_145328_comb;
  wire [9:0] p1_add_145329_comb;
  wire [9:0] p1_add_145330_comb;
  wire [9:0] p1_add_145331_comb;
  wire [9:0] p1_add_145332_comb;
  wire [9:0] p1_add_145333_comb;
  wire [9:0] p1_add_145334_comb;
  wire [9:0] p1_add_145335_comb;
  wire [9:0] p1_add_145336_comb;
  wire [9:0] p1_add_145337_comb;
  wire [9:0] p1_add_145338_comb;
  wire [9:0] p1_add_145339_comb;
  wire [9:0] p1_add_145340_comb;
  wire [9:0] p1_add_145341_comb;
  wire [9:0] p1_add_145342_comb;
  wire [9:0] p1_add_145343_comb;
  wire [9:0] p1_add_145344_comb;
  wire [9:0] p1_add_145345_comb;
  wire [9:0] p1_add_145346_comb;
  wire [9:0] p1_add_145347_comb;
  wire [9:0] p1_add_145348_comb;
  wire [9:0] p1_add_145349_comb;
  wire [9:0] p1_add_145350_comb;
  wire [9:0] p1_add_145351_comb;
  wire [9:0] p1_add_145352_comb;
  wire [9:0] p1_add_145353_comb;
  wire [9:0] p1_add_145354_comb;
  wire [9:0] p1_add_145355_comb;
  wire [9:0] p1_add_145356_comb;
  wire [9:0] p1_add_145357_comb;
  wire [9:0] p1_add_145358_comb;
  wire [9:0] p1_add_145359_comb;
  wire [9:0] p1_add_145360_comb;
  wire [9:0] p1_add_145361_comb;
  wire [9:0] p1_add_145362_comb;
  wire [9:0] p1_add_145363_comb;
  wire [9:0] p1_add_145364_comb;
  wire [9:0] p1_add_145365_comb;
  wire [9:0] p1_add_145366_comb;
  wire [9:0] p1_add_145367_comb;
  wire [9:0] p1_add_145368_comb;
  wire [1:0] p1_bit_slice_145369_comb;
  wire [1:0] p1_bit_slice_145370_comb;
  wire [1:0] p1_bit_slice_145371_comb;
  wire [1:0] p1_bit_slice_145372_comb;
  wire [1:0] p1_bit_slice_145373_comb;
  wire [1:0] p1_bit_slice_145374_comb;
  wire [1:0] p1_bit_slice_145375_comb;
  wire [1:0] p1_bit_slice_145376_comb;
  wire [1:0] p1_bit_slice_145377_comb;
  wire [1:0] p1_bit_slice_145378_comb;
  wire [1:0] p1_bit_slice_145379_comb;
  wire [1:0] p1_bit_slice_145380_comb;
  wire [1:0] p1_bit_slice_145381_comb;
  wire [1:0] p1_bit_slice_145382_comb;
  wire [1:0] p1_bit_slice_145383_comb;
  wire [1:0] p1_bit_slice_145384_comb;
  wire [1:0] p1_bit_slice_145385_comb;
  wire [1:0] p1_bit_slice_145386_comb;
  wire [1:0] p1_bit_slice_145387_comb;
  wire [1:0] p1_bit_slice_145388_comb;
  wire [1:0] p1_bit_slice_145389_comb;
  wire [1:0] p1_bit_slice_145390_comb;
  wire [1:0] p1_bit_slice_145391_comb;
  wire [1:0] p1_bit_slice_145392_comb;
  wire [1:0] p1_bit_slice_145393_comb;
  wire [1:0] p1_bit_slice_145394_comb;
  wire [1:0] p1_bit_slice_145395_comb;
  wire [1:0] p1_bit_slice_145396_comb;
  wire [1:0] p1_bit_slice_145397_comb;
  wire [1:0] p1_bit_slice_145398_comb;
  wire [1:0] p1_bit_slice_145399_comb;
  wire [1:0] p1_bit_slice_145400_comb;
  wire [1:0] p1_bit_slice_145401_comb;
  wire [1:0] p1_bit_slice_145402_comb;
  wire [1:0] p1_bit_slice_145403_comb;
  wire [1:0] p1_bit_slice_145404_comb;
  wire [1:0] p1_bit_slice_145405_comb;
  wire [1:0] p1_bit_slice_145406_comb;
  wire [1:0] p1_bit_slice_145407_comb;
  wire [1:0] p1_bit_slice_145408_comb;
  wire [1:0] p1_bit_slice_145409_comb;
  wire [1:0] p1_bit_slice_145410_comb;
  wire [1:0] p1_bit_slice_145411_comb;
  wire [1:0] p1_bit_slice_145412_comb;
  wire [1:0] p1_bit_slice_145413_comb;
  wire [1:0] p1_bit_slice_145414_comb;
  wire [1:0] p1_bit_slice_145415_comb;
  wire [1:0] p1_bit_slice_145416_comb;
  wire [1:0] p1_bit_slice_145417_comb;
  wire [1:0] p1_bit_slice_145418_comb;
  wire [1:0] p1_bit_slice_145419_comb;
  wire [1:0] p1_bit_slice_145420_comb;
  wire [1:0] p1_bit_slice_145421_comb;
  wire [1:0] p1_bit_slice_145422_comb;
  wire [1:0] p1_bit_slice_145423_comb;
  wire [1:0] p1_bit_slice_145424_comb;
  wire [1:0] p1_bit_slice_145425_comb;
  wire [1:0] p1_bit_slice_145426_comb;
  wire [1:0] p1_bit_slice_145427_comb;
  wire [1:0] p1_bit_slice_145428_comb;
  wire [1:0] p1_bit_slice_145429_comb;
  wire [1:0] p1_bit_slice_145430_comb;
  wire [1:0] p1_bit_slice_145431_comb;
  wire [1:0] p1_bit_slice_145432_comb;
  wire [2:0] p1_add_145561_comb;
  wire [2:0] p1_add_145562_comb;
  wire [2:0] p1_add_145563_comb;
  wire [2:0] p1_add_145564_comb;
  wire [2:0] p1_add_145565_comb;
  wire [2:0] p1_add_145566_comb;
  wire [2:0] p1_add_145567_comb;
  wire [2:0] p1_add_145568_comb;
  wire [2:0] p1_add_145569_comb;
  wire [2:0] p1_add_145570_comb;
  wire [2:0] p1_add_145571_comb;
  wire [2:0] p1_add_145572_comb;
  wire [2:0] p1_add_145573_comb;
  wire [2:0] p1_add_145574_comb;
  wire [2:0] p1_add_145575_comb;
  wire [2:0] p1_add_145576_comb;
  wire [2:0] p1_add_145577_comb;
  wire [2:0] p1_add_145578_comb;
  wire [2:0] p1_add_145579_comb;
  wire [2:0] p1_add_145580_comb;
  wire [2:0] p1_add_145581_comb;
  wire [2:0] p1_add_145582_comb;
  wire [2:0] p1_add_145583_comb;
  wire [2:0] p1_add_145584_comb;
  wire [2:0] p1_add_145585_comb;
  wire [2:0] p1_add_145586_comb;
  wire [2:0] p1_add_145587_comb;
  wire [2:0] p1_add_145588_comb;
  wire [2:0] p1_add_145589_comb;
  wire [2:0] p1_add_145590_comb;
  wire [2:0] p1_add_145591_comb;
  wire [2:0] p1_add_145592_comb;
  wire [2:0] p1_add_145593_comb;
  wire [2:0] p1_add_145594_comb;
  wire [2:0] p1_add_145595_comb;
  wire [2:0] p1_add_145596_comb;
  wire [2:0] p1_add_145597_comb;
  wire [2:0] p1_add_145598_comb;
  wire [2:0] p1_add_145599_comb;
  wire [2:0] p1_add_145600_comb;
  wire [2:0] p1_add_145601_comb;
  wire [2:0] p1_add_145602_comb;
  wire [2:0] p1_add_145603_comb;
  wire [2:0] p1_add_145604_comb;
  wire [2:0] p1_add_145605_comb;
  wire [2:0] p1_add_145606_comb;
  wire [2:0] p1_add_145607_comb;
  wire [2:0] p1_add_145608_comb;
  wire [2:0] p1_add_145609_comb;
  wire [2:0] p1_add_145610_comb;
  wire [2:0] p1_add_145611_comb;
  wire [2:0] p1_add_145612_comb;
  wire [2:0] p1_add_145613_comb;
  wire [2:0] p1_add_145614_comb;
  wire [2:0] p1_add_145615_comb;
  wire [2:0] p1_add_145616_comb;
  wire [2:0] p1_add_145617_comb;
  wire [2:0] p1_add_145618_comb;
  wire [2:0] p1_add_145619_comb;
  wire [2:0] p1_add_145620_comb;
  wire [2:0] p1_add_145621_comb;
  wire [2:0] p1_add_145622_comb;
  wire [2:0] p1_add_145623_comb;
  wire [2:0] p1_add_145624_comb;
  wire [7:0] p1_clipped__136_comb;
  wire [7:0] p1_clipped__152_comb;
  wire [7:0] p1_clipped__168_comb;
  wire [7:0] p1_clipped__184_comb;
  wire [7:0] p1_clipped__200_comb;
  wire [7:0] p1_clipped__216_comb;
  wire [7:0] p1_clipped__232_comb;
  wire [7:0] p1_clipped__248_comb;
  wire [7:0] p1_clipped__137_comb;
  wire [7:0] p1_clipped__153_comb;
  wire [7:0] p1_clipped__169_comb;
  wire [7:0] p1_clipped__185_comb;
  wire [7:0] p1_clipped__201_comb;
  wire [7:0] p1_clipped__217_comb;
  wire [7:0] p1_clipped__233_comb;
  wire [7:0] p1_clipped__249_comb;
  wire [7:0] p1_clipped__138_comb;
  wire [7:0] p1_clipped__154_comb;
  wire [7:0] p1_clipped__170_comb;
  wire [7:0] p1_clipped__186_comb;
  wire [7:0] p1_clipped__202_comb;
  wire [7:0] p1_clipped__218_comb;
  wire [7:0] p1_clipped__234_comb;
  wire [7:0] p1_clipped__250_comb;
  wire [7:0] p1_clipped__139_comb;
  wire [7:0] p1_clipped__155_comb;
  wire [7:0] p1_clipped__171_comb;
  wire [7:0] p1_clipped__187_comb;
  wire [7:0] p1_clipped__203_comb;
  wire [7:0] p1_clipped__219_comb;
  wire [7:0] p1_clipped__235_comb;
  wire [7:0] p1_clipped__251_comb;
  wire [7:0] p1_clipped__140_comb;
  wire [7:0] p1_clipped__156_comb;
  wire [7:0] p1_clipped__172_comb;
  wire [7:0] p1_clipped__188_comb;
  wire [7:0] p1_clipped__204_comb;
  wire [7:0] p1_clipped__220_comb;
  wire [7:0] p1_clipped__236_comb;
  wire [7:0] p1_clipped__252_comb;
  wire [7:0] p1_clipped__141_comb;
  wire [7:0] p1_clipped__157_comb;
  wire [7:0] p1_clipped__173_comb;
  wire [7:0] p1_clipped__189_comb;
  wire [7:0] p1_clipped__205_comb;
  wire [7:0] p1_clipped__221_comb;
  wire [7:0] p1_clipped__237_comb;
  wire [7:0] p1_clipped__253_comb;
  wire [7:0] p1_clipped__142_comb;
  wire [7:0] p1_clipped__158_comb;
  wire [7:0] p1_clipped__174_comb;
  wire [7:0] p1_clipped__190_comb;
  wire [7:0] p1_clipped__206_comb;
  wire [7:0] p1_clipped__222_comb;
  wire [7:0] p1_clipped__238_comb;
  wire [7:0] p1_clipped__254_comb;
  wire [7:0] p1_clipped__143_comb;
  wire [7:0] p1_clipped__159_comb;
  wire [7:0] p1_clipped__175_comb;
  wire [7:0] p1_clipped__191_comb;
  wire [7:0] p1_clipped__207_comb;
  wire [7:0] p1_clipped__223_comb;
  wire [7:0] p1_clipped__239_comb;
  wire [7:0] p1_clipped__255_comb;
  wire [7:0] p1_array_146009_comb[0:7];
  wire [7:0] p1_array_146010_comb[0:7];
  wire [7:0] p1_array_146011_comb[0:7];
  wire [7:0] p1_array_146012_comb[0:7];
  wire [7:0] p1_array_146013_comb[0:7];
  wire [7:0] p1_array_146014_comb[0:7];
  wire [7:0] p1_array_146015_comb[0:7];
  wire [7:0] p1_array_146016_comb[0:7];
  wire [7:0] p1_col_transformed_comb[0:7][0:7];
  assign p1_array_index_130665_comb = p0_x[3'h2][3'h2];
  assign p1_array_index_130666_comb = p0_x[3'h2][3'h3];
  assign p1_array_index_130667_comb = p0_x[3'h2][3'h4];
  assign p1_array_index_130668_comb = p0_x[3'h2][3'h5];
  assign p1_array_index_130669_comb = p0_x[3'h3][3'h2];
  assign p1_array_index_130670_comb = p0_x[3'h3][3'h3];
  assign p1_array_index_130671_comb = p0_x[3'h3][3'h4];
  assign p1_array_index_130672_comb = p0_x[3'h3][3'h5];
  assign p1_array_index_130673_comb = p0_x[3'h4][3'h2];
  assign p1_array_index_130674_comb = p0_x[3'h4][3'h3];
  assign p1_array_index_130675_comb = p0_x[3'h4][3'h4];
  assign p1_array_index_130676_comb = p0_x[3'h4][3'h5];
  assign p1_array_index_130677_comb = p0_x[3'h5][3'h2];
  assign p1_array_index_130678_comb = p0_x[3'h5][3'h3];
  assign p1_array_index_130679_comb = p0_x[3'h5][3'h4];
  assign p1_array_index_130680_comb = p0_x[3'h5][3'h5];
  assign p1_array_index_130681_comb = p0_x[3'h2][3'h0];
  assign p1_array_index_130682_comb = p0_x[3'h2][3'h7];
  assign p1_array_index_130683_comb = p0_x[3'h3][3'h0];
  assign p1_array_index_130684_comb = p0_x[3'h3][3'h7];
  assign p1_array_index_130685_comb = p0_x[3'h4][3'h0];
  assign p1_array_index_130686_comb = p0_x[3'h4][3'h7];
  assign p1_array_index_130687_comb = p0_x[3'h5][3'h0];
  assign p1_array_index_130688_comb = p0_x[3'h5][3'h7];
  assign p1_array_index_130689_comb = p0_x[3'h2][3'h1];
  assign p1_array_index_130690_comb = p0_x[3'h2][3'h6];
  assign p1_array_index_130691_comb = p0_x[3'h3][3'h1];
  assign p1_array_index_130692_comb = p0_x[3'h3][3'h6];
  assign p1_array_index_130693_comb = p0_x[3'h4][3'h1];
  assign p1_array_index_130694_comb = p0_x[3'h4][3'h6];
  assign p1_array_index_130695_comb = p0_x[3'h5][3'h1];
  assign p1_array_index_130696_comb = p0_x[3'h5][3'h6];
  assign p1_array_index_130697_comb = p0_x[3'h0][3'h2];
  assign p1_array_index_130698_comb = p0_x[3'h0][3'h3];
  assign p1_array_index_130699_comb = p0_x[3'h0][3'h4];
  assign p1_array_index_130700_comb = p0_x[3'h0][3'h5];
  assign p1_array_index_130701_comb = p0_x[3'h7][3'h2];
  assign p1_array_index_130702_comb = p0_x[3'h7][3'h3];
  assign p1_array_index_130703_comb = p0_x[3'h7][3'h4];
  assign p1_array_index_130704_comb = p0_x[3'h7][3'h5];
  assign p1_array_index_130705_comb = p0_x[3'h0][3'h0];
  assign p1_array_index_130706_comb = p0_x[3'h0][3'h7];
  assign p1_array_index_130707_comb = p0_x[3'h7][3'h0];
  assign p1_array_index_130708_comb = p0_x[3'h7][3'h7];
  assign p1_array_index_130709_comb = p0_x[3'h0][3'h1];
  assign p1_array_index_130710_comb = p0_x[3'h0][3'h6];
  assign p1_array_index_130711_comb = p0_x[3'h7][3'h1];
  assign p1_array_index_130712_comb = p0_x[3'h7][3'h6];
  assign p1_array_index_130713_comb = p0_x[3'h1][3'h2];
  assign p1_array_index_130714_comb = p0_x[3'h1][3'h3];
  assign p1_array_index_130715_comb = p0_x[3'h1][3'h4];
  assign p1_array_index_130716_comb = p0_x[3'h1][3'h5];
  assign p1_array_index_130717_comb = p0_x[3'h6][3'h2];
  assign p1_array_index_130718_comb = p0_x[3'h6][3'h3];
  assign p1_array_index_130719_comb = p0_x[3'h6][3'h4];
  assign p1_array_index_130720_comb = p0_x[3'h6][3'h5];
  assign p1_array_index_130721_comb = p0_x[3'h1][3'h0];
  assign p1_array_index_130722_comb = p0_x[3'h1][3'h7];
  assign p1_array_index_130723_comb = p0_x[3'h6][3'h0];
  assign p1_array_index_130724_comb = p0_x[3'h6][3'h7];
  assign p1_array_index_130725_comb = p0_x[3'h1][3'h1];
  assign p1_array_index_130726_comb = p0_x[3'h1][3'h6];
  assign p1_array_index_130727_comb = p0_x[3'h6][3'h1];
  assign p1_array_index_130728_comb = p0_x[3'h6][3'h6];
  assign p1_shifted__18_squeezed_comb = {~p1_array_index_130665_comb[7], p1_array_index_130665_comb[6:0]};
  assign p1_shifted__19_squeezed_comb = {~p1_array_index_130666_comb[7], p1_array_index_130666_comb[6:0]};
  assign p1_shifted__20_squeezed_comb = {~p1_array_index_130667_comb[7], p1_array_index_130667_comb[6:0]};
  assign p1_shifted__21_squeezed_comb = {~p1_array_index_130668_comb[7], p1_array_index_130668_comb[6:0]};
  assign p1_shifted__26_squeezed_comb = {~p1_array_index_130669_comb[7], p1_array_index_130669_comb[6:0]};
  assign p1_shifted__27_squeezed_comb = {~p1_array_index_130670_comb[7], p1_array_index_130670_comb[6:0]};
  assign p1_shifted__28_squeezed_comb = {~p1_array_index_130671_comb[7], p1_array_index_130671_comb[6:0]};
  assign p1_shifted__29_squeezed_comb = {~p1_array_index_130672_comb[7], p1_array_index_130672_comb[6:0]};
  assign p1_shifted__34_squeezed_comb = {~p1_array_index_130673_comb[7], p1_array_index_130673_comb[6:0]};
  assign p1_shifted__35_squeezed_comb = {~p1_array_index_130674_comb[7], p1_array_index_130674_comb[6:0]};
  assign p1_shifted__36_squeezed_comb = {~p1_array_index_130675_comb[7], p1_array_index_130675_comb[6:0]};
  assign p1_shifted__37_squeezed_comb = {~p1_array_index_130676_comb[7], p1_array_index_130676_comb[6:0]};
  assign p1_shifted__42_squeezed_comb = {~p1_array_index_130677_comb[7], p1_array_index_130677_comb[6:0]};
  assign p1_shifted__43_squeezed_comb = {~p1_array_index_130678_comb[7], p1_array_index_130678_comb[6:0]};
  assign p1_shifted__44_squeezed_comb = {~p1_array_index_130679_comb[7], p1_array_index_130679_comb[6:0]};
  assign p1_shifted__45_squeezed_comb = {~p1_array_index_130680_comb[7], p1_array_index_130680_comb[6:0]};
  assign p1_shifted__16_squeezed_comb = {~p1_array_index_130681_comb[7], p1_array_index_130681_comb[6:0]};
  assign p1_shifted__23_squeezed_comb = {~p1_array_index_130682_comb[7], p1_array_index_130682_comb[6:0]};
  assign p1_shifted__24_squeezed_comb = {~p1_array_index_130683_comb[7], p1_array_index_130683_comb[6:0]};
  assign p1_shifted__31_squeezed_comb = {~p1_array_index_130684_comb[7], p1_array_index_130684_comb[6:0]};
  assign p1_shifted__32_squeezed_comb = {~p1_array_index_130685_comb[7], p1_array_index_130685_comb[6:0]};
  assign p1_shifted__39_squeezed_comb = {~p1_array_index_130686_comb[7], p1_array_index_130686_comb[6:0]};
  assign p1_shifted__40_squeezed_comb = {~p1_array_index_130687_comb[7], p1_array_index_130687_comb[6:0]};
  assign p1_shifted__47_squeezed_comb = {~p1_array_index_130688_comb[7], p1_array_index_130688_comb[6:0]};
  assign p1_shifted__17_squeezed_comb = {~p1_array_index_130689_comb[7], p1_array_index_130689_comb[6:0]};
  assign p1_shifted__22_squeezed_comb = {~p1_array_index_130690_comb[7], p1_array_index_130690_comb[6:0]};
  assign p1_shifted__25_squeezed_comb = {~p1_array_index_130691_comb[7], p1_array_index_130691_comb[6:0]};
  assign p1_shifted__30_squeezed_comb = {~p1_array_index_130692_comb[7], p1_array_index_130692_comb[6:0]};
  assign p1_shifted__33_squeezed_comb = {~p1_array_index_130693_comb[7], p1_array_index_130693_comb[6:0]};
  assign p1_shifted__38_squeezed_comb = {~p1_array_index_130694_comb[7], p1_array_index_130694_comb[6:0]};
  assign p1_shifted__41_squeezed_comb = {~p1_array_index_130695_comb[7], p1_array_index_130695_comb[6:0]};
  assign p1_shifted__46_squeezed_comb = {~p1_array_index_130696_comb[7], p1_array_index_130696_comb[6:0]};
  assign p1_shifted__2_squeezed_comb = {~p1_array_index_130697_comb[7], p1_array_index_130697_comb[6:0]};
  assign p1_shifted__3_squeezed_comb = {~p1_array_index_130698_comb[7], p1_array_index_130698_comb[6:0]};
  assign p1_shifted__4_squeezed_comb = {~p1_array_index_130699_comb[7], p1_array_index_130699_comb[6:0]};
  assign p1_shifted__5_squeezed_comb = {~p1_array_index_130700_comb[7], p1_array_index_130700_comb[6:0]};
  assign p1_shifted__58_squeezed_comb = {~p1_array_index_130701_comb[7], p1_array_index_130701_comb[6:0]};
  assign p1_shifted__59_squeezed_comb = {~p1_array_index_130702_comb[7], p1_array_index_130702_comb[6:0]};
  assign p1_shifted__60_squeezed_comb = {~p1_array_index_130703_comb[7], p1_array_index_130703_comb[6:0]};
  assign p1_shifted__61_squeezed_comb = {~p1_array_index_130704_comb[7], p1_array_index_130704_comb[6:0]};
  assign p1_shifted_squeezed_comb = {~p1_array_index_130705_comb[7], p1_array_index_130705_comb[6:0]};
  assign p1_shifted__7_squeezed_comb = {~p1_array_index_130706_comb[7], p1_array_index_130706_comb[6:0]};
  assign p1_shifted__56_squeezed_comb = {~p1_array_index_130707_comb[7], p1_array_index_130707_comb[6:0]};
  assign p1_shifted__63_squeezed_comb = {~p1_array_index_130708_comb[7], p1_array_index_130708_comb[6:0]};
  assign p1_shifted__1_squeezed_comb = {~p1_array_index_130709_comb[7], p1_array_index_130709_comb[6:0]};
  assign p1_shifted__6_squeezed_comb = {~p1_array_index_130710_comb[7], p1_array_index_130710_comb[6:0]};
  assign p1_shifted__57_squeezed_comb = {~p1_array_index_130711_comb[7], p1_array_index_130711_comb[6:0]};
  assign p1_shifted__62_squeezed_comb = {~p1_array_index_130712_comb[7], p1_array_index_130712_comb[6:0]};
  assign p1_shifted__10_squeezed_comb = {~p1_array_index_130713_comb[7], p1_array_index_130713_comb[6:0]};
  assign p1_shifted__11_squeezed_comb = {~p1_array_index_130714_comb[7], p1_array_index_130714_comb[6:0]};
  assign p1_shifted__12_squeezed_comb = {~p1_array_index_130715_comb[7], p1_array_index_130715_comb[6:0]};
  assign p1_shifted__13_squeezed_comb = {~p1_array_index_130716_comb[7], p1_array_index_130716_comb[6:0]};
  assign p1_shifted__50_squeezed_comb = {~p1_array_index_130717_comb[7], p1_array_index_130717_comb[6:0]};
  assign p1_shifted__51_squeezed_comb = {~p1_array_index_130718_comb[7], p1_array_index_130718_comb[6:0]};
  assign p1_shifted__52_squeezed_comb = {~p1_array_index_130719_comb[7], p1_array_index_130719_comb[6:0]};
  assign p1_shifted__53_squeezed_comb = {~p1_array_index_130720_comb[7], p1_array_index_130720_comb[6:0]};
  assign p1_shifted__8_squeezed_comb = {~p1_array_index_130721_comb[7], p1_array_index_130721_comb[6:0]};
  assign p1_shifted__15_squeezed_comb = {~p1_array_index_130722_comb[7], p1_array_index_130722_comb[6:0]};
  assign p1_shifted__48_squeezed_comb = {~p1_array_index_130723_comb[7], p1_array_index_130723_comb[6:0]};
  assign p1_shifted__55_squeezed_comb = {~p1_array_index_130724_comb[7], p1_array_index_130724_comb[6:0]};
  assign p1_shifted__9_squeezed_comb = {~p1_array_index_130725_comb[7], p1_array_index_130725_comb[6:0]};
  assign p1_shifted__14_squeezed_comb = {~p1_array_index_130726_comb[7], p1_array_index_130726_comb[6:0]};
  assign p1_shifted__49_squeezed_comb = {~p1_array_index_130727_comb[7], p1_array_index_130727_comb[6:0]};
  assign p1_shifted__54_squeezed_comb = {~p1_array_index_130728_comb[7], p1_array_index_130728_comb[6:0]};
  assign p1_smul_57362_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__18_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___8_comb = 9'h000;
  assign p1_smul_57364_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__19_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___9_comb = 9'h000;
  assign p1_smul_57366_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__20_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___10_comb = 9'h000;
  assign p1_smul_57368_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__21_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___11_comb = 9'h000;
  assign p1_smul_57378_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__26_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___12_comb = 9'h000;
  assign p1_smul_57380_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__27_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___13_comb = 9'h000;
  assign p1_smul_57382_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__28_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___14_comb = 9'h000;
  assign p1_smul_57384_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__29_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___15_comb = 9'h000;
  assign p1_smul_57394_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__34_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___16_comb = 9'h000;
  assign p1_smul_57396_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__35_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___17_comb = 9'h000;
  assign p1_smul_57398_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__36_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___18_comb = 9'h000;
  assign p1_smul_57400_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__37_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___19_comb = 9'h000;
  assign p1_smul_57410_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__42_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___20_comb = 9'h000;
  assign p1_smul_57412_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__43_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___21_comb = 9'h000;
  assign p1_smul_57414_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__44_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___22_comb = 9'h000;
  assign p1_smul_57416_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__45_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___23_comb = 9'h000;
  assign p1_smul_57486_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__16_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___8_comb = 10'h000;
  assign p1_smul_57492_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__19_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___9_comb = 10'h000;
  assign p1_smul_57494_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__20_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___10_comb = 10'h000;
  assign p1_smul_57500_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__23_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___11_comb = 10'h000;
  assign p1_smul_57502_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__24_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___12_comb = 10'h000;
  assign p1_smul_57508_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__27_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___13_comb = 10'h000;
  assign p1_smul_57510_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__28_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___14_comb = 10'h000;
  assign p1_smul_57516_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__31_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___15_comb = 10'h000;
  assign p1_smul_57518_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__32_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___16_comb = 10'h000;
  assign p1_smul_57524_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__35_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___17_comb = 10'h000;
  assign p1_smul_57526_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__36_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___18_comb = 10'h000;
  assign p1_smul_57532_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__39_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___19_comb = 10'h000;
  assign p1_smul_57534_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__40_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___20_comb = 10'h000;
  assign p1_smul_57540_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__43_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___21_comb = 10'h000;
  assign p1_smul_57542_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__44_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___22_comb = 10'h000;
  assign p1_smul_57548_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__47_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___23_comb = 10'h000;
  assign p1_smul_57616_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__17_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___40_comb = 9'h000;
  assign p1_smul_57620_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__19_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___41_comb = 9'h000;
  assign p1_smul_57622_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__20_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___42_comb = 9'h000;
  assign p1_smul_57626_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__22_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___43_comb = 9'h000;
  assign p1_smul_57632_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__25_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___44_comb = 9'h000;
  assign p1_smul_57636_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__27_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___45_comb = 9'h000;
  assign p1_smul_57638_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__28_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___46_comb = 9'h000;
  assign p1_smul_57642_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__30_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___47_comb = 9'h000;
  assign p1_smul_57648_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__33_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___48_comb = 9'h000;
  assign p1_smul_57652_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__35_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___49_comb = 9'h000;
  assign p1_smul_57654_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__36_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___50_comb = 9'h000;
  assign p1_smul_57658_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__38_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___51_comb = 9'h000;
  assign p1_smul_57664_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__41_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___52_comb = 9'h000;
  assign p1_smul_57668_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__43_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___53_comb = 9'h000;
  assign p1_smul_57670_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__44_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___54_comb = 9'h000;
  assign p1_smul_57674_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__46_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___55_comb = 9'h000;
  assign p1_smul_57870_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__16_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___72_comb = 9'h000;
  assign p1_smul_57874_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__18_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___73_comb = 9'h000;
  assign p1_smul_57880_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__21_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___74_comb = 9'h000;
  assign p1_smul_57884_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__23_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___75_comb = 9'h000;
  assign p1_smul_57886_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__24_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___76_comb = 9'h000;
  assign p1_smul_57890_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__26_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___77_comb = 9'h000;
  assign p1_smul_57896_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__29_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___78_comb = 9'h000;
  assign p1_smul_57900_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__31_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___79_comb = 9'h000;
  assign p1_smul_57902_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__32_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___80_comb = 9'h000;
  assign p1_smul_57906_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__34_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___81_comb = 9'h000;
  assign p1_smul_57912_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__37_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___82_comb = 9'h000;
  assign p1_smul_57916_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__39_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___83_comb = 9'h000;
  assign p1_smul_57918_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__40_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___84_comb = 9'h000;
  assign p1_smul_57922_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__42_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___85_comb = 9'h000;
  assign p1_smul_57928_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__45_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___86_comb = 9'h000;
  assign p1_smul_57932_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__47_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___87_comb = 9'h000;
  assign p1_smul_58000_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__17_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___40_comb = 10'h000;
  assign p1_smul_58004_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__19_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___41_comb = 10'h000;
  assign p1_smul_58006_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__20_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___42_comb = 10'h000;
  assign p1_smul_58010_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__22_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___43_comb = 10'h000;
  assign p1_smul_58016_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__25_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___44_comb = 10'h000;
  assign p1_smul_58020_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__27_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___45_comb = 10'h000;
  assign p1_smul_58022_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__28_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___46_comb = 10'h000;
  assign p1_smul_58026_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__30_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___47_comb = 10'h000;
  assign p1_smul_58032_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__33_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___48_comb = 10'h000;
  assign p1_smul_58036_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__35_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___49_comb = 10'h000;
  assign p1_smul_58038_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__36_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___50_comb = 10'h000;
  assign p1_smul_58042_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__38_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___51_comb = 10'h000;
  assign p1_smul_58048_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__41_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___52_comb = 10'h000;
  assign p1_smul_58052_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__43_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___53_comb = 10'h000;
  assign p1_smul_58054_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__44_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___54_comb = 10'h000;
  assign p1_smul_58058_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__46_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___55_comb = 10'h000;
  assign p1_smul_58126_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__16_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___104_comb = 9'h000;
  assign p1_smul_58128_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__17_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___105_comb = 9'h000;
  assign p1_smul_58138_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__22_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___106_comb = 9'h000;
  assign p1_smul_58140_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__23_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___107_comb = 9'h000;
  assign p1_smul_58142_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__24_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___108_comb = 9'h000;
  assign p1_smul_58144_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__25_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___109_comb = 9'h000;
  assign p1_smul_58154_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__30_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___110_comb = 9'h000;
  assign p1_smul_58156_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__31_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___111_comb = 9'h000;
  assign p1_smul_58158_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__32_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___112_comb = 9'h000;
  assign p1_smul_58160_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__33_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___113_comb = 9'h000;
  assign p1_smul_58170_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__38_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___114_comb = 9'h000;
  assign p1_smul_58172_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__39_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___115_comb = 9'h000;
  assign p1_smul_58174_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__40_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___116_comb = 9'h000;
  assign p1_smul_58176_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__41_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___117_comb = 9'h000;
  assign p1_smul_58186_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__46_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___118_comb = 9'h000;
  assign p1_smul_58188_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__47_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___119_comb = 9'h000;
  assign p1_smul_57330_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__2_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits__comb = 9'h000;
  assign p1_smul_57332_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__3_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___1_comb = 9'h000;
  assign p1_smul_57334_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__4_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___2_comb = 9'h000;
  assign p1_smul_57336_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__5_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___3_comb = 9'h000;
  assign p1_smul_57442_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__58_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___28_comb = 9'h000;
  assign p1_smul_57444_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__59_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___29_comb = 9'h000;
  assign p1_smul_57446_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__60_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___30_comb = 9'h000;
  assign p1_smul_57448_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__61_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___31_comb = 9'h000;
  assign p1_smul_57454_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits__comb = 10'h000;
  assign p1_smul_57460_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__3_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___1_comb = 10'h000;
  assign p1_smul_57462_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__4_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___2_comb = 10'h000;
  assign p1_smul_57468_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__7_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___3_comb = 10'h000;
  assign p1_smul_57566_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__56_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___28_comb = 10'h000;
  assign p1_smul_57572_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__59_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___29_comb = 10'h000;
  assign p1_smul_57574_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__60_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___30_comb = 10'h000;
  assign p1_smul_57580_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__63_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___31_comb = 10'h000;
  assign p1_smul_57584_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__1_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___32_comb = 9'h000;
  assign p1_smul_57588_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__3_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___33_comb = 9'h000;
  assign p1_smul_57590_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__4_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___34_comb = 9'h000;
  assign p1_smul_57594_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__6_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___35_comb = 9'h000;
  assign p1_smul_57696_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__57_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___60_comb = 9'h000;
  assign p1_smul_57700_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__59_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___61_comb = 9'h000;
  assign p1_smul_57702_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__60_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___62_comb = 9'h000;
  assign p1_smul_57706_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__62_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___63_comb = 9'h000;
  assign p1_smul_57838_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___64_comb = 9'h000;
  assign p1_smul_57842_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__2_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___65_comb = 9'h000;
  assign p1_smul_57848_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__5_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___66_comb = 9'h000;
  assign p1_smul_57852_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__7_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___67_comb = 9'h000;
  assign p1_smul_57950_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__56_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___92_comb = 9'h000;
  assign p1_smul_57954_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__58_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___93_comb = 9'h000;
  assign p1_smul_57960_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__61_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___94_comb = 9'h000;
  assign p1_smul_57964_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__63_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___95_comb = 9'h000;
  assign p1_smul_57968_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__1_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___32_comb = 10'h000;
  assign p1_smul_57972_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__3_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___33_comb = 10'h000;
  assign p1_smul_57974_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__4_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___34_comb = 10'h000;
  assign p1_smul_57978_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__6_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___35_comb = 10'h000;
  assign p1_smul_58080_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__57_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___60_comb = 10'h000;
  assign p1_smul_58084_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__59_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___61_comb = 10'h000;
  assign p1_smul_58086_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__60_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___62_comb = 10'h000;
  assign p1_smul_58090_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__62_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___63_comb = 10'h000;
  assign p1_smul_58094_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___96_comb = 9'h000;
  assign p1_smul_58096_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__1_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___97_comb = 9'h000;
  assign p1_smul_58106_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__6_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___98_comb = 9'h000;
  assign p1_smul_58108_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__7_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___99_comb = 9'h000;
  assign p1_smul_58206_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__56_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___124_comb = 9'h000;
  assign p1_smul_58208_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__57_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___125_comb = 9'h000;
  assign p1_smul_58218_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__62_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___126_comb = 9'h000;
  assign p1_smul_58220_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__63_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___127_comb = 9'h000;
  assign p1_smul_57346_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__10_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___4_comb = 9'h000;
  assign p1_smul_57348_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__11_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___5_comb = 9'h000;
  assign p1_smul_57350_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__12_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___6_comb = 9'h000;
  assign p1_smul_57352_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__13_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___7_comb = 9'h000;
  assign p1_smul_57426_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__50_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___24_comb = 9'h000;
  assign p1_smul_57428_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__51_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___25_comb = 9'h000;
  assign p1_smul_57430_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__52_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___26_comb = 9'h000;
  assign p1_smul_57432_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__53_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___27_comb = 9'h000;
  assign p1_smul_57470_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__8_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___4_comb = 10'h000;
  assign p1_smul_57476_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__11_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___5_comb = 10'h000;
  assign p1_smul_57478_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__12_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___6_comb = 10'h000;
  assign p1_smul_57484_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__15_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___7_comb = 10'h000;
  assign p1_smul_57550_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__48_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___24_comb = 10'h000;
  assign p1_smul_57556_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__51_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___25_comb = 10'h000;
  assign p1_smul_57558_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__52_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___26_comb = 10'h000;
  assign p1_smul_57564_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__55_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___27_comb = 10'h000;
  assign p1_smul_57600_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__9_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___36_comb = 9'h000;
  assign p1_smul_57604_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__11_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___37_comb = 9'h000;
  assign p1_smul_57606_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__12_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___38_comb = 9'h000;
  assign p1_smul_57610_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__14_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___39_comb = 9'h000;
  assign p1_smul_57680_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__49_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___56_comb = 9'h000;
  assign p1_smul_57684_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__51_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___57_comb = 9'h000;
  assign p1_smul_57686_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__52_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___58_comb = 9'h000;
  assign p1_smul_57690_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__54_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___59_comb = 9'h000;
  assign p1_smul_57854_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__8_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___68_comb = 9'h000;
  assign p1_smul_57858_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__10_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___69_comb = 9'h000;
  assign p1_smul_57864_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__13_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___70_comb = 9'h000;
  assign p1_smul_57868_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__15_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___71_comb = 9'h000;
  assign p1_smul_57934_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__48_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___88_comb = 9'h000;
  assign p1_smul_57938_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__50_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___89_comb = 9'h000;
  assign p1_smul_57944_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__53_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___90_comb = 9'h000;
  assign p1_smul_57948_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__55_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___91_comb = 9'h000;
  assign p1_smul_57984_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__9_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___36_comb = 10'h000;
  assign p1_smul_57988_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__11_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___37_comb = 10'h000;
  assign p1_smul_57990_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__12_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___38_comb = 10'h000;
  assign p1_smul_57994_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__14_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___39_comb = 10'h000;
  assign p1_smul_58064_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__49_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___56_comb = 10'h000;
  assign p1_smul_58068_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__51_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___57_comb = 10'h000;
  assign p1_smul_58070_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__52_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___58_comb = 10'h000;
  assign p1_smul_58074_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__54_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___59_comb = 10'h000;
  assign p1_smul_58110_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__8_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___100_comb = 9'h000;
  assign p1_smul_58112_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__9_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___101_comb = 9'h000;
  assign p1_smul_58122_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__14_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___102_comb = 9'h000;
  assign p1_smul_58124_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__15_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___103_comb = 9'h000;
  assign p1_smul_58190_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__48_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___120_comb = 9'h000;
  assign p1_smul_58192_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__49_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___121_comb = 9'h000;
  assign p1_smul_58202_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__54_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___122_comb = 9'h000;
  assign p1_smul_58204_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__55_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___123_comb = 9'h000;
  assign p1_smul_57326_TrailingBits___144_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___145_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___146_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___147_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___148_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___149_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___150_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___151_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___152_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___153_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___154_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___155_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___156_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___157_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___158_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___159_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___160_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___161_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___162_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___163_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___164_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___165_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___166_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___167_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___168_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___169_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___170_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___171_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___172_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___173_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___174_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___175_comb = 8'h00;
  assign p1_concat_131721_comb = {p1_smul_57362_NarrowedMult__comb, p1_smul_57330_TrailingBits___8_comb};
  assign p1_concat_131722_comb = {p1_smul_57364_NarrowedMult__comb, p1_smul_57330_TrailingBits___9_comb};
  assign p1_concat_131723_comb = {p1_smul_57366_NarrowedMult__comb, p1_smul_57330_TrailingBits___10_comb};
  assign p1_concat_131724_comb = {p1_smul_57368_NarrowedMult__comb, p1_smul_57330_TrailingBits___11_comb};
  assign p1_concat_131725_comb = {p1_smul_57378_NarrowedMult__comb, p1_smul_57330_TrailingBits___12_comb};
  assign p1_concat_131726_comb = {p1_smul_57380_NarrowedMult__comb, p1_smul_57330_TrailingBits___13_comb};
  assign p1_concat_131727_comb = {p1_smul_57382_NarrowedMult__comb, p1_smul_57330_TrailingBits___14_comb};
  assign p1_concat_131728_comb = {p1_smul_57384_NarrowedMult__comb, p1_smul_57330_TrailingBits___15_comb};
  assign p1_concat_131729_comb = {p1_smul_57394_NarrowedMult__comb, p1_smul_57330_TrailingBits___16_comb};
  assign p1_concat_131730_comb = {p1_smul_57396_NarrowedMult__comb, p1_smul_57330_TrailingBits___17_comb};
  assign p1_concat_131731_comb = {p1_smul_57398_NarrowedMult__comb, p1_smul_57330_TrailingBits___18_comb};
  assign p1_concat_131732_comb = {p1_smul_57400_NarrowedMult__comb, p1_smul_57330_TrailingBits___19_comb};
  assign p1_concat_131733_comb = {p1_smul_57410_NarrowedMult__comb, p1_smul_57330_TrailingBits___20_comb};
  assign p1_concat_131734_comb = {p1_smul_57412_NarrowedMult__comb, p1_smul_57330_TrailingBits___21_comb};
  assign p1_concat_131735_comb = {p1_smul_57414_NarrowedMult__comb, p1_smul_57330_TrailingBits___22_comb};
  assign p1_concat_131736_comb = {p1_smul_57416_NarrowedMult__comb, p1_smul_57330_TrailingBits___23_comb};
  assign p1_concat_131737_comb = {p1_smul_57486_NarrowedMult__comb, p1_smul_57454_TrailingBits___8_comb};
  assign p1_concat_131738_comb = {p1_smul_57492_NarrowedMult__comb, p1_smul_57454_TrailingBits___9_comb};
  assign p1_concat_131739_comb = {p1_smul_57494_NarrowedMult__comb, p1_smul_57454_TrailingBits___10_comb};
  assign p1_concat_131740_comb = {p1_smul_57500_NarrowedMult__comb, p1_smul_57454_TrailingBits___11_comb};
  assign p1_concat_131741_comb = {p1_smul_57502_NarrowedMult__comb, p1_smul_57454_TrailingBits___12_comb};
  assign p1_concat_131742_comb = {p1_smul_57508_NarrowedMult__comb, p1_smul_57454_TrailingBits___13_comb};
  assign p1_concat_131743_comb = {p1_smul_57510_NarrowedMult__comb, p1_smul_57454_TrailingBits___14_comb};
  assign p1_concat_131744_comb = {p1_smul_57516_NarrowedMult__comb, p1_smul_57454_TrailingBits___15_comb};
  assign p1_concat_131745_comb = {p1_smul_57518_NarrowedMult__comb, p1_smul_57454_TrailingBits___16_comb};
  assign p1_concat_131746_comb = {p1_smul_57524_NarrowedMult__comb, p1_smul_57454_TrailingBits___17_comb};
  assign p1_concat_131747_comb = {p1_smul_57526_NarrowedMult__comb, p1_smul_57454_TrailingBits___18_comb};
  assign p1_concat_131748_comb = {p1_smul_57532_NarrowedMult__comb, p1_smul_57454_TrailingBits___19_comb};
  assign p1_concat_131749_comb = {p1_smul_57534_NarrowedMult__comb, p1_smul_57454_TrailingBits___20_comb};
  assign p1_concat_131750_comb = {p1_smul_57540_NarrowedMult__comb, p1_smul_57454_TrailingBits___21_comb};
  assign p1_concat_131751_comb = {p1_smul_57542_NarrowedMult__comb, p1_smul_57454_TrailingBits___22_comb};
  assign p1_concat_131752_comb = {p1_smul_57548_NarrowedMult__comb, p1_smul_57454_TrailingBits___23_comb};
  assign p1_concat_131753_comb = {p1_smul_57616_NarrowedMult__comb, p1_smul_57330_TrailingBits___40_comb};
  assign p1_concat_131754_comb = {p1_smul_57620_NarrowedMult__comb, p1_smul_57330_TrailingBits___41_comb};
  assign p1_concat_131755_comb = {p1_smul_57622_NarrowedMult__comb, p1_smul_57330_TrailingBits___42_comb};
  assign p1_concat_131756_comb = {p1_smul_57626_NarrowedMult__comb, p1_smul_57330_TrailingBits___43_comb};
  assign p1_concat_131757_comb = {p1_smul_57632_NarrowedMult__comb, p1_smul_57330_TrailingBits___44_comb};
  assign p1_concat_131758_comb = {p1_smul_57636_NarrowedMult__comb, p1_smul_57330_TrailingBits___45_comb};
  assign p1_concat_131759_comb = {p1_smul_57638_NarrowedMult__comb, p1_smul_57330_TrailingBits___46_comb};
  assign p1_concat_131760_comb = {p1_smul_57642_NarrowedMult__comb, p1_smul_57330_TrailingBits___47_comb};
  assign p1_concat_131761_comb = {p1_smul_57648_NarrowedMult__comb, p1_smul_57330_TrailingBits___48_comb};
  assign p1_concat_131762_comb = {p1_smul_57652_NarrowedMult__comb, p1_smul_57330_TrailingBits___49_comb};
  assign p1_concat_131763_comb = {p1_smul_57654_NarrowedMult__comb, p1_smul_57330_TrailingBits___50_comb};
  assign p1_concat_131764_comb = {p1_smul_57658_NarrowedMult__comb, p1_smul_57330_TrailingBits___51_comb};
  assign p1_concat_131765_comb = {p1_smul_57664_NarrowedMult__comb, p1_smul_57330_TrailingBits___52_comb};
  assign p1_concat_131766_comb = {p1_smul_57668_NarrowedMult__comb, p1_smul_57330_TrailingBits___53_comb};
  assign p1_concat_131767_comb = {p1_smul_57670_NarrowedMult__comb, p1_smul_57330_TrailingBits___54_comb};
  assign p1_concat_131768_comb = {p1_smul_57674_NarrowedMult__comb, p1_smul_57330_TrailingBits___55_comb};
  assign p1_concat_131769_comb = {p1_smul_57870_NarrowedMult__comb, p1_smul_57330_TrailingBits___72_comb};
  assign p1_concat_131770_comb = {p1_smul_57874_NarrowedMult__comb, p1_smul_57330_TrailingBits___73_comb};
  assign p1_concat_131771_comb = {p1_smul_57880_NarrowedMult__comb, p1_smul_57330_TrailingBits___74_comb};
  assign p1_concat_131772_comb = {p1_smul_57884_NarrowedMult__comb, p1_smul_57330_TrailingBits___75_comb};
  assign p1_concat_131773_comb = {p1_smul_57886_NarrowedMult__comb, p1_smul_57330_TrailingBits___76_comb};
  assign p1_concat_131774_comb = {p1_smul_57890_NarrowedMult__comb, p1_smul_57330_TrailingBits___77_comb};
  assign p1_concat_131775_comb = {p1_smul_57896_NarrowedMult__comb, p1_smul_57330_TrailingBits___78_comb};
  assign p1_concat_131776_comb = {p1_smul_57900_NarrowedMult__comb, p1_smul_57330_TrailingBits___79_comb};
  assign p1_concat_131777_comb = {p1_smul_57902_NarrowedMult__comb, p1_smul_57330_TrailingBits___80_comb};
  assign p1_concat_131778_comb = {p1_smul_57906_NarrowedMult__comb, p1_smul_57330_TrailingBits___81_comb};
  assign p1_concat_131779_comb = {p1_smul_57912_NarrowedMult__comb, p1_smul_57330_TrailingBits___82_comb};
  assign p1_concat_131780_comb = {p1_smul_57916_NarrowedMult__comb, p1_smul_57330_TrailingBits___83_comb};
  assign p1_concat_131781_comb = {p1_smul_57918_NarrowedMult__comb, p1_smul_57330_TrailingBits___84_comb};
  assign p1_concat_131782_comb = {p1_smul_57922_NarrowedMult__comb, p1_smul_57330_TrailingBits___85_comb};
  assign p1_concat_131783_comb = {p1_smul_57928_NarrowedMult__comb, p1_smul_57330_TrailingBits___86_comb};
  assign p1_concat_131784_comb = {p1_smul_57932_NarrowedMult__comb, p1_smul_57330_TrailingBits___87_comb};
  assign p1_concat_131785_comb = {p1_smul_58000_NarrowedMult__comb, p1_smul_57454_TrailingBits___40_comb};
  assign p1_concat_131786_comb = {p1_smul_58004_NarrowedMult__comb, p1_smul_57454_TrailingBits___41_comb};
  assign p1_concat_131787_comb = {p1_smul_58006_NarrowedMult__comb, p1_smul_57454_TrailingBits___42_comb};
  assign p1_concat_131788_comb = {p1_smul_58010_NarrowedMult__comb, p1_smul_57454_TrailingBits___43_comb};
  assign p1_concat_131789_comb = {p1_smul_58016_NarrowedMult__comb, p1_smul_57454_TrailingBits___44_comb};
  assign p1_concat_131790_comb = {p1_smul_58020_NarrowedMult__comb, p1_smul_57454_TrailingBits___45_comb};
  assign p1_concat_131791_comb = {p1_smul_58022_NarrowedMult__comb, p1_smul_57454_TrailingBits___46_comb};
  assign p1_concat_131792_comb = {p1_smul_58026_NarrowedMult__comb, p1_smul_57454_TrailingBits___47_comb};
  assign p1_concat_131793_comb = {p1_smul_58032_NarrowedMult__comb, p1_smul_57454_TrailingBits___48_comb};
  assign p1_concat_131794_comb = {p1_smul_58036_NarrowedMult__comb, p1_smul_57454_TrailingBits___49_comb};
  assign p1_concat_131795_comb = {p1_smul_58038_NarrowedMult__comb, p1_smul_57454_TrailingBits___50_comb};
  assign p1_concat_131796_comb = {p1_smul_58042_NarrowedMult__comb, p1_smul_57454_TrailingBits___51_comb};
  assign p1_concat_131797_comb = {p1_smul_58048_NarrowedMult__comb, p1_smul_57454_TrailingBits___52_comb};
  assign p1_concat_131798_comb = {p1_smul_58052_NarrowedMult__comb, p1_smul_57454_TrailingBits___53_comb};
  assign p1_concat_131799_comb = {p1_smul_58054_NarrowedMult__comb, p1_smul_57454_TrailingBits___54_comb};
  assign p1_concat_131800_comb = {p1_smul_58058_NarrowedMult__comb, p1_smul_57454_TrailingBits___55_comb};
  assign p1_concat_131801_comb = {p1_smul_58126_NarrowedMult__comb, p1_smul_57330_TrailingBits___104_comb};
  assign p1_concat_131802_comb = {p1_smul_58128_NarrowedMult__comb, p1_smul_57330_TrailingBits___105_comb};
  assign p1_concat_131803_comb = {p1_smul_58138_NarrowedMult__comb, p1_smul_57330_TrailingBits___106_comb};
  assign p1_concat_131804_comb = {p1_smul_58140_NarrowedMult__comb, p1_smul_57330_TrailingBits___107_comb};
  assign p1_concat_131805_comb = {p1_smul_58142_NarrowedMult__comb, p1_smul_57330_TrailingBits___108_comb};
  assign p1_concat_131806_comb = {p1_smul_58144_NarrowedMult__comb, p1_smul_57330_TrailingBits___109_comb};
  assign p1_concat_131807_comb = {p1_smul_58154_NarrowedMult__comb, p1_smul_57330_TrailingBits___110_comb};
  assign p1_concat_131808_comb = {p1_smul_58156_NarrowedMult__comb, p1_smul_57330_TrailingBits___111_comb};
  assign p1_concat_131809_comb = {p1_smul_58158_NarrowedMult__comb, p1_smul_57330_TrailingBits___112_comb};
  assign p1_concat_131810_comb = {p1_smul_58160_NarrowedMult__comb, p1_smul_57330_TrailingBits___113_comb};
  assign p1_concat_131811_comb = {p1_smul_58170_NarrowedMult__comb, p1_smul_57330_TrailingBits___114_comb};
  assign p1_concat_131812_comb = {p1_smul_58172_NarrowedMult__comb, p1_smul_57330_TrailingBits___115_comb};
  assign p1_concat_131813_comb = {p1_smul_58174_NarrowedMult__comb, p1_smul_57330_TrailingBits___116_comb};
  assign p1_concat_131814_comb = {p1_smul_58176_NarrowedMult__comb, p1_smul_57330_TrailingBits___117_comb};
  assign p1_concat_131815_comb = {p1_smul_58186_NarrowedMult__comb, p1_smul_57330_TrailingBits___118_comb};
  assign p1_concat_131816_comb = {p1_smul_58188_NarrowedMult__comb, p1_smul_57330_TrailingBits___119_comb};
  assign p1_smul_57326_TrailingBits___128_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___129_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___130_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___131_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___132_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___133_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___134_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___135_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___184_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___185_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___186_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___187_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___188_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___189_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___190_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___191_comb = 8'h00;
  assign p1_concat_131865_comb = {p1_smul_57330_NarrowedMult__comb, p1_smul_57330_TrailingBits__comb};
  assign p1_concat_131866_comb = {p1_smul_57332_NarrowedMult__comb, p1_smul_57330_TrailingBits___1_comb};
  assign p1_concat_131867_comb = {p1_smul_57334_NarrowedMult__comb, p1_smul_57330_TrailingBits___2_comb};
  assign p1_concat_131868_comb = {p1_smul_57336_NarrowedMult__comb, p1_smul_57330_TrailingBits___3_comb};
  assign p1_concat_131869_comb = {p1_smul_57442_NarrowedMult__comb, p1_smul_57330_TrailingBits___28_comb};
  assign p1_concat_131870_comb = {p1_smul_57444_NarrowedMult__comb, p1_smul_57330_TrailingBits___29_comb};
  assign p1_concat_131871_comb = {p1_smul_57446_NarrowedMult__comb, p1_smul_57330_TrailingBits___30_comb};
  assign p1_concat_131872_comb = {p1_smul_57448_NarrowedMult__comb, p1_smul_57330_TrailingBits___31_comb};
  assign p1_concat_131873_comb = {p1_smul_57454_NarrowedMult__comb, p1_smul_57454_TrailingBits__comb};
  assign p1_concat_131874_comb = {p1_smul_57460_NarrowedMult__comb, p1_smul_57454_TrailingBits___1_comb};
  assign p1_concat_131875_comb = {p1_smul_57462_NarrowedMult__comb, p1_smul_57454_TrailingBits___2_comb};
  assign p1_concat_131876_comb = {p1_smul_57468_NarrowedMult__comb, p1_smul_57454_TrailingBits___3_comb};
  assign p1_concat_131877_comb = {p1_smul_57566_NarrowedMult__comb, p1_smul_57454_TrailingBits___28_comb};
  assign p1_concat_131878_comb = {p1_smul_57572_NarrowedMult__comb, p1_smul_57454_TrailingBits___29_comb};
  assign p1_concat_131879_comb = {p1_smul_57574_NarrowedMult__comb, p1_smul_57454_TrailingBits___30_comb};
  assign p1_concat_131880_comb = {p1_smul_57580_NarrowedMult__comb, p1_smul_57454_TrailingBits___31_comb};
  assign p1_concat_131881_comb = {p1_smul_57584_NarrowedMult__comb, p1_smul_57330_TrailingBits___32_comb};
  assign p1_concat_131882_comb = {p1_smul_57588_NarrowedMult__comb, p1_smul_57330_TrailingBits___33_comb};
  assign p1_concat_131883_comb = {p1_smul_57590_NarrowedMult__comb, p1_smul_57330_TrailingBits___34_comb};
  assign p1_concat_131884_comb = {p1_smul_57594_NarrowedMult__comb, p1_smul_57330_TrailingBits___35_comb};
  assign p1_concat_131885_comb = {p1_smul_57696_NarrowedMult__comb, p1_smul_57330_TrailingBits___60_comb};
  assign p1_concat_131886_comb = {p1_smul_57700_NarrowedMult__comb, p1_smul_57330_TrailingBits___61_comb};
  assign p1_concat_131887_comb = {p1_smul_57702_NarrowedMult__comb, p1_smul_57330_TrailingBits___62_comb};
  assign p1_concat_131888_comb = {p1_smul_57706_NarrowedMult__comb, p1_smul_57330_TrailingBits___63_comb};
  assign p1_concat_131889_comb = {p1_smul_57838_NarrowedMult__comb, p1_smul_57330_TrailingBits___64_comb};
  assign p1_concat_131890_comb = {p1_smul_57842_NarrowedMult__comb, p1_smul_57330_TrailingBits___65_comb};
  assign p1_concat_131891_comb = {p1_smul_57848_NarrowedMult__comb, p1_smul_57330_TrailingBits___66_comb};
  assign p1_concat_131892_comb = {p1_smul_57852_NarrowedMult__comb, p1_smul_57330_TrailingBits___67_comb};
  assign p1_concat_131893_comb = {p1_smul_57950_NarrowedMult__comb, p1_smul_57330_TrailingBits___92_comb};
  assign p1_concat_131894_comb = {p1_smul_57954_NarrowedMult__comb, p1_smul_57330_TrailingBits___93_comb};
  assign p1_concat_131895_comb = {p1_smul_57960_NarrowedMult__comb, p1_smul_57330_TrailingBits___94_comb};
  assign p1_concat_131896_comb = {p1_smul_57964_NarrowedMult__comb, p1_smul_57330_TrailingBits___95_comb};
  assign p1_concat_131897_comb = {p1_smul_57968_NarrowedMult__comb, p1_smul_57454_TrailingBits___32_comb};
  assign p1_concat_131898_comb = {p1_smul_57972_NarrowedMult__comb, p1_smul_57454_TrailingBits___33_comb};
  assign p1_concat_131899_comb = {p1_smul_57974_NarrowedMult__comb, p1_smul_57454_TrailingBits___34_comb};
  assign p1_concat_131900_comb = {p1_smul_57978_NarrowedMult__comb, p1_smul_57454_TrailingBits___35_comb};
  assign p1_concat_131901_comb = {p1_smul_58080_NarrowedMult__comb, p1_smul_57454_TrailingBits___60_comb};
  assign p1_concat_131902_comb = {p1_smul_58084_NarrowedMult__comb, p1_smul_57454_TrailingBits___61_comb};
  assign p1_concat_131903_comb = {p1_smul_58086_NarrowedMult__comb, p1_smul_57454_TrailingBits___62_comb};
  assign p1_concat_131904_comb = {p1_smul_58090_NarrowedMult__comb, p1_smul_57454_TrailingBits___63_comb};
  assign p1_concat_131905_comb = {p1_smul_58094_NarrowedMult__comb, p1_smul_57330_TrailingBits___96_comb};
  assign p1_concat_131906_comb = {p1_smul_58096_NarrowedMult__comb, p1_smul_57330_TrailingBits___97_comb};
  assign p1_concat_131907_comb = {p1_smul_58106_NarrowedMult__comb, p1_smul_57330_TrailingBits___98_comb};
  assign p1_concat_131908_comb = {p1_smul_58108_NarrowedMult__comb, p1_smul_57330_TrailingBits___99_comb};
  assign p1_concat_131909_comb = {p1_smul_58206_NarrowedMult__comb, p1_smul_57330_TrailingBits___124_comb};
  assign p1_concat_131910_comb = {p1_smul_58208_NarrowedMult__comb, p1_smul_57330_TrailingBits___125_comb};
  assign p1_concat_131911_comb = {p1_smul_58218_NarrowedMult__comb, p1_smul_57330_TrailingBits___126_comb};
  assign p1_concat_131912_comb = {p1_smul_58220_NarrowedMult__comb, p1_smul_57330_TrailingBits___127_comb};
  assign p1_smul_57326_TrailingBits___136_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___137_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___138_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___139_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___140_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___141_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___142_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___143_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___176_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___177_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___178_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___179_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___180_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___181_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___182_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___183_comb = 8'h00;
  assign p1_concat_131961_comb = {p1_smul_57346_NarrowedMult__comb, p1_smul_57330_TrailingBits___4_comb};
  assign p1_concat_131962_comb = {p1_smul_57348_NarrowedMult__comb, p1_smul_57330_TrailingBits___5_comb};
  assign p1_concat_131963_comb = {p1_smul_57350_NarrowedMult__comb, p1_smul_57330_TrailingBits___6_comb};
  assign p1_concat_131964_comb = {p1_smul_57352_NarrowedMult__comb, p1_smul_57330_TrailingBits___7_comb};
  assign p1_concat_131965_comb = {p1_smul_57426_NarrowedMult__comb, p1_smul_57330_TrailingBits___24_comb};
  assign p1_concat_131966_comb = {p1_smul_57428_NarrowedMult__comb, p1_smul_57330_TrailingBits___25_comb};
  assign p1_concat_131967_comb = {p1_smul_57430_NarrowedMult__comb, p1_smul_57330_TrailingBits___26_comb};
  assign p1_concat_131968_comb = {p1_smul_57432_NarrowedMult__comb, p1_smul_57330_TrailingBits___27_comb};
  assign p1_concat_131969_comb = {p1_smul_57470_NarrowedMult__comb, p1_smul_57454_TrailingBits___4_comb};
  assign p1_concat_131970_comb = {p1_smul_57476_NarrowedMult__comb, p1_smul_57454_TrailingBits___5_comb};
  assign p1_concat_131971_comb = {p1_smul_57478_NarrowedMult__comb, p1_smul_57454_TrailingBits___6_comb};
  assign p1_concat_131972_comb = {p1_smul_57484_NarrowedMult__comb, p1_smul_57454_TrailingBits___7_comb};
  assign p1_concat_131973_comb = {p1_smul_57550_NarrowedMult__comb, p1_smul_57454_TrailingBits___24_comb};
  assign p1_concat_131974_comb = {p1_smul_57556_NarrowedMult__comb, p1_smul_57454_TrailingBits___25_comb};
  assign p1_concat_131975_comb = {p1_smul_57558_NarrowedMult__comb, p1_smul_57454_TrailingBits___26_comb};
  assign p1_concat_131976_comb = {p1_smul_57564_NarrowedMult__comb, p1_smul_57454_TrailingBits___27_comb};
  assign p1_concat_131977_comb = {p1_smul_57600_NarrowedMult__comb, p1_smul_57330_TrailingBits___36_comb};
  assign p1_concat_131978_comb = {p1_smul_57604_NarrowedMult__comb, p1_smul_57330_TrailingBits___37_comb};
  assign p1_concat_131979_comb = {p1_smul_57606_NarrowedMult__comb, p1_smul_57330_TrailingBits___38_comb};
  assign p1_concat_131980_comb = {p1_smul_57610_NarrowedMult__comb, p1_smul_57330_TrailingBits___39_comb};
  assign p1_concat_131981_comb = {p1_smul_57680_NarrowedMult__comb, p1_smul_57330_TrailingBits___56_comb};
  assign p1_concat_131982_comb = {p1_smul_57684_NarrowedMult__comb, p1_smul_57330_TrailingBits___57_comb};
  assign p1_concat_131983_comb = {p1_smul_57686_NarrowedMult__comb, p1_smul_57330_TrailingBits___58_comb};
  assign p1_concat_131984_comb = {p1_smul_57690_NarrowedMult__comb, p1_smul_57330_TrailingBits___59_comb};
  assign p1_concat_131985_comb = {p1_smul_57854_NarrowedMult__comb, p1_smul_57330_TrailingBits___68_comb};
  assign p1_concat_131986_comb = {p1_smul_57858_NarrowedMult__comb, p1_smul_57330_TrailingBits___69_comb};
  assign p1_concat_131987_comb = {p1_smul_57864_NarrowedMult__comb, p1_smul_57330_TrailingBits___70_comb};
  assign p1_concat_131988_comb = {p1_smul_57868_NarrowedMult__comb, p1_smul_57330_TrailingBits___71_comb};
  assign p1_concat_131989_comb = {p1_smul_57934_NarrowedMult__comb, p1_smul_57330_TrailingBits___88_comb};
  assign p1_concat_131990_comb = {p1_smul_57938_NarrowedMult__comb, p1_smul_57330_TrailingBits___89_comb};
  assign p1_concat_131991_comb = {p1_smul_57944_NarrowedMult__comb, p1_smul_57330_TrailingBits___90_comb};
  assign p1_concat_131992_comb = {p1_smul_57948_NarrowedMult__comb, p1_smul_57330_TrailingBits___91_comb};
  assign p1_concat_131993_comb = {p1_smul_57984_NarrowedMult__comb, p1_smul_57454_TrailingBits___36_comb};
  assign p1_concat_131994_comb = {p1_smul_57988_NarrowedMult__comb, p1_smul_57454_TrailingBits___37_comb};
  assign p1_concat_131995_comb = {p1_smul_57990_NarrowedMult__comb, p1_smul_57454_TrailingBits___38_comb};
  assign p1_concat_131996_comb = {p1_smul_57994_NarrowedMult__comb, p1_smul_57454_TrailingBits___39_comb};
  assign p1_concat_131997_comb = {p1_smul_58064_NarrowedMult__comb, p1_smul_57454_TrailingBits___56_comb};
  assign p1_concat_131998_comb = {p1_smul_58068_NarrowedMult__comb, p1_smul_57454_TrailingBits___57_comb};
  assign p1_concat_131999_comb = {p1_smul_58070_NarrowedMult__comb, p1_smul_57454_TrailingBits___58_comb};
  assign p1_concat_132000_comb = {p1_smul_58074_NarrowedMult__comb, p1_smul_57454_TrailingBits___59_comb};
  assign p1_concat_132001_comb = {p1_smul_58110_NarrowedMult__comb, p1_smul_57330_TrailingBits___100_comb};
  assign p1_concat_132002_comb = {p1_smul_58112_NarrowedMult__comb, p1_smul_57330_TrailingBits___101_comb};
  assign p1_concat_132003_comb = {p1_smul_58122_NarrowedMult__comb, p1_smul_57330_TrailingBits___102_comb};
  assign p1_concat_132004_comb = {p1_smul_58124_NarrowedMult__comb, p1_smul_57330_TrailingBits___103_comb};
  assign p1_concat_132005_comb = {p1_smul_58190_NarrowedMult__comb, p1_smul_57330_TrailingBits___120_comb};
  assign p1_concat_132006_comb = {p1_smul_58192_NarrowedMult__comb, p1_smul_57330_TrailingBits___121_comb};
  assign p1_concat_132007_comb = {p1_smul_58202_NarrowedMult__comb, p1_smul_57330_TrailingBits___122_comb};
  assign p1_concat_132008_comb = {p1_smul_58204_NarrowedMult__comb, p1_smul_57330_TrailingBits___123_comb};
  assign p1_shifted__16_comb = {~p1_array_index_130681_comb[7], p1_array_index_130681_comb[6:0], p1_smul_57326_TrailingBits___144_comb};
  assign p1_smul_57326_TrailingBits___16_comb = 8'h00;
  assign p1_shifted__17_comb = {~p1_array_index_130689_comb[7], p1_array_index_130689_comb[6:0], p1_smul_57326_TrailingBits___145_comb};
  assign p1_smul_57326_TrailingBits___17_comb = 8'h00;
  assign p1_shifted__18_comb = {~p1_array_index_130665_comb[7], p1_array_index_130665_comb[6:0], p1_smul_57326_TrailingBits___146_comb};
  assign p1_smul_57326_TrailingBits___18_comb = 8'h00;
  assign p1_shifted__19_comb = {~p1_array_index_130666_comb[7], p1_array_index_130666_comb[6:0], p1_smul_57326_TrailingBits___147_comb};
  assign p1_smul_57326_TrailingBits___19_comb = 8'h00;
  assign p1_shifted__20_comb = {~p1_array_index_130667_comb[7], p1_array_index_130667_comb[6:0], p1_smul_57326_TrailingBits___148_comb};
  assign p1_smul_57326_TrailingBits___20_comb = 8'h00;
  assign p1_shifted__21_comb = {~p1_array_index_130668_comb[7], p1_array_index_130668_comb[6:0], p1_smul_57326_TrailingBits___149_comb};
  assign p1_smul_57326_TrailingBits___21_comb = 8'h00;
  assign p1_shifted__22_comb = {~p1_array_index_130690_comb[7], p1_array_index_130690_comb[6:0], p1_smul_57326_TrailingBits___150_comb};
  assign p1_smul_57326_TrailingBits___22_comb = 8'h00;
  assign p1_shifted__23_comb = {~p1_array_index_130682_comb[7], p1_array_index_130682_comb[6:0], p1_smul_57326_TrailingBits___151_comb};
  assign p1_smul_57326_TrailingBits___23_comb = 8'h00;
  assign p1_shifted__24_comb = {~p1_array_index_130683_comb[7], p1_array_index_130683_comb[6:0], p1_smul_57326_TrailingBits___152_comb};
  assign p1_smul_57326_TrailingBits___24_comb = 8'h00;
  assign p1_shifted__25_comb = {~p1_array_index_130691_comb[7], p1_array_index_130691_comb[6:0], p1_smul_57326_TrailingBits___153_comb};
  assign p1_smul_57326_TrailingBits___25_comb = 8'h00;
  assign p1_shifted__26_comb = {~p1_array_index_130669_comb[7], p1_array_index_130669_comb[6:0], p1_smul_57326_TrailingBits___154_comb};
  assign p1_smul_57326_TrailingBits___26_comb = 8'h00;
  assign p1_shifted__27_comb = {~p1_array_index_130670_comb[7], p1_array_index_130670_comb[6:0], p1_smul_57326_TrailingBits___155_comb};
  assign p1_smul_57326_TrailingBits___27_comb = 8'h00;
  assign p1_shifted__28_comb = {~p1_array_index_130671_comb[7], p1_array_index_130671_comb[6:0], p1_smul_57326_TrailingBits___156_comb};
  assign p1_smul_57326_TrailingBits___28_comb = 8'h00;
  assign p1_shifted__29_comb = {~p1_array_index_130672_comb[7], p1_array_index_130672_comb[6:0], p1_smul_57326_TrailingBits___157_comb};
  assign p1_smul_57326_TrailingBits___29_comb = 8'h00;
  assign p1_shifted__30_comb = {~p1_array_index_130692_comb[7], p1_array_index_130692_comb[6:0], p1_smul_57326_TrailingBits___158_comb};
  assign p1_smul_57326_TrailingBits___30_comb = 8'h00;
  assign p1_shifted__31_comb = {~p1_array_index_130684_comb[7], p1_array_index_130684_comb[6:0], p1_smul_57326_TrailingBits___159_comb};
  assign p1_smul_57326_TrailingBits___31_comb = 8'h00;
  assign p1_shifted__32_comb = {~p1_array_index_130685_comb[7], p1_array_index_130685_comb[6:0], p1_smul_57326_TrailingBits___160_comb};
  assign p1_smul_57326_TrailingBits___32_comb = 8'h00;
  assign p1_shifted__33_comb = {~p1_array_index_130693_comb[7], p1_array_index_130693_comb[6:0], p1_smul_57326_TrailingBits___161_comb};
  assign p1_smul_57326_TrailingBits___33_comb = 8'h00;
  assign p1_shifted__34_comb = {~p1_array_index_130673_comb[7], p1_array_index_130673_comb[6:0], p1_smul_57326_TrailingBits___162_comb};
  assign p1_smul_57326_TrailingBits___34_comb = 8'h00;
  assign p1_shifted__35_comb = {~p1_array_index_130674_comb[7], p1_array_index_130674_comb[6:0], p1_smul_57326_TrailingBits___163_comb};
  assign p1_smul_57326_TrailingBits___35_comb = 8'h00;
  assign p1_shifted__36_comb = {~p1_array_index_130675_comb[7], p1_array_index_130675_comb[6:0], p1_smul_57326_TrailingBits___164_comb};
  assign p1_smul_57326_TrailingBits___36_comb = 8'h00;
  assign p1_shifted__37_comb = {~p1_array_index_130676_comb[7], p1_array_index_130676_comb[6:0], p1_smul_57326_TrailingBits___165_comb};
  assign p1_smul_57326_TrailingBits___37_comb = 8'h00;
  assign p1_shifted__38_comb = {~p1_array_index_130694_comb[7], p1_array_index_130694_comb[6:0], p1_smul_57326_TrailingBits___166_comb};
  assign p1_smul_57326_TrailingBits___38_comb = 8'h00;
  assign p1_shifted__39_comb = {~p1_array_index_130686_comb[7], p1_array_index_130686_comb[6:0], p1_smul_57326_TrailingBits___167_comb};
  assign p1_smul_57326_TrailingBits___39_comb = 8'h00;
  assign p1_shifted__40_comb = {~p1_array_index_130687_comb[7], p1_array_index_130687_comb[6:0], p1_smul_57326_TrailingBits___168_comb};
  assign p1_smul_57326_TrailingBits___40_comb = 8'h00;
  assign p1_shifted__41_comb = {~p1_array_index_130695_comb[7], p1_array_index_130695_comb[6:0], p1_smul_57326_TrailingBits___169_comb};
  assign p1_smul_57326_TrailingBits___41_comb = 8'h00;
  assign p1_shifted__42_comb = {~p1_array_index_130677_comb[7], p1_array_index_130677_comb[6:0], p1_smul_57326_TrailingBits___170_comb};
  assign p1_smul_57326_TrailingBits___42_comb = 8'h00;
  assign p1_shifted__43_comb = {~p1_array_index_130678_comb[7], p1_array_index_130678_comb[6:0], p1_smul_57326_TrailingBits___171_comb};
  assign p1_smul_57326_TrailingBits___43_comb = 8'h00;
  assign p1_shifted__44_comb = {~p1_array_index_130679_comb[7], p1_array_index_130679_comb[6:0], p1_smul_57326_TrailingBits___172_comb};
  assign p1_smul_57326_TrailingBits___44_comb = 8'h00;
  assign p1_shifted__45_comb = {~p1_array_index_130680_comb[7], p1_array_index_130680_comb[6:0], p1_smul_57326_TrailingBits___173_comb};
  assign p1_smul_57326_TrailingBits___45_comb = 8'h00;
  assign p1_shifted__46_comb = {~p1_array_index_130696_comb[7], p1_array_index_130696_comb[6:0], p1_smul_57326_TrailingBits___174_comb};
  assign p1_smul_57326_TrailingBits___46_comb = 8'h00;
  assign p1_shifted__47_comb = {~p1_array_index_130688_comb[7], p1_array_index_130688_comb[6:0], p1_smul_57326_TrailingBits___175_comb};
  assign p1_smul_57326_TrailingBits___47_comb = 8'h00;
  assign p1_prod__135_comb = {{7{p1_concat_131721_comb[24]}}, p1_concat_131721_comb};
  assign p1_prod__139_comb = {{9{p1_concat_131722_comb[22]}}, p1_concat_131722_comb};
  assign p1_prod__144_comb = {{9{p1_concat_131723_comb[22]}}, p1_concat_131723_comb};
  assign p1_prod__150_comb = {{7{p1_concat_131724_comb[24]}}, p1_concat_131724_comb};
  assign p1_prod__199_comb = {{7{p1_concat_131725_comb[24]}}, p1_concat_131725_comb};
  assign p1_prod__203_comb = {{9{p1_concat_131726_comb[22]}}, p1_concat_131726_comb};
  assign p1_prod__208_comb = {{9{p1_concat_131727_comb[22]}}, p1_concat_131727_comb};
  assign p1_prod__214_comb = {{7{p1_concat_131728_comb[24]}}, p1_concat_131728_comb};
  assign p1_prod__263_comb = {{7{p1_concat_131729_comb[24]}}, p1_concat_131729_comb};
  assign p1_prod__267_comb = {{9{p1_concat_131730_comb[22]}}, p1_concat_131730_comb};
  assign p1_prod__272_comb = {{9{p1_concat_131731_comb[22]}}, p1_concat_131731_comb};
  assign p1_prod__278_comb = {{7{p1_concat_131732_comb[24]}}, p1_concat_131732_comb};
  assign p1_prod__327_comb = {{7{p1_concat_131733_comb[24]}}, p1_concat_131733_comb};
  assign p1_prod__331_comb = {{9{p1_concat_131734_comb[22]}}, p1_concat_131734_comb};
  assign p1_prod__336_comb = {{9{p1_concat_131735_comb[22]}}, p1_concat_131735_comb};
  assign p1_prod__342_comb = {{7{p1_concat_131736_comb[24]}}, p1_concat_131736_comb};
  assign p1_prod__133_comb = {{7{p1_concat_131737_comb[24]}}, p1_concat_131737_comb};
  assign p1_prod__145_comb = {{7{p1_concat_131738_comb[24]}}, p1_concat_131738_comb};
  assign p1_prod__151_comb = {{7{p1_concat_131739_comb[24]}}, p1_concat_131739_comb};
  assign p1_prod__171_comb = {{7{p1_concat_131740_comb[24]}}, p1_concat_131740_comb};
  assign p1_prod__197_comb = {{7{p1_concat_131741_comb[24]}}, p1_concat_131741_comb};
  assign p1_prod__209_comb = {{7{p1_concat_131742_comb[24]}}, p1_concat_131742_comb};
  assign p1_prod__215_comb = {{7{p1_concat_131743_comb[24]}}, p1_concat_131743_comb};
  assign p1_prod__235_comb = {{7{p1_concat_131744_comb[24]}}, p1_concat_131744_comb};
  assign p1_prod__261_comb = {{7{p1_concat_131745_comb[24]}}, p1_concat_131745_comb};
  assign p1_prod__273_comb = {{7{p1_concat_131746_comb[24]}}, p1_concat_131746_comb};
  assign p1_prod__279_comb = {{7{p1_concat_131747_comb[24]}}, p1_concat_131747_comb};
  assign p1_prod__299_comb = {{7{p1_concat_131748_comb[24]}}, p1_concat_131748_comb};
  assign p1_prod__325_comb = {{7{p1_concat_131749_comb[24]}}, p1_concat_131749_comb};
  assign p1_prod__337_comb = {{7{p1_concat_131750_comb[24]}}, p1_concat_131750_comb};
  assign p1_prod__343_comb = {{7{p1_concat_131751_comb[24]}}, p1_concat_131751_comb};
  assign p1_prod__363_comb = {{7{p1_concat_131752_comb[24]}}, p1_concat_131752_comb};
  assign p1_prod__141_comb = {{9{p1_concat_131753_comb[22]}}, p1_concat_131753_comb};
  assign p1_prod__152_comb = {{7{p1_concat_131754_comb[24]}}, p1_concat_131754_comb};
  assign p1_prod__159_comb = {{7{p1_concat_131755_comb[24]}}, p1_concat_131755_comb};
  assign p1_prod__172_comb = {{9{p1_concat_131756_comb[22]}}, p1_concat_131756_comb};
  assign p1_prod__205_comb = {{9{p1_concat_131757_comb[22]}}, p1_concat_131757_comb};
  assign p1_prod__216_comb = {{7{p1_concat_131758_comb[24]}}, p1_concat_131758_comb};
  assign p1_prod__223_comb = {{7{p1_concat_131759_comb[24]}}, p1_concat_131759_comb};
  assign p1_prod__236_comb = {{9{p1_concat_131760_comb[22]}}, p1_concat_131760_comb};
  assign p1_prod__269_comb = {{9{p1_concat_131761_comb[22]}}, p1_concat_131761_comb};
  assign p1_prod__280_comb = {{7{p1_concat_131762_comb[24]}}, p1_concat_131762_comb};
  assign p1_prod__287_comb = {{7{p1_concat_131763_comb[24]}}, p1_concat_131763_comb};
  assign p1_prod__300_comb = {{9{p1_concat_131764_comb[22]}}, p1_concat_131764_comb};
  assign p1_prod__333_comb = {{9{p1_concat_131765_comb[22]}}, p1_concat_131765_comb};
  assign p1_prod__344_comb = {{7{p1_concat_131766_comb[24]}}, p1_concat_131766_comb};
  assign p1_prod__351_comb = {{7{p1_concat_131767_comb[24]}}, p1_concat_131767_comb};
  assign p1_prod__364_comb = {{9{p1_concat_131768_comb[22]}}, p1_concat_131768_comb};
  assign p1_prod__148_comb = {{7{p1_concat_131769_comb[24]}}, p1_concat_131769_comb};
  assign p1_prod__161_comb = {{9{p1_concat_131770_comb[22]}}, p1_concat_131770_comb};
  assign p1_prod__179_comb = {{9{p1_concat_131771_comb[22]}}, p1_concat_131771_comb};
  assign p1_prod__186_comb = {{7{p1_concat_131772_comb[24]}}, p1_concat_131772_comb};
  assign p1_prod__212_comb = {{7{p1_concat_131773_comb[24]}}, p1_concat_131773_comb};
  assign p1_prod__225_comb = {{9{p1_concat_131774_comb[22]}}, p1_concat_131774_comb};
  assign p1_prod__243_comb = {{9{p1_concat_131775_comb[22]}}, p1_concat_131775_comb};
  assign p1_prod__250_comb = {{7{p1_concat_131776_comb[24]}}, p1_concat_131776_comb};
  assign p1_prod__276_comb = {{7{p1_concat_131777_comb[24]}}, p1_concat_131777_comb};
  assign p1_prod__289_comb = {{9{p1_concat_131778_comb[22]}}, p1_concat_131778_comb};
  assign p1_prod__307_comb = {{9{p1_concat_131779_comb[22]}}, p1_concat_131779_comb};
  assign p1_prod__314_comb = {{7{p1_concat_131780_comb[24]}}, p1_concat_131780_comb};
  assign p1_prod__340_comb = {{7{p1_concat_131781_comb[24]}}, p1_concat_131781_comb};
  assign p1_prod__353_comb = {{9{p1_concat_131782_comb[22]}}, p1_concat_131782_comb};
  assign p1_prod__371_comb = {{9{p1_concat_131783_comb[22]}}, p1_concat_131783_comb};
  assign p1_prod__378_comb = {{7{p1_concat_131784_comb[24]}}, p1_concat_131784_comb};
  assign p1_prod__162_comb = {{7{p1_concat_131785_comb[24]}}, p1_concat_131785_comb};
  assign p1_prod__175_comb = {{7{p1_concat_131786_comb[24]}}, p1_concat_131786_comb};
  assign p1_prod__180_comb = {{7{p1_concat_131787_comb[24]}}, p1_concat_131787_comb};
  assign p1_prod__187_comb = {{7{p1_concat_131788_comb[24]}}, p1_concat_131788_comb};
  assign p1_prod__226_comb = {{7{p1_concat_131789_comb[24]}}, p1_concat_131789_comb};
  assign p1_prod__239_comb = {{7{p1_concat_131790_comb[24]}}, p1_concat_131790_comb};
  assign p1_prod__244_comb = {{7{p1_concat_131791_comb[24]}}, p1_concat_131791_comb};
  assign p1_prod__251_comb = {{7{p1_concat_131792_comb[24]}}, p1_concat_131792_comb};
  assign p1_prod__290_comb = {{7{p1_concat_131793_comb[24]}}, p1_concat_131793_comb};
  assign p1_prod__303_comb = {{7{p1_concat_131794_comb[24]}}, p1_concat_131794_comb};
  assign p1_prod__308_comb = {{7{p1_concat_131795_comb[24]}}, p1_concat_131795_comb};
  assign p1_prod__315_comb = {{7{p1_concat_131796_comb[24]}}, p1_concat_131796_comb};
  assign p1_prod__354_comb = {{7{p1_concat_131797_comb[24]}}, p1_concat_131797_comb};
  assign p1_prod__367_comb = {{7{p1_concat_131798_comb[24]}}, p1_concat_131798_comb};
  assign p1_prod__372_comb = {{7{p1_concat_131799_comb[24]}}, p1_concat_131799_comb};
  assign p1_prod__379_comb = {{7{p1_concat_131800_comb[24]}}, p1_concat_131800_comb};
  assign p1_prod__163_comb = {{9{p1_concat_131801_comb[22]}}, p1_concat_131801_comb};
  assign p1_prod__170_comb = {{7{p1_concat_131802_comb[24]}}, p1_concat_131802_comb};
  assign p1_prod__190_comb = {{7{p1_concat_131803_comb[24]}}, p1_concat_131803_comb};
  assign p1_prod__191_comb = {{9{p1_concat_131804_comb[22]}}, p1_concat_131804_comb};
  assign p1_prod__227_comb = {{9{p1_concat_131805_comb[22]}}, p1_concat_131805_comb};
  assign p1_prod__234_comb = {{7{p1_concat_131806_comb[24]}}, p1_concat_131806_comb};
  assign p1_prod__254_comb = {{7{p1_concat_131807_comb[24]}}, p1_concat_131807_comb};
  assign p1_prod__255_comb = {{9{p1_concat_131808_comb[22]}}, p1_concat_131808_comb};
  assign p1_prod__291_comb = {{9{p1_concat_131809_comb[22]}}, p1_concat_131809_comb};
  assign p1_prod__298_comb = {{7{p1_concat_131810_comb[24]}}, p1_concat_131810_comb};
  assign p1_prod__318_comb = {{7{p1_concat_131811_comb[24]}}, p1_concat_131811_comb};
  assign p1_prod__319_comb = {{9{p1_concat_131812_comb[22]}}, p1_concat_131812_comb};
  assign p1_prod__355_comb = {{9{p1_concat_131813_comb[22]}}, p1_concat_131813_comb};
  assign p1_prod__362_comb = {{7{p1_concat_131814_comb[24]}}, p1_concat_131814_comb};
  assign p1_prod__382_comb = {{7{p1_concat_131815_comb[24]}}, p1_concat_131815_comb};
  assign p1_prod__383_comb = {{9{p1_concat_131816_comb[22]}}, p1_concat_131816_comb};
  assign p1_shifted_comb = {~p1_array_index_130705_comb[7], p1_array_index_130705_comb[6:0], p1_smul_57326_TrailingBits___128_comb};
  assign p1_smul_57326_TrailingBits__comb = 8'h00;
  assign p1_shifted__1_comb = {~p1_array_index_130709_comb[7], p1_array_index_130709_comb[6:0], p1_smul_57326_TrailingBits___129_comb};
  assign p1_smul_57326_TrailingBits___1_comb = 8'h00;
  assign p1_shifted__2_comb = {~p1_array_index_130697_comb[7], p1_array_index_130697_comb[6:0], p1_smul_57326_TrailingBits___130_comb};
  assign p1_smul_57326_TrailingBits___2_comb = 8'h00;
  assign p1_shifted__3_comb = {~p1_array_index_130698_comb[7], p1_array_index_130698_comb[6:0], p1_smul_57326_TrailingBits___131_comb};
  assign p1_smul_57326_TrailingBits___3_comb = 8'h00;
  assign p1_shifted__4_comb = {~p1_array_index_130699_comb[7], p1_array_index_130699_comb[6:0], p1_smul_57326_TrailingBits___132_comb};
  assign p1_smul_57326_TrailingBits___4_comb = 8'h00;
  assign p1_shifted__5_comb = {~p1_array_index_130700_comb[7], p1_array_index_130700_comb[6:0], p1_smul_57326_TrailingBits___133_comb};
  assign p1_smul_57326_TrailingBits___5_comb = 8'h00;
  assign p1_shifted__6_comb = {~p1_array_index_130710_comb[7], p1_array_index_130710_comb[6:0], p1_smul_57326_TrailingBits___134_comb};
  assign p1_smul_57326_TrailingBits___6_comb = 8'h00;
  assign p1_shifted__7_comb = {~p1_array_index_130706_comb[7], p1_array_index_130706_comb[6:0], p1_smul_57326_TrailingBits___135_comb};
  assign p1_smul_57326_TrailingBits___7_comb = 8'h00;
  assign p1_shifted__56_comb = {~p1_array_index_130707_comb[7], p1_array_index_130707_comb[6:0], p1_smul_57326_TrailingBits___184_comb};
  assign p1_smul_57326_TrailingBits___56_comb = 8'h00;
  assign p1_shifted__57_comb = {~p1_array_index_130711_comb[7], p1_array_index_130711_comb[6:0], p1_smul_57326_TrailingBits___185_comb};
  assign p1_smul_57326_TrailingBits___57_comb = 8'h00;
  assign p1_shifted__58_comb = {~p1_array_index_130701_comb[7], p1_array_index_130701_comb[6:0], p1_smul_57326_TrailingBits___186_comb};
  assign p1_smul_57326_TrailingBits___58_comb = 8'h00;
  assign p1_shifted__59_comb = {~p1_array_index_130702_comb[7], p1_array_index_130702_comb[6:0], p1_smul_57326_TrailingBits___187_comb};
  assign p1_smul_57326_TrailingBits___59_comb = 8'h00;
  assign p1_shifted__60_comb = {~p1_array_index_130703_comb[7], p1_array_index_130703_comb[6:0], p1_smul_57326_TrailingBits___188_comb};
  assign p1_smul_57326_TrailingBits___60_comb = 8'h00;
  assign p1_shifted__61_comb = {~p1_array_index_130704_comb[7], p1_array_index_130704_comb[6:0], p1_smul_57326_TrailingBits___189_comb};
  assign p1_smul_57326_TrailingBits___61_comb = 8'h00;
  assign p1_shifted__62_comb = {~p1_array_index_130712_comb[7], p1_array_index_130712_comb[6:0], p1_smul_57326_TrailingBits___190_comb};
  assign p1_smul_57326_TrailingBits___62_comb = 8'h00;
  assign p1_shifted__63_comb = {~p1_array_index_130708_comb[7], p1_array_index_130708_comb[6:0], p1_smul_57326_TrailingBits___191_comb};
  assign p1_smul_57326_TrailingBits___63_comb = 8'h00;
  assign p1_prod__10_comb = {{7{p1_concat_131865_comb[24]}}, p1_concat_131865_comb};
  assign p1_prod__11_comb = {{9{p1_concat_131866_comb[22]}}, p1_concat_131866_comb};
  assign p1_prod__12_comb = {{9{p1_concat_131867_comb[22]}}, p1_concat_131867_comb};
  assign p1_prod__13_comb = {{7{p1_concat_131868_comb[24]}}, p1_concat_131868_comb};
  assign p1_prod__455_comb = {{7{p1_concat_131869_comb[24]}}, p1_concat_131869_comb};
  assign p1_prod__459_comb = {{9{p1_concat_131870_comb[22]}}, p1_concat_131870_comb};
  assign p1_prod__464_comb = {{9{p1_concat_131871_comb[22]}}, p1_concat_131871_comb};
  assign p1_prod__470_comb = {{7{p1_concat_131872_comb[24]}}, p1_concat_131872_comb};
  assign p1_prod__16_comb = {{7{p1_concat_131873_comb[24]}}, p1_concat_131873_comb};
  assign p1_prod__19_comb = {{7{p1_concat_131874_comb[24]}}, p1_concat_131874_comb};
  assign p1_prod__20_comb = {{7{p1_concat_131875_comb[24]}}, p1_concat_131875_comb};
  assign p1_prod__23_comb = {{7{p1_concat_131876_comb[24]}}, p1_concat_131876_comb};
  assign p1_prod__453_comb = {{7{p1_concat_131877_comb[24]}}, p1_concat_131877_comb};
  assign p1_prod__465_comb = {{7{p1_concat_131878_comb[24]}}, p1_concat_131878_comb};
  assign p1_prod__471_comb = {{7{p1_concat_131879_comb[24]}}, p1_concat_131879_comb};
  assign p1_prod__491_comb = {{7{p1_concat_131880_comb[24]}}, p1_concat_131880_comb};
  assign p1_prod__25_comb = {{9{p1_concat_131881_comb[22]}}, p1_concat_131881_comb};
  assign p1_prod__27_comb = {{7{p1_concat_131882_comb[24]}}, p1_concat_131882_comb};
  assign p1_prod__28_comb = {{7{p1_concat_131883_comb[24]}}, p1_concat_131883_comb};
  assign p1_prod__30_comb = {{9{p1_concat_131884_comb[22]}}, p1_concat_131884_comb};
  assign p1_prod__461_comb = {{9{p1_concat_131885_comb[22]}}, p1_concat_131885_comb};
  assign p1_prod__472_comb = {{7{p1_concat_131886_comb[24]}}, p1_concat_131886_comb};
  assign p1_prod__479_comb = {{7{p1_concat_131887_comb[24]}}, p1_concat_131887_comb};
  assign p1_prod__492_comb = {{9{p1_concat_131888_comb[22]}}, p1_concat_131888_comb};
  assign p1_prod__40_comb = {{7{p1_concat_131889_comb[24]}}, p1_concat_131889_comb};
  assign p1_prod__42_comb = {{9{p1_concat_131890_comb[22]}}, p1_concat_131890_comb};
  assign p1_prod__45_comb = {{9{p1_concat_131891_comb[22]}}, p1_concat_131891_comb};
  assign p1_prod__47_comb = {{7{p1_concat_131892_comb[24]}}, p1_concat_131892_comb};
  assign p1_prod__468_comb = {{7{p1_concat_131893_comb[24]}}, p1_concat_131893_comb};
  assign p1_prod__481_comb = {{9{p1_concat_131894_comb[22]}}, p1_concat_131894_comb};
  assign p1_prod__499_comb = {{9{p1_concat_131895_comb[22]}}, p1_concat_131895_comb};
  assign p1_prod__506_comb = {{7{p1_concat_131896_comb[24]}}, p1_concat_131896_comb};
  assign p1_prod__49_comb = {{7{p1_concat_131897_comb[24]}}, p1_concat_131897_comb};
  assign p1_prod__51_comb = {{7{p1_concat_131898_comb[24]}}, p1_concat_131898_comb};
  assign p1_prod__52_comb = {{7{p1_concat_131899_comb[24]}}, p1_concat_131899_comb};
  assign p1_prod__54_comb = {{7{p1_concat_131900_comb[24]}}, p1_concat_131900_comb};
  assign p1_prod__482_comb = {{7{p1_concat_131901_comb[24]}}, p1_concat_131901_comb};
  assign p1_prod__495_comb = {{7{p1_concat_131902_comb[24]}}, p1_concat_131902_comb};
  assign p1_prod__500_comb = {{7{p1_concat_131903_comb[24]}}, p1_concat_131903_comb};
  assign p1_prod__507_comb = {{7{p1_concat_131904_comb[24]}}, p1_concat_131904_comb};
  assign p1_prod__56_comb = {{9{p1_concat_131905_comb[22]}}, p1_concat_131905_comb};
  assign p1_prod__57_comb = {{7{p1_concat_131906_comb[24]}}, p1_concat_131906_comb};
  assign p1_prod__62_comb = {{7{p1_concat_131907_comb[24]}}, p1_concat_131907_comb};
  assign p1_prod__63_comb = {{9{p1_concat_131908_comb[22]}}, p1_concat_131908_comb};
  assign p1_prod__483_comb = {{9{p1_concat_131909_comb[22]}}, p1_concat_131909_comb};
  assign p1_prod__490_comb = {{7{p1_concat_131910_comb[24]}}, p1_concat_131910_comb};
  assign p1_prod__510_comb = {{7{p1_concat_131911_comb[24]}}, p1_concat_131911_comb};
  assign p1_prod__511_comb = {{9{p1_concat_131912_comb[22]}}, p1_concat_131912_comb};
  assign p1_shifted__8_comb = {~p1_array_index_130721_comb[7], p1_array_index_130721_comb[6:0], p1_smul_57326_TrailingBits___136_comb};
  assign p1_smul_57326_TrailingBits___8_comb = 8'h00;
  assign p1_shifted__9_comb = {~p1_array_index_130725_comb[7], p1_array_index_130725_comb[6:0], p1_smul_57326_TrailingBits___137_comb};
  assign p1_smul_57326_TrailingBits___9_comb = 8'h00;
  assign p1_shifted__10_comb = {~p1_array_index_130713_comb[7], p1_array_index_130713_comb[6:0], p1_smul_57326_TrailingBits___138_comb};
  assign p1_smul_57326_TrailingBits___10_comb = 8'h00;
  assign p1_shifted__11_comb = {~p1_array_index_130714_comb[7], p1_array_index_130714_comb[6:0], p1_smul_57326_TrailingBits___139_comb};
  assign p1_smul_57326_TrailingBits___11_comb = 8'h00;
  assign p1_shifted__12_comb = {~p1_array_index_130715_comb[7], p1_array_index_130715_comb[6:0], p1_smul_57326_TrailingBits___140_comb};
  assign p1_smul_57326_TrailingBits___12_comb = 8'h00;
  assign p1_shifted__13_comb = {~p1_array_index_130716_comb[7], p1_array_index_130716_comb[6:0], p1_smul_57326_TrailingBits___141_comb};
  assign p1_smul_57326_TrailingBits___13_comb = 8'h00;
  assign p1_shifted__14_comb = {~p1_array_index_130726_comb[7], p1_array_index_130726_comb[6:0], p1_smul_57326_TrailingBits___142_comb};
  assign p1_smul_57326_TrailingBits___14_comb = 8'h00;
  assign p1_shifted__15_comb = {~p1_array_index_130722_comb[7], p1_array_index_130722_comb[6:0], p1_smul_57326_TrailingBits___143_comb};
  assign p1_smul_57326_TrailingBits___15_comb = 8'h00;
  assign p1_shifted__48_comb = {~p1_array_index_130723_comb[7], p1_array_index_130723_comb[6:0], p1_smul_57326_TrailingBits___176_comb};
  assign p1_smul_57326_TrailingBits___48_comb = 8'h00;
  assign p1_shifted__49_comb = {~p1_array_index_130727_comb[7], p1_array_index_130727_comb[6:0], p1_smul_57326_TrailingBits___177_comb};
  assign p1_smul_57326_TrailingBits___49_comb = 8'h00;
  assign p1_shifted__50_comb = {~p1_array_index_130717_comb[7], p1_array_index_130717_comb[6:0], p1_smul_57326_TrailingBits___178_comb};
  assign p1_smul_57326_TrailingBits___50_comb = 8'h00;
  assign p1_shifted__51_comb = {~p1_array_index_130718_comb[7], p1_array_index_130718_comb[6:0], p1_smul_57326_TrailingBits___179_comb};
  assign p1_smul_57326_TrailingBits___51_comb = 8'h00;
  assign p1_shifted__52_comb = {~p1_array_index_130719_comb[7], p1_array_index_130719_comb[6:0], p1_smul_57326_TrailingBits___180_comb};
  assign p1_smul_57326_TrailingBits___52_comb = 8'h00;
  assign p1_shifted__53_comb = {~p1_array_index_130720_comb[7], p1_array_index_130720_comb[6:0], p1_smul_57326_TrailingBits___181_comb};
  assign p1_smul_57326_TrailingBits___53_comb = 8'h00;
  assign p1_shifted__54_comb = {~p1_array_index_130728_comb[7], p1_array_index_130728_comb[6:0], p1_smul_57326_TrailingBits___182_comb};
  assign p1_smul_57326_TrailingBits___54_comb = 8'h00;
  assign p1_shifted__55_comb = {~p1_array_index_130724_comb[7], p1_array_index_130724_comb[6:0], p1_smul_57326_TrailingBits___183_comb};
  assign p1_smul_57326_TrailingBits___55_comb = 8'h00;
  assign p1_prod__71_comb = {{7{p1_concat_131961_comb[24]}}, p1_concat_131961_comb};
  assign p1_prod__75_comb = {{9{p1_concat_131962_comb[22]}}, p1_concat_131962_comb};
  assign p1_prod__80_comb = {{9{p1_concat_131963_comb[22]}}, p1_concat_131963_comb};
  assign p1_prod__86_comb = {{7{p1_concat_131964_comb[24]}}, p1_concat_131964_comb};
  assign p1_prod__391_comb = {{7{p1_concat_131965_comb[24]}}, p1_concat_131965_comb};
  assign p1_prod__395_comb = {{9{p1_concat_131966_comb[22]}}, p1_concat_131966_comb};
  assign p1_prod__400_comb = {{9{p1_concat_131967_comb[22]}}, p1_concat_131967_comb};
  assign p1_prod__406_comb = {{7{p1_concat_131968_comb[24]}}, p1_concat_131968_comb};
  assign p1_prod__69_comb = {{7{p1_concat_131969_comb[24]}}, p1_concat_131969_comb};
  assign p1_prod__81_comb = {{7{p1_concat_131970_comb[24]}}, p1_concat_131970_comb};
  assign p1_prod__87_comb = {{7{p1_concat_131971_comb[24]}}, p1_concat_131971_comb};
  assign p1_prod__107_comb = {{7{p1_concat_131972_comb[24]}}, p1_concat_131972_comb};
  assign p1_prod__389_comb = {{7{p1_concat_131973_comb[24]}}, p1_concat_131973_comb};
  assign p1_prod__401_comb = {{7{p1_concat_131974_comb[24]}}, p1_concat_131974_comb};
  assign p1_prod__407_comb = {{7{p1_concat_131975_comb[24]}}, p1_concat_131975_comb};
  assign p1_prod__427_comb = {{7{p1_concat_131976_comb[24]}}, p1_concat_131976_comb};
  assign p1_prod__77_comb = {{9{p1_concat_131977_comb[22]}}, p1_concat_131977_comb};
  assign p1_prod__88_comb = {{7{p1_concat_131978_comb[24]}}, p1_concat_131978_comb};
  assign p1_prod__95_comb = {{7{p1_concat_131979_comb[24]}}, p1_concat_131979_comb};
  assign p1_prod__108_comb = {{9{p1_concat_131980_comb[22]}}, p1_concat_131980_comb};
  assign p1_prod__397_comb = {{9{p1_concat_131981_comb[22]}}, p1_concat_131981_comb};
  assign p1_prod__408_comb = {{7{p1_concat_131982_comb[24]}}, p1_concat_131982_comb};
  assign p1_prod__415_comb = {{7{p1_concat_131983_comb[24]}}, p1_concat_131983_comb};
  assign p1_prod__428_comb = {{9{p1_concat_131984_comb[22]}}, p1_concat_131984_comb};
  assign p1_prod__84_comb = {{7{p1_concat_131985_comb[24]}}, p1_concat_131985_comb};
  assign p1_prod__97_comb = {{9{p1_concat_131986_comb[22]}}, p1_concat_131986_comb};
  assign p1_prod__115_comb = {{9{p1_concat_131987_comb[22]}}, p1_concat_131987_comb};
  assign p1_prod__122_comb = {{7{p1_concat_131988_comb[24]}}, p1_concat_131988_comb};
  assign p1_prod__404_comb = {{7{p1_concat_131989_comb[24]}}, p1_concat_131989_comb};
  assign p1_prod__417_comb = {{9{p1_concat_131990_comb[22]}}, p1_concat_131990_comb};
  assign p1_prod__435_comb = {{9{p1_concat_131991_comb[22]}}, p1_concat_131991_comb};
  assign p1_prod__442_comb = {{7{p1_concat_131992_comb[24]}}, p1_concat_131992_comb};
  assign p1_prod__98_comb = {{7{p1_concat_131993_comb[24]}}, p1_concat_131993_comb};
  assign p1_prod__111_comb = {{7{p1_concat_131994_comb[24]}}, p1_concat_131994_comb};
  assign p1_prod__116_comb = {{7{p1_concat_131995_comb[24]}}, p1_concat_131995_comb};
  assign p1_prod__123_comb = {{7{p1_concat_131996_comb[24]}}, p1_concat_131996_comb};
  assign p1_prod__418_comb = {{7{p1_concat_131997_comb[24]}}, p1_concat_131997_comb};
  assign p1_prod__431_comb = {{7{p1_concat_131998_comb[24]}}, p1_concat_131998_comb};
  assign p1_prod__436_comb = {{7{p1_concat_131999_comb[24]}}, p1_concat_131999_comb};
  assign p1_prod__443_comb = {{7{p1_concat_132000_comb[24]}}, p1_concat_132000_comb};
  assign p1_prod__99_comb = {{9{p1_concat_132001_comb[22]}}, p1_concat_132001_comb};
  assign p1_prod__106_comb = {{7{p1_concat_132002_comb[24]}}, p1_concat_132002_comb};
  assign p1_prod__126_comb = {{7{p1_concat_132003_comb[24]}}, p1_concat_132003_comb};
  assign p1_prod__127_comb = {{9{p1_concat_132004_comb[22]}}, p1_concat_132004_comb};
  assign p1_prod__419_comb = {{9{p1_concat_132005_comb[22]}}, p1_concat_132005_comb};
  assign p1_prod__426_comb = {{7{p1_concat_132006_comb[24]}}, p1_concat_132006_comb};
  assign p1_prod__446_comb = {{7{p1_concat_132007_comb[24]}}, p1_concat_132007_comb};
  assign p1_prod__447_comb = {{9{p1_concat_132008_comb[22]}}, p1_concat_132008_comb};
  assign p1_or_132809_comb = p1_prod__135_comb | 32'h0000_0080;
  assign p1_or_132810_comb = p1_prod__139_comb | 32'h0000_0080;
  assign p1_or_132811_comb = p1_prod__144_comb | 32'h0000_0080;
  assign p1_or_132812_comb = p1_prod__150_comb | 32'h0000_0080;
  assign p1_or_132813_comb = p1_prod__199_comb | 32'h0000_0080;
  assign p1_or_132814_comb = p1_prod__203_comb | 32'h0000_0080;
  assign p1_or_132815_comb = p1_prod__208_comb | 32'h0000_0080;
  assign p1_or_132816_comb = p1_prod__214_comb | 32'h0000_0080;
  assign p1_or_132817_comb = p1_prod__263_comb | 32'h0000_0080;
  assign p1_or_132818_comb = p1_prod__267_comb | 32'h0000_0080;
  assign p1_or_132819_comb = p1_prod__272_comb | 32'h0000_0080;
  assign p1_or_132820_comb = p1_prod__278_comb | 32'h0000_0080;
  assign p1_or_132821_comb = p1_prod__327_comb | 32'h0000_0080;
  assign p1_or_132822_comb = p1_prod__331_comb | 32'h0000_0080;
  assign p1_or_132823_comb = p1_prod__336_comb | 32'h0000_0080;
  assign p1_or_132824_comb = p1_prod__342_comb | 32'h0000_0080;
  assign p1_or_132825_comb = p1_prod__133_comb | 32'h0000_0080;
  assign p1_smul_57488_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__17_squeezed_comb, 7'h31);
  assign p1_smul_57490_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__18_squeezed_comb, 7'h4f);
  assign p1_or_132830_comb = p1_prod__145_comb | 32'h0000_0080;
  assign p1_or_132831_comb = p1_prod__151_comb | 32'h0000_0080;
  assign p1_smul_57496_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__21_squeezed_comb, 7'h4f);
  assign p1_smul_57498_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__22_squeezed_comb, 7'h31);
  assign p1_or_132836_comb = p1_prod__171_comb | 32'h0000_0080;
  assign p1_or_132837_comb = p1_prod__197_comb | 32'h0000_0080;
  assign p1_smul_57504_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__25_squeezed_comb, 7'h31);
  assign p1_smul_57506_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__26_squeezed_comb, 7'h4f);
  assign p1_or_132842_comb = p1_prod__209_comb | 32'h0000_0080;
  assign p1_or_132843_comb = p1_prod__215_comb | 32'h0000_0080;
  assign p1_smul_57512_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__29_squeezed_comb, 7'h4f);
  assign p1_smul_57514_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__30_squeezed_comb, 7'h31);
  assign p1_or_132848_comb = p1_prod__235_comb | 32'h0000_0080;
  assign p1_or_132849_comb = p1_prod__261_comb | 32'h0000_0080;
  assign p1_smul_57520_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__33_squeezed_comb, 7'h31);
  assign p1_smul_57522_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__34_squeezed_comb, 7'h4f);
  assign p1_or_132854_comb = p1_prod__273_comb | 32'h0000_0080;
  assign p1_or_132855_comb = p1_prod__279_comb | 32'h0000_0080;
  assign p1_smul_57528_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__37_squeezed_comb, 7'h4f);
  assign p1_smul_57530_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__38_squeezed_comb, 7'h31);
  assign p1_or_132860_comb = p1_prod__299_comb | 32'h0000_0080;
  assign p1_or_132861_comb = p1_prod__325_comb | 32'h0000_0080;
  assign p1_smul_57536_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__41_squeezed_comb, 7'h31);
  assign p1_smul_57538_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__42_squeezed_comb, 7'h4f);
  assign p1_or_132866_comb = p1_prod__337_comb | 32'h0000_0080;
  assign p1_or_132867_comb = p1_prod__343_comb | 32'h0000_0080;
  assign p1_smul_57544_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__45_squeezed_comb, 7'h4f);
  assign p1_smul_57546_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__46_squeezed_comb, 7'h31);
  assign p1_or_132872_comb = p1_prod__363_comb | 32'h0000_0080;
  assign p1_or_132873_comb = p1_prod__141_comb | 32'h0000_0080;
  assign p1_or_132874_comb = p1_prod__152_comb | 32'h0000_0080;
  assign p1_or_132875_comb = p1_prod__159_comb | 32'h0000_0080;
  assign p1_or_132876_comb = p1_prod__172_comb | 32'h0000_0080;
  assign p1_or_132877_comb = p1_prod__205_comb | 32'h0000_0080;
  assign p1_or_132878_comb = p1_prod__216_comb | 32'h0000_0080;
  assign p1_or_132879_comb = p1_prod__223_comb | 32'h0000_0080;
  assign p1_or_132880_comb = p1_prod__236_comb | 32'h0000_0080;
  assign p1_or_132881_comb = p1_prod__269_comb | 32'h0000_0080;
  assign p1_or_132882_comb = p1_prod__280_comb | 32'h0000_0080;
  assign p1_or_132883_comb = p1_prod__287_comb | 32'h0000_0080;
  assign p1_or_132884_comb = p1_prod__300_comb | 32'h0000_0080;
  assign p1_or_132885_comb = p1_prod__333_comb | 32'h0000_0080;
  assign p1_or_132886_comb = p1_prod__344_comb | 32'h0000_0080;
  assign p1_or_132887_comb = p1_prod__351_comb | 32'h0000_0080;
  assign p1_or_132888_comb = p1_prod__364_comb | 32'h0000_0080;
  assign p1_or_132889_comb = p1_prod__148_comb | 32'h0000_0080;
  assign p1_or_132890_comb = p1_prod__161_comb | 32'h0000_0080;
  assign p1_or_132891_comb = p1_prod__179_comb | 32'h0000_0080;
  assign p1_or_132892_comb = p1_prod__186_comb | 32'h0000_0080;
  assign p1_or_132893_comb = p1_prod__212_comb | 32'h0000_0080;
  assign p1_or_132894_comb = p1_prod__225_comb | 32'h0000_0080;
  assign p1_or_132895_comb = p1_prod__243_comb | 32'h0000_0080;
  assign p1_or_132896_comb = p1_prod__250_comb | 32'h0000_0080;
  assign p1_or_132897_comb = p1_prod__276_comb | 32'h0000_0080;
  assign p1_or_132898_comb = p1_prod__289_comb | 32'h0000_0080;
  assign p1_or_132899_comb = p1_prod__307_comb | 32'h0000_0080;
  assign p1_or_132900_comb = p1_prod__314_comb | 32'h0000_0080;
  assign p1_or_132901_comb = p1_prod__340_comb | 32'h0000_0080;
  assign p1_or_132902_comb = p1_prod__353_comb | 32'h0000_0080;
  assign p1_or_132903_comb = p1_prod__371_comb | 32'h0000_0080;
  assign p1_or_132904_comb = p1_prod__378_comb | 32'h0000_0080;
  assign p1_smul_57998_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__16_squeezed_comb, 7'h31);
  assign p1_or_132907_comb = p1_prod__162_comb | 32'h0000_0080;
  assign p1_smul_58002_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__18_squeezed_comb, 7'h31);
  assign p1_or_132910_comb = p1_prod__175_comb | 32'h0000_0080;
  assign p1_or_132911_comb = p1_prod__180_comb | 32'h0000_0080;
  assign p1_smul_58008_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__21_squeezed_comb, 7'h31);
  assign p1_or_132914_comb = p1_prod__187_comb | 32'h0000_0080;
  assign p1_smul_58012_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__23_squeezed_comb, 7'h31);
  assign p1_smul_58014_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__24_squeezed_comb, 7'h31);
  assign p1_or_132919_comb = p1_prod__226_comb | 32'h0000_0080;
  assign p1_smul_58018_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__26_squeezed_comb, 7'h31);
  assign p1_or_132922_comb = p1_prod__239_comb | 32'h0000_0080;
  assign p1_or_132923_comb = p1_prod__244_comb | 32'h0000_0080;
  assign p1_smul_58024_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__29_squeezed_comb, 7'h31);
  assign p1_or_132926_comb = p1_prod__251_comb | 32'h0000_0080;
  assign p1_smul_58028_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__31_squeezed_comb, 7'h31);
  assign p1_smul_58030_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__32_squeezed_comb, 7'h31);
  assign p1_or_132931_comb = p1_prod__290_comb | 32'h0000_0080;
  assign p1_smul_58034_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__34_squeezed_comb, 7'h31);
  assign p1_or_132934_comb = p1_prod__303_comb | 32'h0000_0080;
  assign p1_or_132935_comb = p1_prod__308_comb | 32'h0000_0080;
  assign p1_smul_58040_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__37_squeezed_comb, 7'h31);
  assign p1_or_132938_comb = p1_prod__315_comb | 32'h0000_0080;
  assign p1_smul_58044_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__39_squeezed_comb, 7'h31);
  assign p1_smul_58046_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__40_squeezed_comb, 7'h31);
  assign p1_or_132943_comb = p1_prod__354_comb | 32'h0000_0080;
  assign p1_smul_58050_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__42_squeezed_comb, 7'h31);
  assign p1_or_132946_comb = p1_prod__367_comb | 32'h0000_0080;
  assign p1_or_132947_comb = p1_prod__372_comb | 32'h0000_0080;
  assign p1_smul_58056_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__45_squeezed_comb, 7'h31);
  assign p1_or_132950_comb = p1_prod__379_comb | 32'h0000_0080;
  assign p1_smul_58060_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__47_squeezed_comb, 7'h31);
  assign p1_or_132953_comb = p1_prod__163_comb | 32'h0000_0080;
  assign p1_or_132954_comb = p1_prod__170_comb | 32'h0000_0080;
  assign p1_or_132955_comb = p1_prod__190_comb | 32'h0000_0080;
  assign p1_or_132956_comb = p1_prod__191_comb | 32'h0000_0080;
  assign p1_or_132957_comb = p1_prod__227_comb | 32'h0000_0080;
  assign p1_or_132958_comb = p1_prod__234_comb | 32'h0000_0080;
  assign p1_or_132959_comb = p1_prod__254_comb | 32'h0000_0080;
  assign p1_or_132960_comb = p1_prod__255_comb | 32'h0000_0080;
  assign p1_or_132961_comb = p1_prod__291_comb | 32'h0000_0080;
  assign p1_or_132962_comb = p1_prod__298_comb | 32'h0000_0080;
  assign p1_or_132963_comb = p1_prod__318_comb | 32'h0000_0080;
  assign p1_or_132964_comb = p1_prod__319_comb | 32'h0000_0080;
  assign p1_or_132965_comb = p1_prod__355_comb | 32'h0000_0080;
  assign p1_or_132966_comb = p1_prod__362_comb | 32'h0000_0080;
  assign p1_or_132967_comb = p1_prod__382_comb | 32'h0000_0080;
  assign p1_or_132968_comb = p1_prod__383_comb | 32'h0000_0080;
  assign p1_or_133017_comb = p1_prod__10_comb | 32'h0000_0080;
  assign p1_or_133018_comb = p1_prod__11_comb | 32'h0000_0080;
  assign p1_or_133019_comb = p1_prod__12_comb | 32'h0000_0080;
  assign p1_or_133020_comb = p1_prod__13_comb | 32'h0000_0080;
  assign p1_or_133021_comb = p1_prod__455_comb | 32'h0000_0080;
  assign p1_or_133022_comb = p1_prod__459_comb | 32'h0000_0080;
  assign p1_or_133023_comb = p1_prod__464_comb | 32'h0000_0080;
  assign p1_or_133024_comb = p1_prod__470_comb | 32'h0000_0080;
  assign p1_or_133025_comb = p1_prod__16_comb | 32'h0000_0080;
  assign p1_smul_57456_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__1_squeezed_comb, 7'h31);
  assign p1_smul_57458_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__2_squeezed_comb, 7'h4f);
  assign p1_or_133030_comb = p1_prod__19_comb | 32'h0000_0080;
  assign p1_or_133031_comb = p1_prod__20_comb | 32'h0000_0080;
  assign p1_smul_57464_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__5_squeezed_comb, 7'h4f);
  assign p1_smul_57466_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__6_squeezed_comb, 7'h31);
  assign p1_or_133036_comb = p1_prod__23_comb | 32'h0000_0080;
  assign p1_or_133037_comb = p1_prod__453_comb | 32'h0000_0080;
  assign p1_smul_57568_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__57_squeezed_comb, 7'h31);
  assign p1_smul_57570_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__58_squeezed_comb, 7'h4f);
  assign p1_or_133042_comb = p1_prod__465_comb | 32'h0000_0080;
  assign p1_or_133043_comb = p1_prod__471_comb | 32'h0000_0080;
  assign p1_smul_57576_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__61_squeezed_comb, 7'h4f);
  assign p1_smul_57578_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__62_squeezed_comb, 7'h31);
  assign p1_or_133048_comb = p1_prod__491_comb | 32'h0000_0080;
  assign p1_or_133049_comb = p1_prod__25_comb | 32'h0000_0080;
  assign p1_or_133050_comb = p1_prod__27_comb | 32'h0000_0080;
  assign p1_or_133051_comb = p1_prod__28_comb | 32'h0000_0080;
  assign p1_or_133052_comb = p1_prod__30_comb | 32'h0000_0080;
  assign p1_or_133053_comb = p1_prod__461_comb | 32'h0000_0080;
  assign p1_or_133054_comb = p1_prod__472_comb | 32'h0000_0080;
  assign p1_or_133055_comb = p1_prod__479_comb | 32'h0000_0080;
  assign p1_or_133056_comb = p1_prod__492_comb | 32'h0000_0080;
  assign p1_or_133057_comb = p1_prod__40_comb | 32'h0000_0080;
  assign p1_or_133058_comb = p1_prod__42_comb | 32'h0000_0080;
  assign p1_or_133059_comb = p1_prod__45_comb | 32'h0000_0080;
  assign p1_or_133060_comb = p1_prod__47_comb | 32'h0000_0080;
  assign p1_or_133061_comb = p1_prod__468_comb | 32'h0000_0080;
  assign p1_or_133062_comb = p1_prod__481_comb | 32'h0000_0080;
  assign p1_or_133063_comb = p1_prod__499_comb | 32'h0000_0080;
  assign p1_or_133064_comb = p1_prod__506_comb | 32'h0000_0080;
  assign p1_smul_57966_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted_squeezed_comb, 7'h31);
  assign p1_or_133067_comb = p1_prod__49_comb | 32'h0000_0080;
  assign p1_smul_57970_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__2_squeezed_comb, 7'h31);
  assign p1_or_133070_comb = p1_prod__51_comb | 32'h0000_0080;
  assign p1_or_133071_comb = p1_prod__52_comb | 32'h0000_0080;
  assign p1_smul_57976_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__5_squeezed_comb, 7'h31);
  assign p1_or_133074_comb = p1_prod__54_comb | 32'h0000_0080;
  assign p1_smul_57980_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__7_squeezed_comb, 7'h31);
  assign p1_smul_58078_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__56_squeezed_comb, 7'h31);
  assign p1_or_133079_comb = p1_prod__482_comb | 32'h0000_0080;
  assign p1_smul_58082_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__58_squeezed_comb, 7'h31);
  assign p1_or_133082_comb = p1_prod__495_comb | 32'h0000_0080;
  assign p1_or_133083_comb = p1_prod__500_comb | 32'h0000_0080;
  assign p1_smul_58088_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__61_squeezed_comb, 7'h31);
  assign p1_or_133086_comb = p1_prod__507_comb | 32'h0000_0080;
  assign p1_smul_58092_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__63_squeezed_comb, 7'h31);
  assign p1_or_133089_comb = p1_prod__56_comb | 32'h0000_0080;
  assign p1_or_133090_comb = p1_prod__57_comb | 32'h0000_0080;
  assign p1_or_133091_comb = p1_prod__62_comb | 32'h0000_0080;
  assign p1_or_133092_comb = p1_prod__63_comb | 32'h0000_0080;
  assign p1_or_133093_comb = p1_prod__483_comb | 32'h0000_0080;
  assign p1_or_133094_comb = p1_prod__490_comb | 32'h0000_0080;
  assign p1_or_133095_comb = p1_prod__510_comb | 32'h0000_0080;
  assign p1_or_133096_comb = p1_prod__511_comb | 32'h0000_0080;
  assign p1_or_133145_comb = p1_prod__71_comb | 32'h0000_0080;
  assign p1_or_133146_comb = p1_prod__75_comb | 32'h0000_0080;
  assign p1_or_133147_comb = p1_prod__80_comb | 32'h0000_0080;
  assign p1_or_133148_comb = p1_prod__86_comb | 32'h0000_0080;
  assign p1_or_133149_comb = p1_prod__391_comb | 32'h0000_0080;
  assign p1_or_133150_comb = p1_prod__395_comb | 32'h0000_0080;
  assign p1_or_133151_comb = p1_prod__400_comb | 32'h0000_0080;
  assign p1_or_133152_comb = p1_prod__406_comb | 32'h0000_0080;
  assign p1_or_133153_comb = p1_prod__69_comb | 32'h0000_0080;
  assign p1_smul_57472_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__9_squeezed_comb, 7'h31);
  assign p1_smul_57474_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__10_squeezed_comb, 7'h4f);
  assign p1_or_133158_comb = p1_prod__81_comb | 32'h0000_0080;
  assign p1_or_133159_comb = p1_prod__87_comb | 32'h0000_0080;
  assign p1_smul_57480_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__13_squeezed_comb, 7'h4f);
  assign p1_smul_57482_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__14_squeezed_comb, 7'h31);
  assign p1_or_133164_comb = p1_prod__107_comb | 32'h0000_0080;
  assign p1_or_133165_comb = p1_prod__389_comb | 32'h0000_0080;
  assign p1_smul_57552_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__49_squeezed_comb, 7'h31);
  assign p1_smul_57554_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__50_squeezed_comb, 7'h4f);
  assign p1_or_133170_comb = p1_prod__401_comb | 32'h0000_0080;
  assign p1_or_133171_comb = p1_prod__407_comb | 32'h0000_0080;
  assign p1_smul_57560_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__53_squeezed_comb, 7'h4f);
  assign p1_smul_57562_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__54_squeezed_comb, 7'h31);
  assign p1_or_133176_comb = p1_prod__427_comb | 32'h0000_0080;
  assign p1_or_133177_comb = p1_prod__77_comb | 32'h0000_0080;
  assign p1_or_133178_comb = p1_prod__88_comb | 32'h0000_0080;
  assign p1_or_133179_comb = p1_prod__95_comb | 32'h0000_0080;
  assign p1_or_133180_comb = p1_prod__108_comb | 32'h0000_0080;
  assign p1_or_133181_comb = p1_prod__397_comb | 32'h0000_0080;
  assign p1_or_133182_comb = p1_prod__408_comb | 32'h0000_0080;
  assign p1_or_133183_comb = p1_prod__415_comb | 32'h0000_0080;
  assign p1_or_133184_comb = p1_prod__428_comb | 32'h0000_0080;
  assign p1_or_133185_comb = p1_prod__84_comb | 32'h0000_0080;
  assign p1_or_133186_comb = p1_prod__97_comb | 32'h0000_0080;
  assign p1_or_133187_comb = p1_prod__115_comb | 32'h0000_0080;
  assign p1_or_133188_comb = p1_prod__122_comb | 32'h0000_0080;
  assign p1_or_133189_comb = p1_prod__404_comb | 32'h0000_0080;
  assign p1_or_133190_comb = p1_prod__417_comb | 32'h0000_0080;
  assign p1_or_133191_comb = p1_prod__435_comb | 32'h0000_0080;
  assign p1_or_133192_comb = p1_prod__442_comb | 32'h0000_0080;
  assign p1_smul_57982_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__8_squeezed_comb, 7'h31);
  assign p1_or_133195_comb = p1_prod__98_comb | 32'h0000_0080;
  assign p1_smul_57986_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__10_squeezed_comb, 7'h31);
  assign p1_or_133198_comb = p1_prod__111_comb | 32'h0000_0080;
  assign p1_or_133199_comb = p1_prod__116_comb | 32'h0000_0080;
  assign p1_smul_57992_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__13_squeezed_comb, 7'h31);
  assign p1_or_133202_comb = p1_prod__123_comb | 32'h0000_0080;
  assign p1_smul_57996_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__15_squeezed_comb, 7'h31);
  assign p1_smul_58062_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__48_squeezed_comb, 7'h31);
  assign p1_or_133207_comb = p1_prod__418_comb | 32'h0000_0080;
  assign p1_smul_58066_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__50_squeezed_comb, 7'h31);
  assign p1_or_133210_comb = p1_prod__431_comb | 32'h0000_0080;
  assign p1_or_133211_comb = p1_prod__436_comb | 32'h0000_0080;
  assign p1_smul_58072_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__53_squeezed_comb, 7'h31);
  assign p1_or_133214_comb = p1_prod__443_comb | 32'h0000_0080;
  assign p1_smul_58076_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__55_squeezed_comb, 7'h31);
  assign p1_or_133217_comb = p1_prod__99_comb | 32'h0000_0080;
  assign p1_or_133218_comb = p1_prod__106_comb | 32'h0000_0080;
  assign p1_or_133219_comb = p1_prod__126_comb | 32'h0000_0080;
  assign p1_or_133220_comb = p1_prod__127_comb | 32'h0000_0080;
  assign p1_or_133221_comb = p1_prod__419_comb | 32'h0000_0080;
  assign p1_or_133222_comb = p1_prod__426_comb | 32'h0000_0080;
  assign p1_or_133223_comb = p1_prod__446_comb | 32'h0000_0080;
  assign p1_or_133224_comb = p1_prod__447_comb | 32'h0000_0080;
  assign p1_sel_133225_comb = $signed(p1_shifted__16_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__16_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__16_squeezed_comb, p1_smul_57326_TrailingBits___16_comb};
  assign p1_sel_133226_comb = $signed(p1_shifted__17_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__17_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__17_squeezed_comb, p1_smul_57326_TrailingBits___17_comb};
  assign p1_sel_133227_comb = $signed(p1_shifted__18_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__18_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__18_squeezed_comb, p1_smul_57326_TrailingBits___18_comb};
  assign p1_sel_133228_comb = $signed(p1_shifted__19_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__19_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__19_squeezed_comb, p1_smul_57326_TrailingBits___19_comb};
  assign p1_sel_133229_comb = $signed(p1_shifted__20_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__20_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__20_squeezed_comb, p1_smul_57326_TrailingBits___20_comb};
  assign p1_sel_133230_comb = $signed(p1_shifted__21_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__21_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__21_squeezed_comb, p1_smul_57326_TrailingBits___21_comb};
  assign p1_sel_133231_comb = $signed(p1_shifted__22_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__22_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__22_squeezed_comb, p1_smul_57326_TrailingBits___22_comb};
  assign p1_sel_133232_comb = $signed(p1_shifted__23_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__23_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__23_squeezed_comb, p1_smul_57326_TrailingBits___23_comb};
  assign p1_sel_133233_comb = $signed(p1_shifted__24_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__24_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__24_squeezed_comb, p1_smul_57326_TrailingBits___24_comb};
  assign p1_sel_133234_comb = $signed(p1_shifted__25_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__25_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__25_squeezed_comb, p1_smul_57326_TrailingBits___25_comb};
  assign p1_sel_133235_comb = $signed(p1_shifted__26_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__26_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__26_squeezed_comb, p1_smul_57326_TrailingBits___26_comb};
  assign p1_sel_133236_comb = $signed(p1_shifted__27_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__27_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__27_squeezed_comb, p1_smul_57326_TrailingBits___27_comb};
  assign p1_sel_133237_comb = $signed(p1_shifted__28_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__28_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__28_squeezed_comb, p1_smul_57326_TrailingBits___28_comb};
  assign p1_sel_133238_comb = $signed(p1_shifted__29_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__29_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__29_squeezed_comb, p1_smul_57326_TrailingBits___29_comb};
  assign p1_sel_133239_comb = $signed(p1_shifted__30_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__30_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__30_squeezed_comb, p1_smul_57326_TrailingBits___30_comb};
  assign p1_sel_133240_comb = $signed(p1_shifted__31_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__31_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__31_squeezed_comb, p1_smul_57326_TrailingBits___31_comb};
  assign p1_sel_133241_comb = $signed(p1_shifted__32_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__32_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__32_squeezed_comb, p1_smul_57326_TrailingBits___32_comb};
  assign p1_sel_133242_comb = $signed(p1_shifted__33_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__33_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__33_squeezed_comb, p1_smul_57326_TrailingBits___33_comb};
  assign p1_sel_133243_comb = $signed(p1_shifted__34_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__34_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__34_squeezed_comb, p1_smul_57326_TrailingBits___34_comb};
  assign p1_sel_133244_comb = $signed(p1_shifted__35_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__35_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__35_squeezed_comb, p1_smul_57326_TrailingBits___35_comb};
  assign p1_sel_133245_comb = $signed(p1_shifted__36_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__36_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__36_squeezed_comb, p1_smul_57326_TrailingBits___36_comb};
  assign p1_sel_133246_comb = $signed(p1_shifted__37_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__37_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__37_squeezed_comb, p1_smul_57326_TrailingBits___37_comb};
  assign p1_sel_133247_comb = $signed(p1_shifted__38_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__38_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__38_squeezed_comb, p1_smul_57326_TrailingBits___38_comb};
  assign p1_sel_133248_comb = $signed(p1_shifted__39_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__39_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__39_squeezed_comb, p1_smul_57326_TrailingBits___39_comb};
  assign p1_sel_133249_comb = $signed(p1_shifted__40_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__40_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__40_squeezed_comb, p1_smul_57326_TrailingBits___40_comb};
  assign p1_sel_133250_comb = $signed(p1_shifted__41_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__41_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__41_squeezed_comb, p1_smul_57326_TrailingBits___41_comb};
  assign p1_sel_133251_comb = $signed(p1_shifted__42_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__42_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__42_squeezed_comb, p1_smul_57326_TrailingBits___42_comb};
  assign p1_sel_133252_comb = $signed(p1_shifted__43_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__43_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__43_squeezed_comb, p1_smul_57326_TrailingBits___43_comb};
  assign p1_sel_133253_comb = $signed(p1_shifted__44_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__44_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__44_squeezed_comb, p1_smul_57326_TrailingBits___44_comb};
  assign p1_sel_133254_comb = $signed(p1_shifted__45_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__45_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__45_squeezed_comb, p1_smul_57326_TrailingBits___45_comb};
  assign p1_sel_133255_comb = $signed(p1_shifted__46_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__46_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__46_squeezed_comb, p1_smul_57326_TrailingBits___46_comb};
  assign p1_sel_133256_comb = $signed(p1_shifted__47_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__47_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__47_squeezed_comb, p1_smul_57326_TrailingBits___47_comb};
  assign p1_concat_133325_comb = {p1_smul_57488_NarrowedMult__comb, 1'h0};
  assign p1_concat_133327_comb = {p1_smul_57490_NarrowedMult__comb, 1'h0};
  assign p1_concat_133337_comb = {p1_smul_57496_NarrowedMult__comb, 1'h0};
  assign p1_concat_133339_comb = {p1_smul_57498_NarrowedMult__comb, 1'h0};
  assign p1_concat_133349_comb = {p1_smul_57504_NarrowedMult__comb, 1'h0};
  assign p1_concat_133351_comb = {p1_smul_57506_NarrowedMult__comb, 1'h0};
  assign p1_concat_133361_comb = {p1_smul_57512_NarrowedMult__comb, 1'h0};
  assign p1_concat_133363_comb = {p1_smul_57514_NarrowedMult__comb, 1'h0};
  assign p1_concat_133373_comb = {p1_smul_57520_NarrowedMult__comb, 1'h0};
  assign p1_concat_133375_comb = {p1_smul_57522_NarrowedMult__comb, 1'h0};
  assign p1_concat_133385_comb = {p1_smul_57528_NarrowedMult__comb, 1'h0};
  assign p1_concat_133387_comb = {p1_smul_57530_NarrowedMult__comb, 1'h0};
  assign p1_concat_133397_comb = {p1_smul_57536_NarrowedMult__comb, 1'h0};
  assign p1_concat_133399_comb = {p1_smul_57538_NarrowedMult__comb, 1'h0};
  assign p1_concat_133409_comb = {p1_smul_57544_NarrowedMult__comb, 1'h0};
  assign p1_concat_133411_comb = {p1_smul_57546_NarrowedMult__comb, 1'h0};
  assign p1_concat_133545_comb = {p1_smul_57998_NarrowedMult__comb, 1'h0};
  assign p1_concat_133551_comb = {p1_smul_58002_NarrowedMult__comb, 1'h0};
  assign p1_concat_133561_comb = {p1_smul_58008_NarrowedMult__comb, 1'h0};
  assign p1_concat_133567_comb = {p1_smul_58012_NarrowedMult__comb, 1'h0};
  assign p1_concat_133569_comb = {p1_smul_58014_NarrowedMult__comb, 1'h0};
  assign p1_concat_133575_comb = {p1_smul_58018_NarrowedMult__comb, 1'h0};
  assign p1_concat_133585_comb = {p1_smul_58024_NarrowedMult__comb, 1'h0};
  assign p1_concat_133591_comb = {p1_smul_58028_NarrowedMult__comb, 1'h0};
  assign p1_concat_133593_comb = {p1_smul_58030_NarrowedMult__comb, 1'h0};
  assign p1_concat_133599_comb = {p1_smul_58034_NarrowedMult__comb, 1'h0};
  assign p1_concat_133609_comb = {p1_smul_58040_NarrowedMult__comb, 1'h0};
  assign p1_concat_133615_comb = {p1_smul_58044_NarrowedMult__comb, 1'h0};
  assign p1_concat_133617_comb = {p1_smul_58046_NarrowedMult__comb, 1'h0};
  assign p1_concat_133623_comb = {p1_smul_58050_NarrowedMult__comb, 1'h0};
  assign p1_concat_133633_comb = {p1_smul_58056_NarrowedMult__comb, 1'h0};
  assign p1_concat_133639_comb = {p1_smul_58060_NarrowedMult__comb, 1'h0};
  assign p1_sel_133705_comb = $signed(p1_shifted_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted_squeezed_comb, p1_smul_57326_TrailingBits__comb};
  assign p1_sel_133706_comb = $signed(p1_shifted__1_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__1_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__1_squeezed_comb, p1_smul_57326_TrailingBits___1_comb};
  assign p1_sel_133707_comb = $signed(p1_shifted__2_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__2_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__2_squeezed_comb, p1_smul_57326_TrailingBits___2_comb};
  assign p1_sel_133708_comb = $signed(p1_shifted__3_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__3_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__3_squeezed_comb, p1_smul_57326_TrailingBits___3_comb};
  assign p1_sel_133709_comb = $signed(p1_shifted__4_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__4_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__4_squeezed_comb, p1_smul_57326_TrailingBits___4_comb};
  assign p1_sel_133710_comb = $signed(p1_shifted__5_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__5_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__5_squeezed_comb, p1_smul_57326_TrailingBits___5_comb};
  assign p1_sel_133711_comb = $signed(p1_shifted__6_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__6_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__6_squeezed_comb, p1_smul_57326_TrailingBits___6_comb};
  assign p1_sel_133712_comb = $signed(p1_shifted__7_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__7_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__7_squeezed_comb, p1_smul_57326_TrailingBits___7_comb};
  assign p1_sel_133713_comb = $signed(p1_shifted__56_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__56_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__56_squeezed_comb, p1_smul_57326_TrailingBits___56_comb};
  assign p1_sel_133714_comb = $signed(p1_shifted__57_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__57_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__57_squeezed_comb, p1_smul_57326_TrailingBits___57_comb};
  assign p1_sel_133715_comb = $signed(p1_shifted__58_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__58_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__58_squeezed_comb, p1_smul_57326_TrailingBits___58_comb};
  assign p1_sel_133716_comb = $signed(p1_shifted__59_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__59_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__59_squeezed_comb, p1_smul_57326_TrailingBits___59_comb};
  assign p1_sel_133717_comb = $signed(p1_shifted__60_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__60_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__60_squeezed_comb, p1_smul_57326_TrailingBits___60_comb};
  assign p1_sel_133718_comb = $signed(p1_shifted__61_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__61_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__61_squeezed_comb, p1_smul_57326_TrailingBits___61_comb};
  assign p1_sel_133719_comb = $signed(p1_shifted__62_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__62_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__62_squeezed_comb, p1_smul_57326_TrailingBits___62_comb};
  assign p1_sel_133720_comb = $signed(p1_shifted__63_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__63_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__63_squeezed_comb, p1_smul_57326_TrailingBits___63_comb};
  assign p1_concat_133757_comb = {p1_smul_57456_NarrowedMult__comb, 1'h0};
  assign p1_concat_133759_comb = {p1_smul_57458_NarrowedMult__comb, 1'h0};
  assign p1_concat_133769_comb = {p1_smul_57464_NarrowedMult__comb, 1'h0};
  assign p1_concat_133771_comb = {p1_smul_57466_NarrowedMult__comb, 1'h0};
  assign p1_concat_133781_comb = {p1_smul_57568_NarrowedMult__comb, 1'h0};
  assign p1_concat_133783_comb = {p1_smul_57570_NarrowedMult__comb, 1'h0};
  assign p1_concat_133793_comb = {p1_smul_57576_NarrowedMult__comb, 1'h0};
  assign p1_concat_133795_comb = {p1_smul_57578_NarrowedMult__comb, 1'h0};
  assign p1_concat_133865_comb = {p1_smul_57966_NarrowedMult__comb, 1'h0};
  assign p1_concat_133871_comb = {p1_smul_57970_NarrowedMult__comb, 1'h0};
  assign p1_concat_133881_comb = {p1_smul_57976_NarrowedMult__comb, 1'h0};
  assign p1_concat_133887_comb = {p1_smul_57980_NarrowedMult__comb, 1'h0};
  assign p1_concat_133889_comb = {p1_smul_58078_NarrowedMult__comb, 1'h0};
  assign p1_concat_133895_comb = {p1_smul_58082_NarrowedMult__comb, 1'h0};
  assign p1_concat_133905_comb = {p1_smul_58088_NarrowedMult__comb, 1'h0};
  assign p1_concat_133911_comb = {p1_smul_58092_NarrowedMult__comb, 1'h0};
  assign p1_sel_133945_comb = $signed(p1_shifted__8_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__8_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__8_squeezed_comb, p1_smul_57326_TrailingBits___8_comb};
  assign p1_sel_133946_comb = $signed(p1_shifted__9_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__9_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__9_squeezed_comb, p1_smul_57326_TrailingBits___9_comb};
  assign p1_sel_133947_comb = $signed(p1_shifted__10_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__10_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__10_squeezed_comb, p1_smul_57326_TrailingBits___10_comb};
  assign p1_sel_133948_comb = $signed(p1_shifted__11_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__11_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__11_squeezed_comb, p1_smul_57326_TrailingBits___11_comb};
  assign p1_sel_133949_comb = $signed(p1_shifted__12_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__12_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__12_squeezed_comb, p1_smul_57326_TrailingBits___12_comb};
  assign p1_sel_133950_comb = $signed(p1_shifted__13_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__13_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__13_squeezed_comb, p1_smul_57326_TrailingBits___13_comb};
  assign p1_sel_133951_comb = $signed(p1_shifted__14_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__14_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__14_squeezed_comb, p1_smul_57326_TrailingBits___14_comb};
  assign p1_sel_133952_comb = $signed(p1_shifted__15_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__15_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__15_squeezed_comb, p1_smul_57326_TrailingBits___15_comb};
  assign p1_sel_133953_comb = $signed(p1_shifted__48_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__48_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__48_squeezed_comb, p1_smul_57326_TrailingBits___48_comb};
  assign p1_sel_133954_comb = $signed(p1_shifted__49_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__49_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__49_squeezed_comb, p1_smul_57326_TrailingBits___49_comb};
  assign p1_sel_133955_comb = $signed(p1_shifted__50_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__50_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__50_squeezed_comb, p1_smul_57326_TrailingBits___50_comb};
  assign p1_sel_133956_comb = $signed(p1_shifted__51_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__51_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__51_squeezed_comb, p1_smul_57326_TrailingBits___51_comb};
  assign p1_sel_133957_comb = $signed(p1_shifted__52_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__52_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__52_squeezed_comb, p1_smul_57326_TrailingBits___52_comb};
  assign p1_sel_133958_comb = $signed(p1_shifted__53_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__53_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__53_squeezed_comb, p1_smul_57326_TrailingBits___53_comb};
  assign p1_sel_133959_comb = $signed(p1_shifted__54_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__54_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__54_squeezed_comb, p1_smul_57326_TrailingBits___54_comb};
  assign p1_sel_133960_comb = $signed(p1_shifted__55_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__55_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__55_squeezed_comb, p1_smul_57326_TrailingBits___55_comb};
  assign p1_concat_133997_comb = {p1_smul_57472_NarrowedMult__comb, 1'h0};
  assign p1_concat_133999_comb = {p1_smul_57474_NarrowedMult__comb, 1'h0};
  assign p1_concat_134009_comb = {p1_smul_57480_NarrowedMult__comb, 1'h0};
  assign p1_concat_134011_comb = {p1_smul_57482_NarrowedMult__comb, 1'h0};
  assign p1_concat_134021_comb = {p1_smul_57552_NarrowedMult__comb, 1'h0};
  assign p1_concat_134023_comb = {p1_smul_57554_NarrowedMult__comb, 1'h0};
  assign p1_concat_134033_comb = {p1_smul_57560_NarrowedMult__comb, 1'h0};
  assign p1_concat_134035_comb = {p1_smul_57562_NarrowedMult__comb, 1'h0};
  assign p1_concat_134105_comb = {p1_smul_57982_NarrowedMult__comb, 1'h0};
  assign p1_concat_134111_comb = {p1_smul_57986_NarrowedMult__comb, 1'h0};
  assign p1_concat_134121_comb = {p1_smul_57992_NarrowedMult__comb, 1'h0};
  assign p1_concat_134127_comb = {p1_smul_57996_NarrowedMult__comb, 1'h0};
  assign p1_concat_134129_comb = {p1_smul_58062_NarrowedMult__comb, 1'h0};
  assign p1_concat_134135_comb = {p1_smul_58066_NarrowedMult__comb, 1'h0};
  assign p1_concat_134145_comb = {p1_smul_58072_NarrowedMult__comb, 1'h0};
  assign p1_concat_134151_comb = {p1_smul_58076_NarrowedMult__comb, 1'h0};
  assign p1_add_135145_comb = {{1{p1_sel_133225_comb[15]}}, p1_sel_133225_comb} + {{1{p1_sel_133226_comb[15]}}, p1_sel_133226_comb};
  assign p1_add_135146_comb = {{1{p1_sel_133227_comb[15]}}, p1_sel_133227_comb} + {{1{p1_sel_133228_comb[15]}}, p1_sel_133228_comb};
  assign p1_add_135147_comb = {{1{p1_sel_133229_comb[15]}}, p1_sel_133229_comb} + {{1{p1_sel_133230_comb[15]}}, p1_sel_133230_comb};
  assign p1_add_135148_comb = {{1{p1_sel_133231_comb[15]}}, p1_sel_133231_comb} + {{1{p1_sel_133232_comb[15]}}, p1_sel_133232_comb};
  assign p1_add_135149_comb = {{1{p1_sel_133233_comb[15]}}, p1_sel_133233_comb} + {{1{p1_sel_133234_comb[15]}}, p1_sel_133234_comb};
  assign p1_add_135150_comb = {{1{p1_sel_133235_comb[15]}}, p1_sel_133235_comb} + {{1{p1_sel_133236_comb[15]}}, p1_sel_133236_comb};
  assign p1_add_135151_comb = {{1{p1_sel_133237_comb[15]}}, p1_sel_133237_comb} + {{1{p1_sel_133238_comb[15]}}, p1_sel_133238_comb};
  assign p1_add_135152_comb = {{1{p1_sel_133239_comb[15]}}, p1_sel_133239_comb} + {{1{p1_sel_133240_comb[15]}}, p1_sel_133240_comb};
  assign p1_add_135153_comb = {{1{p1_sel_133241_comb[15]}}, p1_sel_133241_comb} + {{1{p1_sel_133242_comb[15]}}, p1_sel_133242_comb};
  assign p1_add_135154_comb = {{1{p1_sel_133243_comb[15]}}, p1_sel_133243_comb} + {{1{p1_sel_133244_comb[15]}}, p1_sel_133244_comb};
  assign p1_add_135155_comb = {{1{p1_sel_133245_comb[15]}}, p1_sel_133245_comb} + {{1{p1_sel_133246_comb[15]}}, p1_sel_133246_comb};
  assign p1_add_135156_comb = {{1{p1_sel_133247_comb[15]}}, p1_sel_133247_comb} + {{1{p1_sel_133248_comb[15]}}, p1_sel_133248_comb};
  assign p1_add_135157_comb = {{1{p1_sel_133249_comb[15]}}, p1_sel_133249_comb} + {{1{p1_sel_133250_comb[15]}}, p1_sel_133250_comb};
  assign p1_add_135158_comb = {{1{p1_sel_133251_comb[15]}}, p1_sel_133251_comb} + {{1{p1_sel_133252_comb[15]}}, p1_sel_133252_comb};
  assign p1_add_135159_comb = {{1{p1_sel_133253_comb[15]}}, p1_sel_133253_comb} + {{1{p1_sel_133254_comb[15]}}, p1_sel_133254_comb};
  assign p1_add_135160_comb = {{1{p1_sel_133255_comb[15]}}, p1_sel_133255_comb} + {{1{p1_sel_133256_comb[15]}}, p1_sel_133256_comb};
  assign p1_smul_135161_comb = smul16b_8b_x_9b(p1_shifted__16_squeezed_comb, 9'h0fb);
  assign p1_smul_135162_comb = smul16b_8b_x_9b(p1_shifted__17_squeezed_comb, 9'h0d5);
  assign p1_sel_135163_comb = $signed(p1_or_132809_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132809_comb[23:9], 1'h0};
  assign p1_sel_135164_comb = $signed(p1_or_132810_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132810_comb[23:9], 1'h0};
  assign p1_sel_135165_comb = $signed(p1_or_132811_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132811_comb[23:9], 1'h0};
  assign p1_sel_135166_comb = $signed(p1_or_132812_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132812_comb[23:9], 1'h0};
  assign p1_smul_135167_comb = smul16b_8b_x_9b(p1_shifted__22_squeezed_comb, 9'h12b);
  assign p1_smul_135168_comb = smul16b_8b_x_9b(p1_shifted__23_squeezed_comb, 9'h105);
  assign p1_smul_135169_comb = smul16b_8b_x_9b(p1_shifted__24_squeezed_comb, 9'h0fb);
  assign p1_smul_135170_comb = smul16b_8b_x_9b(p1_shifted__25_squeezed_comb, 9'h0d5);
  assign p1_sel_135171_comb = $signed(p1_or_132813_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132813_comb[23:9], 1'h0};
  assign p1_sel_135172_comb = $signed(p1_or_132814_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132814_comb[23:9], 1'h0};
  assign p1_sel_135173_comb = $signed(p1_or_132815_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132815_comb[23:9], 1'h0};
  assign p1_sel_135174_comb = $signed(p1_or_132816_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132816_comb[23:9], 1'h0};
  assign p1_smul_135175_comb = smul16b_8b_x_9b(p1_shifted__30_squeezed_comb, 9'h12b);
  assign p1_smul_135176_comb = smul16b_8b_x_9b(p1_shifted__31_squeezed_comb, 9'h105);
  assign p1_smul_135177_comb = smul16b_8b_x_9b(p1_shifted__32_squeezed_comb, 9'h0fb);
  assign p1_smul_135178_comb = smul16b_8b_x_9b(p1_shifted__33_squeezed_comb, 9'h0d5);
  assign p1_sel_135179_comb = $signed(p1_or_132817_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132817_comb[23:9], 1'h0};
  assign p1_sel_135180_comb = $signed(p1_or_132818_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132818_comb[23:9], 1'h0};
  assign p1_sel_135181_comb = $signed(p1_or_132819_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132819_comb[23:9], 1'h0};
  assign p1_sel_135182_comb = $signed(p1_or_132820_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132820_comb[23:9], 1'h0};
  assign p1_smul_135183_comb = smul16b_8b_x_9b(p1_shifted__38_squeezed_comb, 9'h12b);
  assign p1_smul_135184_comb = smul16b_8b_x_9b(p1_shifted__39_squeezed_comb, 9'h105);
  assign p1_smul_135185_comb = smul16b_8b_x_9b(p1_shifted__40_squeezed_comb, 9'h0fb);
  assign p1_smul_135186_comb = smul16b_8b_x_9b(p1_shifted__41_squeezed_comb, 9'h0d5);
  assign p1_sel_135187_comb = $signed(p1_or_132821_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132821_comb[23:9], 1'h0};
  assign p1_sel_135188_comb = $signed(p1_or_132822_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132822_comb[23:9], 1'h0};
  assign p1_sel_135189_comb = $signed(p1_or_132823_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132823_comb[23:9], 1'h0};
  assign p1_sel_135190_comb = $signed(p1_or_132824_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132824_comb[23:9], 1'h0};
  assign p1_smul_135191_comb = smul16b_8b_x_9b(p1_shifted__46_squeezed_comb, 9'h12b);
  assign p1_smul_135192_comb = smul16b_8b_x_9b(p1_shifted__47_squeezed_comb, 9'h105);
  assign p1_sel_135193_comb = $signed(p1_or_132825_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132825_comb[23:10], 2'h0};
  assign p1_sel_135194_comb = $signed(p1_concat_133325_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133325_comb;
  assign p1_sel_135195_comb = $signed(p1_concat_133327_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133327_comb;
  assign p1_sel_135196_comb = $signed(p1_or_132830_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132830_comb[23:10], 2'h0};
  assign p1_sel_135197_comb = $signed(p1_or_132831_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132831_comb[23:10], 2'h0};
  assign p1_sel_135198_comb = $signed(p1_concat_133337_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133337_comb;
  assign p1_sel_135199_comb = $signed(p1_concat_133339_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133339_comb;
  assign p1_sel_135200_comb = $signed(p1_or_132836_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132836_comb[23:10], 2'h0};
  assign p1_sel_135201_comb = $signed(p1_or_132837_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132837_comb[23:10], 2'h0};
  assign p1_sel_135202_comb = $signed(p1_concat_133349_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133349_comb;
  assign p1_sel_135203_comb = $signed(p1_concat_133351_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133351_comb;
  assign p1_sel_135204_comb = $signed(p1_or_132842_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132842_comb[23:10], 2'h0};
  assign p1_sel_135205_comb = $signed(p1_or_132843_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132843_comb[23:10], 2'h0};
  assign p1_sel_135206_comb = $signed(p1_concat_133361_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133361_comb;
  assign p1_sel_135207_comb = $signed(p1_concat_133363_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133363_comb;
  assign p1_sel_135208_comb = $signed(p1_or_132848_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132848_comb[23:10], 2'h0};
  assign p1_sel_135209_comb = $signed(p1_or_132849_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132849_comb[23:10], 2'h0};
  assign p1_sel_135210_comb = $signed(p1_concat_133373_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133373_comb;
  assign p1_sel_135211_comb = $signed(p1_concat_133375_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133375_comb;
  assign p1_sel_135212_comb = $signed(p1_or_132854_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132854_comb[23:10], 2'h0};
  assign p1_sel_135213_comb = $signed(p1_or_132855_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132855_comb[23:10], 2'h0};
  assign p1_sel_135214_comb = $signed(p1_concat_133385_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133385_comb;
  assign p1_sel_135215_comb = $signed(p1_concat_133387_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133387_comb;
  assign p1_sel_135216_comb = $signed(p1_or_132860_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132860_comb[23:10], 2'h0};
  assign p1_sel_135217_comb = $signed(p1_or_132861_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132861_comb[23:10], 2'h0};
  assign p1_sel_135218_comb = $signed(p1_concat_133397_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133397_comb;
  assign p1_sel_135219_comb = $signed(p1_concat_133399_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133399_comb;
  assign p1_sel_135220_comb = $signed(p1_or_132866_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132866_comb[23:10], 2'h0};
  assign p1_sel_135221_comb = $signed(p1_or_132867_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132867_comb[23:10], 2'h0};
  assign p1_sel_135222_comb = $signed(p1_concat_133409_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133409_comb;
  assign p1_sel_135223_comb = $signed(p1_concat_133411_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133411_comb;
  assign p1_sel_135224_comb = $signed(p1_or_132872_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132872_comb[23:10], 2'h0};
  assign p1_smul_135225_comb = smul16b_8b_x_9b(p1_shifted__16_squeezed_comb, 9'h0d5);
  assign p1_sel_135226_comb = $signed(p1_or_132873_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132873_comb[23:9], 1'h0};
  assign p1_smul_135227_comb = smul16b_8b_x_9b(p1_shifted__18_squeezed_comb, 9'h105);
  assign p1_sel_135228_comb = $signed(p1_or_132874_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132874_comb[23:9], 1'h0};
  assign p1_sel_135229_comb = $signed(p1_or_132875_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132875_comb[23:9], 1'h0};
  assign p1_smul_135230_comb = smul16b_8b_x_9b(p1_shifted__21_squeezed_comb, 9'h0fb);
  assign p1_sel_135231_comb = $signed(p1_or_132876_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132876_comb[23:9], 1'h0};
  assign p1_smul_135232_comb = smul16b_8b_x_9b(p1_shifted__23_squeezed_comb, 9'h12b);
  assign p1_smul_135233_comb = smul16b_8b_x_9b(p1_shifted__24_squeezed_comb, 9'h0d5);
  assign p1_sel_135234_comb = $signed(p1_or_132877_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132877_comb[23:9], 1'h0};
  assign p1_smul_135235_comb = smul16b_8b_x_9b(p1_shifted__26_squeezed_comb, 9'h105);
  assign p1_sel_135236_comb = $signed(p1_or_132878_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132878_comb[23:9], 1'h0};
  assign p1_sel_135237_comb = $signed(p1_or_132879_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132879_comb[23:9], 1'h0};
  assign p1_smul_135238_comb = smul16b_8b_x_9b(p1_shifted__29_squeezed_comb, 9'h0fb);
  assign p1_sel_135239_comb = $signed(p1_or_132880_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132880_comb[23:9], 1'h0};
  assign p1_smul_135240_comb = smul16b_8b_x_9b(p1_shifted__31_squeezed_comb, 9'h12b);
  assign p1_smul_135241_comb = smul16b_8b_x_9b(p1_shifted__32_squeezed_comb, 9'h0d5);
  assign p1_sel_135242_comb = $signed(p1_or_132881_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132881_comb[23:9], 1'h0};
  assign p1_smul_135243_comb = smul16b_8b_x_9b(p1_shifted__34_squeezed_comb, 9'h105);
  assign p1_sel_135244_comb = $signed(p1_or_132882_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132882_comb[23:9], 1'h0};
  assign p1_sel_135245_comb = $signed(p1_or_132883_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132883_comb[23:9], 1'h0};
  assign p1_smul_135246_comb = smul16b_8b_x_9b(p1_shifted__37_squeezed_comb, 9'h0fb);
  assign p1_sel_135247_comb = $signed(p1_or_132884_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132884_comb[23:9], 1'h0};
  assign p1_smul_135248_comb = smul16b_8b_x_9b(p1_shifted__39_squeezed_comb, 9'h12b);
  assign p1_smul_135249_comb = smul16b_8b_x_9b(p1_shifted__40_squeezed_comb, 9'h0d5);
  assign p1_sel_135250_comb = $signed(p1_or_132885_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132885_comb[23:9], 1'h0};
  assign p1_smul_135251_comb = smul16b_8b_x_9b(p1_shifted__42_squeezed_comb, 9'h105);
  assign p1_sel_135252_comb = $signed(p1_or_132886_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132886_comb[23:9], 1'h0};
  assign p1_sel_135253_comb = $signed(p1_or_132887_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132887_comb[23:9], 1'h0};
  assign p1_smul_135254_comb = smul16b_8b_x_9b(p1_shifted__45_squeezed_comb, 9'h0fb);
  assign p1_sel_135255_comb = $signed(p1_or_132888_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132888_comb[23:9], 1'h0};
  assign p1_smul_135256_comb = smul16b_8b_x_9b(p1_shifted__47_squeezed_comb, 9'h12b);
  assign p1_smul_135257_comb = smul16b_8b_x_9b(p1_shifted__16_squeezed_comb, 9'h0b5);
  assign p1_smul_135258_comb = smul16b_8b_x_9b(p1_shifted__17_squeezed_comb, 9'h14b);
  assign p1_smul_135259_comb = smul16b_8b_x_9b(p1_shifted__18_squeezed_comb, 9'h14b);
  assign p1_smul_135260_comb = smul16b_8b_x_9b(p1_shifted__19_squeezed_comb, 9'h0b5);
  assign p1_smul_135261_comb = smul16b_8b_x_9b(p1_shifted__20_squeezed_comb, 9'h0b5);
  assign p1_smul_135262_comb = smul16b_8b_x_9b(p1_shifted__21_squeezed_comb, 9'h14b);
  assign p1_smul_135263_comb = smul16b_8b_x_9b(p1_shifted__22_squeezed_comb, 9'h14b);
  assign p1_smul_135264_comb = smul16b_8b_x_9b(p1_shifted__23_squeezed_comb, 9'h0b5);
  assign p1_smul_135265_comb = smul16b_8b_x_9b(p1_shifted__24_squeezed_comb, 9'h0b5);
  assign p1_smul_135266_comb = smul16b_8b_x_9b(p1_shifted__25_squeezed_comb, 9'h14b);
  assign p1_smul_135267_comb = smul16b_8b_x_9b(p1_shifted__26_squeezed_comb, 9'h14b);
  assign p1_smul_135268_comb = smul16b_8b_x_9b(p1_shifted__27_squeezed_comb, 9'h0b5);
  assign p1_smul_135269_comb = smul16b_8b_x_9b(p1_shifted__28_squeezed_comb, 9'h0b5);
  assign p1_smul_135270_comb = smul16b_8b_x_9b(p1_shifted__29_squeezed_comb, 9'h14b);
  assign p1_smul_135271_comb = smul16b_8b_x_9b(p1_shifted__30_squeezed_comb, 9'h14b);
  assign p1_smul_135272_comb = smul16b_8b_x_9b(p1_shifted__31_squeezed_comb, 9'h0b5);
  assign p1_smul_135273_comb = smul16b_8b_x_9b(p1_shifted__32_squeezed_comb, 9'h0b5);
  assign p1_smul_135274_comb = smul16b_8b_x_9b(p1_shifted__33_squeezed_comb, 9'h14b);
  assign p1_smul_135275_comb = smul16b_8b_x_9b(p1_shifted__34_squeezed_comb, 9'h14b);
  assign p1_smul_135276_comb = smul16b_8b_x_9b(p1_shifted__35_squeezed_comb, 9'h0b5);
  assign p1_smul_135277_comb = smul16b_8b_x_9b(p1_shifted__36_squeezed_comb, 9'h0b5);
  assign p1_smul_135278_comb = smul16b_8b_x_9b(p1_shifted__37_squeezed_comb, 9'h14b);
  assign p1_smul_135279_comb = smul16b_8b_x_9b(p1_shifted__38_squeezed_comb, 9'h14b);
  assign p1_smul_135280_comb = smul16b_8b_x_9b(p1_shifted__39_squeezed_comb, 9'h0b5);
  assign p1_smul_135281_comb = smul16b_8b_x_9b(p1_shifted__40_squeezed_comb, 9'h0b5);
  assign p1_smul_135282_comb = smul16b_8b_x_9b(p1_shifted__41_squeezed_comb, 9'h14b);
  assign p1_smul_135283_comb = smul16b_8b_x_9b(p1_shifted__42_squeezed_comb, 9'h14b);
  assign p1_smul_135284_comb = smul16b_8b_x_9b(p1_shifted__43_squeezed_comb, 9'h0b5);
  assign p1_smul_135285_comb = smul16b_8b_x_9b(p1_shifted__44_squeezed_comb, 9'h0b5);
  assign p1_smul_135286_comb = smul16b_8b_x_9b(p1_shifted__45_squeezed_comb, 9'h14b);
  assign p1_smul_135287_comb = smul16b_8b_x_9b(p1_shifted__46_squeezed_comb, 9'h14b);
  assign p1_smul_135288_comb = smul16b_8b_x_9b(p1_shifted__47_squeezed_comb, 9'h0b5);
  assign p1_sel_135289_comb = $signed(p1_or_132889_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132889_comb[23:9], 1'h0};
  assign p1_smul_135290_comb = smul16b_8b_x_9b(p1_shifted__17_squeezed_comb, 9'h105);
  assign p1_sel_135291_comb = $signed(p1_or_132890_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132890_comb[23:9], 1'h0};
  assign p1_smul_135292_comb = smul16b_8b_x_9b(p1_shifted__19_squeezed_comb, 9'h0d5);
  assign p1_smul_135293_comb = smul16b_8b_x_9b(p1_shifted__20_squeezed_comb, 9'h0d5);
  assign p1_sel_135294_comb = $signed(p1_or_132891_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132891_comb[23:9], 1'h0};
  assign p1_smul_135295_comb = smul16b_8b_x_9b(p1_shifted__22_squeezed_comb, 9'h105);
  assign p1_sel_135296_comb = $signed(p1_or_132892_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132892_comb[23:9], 1'h0};
  assign p1_sel_135297_comb = $signed(p1_or_132893_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132893_comb[23:9], 1'h0};
  assign p1_smul_135298_comb = smul16b_8b_x_9b(p1_shifted__25_squeezed_comb, 9'h105);
  assign p1_sel_135299_comb = $signed(p1_or_132894_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132894_comb[23:9], 1'h0};
  assign p1_smul_135300_comb = smul16b_8b_x_9b(p1_shifted__27_squeezed_comb, 9'h0d5);
  assign p1_smul_135301_comb = smul16b_8b_x_9b(p1_shifted__28_squeezed_comb, 9'h0d5);
  assign p1_sel_135302_comb = $signed(p1_or_132895_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132895_comb[23:9], 1'h0};
  assign p1_smul_135303_comb = smul16b_8b_x_9b(p1_shifted__30_squeezed_comb, 9'h105);
  assign p1_sel_135304_comb = $signed(p1_or_132896_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132896_comb[23:9], 1'h0};
  assign p1_sel_135305_comb = $signed(p1_or_132897_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132897_comb[23:9], 1'h0};
  assign p1_smul_135306_comb = smul16b_8b_x_9b(p1_shifted__33_squeezed_comb, 9'h105);
  assign p1_sel_135307_comb = $signed(p1_or_132898_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132898_comb[23:9], 1'h0};
  assign p1_smul_135308_comb = smul16b_8b_x_9b(p1_shifted__35_squeezed_comb, 9'h0d5);
  assign p1_smul_135309_comb = smul16b_8b_x_9b(p1_shifted__36_squeezed_comb, 9'h0d5);
  assign p1_sel_135310_comb = $signed(p1_or_132899_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132899_comb[23:9], 1'h0};
  assign p1_smul_135311_comb = smul16b_8b_x_9b(p1_shifted__38_squeezed_comb, 9'h105);
  assign p1_sel_135312_comb = $signed(p1_or_132900_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132900_comb[23:9], 1'h0};
  assign p1_sel_135313_comb = $signed(p1_or_132901_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132901_comb[23:9], 1'h0};
  assign p1_smul_135314_comb = smul16b_8b_x_9b(p1_shifted__41_squeezed_comb, 9'h105);
  assign p1_sel_135315_comb = $signed(p1_or_132902_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132902_comb[23:9], 1'h0};
  assign p1_smul_135316_comb = smul16b_8b_x_9b(p1_shifted__43_squeezed_comb, 9'h0d5);
  assign p1_smul_135317_comb = smul16b_8b_x_9b(p1_shifted__44_squeezed_comb, 9'h0d5);
  assign p1_sel_135318_comb = $signed(p1_or_132903_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132903_comb[23:9], 1'h0};
  assign p1_smul_135319_comb = smul16b_8b_x_9b(p1_shifted__46_squeezed_comb, 9'h105);
  assign p1_sel_135320_comb = $signed(p1_or_132904_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132904_comb[23:9], 1'h0};
  assign p1_sel_135321_comb = $signed(p1_concat_133545_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133545_comb;
  assign p1_sel_135322_comb = $signed(p1_or_132907_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132907_comb[23:10], 2'h0};
  assign p1_sel_135323_comb = $signed(p1_concat_133551_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133551_comb;
  assign p1_sel_135324_comb = $signed(p1_or_132910_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132910_comb[23:10], 2'h0};
  assign p1_sel_135325_comb = $signed(p1_or_132911_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132911_comb[23:10], 2'h0};
  assign p1_sel_135326_comb = $signed(p1_concat_133561_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133561_comb;
  assign p1_sel_135327_comb = $signed(p1_or_132914_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132914_comb[23:10], 2'h0};
  assign p1_sel_135328_comb = $signed(p1_concat_133567_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133567_comb;
  assign p1_sel_135329_comb = $signed(p1_concat_133569_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133569_comb;
  assign p1_sel_135330_comb = $signed(p1_or_132919_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132919_comb[23:10], 2'h0};
  assign p1_sel_135331_comb = $signed(p1_concat_133575_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133575_comb;
  assign p1_sel_135332_comb = $signed(p1_or_132922_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132922_comb[23:10], 2'h0};
  assign p1_sel_135333_comb = $signed(p1_or_132923_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132923_comb[23:10], 2'h0};
  assign p1_sel_135334_comb = $signed(p1_concat_133585_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133585_comb;
  assign p1_sel_135335_comb = $signed(p1_or_132926_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132926_comb[23:10], 2'h0};
  assign p1_sel_135336_comb = $signed(p1_concat_133591_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133591_comb;
  assign p1_sel_135337_comb = $signed(p1_concat_133593_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133593_comb;
  assign p1_sel_135338_comb = $signed(p1_or_132931_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132931_comb[23:10], 2'h0};
  assign p1_sel_135339_comb = $signed(p1_concat_133599_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133599_comb;
  assign p1_sel_135340_comb = $signed(p1_or_132934_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132934_comb[23:10], 2'h0};
  assign p1_sel_135341_comb = $signed(p1_or_132935_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132935_comb[23:10], 2'h0};
  assign p1_sel_135342_comb = $signed(p1_concat_133609_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133609_comb;
  assign p1_sel_135343_comb = $signed(p1_or_132938_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132938_comb[23:10], 2'h0};
  assign p1_sel_135344_comb = $signed(p1_concat_133615_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133615_comb;
  assign p1_sel_135345_comb = $signed(p1_concat_133617_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133617_comb;
  assign p1_sel_135346_comb = $signed(p1_or_132943_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132943_comb[23:10], 2'h0};
  assign p1_sel_135347_comb = $signed(p1_concat_133623_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133623_comb;
  assign p1_sel_135348_comb = $signed(p1_or_132946_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132946_comb[23:10], 2'h0};
  assign p1_sel_135349_comb = $signed(p1_or_132947_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132947_comb[23:10], 2'h0};
  assign p1_sel_135350_comb = $signed(p1_concat_133633_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133633_comb;
  assign p1_sel_135351_comb = $signed(p1_or_132950_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132950_comb[23:10], 2'h0};
  assign p1_sel_135352_comb = $signed(p1_concat_133639_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133639_comb;
  assign p1_sel_135353_comb = $signed(p1_or_132953_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132953_comb[23:9], 1'h0};
  assign p1_sel_135354_comb = $signed(p1_or_132954_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132954_comb[23:9], 1'h0};
  assign p1_smul_135355_comb = smul16b_8b_x_9b(p1_shifted__18_squeezed_comb, 9'h0d5);
  assign p1_smul_135356_comb = smul16b_8b_x_9b(p1_shifted__19_squeezed_comb, 9'h105);
  assign p1_smul_135357_comb = smul16b_8b_x_9b(p1_shifted__20_squeezed_comb, 9'h105);
  assign p1_smul_135358_comb = smul16b_8b_x_9b(p1_shifted__21_squeezed_comb, 9'h0d5);
  assign p1_sel_135359_comb = $signed(p1_or_132955_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132955_comb[23:9], 1'h0};
  assign p1_sel_135360_comb = $signed(p1_or_132956_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132956_comb[23:9], 1'h0};
  assign p1_sel_135361_comb = $signed(p1_or_132957_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132957_comb[23:9], 1'h0};
  assign p1_sel_135362_comb = $signed(p1_or_132958_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132958_comb[23:9], 1'h0};
  assign p1_smul_135363_comb = smul16b_8b_x_9b(p1_shifted__26_squeezed_comb, 9'h0d5);
  assign p1_smul_135364_comb = smul16b_8b_x_9b(p1_shifted__27_squeezed_comb, 9'h105);
  assign p1_smul_135365_comb = smul16b_8b_x_9b(p1_shifted__28_squeezed_comb, 9'h105);
  assign p1_smul_135366_comb = smul16b_8b_x_9b(p1_shifted__29_squeezed_comb, 9'h0d5);
  assign p1_sel_135367_comb = $signed(p1_or_132959_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132959_comb[23:9], 1'h0};
  assign p1_sel_135368_comb = $signed(p1_or_132960_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132960_comb[23:9], 1'h0};
  assign p1_sel_135369_comb = $signed(p1_or_132961_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132961_comb[23:9], 1'h0};
  assign p1_sel_135370_comb = $signed(p1_or_132962_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132962_comb[23:9], 1'h0};
  assign p1_smul_135371_comb = smul16b_8b_x_9b(p1_shifted__34_squeezed_comb, 9'h0d5);
  assign p1_smul_135372_comb = smul16b_8b_x_9b(p1_shifted__35_squeezed_comb, 9'h105);
  assign p1_smul_135373_comb = smul16b_8b_x_9b(p1_shifted__36_squeezed_comb, 9'h105);
  assign p1_smul_135374_comb = smul16b_8b_x_9b(p1_shifted__37_squeezed_comb, 9'h0d5);
  assign p1_sel_135375_comb = $signed(p1_or_132963_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132963_comb[23:9], 1'h0};
  assign p1_sel_135376_comb = $signed(p1_or_132964_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132964_comb[23:9], 1'h0};
  assign p1_sel_135377_comb = $signed(p1_or_132965_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132965_comb[23:9], 1'h0};
  assign p1_sel_135378_comb = $signed(p1_or_132966_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132966_comb[23:9], 1'h0};
  assign p1_smul_135379_comb = smul16b_8b_x_9b(p1_shifted__42_squeezed_comb, 9'h0d5);
  assign p1_smul_135380_comb = smul16b_8b_x_9b(p1_shifted__43_squeezed_comb, 9'h105);
  assign p1_smul_135381_comb = smul16b_8b_x_9b(p1_shifted__44_squeezed_comb, 9'h105);
  assign p1_smul_135382_comb = smul16b_8b_x_9b(p1_shifted__45_squeezed_comb, 9'h0d5);
  assign p1_sel_135383_comb = $signed(p1_or_132967_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132967_comb[23:9], 1'h0};
  assign p1_sel_135384_comb = $signed(p1_or_132968_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_132968_comb[23:9], 1'h0};
  assign p1_add_135385_comb = {{1{p1_sel_133705_comb[15]}}, p1_sel_133705_comb} + {{1{p1_sel_133706_comb[15]}}, p1_sel_133706_comb};
  assign p1_add_135386_comb = {{1{p1_sel_133707_comb[15]}}, p1_sel_133707_comb} + {{1{p1_sel_133708_comb[15]}}, p1_sel_133708_comb};
  assign p1_add_135387_comb = {{1{p1_sel_133709_comb[15]}}, p1_sel_133709_comb} + {{1{p1_sel_133710_comb[15]}}, p1_sel_133710_comb};
  assign p1_add_135388_comb = {{1{p1_sel_133711_comb[15]}}, p1_sel_133711_comb} + {{1{p1_sel_133712_comb[15]}}, p1_sel_133712_comb};
  assign p1_add_135389_comb = {{1{p1_sel_133713_comb[15]}}, p1_sel_133713_comb} + {{1{p1_sel_133714_comb[15]}}, p1_sel_133714_comb};
  assign p1_add_135390_comb = {{1{p1_sel_133715_comb[15]}}, p1_sel_133715_comb} + {{1{p1_sel_133716_comb[15]}}, p1_sel_133716_comb};
  assign p1_add_135391_comb = {{1{p1_sel_133717_comb[15]}}, p1_sel_133717_comb} + {{1{p1_sel_133718_comb[15]}}, p1_sel_133718_comb};
  assign p1_add_135392_comb = {{1{p1_sel_133719_comb[15]}}, p1_sel_133719_comb} + {{1{p1_sel_133720_comb[15]}}, p1_sel_133720_comb};
  assign p1_smul_135393_comb = smul16b_8b_x_9b(p1_shifted_squeezed_comb, 9'h0fb);
  assign p1_smul_135394_comb = smul16b_8b_x_9b(p1_shifted__1_squeezed_comb, 9'h0d5);
  assign p1_sel_135395_comb = $signed(p1_or_133017_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133017_comb[23:9], 1'h0};
  assign p1_sel_135396_comb = $signed(p1_or_133018_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133018_comb[23:9], 1'h0};
  assign p1_sel_135397_comb = $signed(p1_or_133019_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133019_comb[23:9], 1'h0};
  assign p1_sel_135398_comb = $signed(p1_or_133020_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133020_comb[23:9], 1'h0};
  assign p1_smul_135399_comb = smul16b_8b_x_9b(p1_shifted__6_squeezed_comb, 9'h12b);
  assign p1_smul_135400_comb = smul16b_8b_x_9b(p1_shifted__7_squeezed_comb, 9'h105);
  assign p1_smul_135401_comb = smul16b_8b_x_9b(p1_shifted__56_squeezed_comb, 9'h0fb);
  assign p1_smul_135402_comb = smul16b_8b_x_9b(p1_shifted__57_squeezed_comb, 9'h0d5);
  assign p1_sel_135403_comb = $signed(p1_or_133021_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133021_comb[23:9], 1'h0};
  assign p1_sel_135404_comb = $signed(p1_or_133022_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133022_comb[23:9], 1'h0};
  assign p1_sel_135405_comb = $signed(p1_or_133023_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133023_comb[23:9], 1'h0};
  assign p1_sel_135406_comb = $signed(p1_or_133024_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133024_comb[23:9], 1'h0};
  assign p1_smul_135407_comb = smul16b_8b_x_9b(p1_shifted__62_squeezed_comb, 9'h12b);
  assign p1_smul_135408_comb = smul16b_8b_x_9b(p1_shifted__63_squeezed_comb, 9'h105);
  assign p1_sel_135409_comb = $signed(p1_or_133025_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133025_comb[23:10], 2'h0};
  assign p1_sel_135410_comb = $signed(p1_concat_133757_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133757_comb;
  assign p1_sel_135411_comb = $signed(p1_concat_133759_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133759_comb;
  assign p1_sel_135412_comb = $signed(p1_or_133030_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133030_comb[23:10], 2'h0};
  assign p1_sel_135413_comb = $signed(p1_or_133031_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133031_comb[23:10], 2'h0};
  assign p1_sel_135414_comb = $signed(p1_concat_133769_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133769_comb;
  assign p1_sel_135415_comb = $signed(p1_concat_133771_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133771_comb;
  assign p1_sel_135416_comb = $signed(p1_or_133036_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133036_comb[23:10], 2'h0};
  assign p1_sel_135417_comb = $signed(p1_or_133037_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133037_comb[23:10], 2'h0};
  assign p1_sel_135418_comb = $signed(p1_concat_133781_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133781_comb;
  assign p1_sel_135419_comb = $signed(p1_concat_133783_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133783_comb;
  assign p1_sel_135420_comb = $signed(p1_or_133042_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133042_comb[23:10], 2'h0};
  assign p1_sel_135421_comb = $signed(p1_or_133043_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133043_comb[23:10], 2'h0};
  assign p1_sel_135422_comb = $signed(p1_concat_133793_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133793_comb;
  assign p1_sel_135423_comb = $signed(p1_concat_133795_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133795_comb;
  assign p1_sel_135424_comb = $signed(p1_or_133048_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133048_comb[23:10], 2'h0};
  assign p1_smul_135425_comb = smul16b_8b_x_9b(p1_shifted_squeezed_comb, 9'h0d5);
  assign p1_sel_135426_comb = $signed(p1_or_133049_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133049_comb[23:9], 1'h0};
  assign p1_smul_135427_comb = smul16b_8b_x_9b(p1_shifted__2_squeezed_comb, 9'h105);
  assign p1_sel_135428_comb = $signed(p1_or_133050_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133050_comb[23:9], 1'h0};
  assign p1_sel_135429_comb = $signed(p1_or_133051_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133051_comb[23:9], 1'h0};
  assign p1_smul_135430_comb = smul16b_8b_x_9b(p1_shifted__5_squeezed_comb, 9'h0fb);
  assign p1_sel_135431_comb = $signed(p1_or_133052_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133052_comb[23:9], 1'h0};
  assign p1_smul_135432_comb = smul16b_8b_x_9b(p1_shifted__7_squeezed_comb, 9'h12b);
  assign p1_smul_135433_comb = smul16b_8b_x_9b(p1_shifted__56_squeezed_comb, 9'h0d5);
  assign p1_sel_135434_comb = $signed(p1_or_133053_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133053_comb[23:9], 1'h0};
  assign p1_smul_135435_comb = smul16b_8b_x_9b(p1_shifted__58_squeezed_comb, 9'h105);
  assign p1_sel_135436_comb = $signed(p1_or_133054_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133054_comb[23:9], 1'h0};
  assign p1_sel_135437_comb = $signed(p1_or_133055_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133055_comb[23:9], 1'h0};
  assign p1_smul_135438_comb = smul16b_8b_x_9b(p1_shifted__61_squeezed_comb, 9'h0fb);
  assign p1_sel_135439_comb = $signed(p1_or_133056_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133056_comb[23:9], 1'h0};
  assign p1_smul_135440_comb = smul16b_8b_x_9b(p1_shifted__63_squeezed_comb, 9'h12b);
  assign p1_smul_135441_comb = smul16b_8b_x_9b(p1_shifted_squeezed_comb, 9'h0b5);
  assign p1_smul_135442_comb = smul16b_8b_x_9b(p1_shifted__1_squeezed_comb, 9'h14b);
  assign p1_smul_135443_comb = smul16b_8b_x_9b(p1_shifted__2_squeezed_comb, 9'h14b);
  assign p1_smul_135444_comb = smul16b_8b_x_9b(p1_shifted__3_squeezed_comb, 9'h0b5);
  assign p1_smul_135445_comb = smul16b_8b_x_9b(p1_shifted__4_squeezed_comb, 9'h0b5);
  assign p1_smul_135446_comb = smul16b_8b_x_9b(p1_shifted__5_squeezed_comb, 9'h14b);
  assign p1_smul_135447_comb = smul16b_8b_x_9b(p1_shifted__6_squeezed_comb, 9'h14b);
  assign p1_smul_135448_comb = smul16b_8b_x_9b(p1_shifted__7_squeezed_comb, 9'h0b5);
  assign p1_smul_135449_comb = smul16b_8b_x_9b(p1_shifted__56_squeezed_comb, 9'h0b5);
  assign p1_smul_135450_comb = smul16b_8b_x_9b(p1_shifted__57_squeezed_comb, 9'h14b);
  assign p1_smul_135451_comb = smul16b_8b_x_9b(p1_shifted__58_squeezed_comb, 9'h14b);
  assign p1_smul_135452_comb = smul16b_8b_x_9b(p1_shifted__59_squeezed_comb, 9'h0b5);
  assign p1_smul_135453_comb = smul16b_8b_x_9b(p1_shifted__60_squeezed_comb, 9'h0b5);
  assign p1_smul_135454_comb = smul16b_8b_x_9b(p1_shifted__61_squeezed_comb, 9'h14b);
  assign p1_smul_135455_comb = smul16b_8b_x_9b(p1_shifted__62_squeezed_comb, 9'h14b);
  assign p1_smul_135456_comb = smul16b_8b_x_9b(p1_shifted__63_squeezed_comb, 9'h0b5);
  assign p1_sel_135457_comb = $signed(p1_or_133057_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133057_comb[23:9], 1'h0};
  assign p1_smul_135458_comb = smul16b_8b_x_9b(p1_shifted__1_squeezed_comb, 9'h105);
  assign p1_sel_135459_comb = $signed(p1_or_133058_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133058_comb[23:9], 1'h0};
  assign p1_smul_135460_comb = smul16b_8b_x_9b(p1_shifted__3_squeezed_comb, 9'h0d5);
  assign p1_smul_135461_comb = smul16b_8b_x_9b(p1_shifted__4_squeezed_comb, 9'h0d5);
  assign p1_sel_135462_comb = $signed(p1_or_133059_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133059_comb[23:9], 1'h0};
  assign p1_smul_135463_comb = smul16b_8b_x_9b(p1_shifted__6_squeezed_comb, 9'h105);
  assign p1_sel_135464_comb = $signed(p1_or_133060_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133060_comb[23:9], 1'h0};
  assign p1_sel_135465_comb = $signed(p1_or_133061_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133061_comb[23:9], 1'h0};
  assign p1_smul_135466_comb = smul16b_8b_x_9b(p1_shifted__57_squeezed_comb, 9'h105);
  assign p1_sel_135467_comb = $signed(p1_or_133062_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133062_comb[23:9], 1'h0};
  assign p1_smul_135468_comb = smul16b_8b_x_9b(p1_shifted__59_squeezed_comb, 9'h0d5);
  assign p1_smul_135469_comb = smul16b_8b_x_9b(p1_shifted__60_squeezed_comb, 9'h0d5);
  assign p1_sel_135470_comb = $signed(p1_or_133063_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133063_comb[23:9], 1'h0};
  assign p1_smul_135471_comb = smul16b_8b_x_9b(p1_shifted__62_squeezed_comb, 9'h105);
  assign p1_sel_135472_comb = $signed(p1_or_133064_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133064_comb[23:9], 1'h0};
  assign p1_sel_135473_comb = $signed(p1_concat_133865_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133865_comb;
  assign p1_sel_135474_comb = $signed(p1_or_133067_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133067_comb[23:10], 2'h0};
  assign p1_sel_135475_comb = $signed(p1_concat_133871_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133871_comb;
  assign p1_sel_135476_comb = $signed(p1_or_133070_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133070_comb[23:10], 2'h0};
  assign p1_sel_135477_comb = $signed(p1_or_133071_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133071_comb[23:10], 2'h0};
  assign p1_sel_135478_comb = $signed(p1_concat_133881_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133881_comb;
  assign p1_sel_135479_comb = $signed(p1_or_133074_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133074_comb[23:10], 2'h0};
  assign p1_sel_135480_comb = $signed(p1_concat_133887_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133887_comb;
  assign p1_sel_135481_comb = $signed(p1_concat_133889_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133889_comb;
  assign p1_sel_135482_comb = $signed(p1_or_133079_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133079_comb[23:10], 2'h0};
  assign p1_sel_135483_comb = $signed(p1_concat_133895_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133895_comb;
  assign p1_sel_135484_comb = $signed(p1_or_133082_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133082_comb[23:10], 2'h0};
  assign p1_sel_135485_comb = $signed(p1_or_133083_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133083_comb[23:10], 2'h0};
  assign p1_sel_135486_comb = $signed(p1_concat_133905_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133905_comb;
  assign p1_sel_135487_comb = $signed(p1_or_133086_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133086_comb[23:10], 2'h0};
  assign p1_sel_135488_comb = $signed(p1_concat_133911_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133911_comb;
  assign p1_sel_135489_comb = $signed(p1_or_133089_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133089_comb[23:9], 1'h0};
  assign p1_sel_135490_comb = $signed(p1_or_133090_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133090_comb[23:9], 1'h0};
  assign p1_smul_135491_comb = smul16b_8b_x_9b(p1_shifted__2_squeezed_comb, 9'h0d5);
  assign p1_smul_135492_comb = smul16b_8b_x_9b(p1_shifted__3_squeezed_comb, 9'h105);
  assign p1_smul_135493_comb = smul16b_8b_x_9b(p1_shifted__4_squeezed_comb, 9'h105);
  assign p1_smul_135494_comb = smul16b_8b_x_9b(p1_shifted__5_squeezed_comb, 9'h0d5);
  assign p1_sel_135495_comb = $signed(p1_or_133091_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133091_comb[23:9], 1'h0};
  assign p1_sel_135496_comb = $signed(p1_or_133092_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133092_comb[23:9], 1'h0};
  assign p1_sel_135497_comb = $signed(p1_or_133093_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133093_comb[23:9], 1'h0};
  assign p1_sel_135498_comb = $signed(p1_or_133094_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133094_comb[23:9], 1'h0};
  assign p1_smul_135499_comb = smul16b_8b_x_9b(p1_shifted__58_squeezed_comb, 9'h0d5);
  assign p1_smul_135500_comb = smul16b_8b_x_9b(p1_shifted__59_squeezed_comb, 9'h105);
  assign p1_smul_135501_comb = smul16b_8b_x_9b(p1_shifted__60_squeezed_comb, 9'h105);
  assign p1_smul_135502_comb = smul16b_8b_x_9b(p1_shifted__61_squeezed_comb, 9'h0d5);
  assign p1_sel_135503_comb = $signed(p1_or_133095_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133095_comb[23:9], 1'h0};
  assign p1_sel_135504_comb = $signed(p1_or_133096_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133096_comb[23:9], 1'h0};
  assign p1_add_135505_comb = {{1{p1_sel_133945_comb[15]}}, p1_sel_133945_comb} + {{1{p1_sel_133946_comb[15]}}, p1_sel_133946_comb};
  assign p1_add_135506_comb = {{1{p1_sel_133947_comb[15]}}, p1_sel_133947_comb} + {{1{p1_sel_133948_comb[15]}}, p1_sel_133948_comb};
  assign p1_add_135507_comb = {{1{p1_sel_133949_comb[15]}}, p1_sel_133949_comb} + {{1{p1_sel_133950_comb[15]}}, p1_sel_133950_comb};
  assign p1_add_135508_comb = {{1{p1_sel_133951_comb[15]}}, p1_sel_133951_comb} + {{1{p1_sel_133952_comb[15]}}, p1_sel_133952_comb};
  assign p1_add_135509_comb = {{1{p1_sel_133953_comb[15]}}, p1_sel_133953_comb} + {{1{p1_sel_133954_comb[15]}}, p1_sel_133954_comb};
  assign p1_add_135510_comb = {{1{p1_sel_133955_comb[15]}}, p1_sel_133955_comb} + {{1{p1_sel_133956_comb[15]}}, p1_sel_133956_comb};
  assign p1_add_135511_comb = {{1{p1_sel_133957_comb[15]}}, p1_sel_133957_comb} + {{1{p1_sel_133958_comb[15]}}, p1_sel_133958_comb};
  assign p1_add_135512_comb = {{1{p1_sel_133959_comb[15]}}, p1_sel_133959_comb} + {{1{p1_sel_133960_comb[15]}}, p1_sel_133960_comb};
  assign p1_smul_135513_comb = smul16b_8b_x_9b(p1_shifted__8_squeezed_comb, 9'h0fb);
  assign p1_smul_135514_comb = smul16b_8b_x_9b(p1_shifted__9_squeezed_comb, 9'h0d5);
  assign p1_sel_135515_comb = $signed(p1_or_133145_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133145_comb[23:9], 1'h0};
  assign p1_sel_135516_comb = $signed(p1_or_133146_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133146_comb[23:9], 1'h0};
  assign p1_sel_135517_comb = $signed(p1_or_133147_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133147_comb[23:9], 1'h0};
  assign p1_sel_135518_comb = $signed(p1_or_133148_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133148_comb[23:9], 1'h0};
  assign p1_smul_135519_comb = smul16b_8b_x_9b(p1_shifted__14_squeezed_comb, 9'h12b);
  assign p1_smul_135520_comb = smul16b_8b_x_9b(p1_shifted__15_squeezed_comb, 9'h105);
  assign p1_smul_135521_comb = smul16b_8b_x_9b(p1_shifted__48_squeezed_comb, 9'h0fb);
  assign p1_smul_135522_comb = smul16b_8b_x_9b(p1_shifted__49_squeezed_comb, 9'h0d5);
  assign p1_sel_135523_comb = $signed(p1_or_133149_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133149_comb[23:9], 1'h0};
  assign p1_sel_135524_comb = $signed(p1_or_133150_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133150_comb[23:9], 1'h0};
  assign p1_sel_135525_comb = $signed(p1_or_133151_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133151_comb[23:9], 1'h0};
  assign p1_sel_135526_comb = $signed(p1_or_133152_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133152_comb[23:9], 1'h0};
  assign p1_smul_135527_comb = smul16b_8b_x_9b(p1_shifted__54_squeezed_comb, 9'h12b);
  assign p1_smul_135528_comb = smul16b_8b_x_9b(p1_shifted__55_squeezed_comb, 9'h105);
  assign p1_sel_135529_comb = $signed(p1_or_133153_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133153_comb[23:10], 2'h0};
  assign p1_sel_135530_comb = $signed(p1_concat_133997_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133997_comb;
  assign p1_sel_135531_comb = $signed(p1_concat_133999_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_133999_comb;
  assign p1_sel_135532_comb = $signed(p1_or_133158_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133158_comb[23:10], 2'h0};
  assign p1_sel_135533_comb = $signed(p1_or_133159_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133159_comb[23:10], 2'h0};
  assign p1_sel_135534_comb = $signed(p1_concat_134009_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134009_comb;
  assign p1_sel_135535_comb = $signed(p1_concat_134011_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134011_comb;
  assign p1_sel_135536_comb = $signed(p1_or_133164_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133164_comb[23:10], 2'h0};
  assign p1_sel_135537_comb = $signed(p1_or_133165_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133165_comb[23:10], 2'h0};
  assign p1_sel_135538_comb = $signed(p1_concat_134021_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134021_comb;
  assign p1_sel_135539_comb = $signed(p1_concat_134023_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134023_comb;
  assign p1_sel_135540_comb = $signed(p1_or_133170_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133170_comb[23:10], 2'h0};
  assign p1_sel_135541_comb = $signed(p1_or_133171_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133171_comb[23:10], 2'h0};
  assign p1_sel_135542_comb = $signed(p1_concat_134033_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134033_comb;
  assign p1_sel_135543_comb = $signed(p1_concat_134035_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134035_comb;
  assign p1_sel_135544_comb = $signed(p1_or_133176_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133176_comb[23:10], 2'h0};
  assign p1_smul_135545_comb = smul16b_8b_x_9b(p1_shifted__8_squeezed_comb, 9'h0d5);
  assign p1_sel_135546_comb = $signed(p1_or_133177_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133177_comb[23:9], 1'h0};
  assign p1_smul_135547_comb = smul16b_8b_x_9b(p1_shifted__10_squeezed_comb, 9'h105);
  assign p1_sel_135548_comb = $signed(p1_or_133178_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133178_comb[23:9], 1'h0};
  assign p1_sel_135549_comb = $signed(p1_or_133179_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133179_comb[23:9], 1'h0};
  assign p1_smul_135550_comb = smul16b_8b_x_9b(p1_shifted__13_squeezed_comb, 9'h0fb);
  assign p1_sel_135551_comb = $signed(p1_or_133180_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133180_comb[23:9], 1'h0};
  assign p1_smul_135552_comb = smul16b_8b_x_9b(p1_shifted__15_squeezed_comb, 9'h12b);
  assign p1_smul_135553_comb = smul16b_8b_x_9b(p1_shifted__48_squeezed_comb, 9'h0d5);
  assign p1_sel_135554_comb = $signed(p1_or_133181_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133181_comb[23:9], 1'h0};
  assign p1_smul_135555_comb = smul16b_8b_x_9b(p1_shifted__50_squeezed_comb, 9'h105);
  assign p1_sel_135556_comb = $signed(p1_or_133182_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133182_comb[23:9], 1'h0};
  assign p1_sel_135557_comb = $signed(p1_or_133183_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133183_comb[23:9], 1'h0};
  assign p1_smul_135558_comb = smul16b_8b_x_9b(p1_shifted__53_squeezed_comb, 9'h0fb);
  assign p1_sel_135559_comb = $signed(p1_or_133184_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133184_comb[23:9], 1'h0};
  assign p1_smul_135560_comb = smul16b_8b_x_9b(p1_shifted__55_squeezed_comb, 9'h12b);
  assign p1_smul_135561_comb = smul16b_8b_x_9b(p1_shifted__8_squeezed_comb, 9'h0b5);
  assign p1_smul_135562_comb = smul16b_8b_x_9b(p1_shifted__9_squeezed_comb, 9'h14b);
  assign p1_smul_135563_comb = smul16b_8b_x_9b(p1_shifted__10_squeezed_comb, 9'h14b);
  assign p1_smul_135564_comb = smul16b_8b_x_9b(p1_shifted__11_squeezed_comb, 9'h0b5);
  assign p1_smul_135565_comb = smul16b_8b_x_9b(p1_shifted__12_squeezed_comb, 9'h0b5);
  assign p1_smul_135566_comb = smul16b_8b_x_9b(p1_shifted__13_squeezed_comb, 9'h14b);
  assign p1_smul_135567_comb = smul16b_8b_x_9b(p1_shifted__14_squeezed_comb, 9'h14b);
  assign p1_smul_135568_comb = smul16b_8b_x_9b(p1_shifted__15_squeezed_comb, 9'h0b5);
  assign p1_smul_135569_comb = smul16b_8b_x_9b(p1_shifted__48_squeezed_comb, 9'h0b5);
  assign p1_smul_135570_comb = smul16b_8b_x_9b(p1_shifted__49_squeezed_comb, 9'h14b);
  assign p1_smul_135571_comb = smul16b_8b_x_9b(p1_shifted__50_squeezed_comb, 9'h14b);
  assign p1_smul_135572_comb = smul16b_8b_x_9b(p1_shifted__51_squeezed_comb, 9'h0b5);
  assign p1_smul_135573_comb = smul16b_8b_x_9b(p1_shifted__52_squeezed_comb, 9'h0b5);
  assign p1_smul_135574_comb = smul16b_8b_x_9b(p1_shifted__53_squeezed_comb, 9'h14b);
  assign p1_smul_135575_comb = smul16b_8b_x_9b(p1_shifted__54_squeezed_comb, 9'h14b);
  assign p1_smul_135576_comb = smul16b_8b_x_9b(p1_shifted__55_squeezed_comb, 9'h0b5);
  assign p1_sel_135577_comb = $signed(p1_or_133185_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133185_comb[23:9], 1'h0};
  assign p1_smul_135578_comb = smul16b_8b_x_9b(p1_shifted__9_squeezed_comb, 9'h105);
  assign p1_sel_135579_comb = $signed(p1_or_133186_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133186_comb[23:9], 1'h0};
  assign p1_smul_135580_comb = smul16b_8b_x_9b(p1_shifted__11_squeezed_comb, 9'h0d5);
  assign p1_smul_135581_comb = smul16b_8b_x_9b(p1_shifted__12_squeezed_comb, 9'h0d5);
  assign p1_sel_135582_comb = $signed(p1_or_133187_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133187_comb[23:9], 1'h0};
  assign p1_smul_135583_comb = smul16b_8b_x_9b(p1_shifted__14_squeezed_comb, 9'h105);
  assign p1_sel_135584_comb = $signed(p1_or_133188_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133188_comb[23:9], 1'h0};
  assign p1_sel_135585_comb = $signed(p1_or_133189_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133189_comb[23:9], 1'h0};
  assign p1_smul_135586_comb = smul16b_8b_x_9b(p1_shifted__49_squeezed_comb, 9'h105);
  assign p1_sel_135587_comb = $signed(p1_or_133190_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133190_comb[23:9], 1'h0};
  assign p1_smul_135588_comb = smul16b_8b_x_9b(p1_shifted__51_squeezed_comb, 9'h0d5);
  assign p1_smul_135589_comb = smul16b_8b_x_9b(p1_shifted__52_squeezed_comb, 9'h0d5);
  assign p1_sel_135590_comb = $signed(p1_or_133191_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133191_comb[23:9], 1'h0};
  assign p1_smul_135591_comb = smul16b_8b_x_9b(p1_shifted__54_squeezed_comb, 9'h105);
  assign p1_sel_135592_comb = $signed(p1_or_133192_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133192_comb[23:9], 1'h0};
  assign p1_sel_135593_comb = $signed(p1_concat_134105_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134105_comb;
  assign p1_sel_135594_comb = $signed(p1_or_133195_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133195_comb[23:10], 2'h0};
  assign p1_sel_135595_comb = $signed(p1_concat_134111_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134111_comb;
  assign p1_sel_135596_comb = $signed(p1_or_133198_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133198_comb[23:10], 2'h0};
  assign p1_sel_135597_comb = $signed(p1_or_133199_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133199_comb[23:10], 2'h0};
  assign p1_sel_135598_comb = $signed(p1_concat_134121_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134121_comb;
  assign p1_sel_135599_comb = $signed(p1_or_133202_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133202_comb[23:10], 2'h0};
  assign p1_sel_135600_comb = $signed(p1_concat_134127_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134127_comb;
  assign p1_sel_135601_comb = $signed(p1_concat_134129_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134129_comb;
  assign p1_sel_135602_comb = $signed(p1_or_133207_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133207_comb[23:10], 2'h0};
  assign p1_sel_135603_comb = $signed(p1_concat_134135_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134135_comb;
  assign p1_sel_135604_comb = $signed(p1_or_133210_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133210_comb[23:10], 2'h0};
  assign p1_sel_135605_comb = $signed(p1_or_133211_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133211_comb[23:10], 2'h0};
  assign p1_sel_135606_comb = $signed(p1_concat_134145_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134145_comb;
  assign p1_sel_135607_comb = $signed(p1_or_133214_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133214_comb[23:10], 2'h0};
  assign p1_sel_135608_comb = $signed(p1_concat_134151_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_134151_comb;
  assign p1_sel_135609_comb = $signed(p1_or_133217_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133217_comb[23:9], 1'h0};
  assign p1_sel_135610_comb = $signed(p1_or_133218_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133218_comb[23:9], 1'h0};
  assign p1_smul_135611_comb = smul16b_8b_x_9b(p1_shifted__10_squeezed_comb, 9'h0d5);
  assign p1_smul_135612_comb = smul16b_8b_x_9b(p1_shifted__11_squeezed_comb, 9'h105);
  assign p1_smul_135613_comb = smul16b_8b_x_9b(p1_shifted__12_squeezed_comb, 9'h105);
  assign p1_smul_135614_comb = smul16b_8b_x_9b(p1_shifted__13_squeezed_comb, 9'h0d5);
  assign p1_sel_135615_comb = $signed(p1_or_133219_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133219_comb[23:9], 1'h0};
  assign p1_sel_135616_comb = $signed(p1_or_133220_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133220_comb[23:9], 1'h0};
  assign p1_sel_135617_comb = $signed(p1_or_133221_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133221_comb[23:9], 1'h0};
  assign p1_sel_135618_comb = $signed(p1_or_133222_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133222_comb[23:9], 1'h0};
  assign p1_smul_135619_comb = smul16b_8b_x_9b(p1_shifted__50_squeezed_comb, 9'h0d5);
  assign p1_smul_135620_comb = smul16b_8b_x_9b(p1_shifted__51_squeezed_comb, 9'h105);
  assign p1_smul_135621_comb = smul16b_8b_x_9b(p1_shifted__52_squeezed_comb, 9'h105);
  assign p1_smul_135622_comb = smul16b_8b_x_9b(p1_shifted__53_squeezed_comb, 9'h0d5);
  assign p1_sel_135623_comb = $signed(p1_or_133223_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133223_comb[23:9], 1'h0};
  assign p1_sel_135624_comb = $signed(p1_or_133224_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_133224_comb[23:9], 1'h0};
  assign p1_sum__989_comb = {{15{p1_add_135145_comb[16]}}, p1_add_135145_comb};
  assign p1_sum__990_comb = {{15{p1_add_135146_comb[16]}}, p1_add_135146_comb};
  assign p1_sum__991_comb = {{15{p1_add_135147_comb[16]}}, p1_add_135147_comb};
  assign p1_sum__992_comb = {{15{p1_add_135148_comb[16]}}, p1_add_135148_comb};
  assign p1_sum__961_comb = {{15{p1_add_135149_comb[16]}}, p1_add_135149_comb};
  assign p1_sum__962_comb = {{15{p1_add_135150_comb[16]}}, p1_add_135150_comb};
  assign p1_sum__963_comb = {{15{p1_add_135151_comb[16]}}, p1_add_135151_comb};
  assign p1_sum__964_comb = {{15{p1_add_135152_comb[16]}}, p1_add_135152_comb};
  assign p1_sum__926_comb = {{15{p1_add_135153_comb[16]}}, p1_add_135153_comb};
  assign p1_sum__927_comb = {{15{p1_add_135154_comb[16]}}, p1_add_135154_comb};
  assign p1_sum__928_comb = {{15{p1_add_135155_comb[16]}}, p1_add_135155_comb};
  assign p1_sum__929_comb = {{15{p1_add_135156_comb[16]}}, p1_add_135156_comb};
  assign p1_sum__884_comb = {{15{p1_add_135157_comb[16]}}, p1_add_135157_comb};
  assign p1_sum__885_comb = {{15{p1_add_135158_comb[16]}}, p1_add_135158_comb};
  assign p1_sum__886_comb = {{15{p1_add_135159_comb[16]}}, p1_add_135159_comb};
  assign p1_sum__887_comb = {{15{p1_add_135160_comb[16]}}, p1_add_135160_comb};
  assign p1_sum__1017_comb = {{15{p1_add_135385_comb[16]}}, p1_add_135385_comb};
  assign p1_sum__1018_comb = {{15{p1_add_135386_comb[16]}}, p1_add_135386_comb};
  assign p1_sum__1019_comb = {{15{p1_add_135387_comb[16]}}, p1_add_135387_comb};
  assign p1_sum__1020_comb = {{15{p1_add_135388_comb[16]}}, p1_add_135388_comb};
  assign p1_sum__779_comb = {{15{p1_add_135389_comb[16]}}, p1_add_135389_comb};
  assign p1_sum__780_comb = {{15{p1_add_135390_comb[16]}}, p1_add_135390_comb};
  assign p1_sum__781_comb = {{15{p1_add_135391_comb[16]}}, p1_add_135391_comb};
  assign p1_sum__782_comb = {{15{p1_add_135392_comb[16]}}, p1_add_135392_comb};
  assign p1_sum__1010_comb = {{15{p1_add_135505_comb[16]}}, p1_add_135505_comb};
  assign p1_sum__1011_comb = {{15{p1_add_135506_comb[16]}}, p1_add_135506_comb};
  assign p1_sum__1012_comb = {{15{p1_add_135507_comb[16]}}, p1_add_135507_comb};
  assign p1_sum__1013_comb = {{15{p1_add_135508_comb[16]}}, p1_add_135508_comb};
  assign p1_sum__835_comb = {{15{p1_add_135509_comb[16]}}, p1_add_135509_comb};
  assign p1_sum__836_comb = {{15{p1_add_135510_comb[16]}}, p1_add_135510_comb};
  assign p1_sum__837_comb = {{15{p1_add_135511_comb[16]}}, p1_add_135511_comb};
  assign p1_sum__838_comb = {{15{p1_add_135512_comb[16]}}, p1_add_135512_comb};
  assign p1_sum__993_comb = p1_sum__989_comb + p1_sum__990_comb;
  assign p1_sum__994_comb = p1_sum__991_comb + p1_sum__992_comb;
  assign p1_sum__965_comb = p1_sum__961_comb + p1_sum__962_comb;
  assign p1_sum__966_comb = p1_sum__963_comb + p1_sum__964_comb;
  assign p1_sum__930_comb = p1_sum__926_comb + p1_sum__927_comb;
  assign p1_sum__931_comb = p1_sum__928_comb + p1_sum__929_comb;
  assign p1_sum__888_comb = p1_sum__884_comb + p1_sum__885_comb;
  assign p1_sum__889_comb = p1_sum__886_comb + p1_sum__887_comb;
  assign p1_add_136113_comb = {{1{p1_smul_135161_comb[15]}}, p1_smul_135161_comb} + {{1{p1_smul_135162_comb[15]}}, p1_smul_135162_comb};
  assign p1_add_136114_comb = {{1{p1_sel_135163_comb[15]}}, p1_sel_135163_comb} + {{1{p1_sel_135164_comb[15]}}, p1_sel_135164_comb};
  assign p1_add_136115_comb = {{1{p1_sel_135165_comb[15]}}, p1_sel_135165_comb} + {{1{p1_sel_135166_comb[15]}}, p1_sel_135166_comb};
  assign p1_add_136116_comb = {{1{p1_smul_135167_comb[15]}}, p1_smul_135167_comb} + {{1{p1_smul_135168_comb[15]}}, p1_smul_135168_comb};
  assign p1_add_136117_comb = {{1{p1_smul_135169_comb[15]}}, p1_smul_135169_comb} + {{1{p1_smul_135170_comb[15]}}, p1_smul_135170_comb};
  assign p1_add_136118_comb = {{1{p1_sel_135171_comb[15]}}, p1_sel_135171_comb} + {{1{p1_sel_135172_comb[15]}}, p1_sel_135172_comb};
  assign p1_add_136119_comb = {{1{p1_sel_135173_comb[15]}}, p1_sel_135173_comb} + {{1{p1_sel_135174_comb[15]}}, p1_sel_135174_comb};
  assign p1_add_136120_comb = {{1{p1_smul_135175_comb[15]}}, p1_smul_135175_comb} + {{1{p1_smul_135176_comb[15]}}, p1_smul_135176_comb};
  assign p1_add_136121_comb = {{1{p1_smul_135177_comb[15]}}, p1_smul_135177_comb} + {{1{p1_smul_135178_comb[15]}}, p1_smul_135178_comb};
  assign p1_add_136122_comb = {{1{p1_sel_135179_comb[15]}}, p1_sel_135179_comb} + {{1{p1_sel_135180_comb[15]}}, p1_sel_135180_comb};
  assign p1_add_136123_comb = {{1{p1_sel_135181_comb[15]}}, p1_sel_135181_comb} + {{1{p1_sel_135182_comb[15]}}, p1_sel_135182_comb};
  assign p1_add_136124_comb = {{1{p1_smul_135183_comb[15]}}, p1_smul_135183_comb} + {{1{p1_smul_135184_comb[15]}}, p1_smul_135184_comb};
  assign p1_add_136125_comb = {{1{p1_smul_135185_comb[15]}}, p1_smul_135185_comb} + {{1{p1_smul_135186_comb[15]}}, p1_smul_135186_comb};
  assign p1_add_136126_comb = {{1{p1_sel_135187_comb[15]}}, p1_sel_135187_comb} + {{1{p1_sel_135188_comb[15]}}, p1_sel_135188_comb};
  assign p1_add_136127_comb = {{1{p1_sel_135189_comb[15]}}, p1_sel_135189_comb} + {{1{p1_sel_135190_comb[15]}}, p1_sel_135190_comb};
  assign p1_add_136128_comb = {{1{p1_smul_135191_comb[15]}}, p1_smul_135191_comb} + {{1{p1_smul_135192_comb[15]}}, p1_smul_135192_comb};
  assign p1_add_136129_comb = {{1{p1_sel_135193_comb[15]}}, p1_sel_135193_comb} + {{1{p1_sel_135194_comb[15]}}, p1_sel_135194_comb};
  assign p1_add_136130_comb = {{1{p1_sel_135195_comb[15]}}, p1_sel_135195_comb} + {{1{p1_sel_135196_comb[15]}}, p1_sel_135196_comb};
  assign p1_add_136131_comb = {{1{p1_sel_135197_comb[15]}}, p1_sel_135197_comb} + {{1{p1_sel_135198_comb[15]}}, p1_sel_135198_comb};
  assign p1_add_136132_comb = {{1{p1_sel_135199_comb[15]}}, p1_sel_135199_comb} + {{1{p1_sel_135200_comb[15]}}, p1_sel_135200_comb};
  assign p1_add_136133_comb = {{1{p1_sel_135201_comb[15]}}, p1_sel_135201_comb} + {{1{p1_sel_135202_comb[15]}}, p1_sel_135202_comb};
  assign p1_add_136134_comb = {{1{p1_sel_135203_comb[15]}}, p1_sel_135203_comb} + {{1{p1_sel_135204_comb[15]}}, p1_sel_135204_comb};
  assign p1_add_136135_comb = {{1{p1_sel_135205_comb[15]}}, p1_sel_135205_comb} + {{1{p1_sel_135206_comb[15]}}, p1_sel_135206_comb};
  assign p1_add_136136_comb = {{1{p1_sel_135207_comb[15]}}, p1_sel_135207_comb} + {{1{p1_sel_135208_comb[15]}}, p1_sel_135208_comb};
  assign p1_add_136137_comb = {{1{p1_sel_135209_comb[15]}}, p1_sel_135209_comb} + {{1{p1_sel_135210_comb[15]}}, p1_sel_135210_comb};
  assign p1_add_136138_comb = {{1{p1_sel_135211_comb[15]}}, p1_sel_135211_comb} + {{1{p1_sel_135212_comb[15]}}, p1_sel_135212_comb};
  assign p1_add_136139_comb = {{1{p1_sel_135213_comb[15]}}, p1_sel_135213_comb} + {{1{p1_sel_135214_comb[15]}}, p1_sel_135214_comb};
  assign p1_add_136140_comb = {{1{p1_sel_135215_comb[15]}}, p1_sel_135215_comb} + {{1{p1_sel_135216_comb[15]}}, p1_sel_135216_comb};
  assign p1_add_136141_comb = {{1{p1_sel_135217_comb[15]}}, p1_sel_135217_comb} + {{1{p1_sel_135218_comb[15]}}, p1_sel_135218_comb};
  assign p1_add_136142_comb = {{1{p1_sel_135219_comb[15]}}, p1_sel_135219_comb} + {{1{p1_sel_135220_comb[15]}}, p1_sel_135220_comb};
  assign p1_add_136143_comb = {{1{p1_sel_135221_comb[15]}}, p1_sel_135221_comb} + {{1{p1_sel_135222_comb[15]}}, p1_sel_135222_comb};
  assign p1_add_136144_comb = {{1{p1_sel_135223_comb[15]}}, p1_sel_135223_comb} + {{1{p1_sel_135224_comb[15]}}, p1_sel_135224_comb};
  assign p1_add_136145_comb = {{1{p1_smul_135225_comb[15]}}, p1_smul_135225_comb} + {{1{p1_sel_135226_comb[15]}}, p1_sel_135226_comb};
  assign p1_add_136146_comb = {{1{p1_smul_135227_comb[15]}}, p1_smul_135227_comb} + {{1{p1_sel_135228_comb[15]}}, p1_sel_135228_comb};
  assign p1_add_136147_comb = {{1{p1_sel_135229_comb[15]}}, p1_sel_135229_comb} + {{1{p1_smul_135230_comb[15]}}, p1_smul_135230_comb};
  assign p1_add_136148_comb = {{1{p1_sel_135231_comb[15]}}, p1_sel_135231_comb} + {{1{p1_smul_135232_comb[15]}}, p1_smul_135232_comb};
  assign p1_add_136149_comb = {{1{p1_smul_135233_comb[15]}}, p1_smul_135233_comb} + {{1{p1_sel_135234_comb[15]}}, p1_sel_135234_comb};
  assign p1_add_136150_comb = {{1{p1_smul_135235_comb[15]}}, p1_smul_135235_comb} + {{1{p1_sel_135236_comb[15]}}, p1_sel_135236_comb};
  assign p1_add_136151_comb = {{1{p1_sel_135237_comb[15]}}, p1_sel_135237_comb} + {{1{p1_smul_135238_comb[15]}}, p1_smul_135238_comb};
  assign p1_add_136152_comb = {{1{p1_sel_135239_comb[15]}}, p1_sel_135239_comb} + {{1{p1_smul_135240_comb[15]}}, p1_smul_135240_comb};
  assign p1_add_136153_comb = {{1{p1_smul_135241_comb[15]}}, p1_smul_135241_comb} + {{1{p1_sel_135242_comb[15]}}, p1_sel_135242_comb};
  assign p1_add_136154_comb = {{1{p1_smul_135243_comb[15]}}, p1_smul_135243_comb} + {{1{p1_sel_135244_comb[15]}}, p1_sel_135244_comb};
  assign p1_add_136155_comb = {{1{p1_sel_135245_comb[15]}}, p1_sel_135245_comb} + {{1{p1_smul_135246_comb[15]}}, p1_smul_135246_comb};
  assign p1_add_136156_comb = {{1{p1_sel_135247_comb[15]}}, p1_sel_135247_comb} + {{1{p1_smul_135248_comb[15]}}, p1_smul_135248_comb};
  assign p1_add_136157_comb = {{1{p1_smul_135249_comb[15]}}, p1_smul_135249_comb} + {{1{p1_sel_135250_comb[15]}}, p1_sel_135250_comb};
  assign p1_add_136158_comb = {{1{p1_smul_135251_comb[15]}}, p1_smul_135251_comb} + {{1{p1_sel_135252_comb[15]}}, p1_sel_135252_comb};
  assign p1_add_136159_comb = {{1{p1_sel_135253_comb[15]}}, p1_sel_135253_comb} + {{1{p1_smul_135254_comb[15]}}, p1_smul_135254_comb};
  assign p1_add_136160_comb = {{1{p1_sel_135255_comb[15]}}, p1_sel_135255_comb} + {{1{p1_smul_135256_comb[15]}}, p1_smul_135256_comb};
  assign p1_add_136161_comb = {{1{p1_smul_135257_comb[15]}}, p1_smul_135257_comb} + {{1{p1_smul_135258_comb[15]}}, p1_smul_135258_comb};
  assign p1_add_136162_comb = {{1{p1_smul_135259_comb[15]}}, p1_smul_135259_comb} + {{1{p1_smul_135260_comb[15]}}, p1_smul_135260_comb};
  assign p1_add_136163_comb = {{1{p1_smul_135261_comb[15]}}, p1_smul_135261_comb} + {{1{p1_smul_135262_comb[15]}}, p1_smul_135262_comb};
  assign p1_add_136164_comb = {{1{p1_smul_135263_comb[15]}}, p1_smul_135263_comb} + {{1{p1_smul_135264_comb[15]}}, p1_smul_135264_comb};
  assign p1_add_136165_comb = {{1{p1_smul_135265_comb[15]}}, p1_smul_135265_comb} + {{1{p1_smul_135266_comb[15]}}, p1_smul_135266_comb};
  assign p1_add_136166_comb = {{1{p1_smul_135267_comb[15]}}, p1_smul_135267_comb} + {{1{p1_smul_135268_comb[15]}}, p1_smul_135268_comb};
  assign p1_add_136167_comb = {{1{p1_smul_135269_comb[15]}}, p1_smul_135269_comb} + {{1{p1_smul_135270_comb[15]}}, p1_smul_135270_comb};
  assign p1_add_136168_comb = {{1{p1_smul_135271_comb[15]}}, p1_smul_135271_comb} + {{1{p1_smul_135272_comb[15]}}, p1_smul_135272_comb};
  assign p1_add_136169_comb = {{1{p1_smul_135273_comb[15]}}, p1_smul_135273_comb} + {{1{p1_smul_135274_comb[15]}}, p1_smul_135274_comb};
  assign p1_add_136170_comb = {{1{p1_smul_135275_comb[15]}}, p1_smul_135275_comb} + {{1{p1_smul_135276_comb[15]}}, p1_smul_135276_comb};
  assign p1_add_136171_comb = {{1{p1_smul_135277_comb[15]}}, p1_smul_135277_comb} + {{1{p1_smul_135278_comb[15]}}, p1_smul_135278_comb};
  assign p1_add_136172_comb = {{1{p1_smul_135279_comb[15]}}, p1_smul_135279_comb} + {{1{p1_smul_135280_comb[15]}}, p1_smul_135280_comb};
  assign p1_add_136173_comb = {{1{p1_smul_135281_comb[15]}}, p1_smul_135281_comb} + {{1{p1_smul_135282_comb[15]}}, p1_smul_135282_comb};
  assign p1_add_136174_comb = {{1{p1_smul_135283_comb[15]}}, p1_smul_135283_comb} + {{1{p1_smul_135284_comb[15]}}, p1_smul_135284_comb};
  assign p1_add_136175_comb = {{1{p1_smul_135285_comb[15]}}, p1_smul_135285_comb} + {{1{p1_smul_135286_comb[15]}}, p1_smul_135286_comb};
  assign p1_add_136176_comb = {{1{p1_smul_135287_comb[15]}}, p1_smul_135287_comb} + {{1{p1_smul_135288_comb[15]}}, p1_smul_135288_comb};
  assign p1_add_136177_comb = {{1{p1_sel_135289_comb[15]}}, p1_sel_135289_comb} + {{1{p1_smul_135290_comb[15]}}, p1_smul_135290_comb};
  assign p1_add_136178_comb = {{1{p1_sel_135291_comb[15]}}, p1_sel_135291_comb} + {{1{p1_smul_135292_comb[15]}}, p1_smul_135292_comb};
  assign p1_add_136179_comb = {{1{p1_smul_135293_comb[15]}}, p1_smul_135293_comb} + {{1{p1_sel_135294_comb[15]}}, p1_sel_135294_comb};
  assign p1_add_136180_comb = {{1{p1_smul_135295_comb[15]}}, p1_smul_135295_comb} + {{1{p1_sel_135296_comb[15]}}, p1_sel_135296_comb};
  assign p1_add_136181_comb = {{1{p1_sel_135297_comb[15]}}, p1_sel_135297_comb} + {{1{p1_smul_135298_comb[15]}}, p1_smul_135298_comb};
  assign p1_add_136182_comb = {{1{p1_sel_135299_comb[15]}}, p1_sel_135299_comb} + {{1{p1_smul_135300_comb[15]}}, p1_smul_135300_comb};
  assign p1_add_136183_comb = {{1{p1_smul_135301_comb[15]}}, p1_smul_135301_comb} + {{1{p1_sel_135302_comb[15]}}, p1_sel_135302_comb};
  assign p1_add_136184_comb = {{1{p1_smul_135303_comb[15]}}, p1_smul_135303_comb} + {{1{p1_sel_135304_comb[15]}}, p1_sel_135304_comb};
  assign p1_add_136185_comb = {{1{p1_sel_135305_comb[15]}}, p1_sel_135305_comb} + {{1{p1_smul_135306_comb[15]}}, p1_smul_135306_comb};
  assign p1_add_136186_comb = {{1{p1_sel_135307_comb[15]}}, p1_sel_135307_comb} + {{1{p1_smul_135308_comb[15]}}, p1_smul_135308_comb};
  assign p1_add_136187_comb = {{1{p1_smul_135309_comb[15]}}, p1_smul_135309_comb} + {{1{p1_sel_135310_comb[15]}}, p1_sel_135310_comb};
  assign p1_add_136188_comb = {{1{p1_smul_135311_comb[15]}}, p1_smul_135311_comb} + {{1{p1_sel_135312_comb[15]}}, p1_sel_135312_comb};
  assign p1_add_136189_comb = {{1{p1_sel_135313_comb[15]}}, p1_sel_135313_comb} + {{1{p1_smul_135314_comb[15]}}, p1_smul_135314_comb};
  assign p1_add_136190_comb = {{1{p1_sel_135315_comb[15]}}, p1_sel_135315_comb} + {{1{p1_smul_135316_comb[15]}}, p1_smul_135316_comb};
  assign p1_add_136191_comb = {{1{p1_smul_135317_comb[15]}}, p1_smul_135317_comb} + {{1{p1_sel_135318_comb[15]}}, p1_sel_135318_comb};
  assign p1_add_136192_comb = {{1{p1_smul_135319_comb[15]}}, p1_smul_135319_comb} + {{1{p1_sel_135320_comb[15]}}, p1_sel_135320_comb};
  assign p1_add_136193_comb = {{1{p1_sel_135321_comb[15]}}, p1_sel_135321_comb} + {{1{p1_sel_135322_comb[15]}}, p1_sel_135322_comb};
  assign p1_add_136194_comb = {{1{p1_sel_135323_comb[15]}}, p1_sel_135323_comb} + {{1{p1_sel_135324_comb[15]}}, p1_sel_135324_comb};
  assign p1_add_136195_comb = {{1{p1_sel_135325_comb[15]}}, p1_sel_135325_comb} + {{1{p1_sel_135326_comb[15]}}, p1_sel_135326_comb};
  assign p1_add_136196_comb = {{1{p1_sel_135327_comb[15]}}, p1_sel_135327_comb} + {{1{p1_sel_135328_comb[15]}}, p1_sel_135328_comb};
  assign p1_add_136197_comb = {{1{p1_sel_135329_comb[15]}}, p1_sel_135329_comb} + {{1{p1_sel_135330_comb[15]}}, p1_sel_135330_comb};
  assign p1_add_136198_comb = {{1{p1_sel_135331_comb[15]}}, p1_sel_135331_comb} + {{1{p1_sel_135332_comb[15]}}, p1_sel_135332_comb};
  assign p1_add_136199_comb = {{1{p1_sel_135333_comb[15]}}, p1_sel_135333_comb} + {{1{p1_sel_135334_comb[15]}}, p1_sel_135334_comb};
  assign p1_add_136200_comb = {{1{p1_sel_135335_comb[15]}}, p1_sel_135335_comb} + {{1{p1_sel_135336_comb[15]}}, p1_sel_135336_comb};
  assign p1_add_136201_comb = {{1{p1_sel_135337_comb[15]}}, p1_sel_135337_comb} + {{1{p1_sel_135338_comb[15]}}, p1_sel_135338_comb};
  assign p1_add_136202_comb = {{1{p1_sel_135339_comb[15]}}, p1_sel_135339_comb} + {{1{p1_sel_135340_comb[15]}}, p1_sel_135340_comb};
  assign p1_add_136203_comb = {{1{p1_sel_135341_comb[15]}}, p1_sel_135341_comb} + {{1{p1_sel_135342_comb[15]}}, p1_sel_135342_comb};
  assign p1_add_136204_comb = {{1{p1_sel_135343_comb[15]}}, p1_sel_135343_comb} + {{1{p1_sel_135344_comb[15]}}, p1_sel_135344_comb};
  assign p1_add_136205_comb = {{1{p1_sel_135345_comb[15]}}, p1_sel_135345_comb} + {{1{p1_sel_135346_comb[15]}}, p1_sel_135346_comb};
  assign p1_add_136206_comb = {{1{p1_sel_135347_comb[15]}}, p1_sel_135347_comb} + {{1{p1_sel_135348_comb[15]}}, p1_sel_135348_comb};
  assign p1_add_136207_comb = {{1{p1_sel_135349_comb[15]}}, p1_sel_135349_comb} + {{1{p1_sel_135350_comb[15]}}, p1_sel_135350_comb};
  assign p1_add_136208_comb = {{1{p1_sel_135351_comb[15]}}, p1_sel_135351_comb} + {{1{p1_sel_135352_comb[15]}}, p1_sel_135352_comb};
  assign p1_add_136209_comb = {{1{p1_sel_135353_comb[15]}}, p1_sel_135353_comb} + {{1{p1_sel_135354_comb[15]}}, p1_sel_135354_comb};
  assign p1_add_136210_comb = {{1{p1_smul_135355_comb[15]}}, p1_smul_135355_comb} + {{1{p1_smul_135356_comb[15]}}, p1_smul_135356_comb};
  assign p1_add_136211_comb = {{1{p1_smul_135357_comb[15]}}, p1_smul_135357_comb} + {{1{p1_smul_135358_comb[15]}}, p1_smul_135358_comb};
  assign p1_add_136212_comb = {{1{p1_sel_135359_comb[15]}}, p1_sel_135359_comb} + {{1{p1_sel_135360_comb[15]}}, p1_sel_135360_comb};
  assign p1_add_136213_comb = {{1{p1_sel_135361_comb[15]}}, p1_sel_135361_comb} + {{1{p1_sel_135362_comb[15]}}, p1_sel_135362_comb};
  assign p1_add_136214_comb = {{1{p1_smul_135363_comb[15]}}, p1_smul_135363_comb} + {{1{p1_smul_135364_comb[15]}}, p1_smul_135364_comb};
  assign p1_add_136215_comb = {{1{p1_smul_135365_comb[15]}}, p1_smul_135365_comb} + {{1{p1_smul_135366_comb[15]}}, p1_smul_135366_comb};
  assign p1_add_136216_comb = {{1{p1_sel_135367_comb[15]}}, p1_sel_135367_comb} + {{1{p1_sel_135368_comb[15]}}, p1_sel_135368_comb};
  assign p1_add_136217_comb = {{1{p1_sel_135369_comb[15]}}, p1_sel_135369_comb} + {{1{p1_sel_135370_comb[15]}}, p1_sel_135370_comb};
  assign p1_add_136218_comb = {{1{p1_smul_135371_comb[15]}}, p1_smul_135371_comb} + {{1{p1_smul_135372_comb[15]}}, p1_smul_135372_comb};
  assign p1_add_136219_comb = {{1{p1_smul_135373_comb[15]}}, p1_smul_135373_comb} + {{1{p1_smul_135374_comb[15]}}, p1_smul_135374_comb};
  assign p1_add_136220_comb = {{1{p1_sel_135375_comb[15]}}, p1_sel_135375_comb} + {{1{p1_sel_135376_comb[15]}}, p1_sel_135376_comb};
  assign p1_add_136221_comb = {{1{p1_sel_135377_comb[15]}}, p1_sel_135377_comb} + {{1{p1_sel_135378_comb[15]}}, p1_sel_135378_comb};
  assign p1_add_136222_comb = {{1{p1_smul_135379_comb[15]}}, p1_smul_135379_comb} + {{1{p1_smul_135380_comb[15]}}, p1_smul_135380_comb};
  assign p1_add_136223_comb = {{1{p1_smul_135381_comb[15]}}, p1_smul_135381_comb} + {{1{p1_smul_135382_comb[15]}}, p1_smul_135382_comb};
  assign p1_add_136224_comb = {{1{p1_sel_135383_comb[15]}}, p1_sel_135383_comb} + {{1{p1_sel_135384_comb[15]}}, p1_sel_135384_comb};
  assign p1_sum__1021_comb = p1_sum__1017_comb + p1_sum__1018_comb;
  assign p1_sum__1022_comb = p1_sum__1019_comb + p1_sum__1020_comb;
  assign p1_sum__783_comb = p1_sum__779_comb + p1_sum__780_comb;
  assign p1_sum__784_comb = p1_sum__781_comb + p1_sum__782_comb;
  assign p1_add_136229_comb = {{1{p1_smul_135393_comb[15]}}, p1_smul_135393_comb} + {{1{p1_smul_135394_comb[15]}}, p1_smul_135394_comb};
  assign p1_add_136230_comb = {{1{p1_sel_135395_comb[15]}}, p1_sel_135395_comb} + {{1{p1_sel_135396_comb[15]}}, p1_sel_135396_comb};
  assign p1_add_136231_comb = {{1{p1_sel_135397_comb[15]}}, p1_sel_135397_comb} + {{1{p1_sel_135398_comb[15]}}, p1_sel_135398_comb};
  assign p1_add_136232_comb = {{1{p1_smul_135399_comb[15]}}, p1_smul_135399_comb} + {{1{p1_smul_135400_comb[15]}}, p1_smul_135400_comb};
  assign p1_add_136233_comb = {{1{p1_smul_135401_comb[15]}}, p1_smul_135401_comb} + {{1{p1_smul_135402_comb[15]}}, p1_smul_135402_comb};
  assign p1_add_136234_comb = {{1{p1_sel_135403_comb[15]}}, p1_sel_135403_comb} + {{1{p1_sel_135404_comb[15]}}, p1_sel_135404_comb};
  assign p1_add_136235_comb = {{1{p1_sel_135405_comb[15]}}, p1_sel_135405_comb} + {{1{p1_sel_135406_comb[15]}}, p1_sel_135406_comb};
  assign p1_add_136236_comb = {{1{p1_smul_135407_comb[15]}}, p1_smul_135407_comb} + {{1{p1_smul_135408_comb[15]}}, p1_smul_135408_comb};
  assign p1_add_136237_comb = {{1{p1_sel_135409_comb[15]}}, p1_sel_135409_comb} + {{1{p1_sel_135410_comb[15]}}, p1_sel_135410_comb};
  assign p1_add_136238_comb = {{1{p1_sel_135411_comb[15]}}, p1_sel_135411_comb} + {{1{p1_sel_135412_comb[15]}}, p1_sel_135412_comb};
  assign p1_add_136239_comb = {{1{p1_sel_135413_comb[15]}}, p1_sel_135413_comb} + {{1{p1_sel_135414_comb[15]}}, p1_sel_135414_comb};
  assign p1_add_136240_comb = {{1{p1_sel_135415_comb[15]}}, p1_sel_135415_comb} + {{1{p1_sel_135416_comb[15]}}, p1_sel_135416_comb};
  assign p1_add_136241_comb = {{1{p1_sel_135417_comb[15]}}, p1_sel_135417_comb} + {{1{p1_sel_135418_comb[15]}}, p1_sel_135418_comb};
  assign p1_add_136242_comb = {{1{p1_sel_135419_comb[15]}}, p1_sel_135419_comb} + {{1{p1_sel_135420_comb[15]}}, p1_sel_135420_comb};
  assign p1_add_136243_comb = {{1{p1_sel_135421_comb[15]}}, p1_sel_135421_comb} + {{1{p1_sel_135422_comb[15]}}, p1_sel_135422_comb};
  assign p1_add_136244_comb = {{1{p1_sel_135423_comb[15]}}, p1_sel_135423_comb} + {{1{p1_sel_135424_comb[15]}}, p1_sel_135424_comb};
  assign p1_add_136245_comb = {{1{p1_smul_135425_comb[15]}}, p1_smul_135425_comb} + {{1{p1_sel_135426_comb[15]}}, p1_sel_135426_comb};
  assign p1_add_136246_comb = {{1{p1_smul_135427_comb[15]}}, p1_smul_135427_comb} + {{1{p1_sel_135428_comb[15]}}, p1_sel_135428_comb};
  assign p1_add_136247_comb = {{1{p1_sel_135429_comb[15]}}, p1_sel_135429_comb} + {{1{p1_smul_135430_comb[15]}}, p1_smul_135430_comb};
  assign p1_add_136248_comb = {{1{p1_sel_135431_comb[15]}}, p1_sel_135431_comb} + {{1{p1_smul_135432_comb[15]}}, p1_smul_135432_comb};
  assign p1_add_136249_comb = {{1{p1_smul_135433_comb[15]}}, p1_smul_135433_comb} + {{1{p1_sel_135434_comb[15]}}, p1_sel_135434_comb};
  assign p1_add_136250_comb = {{1{p1_smul_135435_comb[15]}}, p1_smul_135435_comb} + {{1{p1_sel_135436_comb[15]}}, p1_sel_135436_comb};
  assign p1_add_136251_comb = {{1{p1_sel_135437_comb[15]}}, p1_sel_135437_comb} + {{1{p1_smul_135438_comb[15]}}, p1_smul_135438_comb};
  assign p1_add_136252_comb = {{1{p1_sel_135439_comb[15]}}, p1_sel_135439_comb} + {{1{p1_smul_135440_comb[15]}}, p1_smul_135440_comb};
  assign p1_add_136253_comb = {{1{p1_smul_135441_comb[15]}}, p1_smul_135441_comb} + {{1{p1_smul_135442_comb[15]}}, p1_smul_135442_comb};
  assign p1_add_136254_comb = {{1{p1_smul_135443_comb[15]}}, p1_smul_135443_comb} + {{1{p1_smul_135444_comb[15]}}, p1_smul_135444_comb};
  assign p1_add_136255_comb = {{1{p1_smul_135445_comb[15]}}, p1_smul_135445_comb} + {{1{p1_smul_135446_comb[15]}}, p1_smul_135446_comb};
  assign p1_add_136256_comb = {{1{p1_smul_135447_comb[15]}}, p1_smul_135447_comb} + {{1{p1_smul_135448_comb[15]}}, p1_smul_135448_comb};
  assign p1_add_136257_comb = {{1{p1_smul_135449_comb[15]}}, p1_smul_135449_comb} + {{1{p1_smul_135450_comb[15]}}, p1_smul_135450_comb};
  assign p1_add_136258_comb = {{1{p1_smul_135451_comb[15]}}, p1_smul_135451_comb} + {{1{p1_smul_135452_comb[15]}}, p1_smul_135452_comb};
  assign p1_add_136259_comb = {{1{p1_smul_135453_comb[15]}}, p1_smul_135453_comb} + {{1{p1_smul_135454_comb[15]}}, p1_smul_135454_comb};
  assign p1_add_136260_comb = {{1{p1_smul_135455_comb[15]}}, p1_smul_135455_comb} + {{1{p1_smul_135456_comb[15]}}, p1_smul_135456_comb};
  assign p1_add_136261_comb = {{1{p1_sel_135457_comb[15]}}, p1_sel_135457_comb} + {{1{p1_smul_135458_comb[15]}}, p1_smul_135458_comb};
  assign p1_add_136262_comb = {{1{p1_sel_135459_comb[15]}}, p1_sel_135459_comb} + {{1{p1_smul_135460_comb[15]}}, p1_smul_135460_comb};
  assign p1_add_136263_comb = {{1{p1_smul_135461_comb[15]}}, p1_smul_135461_comb} + {{1{p1_sel_135462_comb[15]}}, p1_sel_135462_comb};
  assign p1_add_136264_comb = {{1{p1_smul_135463_comb[15]}}, p1_smul_135463_comb} + {{1{p1_sel_135464_comb[15]}}, p1_sel_135464_comb};
  assign p1_add_136265_comb = {{1{p1_sel_135465_comb[15]}}, p1_sel_135465_comb} + {{1{p1_smul_135466_comb[15]}}, p1_smul_135466_comb};
  assign p1_add_136266_comb = {{1{p1_sel_135467_comb[15]}}, p1_sel_135467_comb} + {{1{p1_smul_135468_comb[15]}}, p1_smul_135468_comb};
  assign p1_add_136267_comb = {{1{p1_smul_135469_comb[15]}}, p1_smul_135469_comb} + {{1{p1_sel_135470_comb[15]}}, p1_sel_135470_comb};
  assign p1_add_136268_comb = {{1{p1_smul_135471_comb[15]}}, p1_smul_135471_comb} + {{1{p1_sel_135472_comb[15]}}, p1_sel_135472_comb};
  assign p1_add_136269_comb = {{1{p1_sel_135473_comb[15]}}, p1_sel_135473_comb} + {{1{p1_sel_135474_comb[15]}}, p1_sel_135474_comb};
  assign p1_add_136270_comb = {{1{p1_sel_135475_comb[15]}}, p1_sel_135475_comb} + {{1{p1_sel_135476_comb[15]}}, p1_sel_135476_comb};
  assign p1_add_136271_comb = {{1{p1_sel_135477_comb[15]}}, p1_sel_135477_comb} + {{1{p1_sel_135478_comb[15]}}, p1_sel_135478_comb};
  assign p1_add_136272_comb = {{1{p1_sel_135479_comb[15]}}, p1_sel_135479_comb} + {{1{p1_sel_135480_comb[15]}}, p1_sel_135480_comb};
  assign p1_add_136273_comb = {{1{p1_sel_135481_comb[15]}}, p1_sel_135481_comb} + {{1{p1_sel_135482_comb[15]}}, p1_sel_135482_comb};
  assign p1_add_136274_comb = {{1{p1_sel_135483_comb[15]}}, p1_sel_135483_comb} + {{1{p1_sel_135484_comb[15]}}, p1_sel_135484_comb};
  assign p1_add_136275_comb = {{1{p1_sel_135485_comb[15]}}, p1_sel_135485_comb} + {{1{p1_sel_135486_comb[15]}}, p1_sel_135486_comb};
  assign p1_add_136276_comb = {{1{p1_sel_135487_comb[15]}}, p1_sel_135487_comb} + {{1{p1_sel_135488_comb[15]}}, p1_sel_135488_comb};
  assign p1_add_136277_comb = {{1{p1_sel_135489_comb[15]}}, p1_sel_135489_comb} + {{1{p1_sel_135490_comb[15]}}, p1_sel_135490_comb};
  assign p1_add_136278_comb = {{1{p1_smul_135491_comb[15]}}, p1_smul_135491_comb} + {{1{p1_smul_135492_comb[15]}}, p1_smul_135492_comb};
  assign p1_add_136279_comb = {{1{p1_smul_135493_comb[15]}}, p1_smul_135493_comb} + {{1{p1_smul_135494_comb[15]}}, p1_smul_135494_comb};
  assign p1_add_136280_comb = {{1{p1_sel_135495_comb[15]}}, p1_sel_135495_comb} + {{1{p1_sel_135496_comb[15]}}, p1_sel_135496_comb};
  assign p1_add_136281_comb = {{1{p1_sel_135497_comb[15]}}, p1_sel_135497_comb} + {{1{p1_sel_135498_comb[15]}}, p1_sel_135498_comb};
  assign p1_add_136282_comb = {{1{p1_smul_135499_comb[15]}}, p1_smul_135499_comb} + {{1{p1_smul_135500_comb[15]}}, p1_smul_135500_comb};
  assign p1_add_136283_comb = {{1{p1_smul_135501_comb[15]}}, p1_smul_135501_comb} + {{1{p1_smul_135502_comb[15]}}, p1_smul_135502_comb};
  assign p1_add_136284_comb = {{1{p1_sel_135503_comb[15]}}, p1_sel_135503_comb} + {{1{p1_sel_135504_comb[15]}}, p1_sel_135504_comb};
  assign p1_sum__1014_comb = p1_sum__1010_comb + p1_sum__1011_comb;
  assign p1_sum__1015_comb = p1_sum__1012_comb + p1_sum__1013_comb;
  assign p1_sum__839_comb = p1_sum__835_comb + p1_sum__836_comb;
  assign p1_sum__840_comb = p1_sum__837_comb + p1_sum__838_comb;
  assign p1_add_136289_comb = {{1{p1_smul_135513_comb[15]}}, p1_smul_135513_comb} + {{1{p1_smul_135514_comb[15]}}, p1_smul_135514_comb};
  assign p1_add_136290_comb = {{1{p1_sel_135515_comb[15]}}, p1_sel_135515_comb} + {{1{p1_sel_135516_comb[15]}}, p1_sel_135516_comb};
  assign p1_add_136291_comb = {{1{p1_sel_135517_comb[15]}}, p1_sel_135517_comb} + {{1{p1_sel_135518_comb[15]}}, p1_sel_135518_comb};
  assign p1_add_136292_comb = {{1{p1_smul_135519_comb[15]}}, p1_smul_135519_comb} + {{1{p1_smul_135520_comb[15]}}, p1_smul_135520_comb};
  assign p1_add_136293_comb = {{1{p1_smul_135521_comb[15]}}, p1_smul_135521_comb} + {{1{p1_smul_135522_comb[15]}}, p1_smul_135522_comb};
  assign p1_add_136294_comb = {{1{p1_sel_135523_comb[15]}}, p1_sel_135523_comb} + {{1{p1_sel_135524_comb[15]}}, p1_sel_135524_comb};
  assign p1_add_136295_comb = {{1{p1_sel_135525_comb[15]}}, p1_sel_135525_comb} + {{1{p1_sel_135526_comb[15]}}, p1_sel_135526_comb};
  assign p1_add_136296_comb = {{1{p1_smul_135527_comb[15]}}, p1_smul_135527_comb} + {{1{p1_smul_135528_comb[15]}}, p1_smul_135528_comb};
  assign p1_add_136297_comb = {{1{p1_sel_135529_comb[15]}}, p1_sel_135529_comb} + {{1{p1_sel_135530_comb[15]}}, p1_sel_135530_comb};
  assign p1_add_136298_comb = {{1{p1_sel_135531_comb[15]}}, p1_sel_135531_comb} + {{1{p1_sel_135532_comb[15]}}, p1_sel_135532_comb};
  assign p1_add_136299_comb = {{1{p1_sel_135533_comb[15]}}, p1_sel_135533_comb} + {{1{p1_sel_135534_comb[15]}}, p1_sel_135534_comb};
  assign p1_add_136300_comb = {{1{p1_sel_135535_comb[15]}}, p1_sel_135535_comb} + {{1{p1_sel_135536_comb[15]}}, p1_sel_135536_comb};
  assign p1_add_136301_comb = {{1{p1_sel_135537_comb[15]}}, p1_sel_135537_comb} + {{1{p1_sel_135538_comb[15]}}, p1_sel_135538_comb};
  assign p1_add_136302_comb = {{1{p1_sel_135539_comb[15]}}, p1_sel_135539_comb} + {{1{p1_sel_135540_comb[15]}}, p1_sel_135540_comb};
  assign p1_add_136303_comb = {{1{p1_sel_135541_comb[15]}}, p1_sel_135541_comb} + {{1{p1_sel_135542_comb[15]}}, p1_sel_135542_comb};
  assign p1_add_136304_comb = {{1{p1_sel_135543_comb[15]}}, p1_sel_135543_comb} + {{1{p1_sel_135544_comb[15]}}, p1_sel_135544_comb};
  assign p1_add_136305_comb = {{1{p1_smul_135545_comb[15]}}, p1_smul_135545_comb} + {{1{p1_sel_135546_comb[15]}}, p1_sel_135546_comb};
  assign p1_add_136306_comb = {{1{p1_smul_135547_comb[15]}}, p1_smul_135547_comb} + {{1{p1_sel_135548_comb[15]}}, p1_sel_135548_comb};
  assign p1_add_136307_comb = {{1{p1_sel_135549_comb[15]}}, p1_sel_135549_comb} + {{1{p1_smul_135550_comb[15]}}, p1_smul_135550_comb};
  assign p1_add_136308_comb = {{1{p1_sel_135551_comb[15]}}, p1_sel_135551_comb} + {{1{p1_smul_135552_comb[15]}}, p1_smul_135552_comb};
  assign p1_add_136309_comb = {{1{p1_smul_135553_comb[15]}}, p1_smul_135553_comb} + {{1{p1_sel_135554_comb[15]}}, p1_sel_135554_comb};
  assign p1_add_136310_comb = {{1{p1_smul_135555_comb[15]}}, p1_smul_135555_comb} + {{1{p1_sel_135556_comb[15]}}, p1_sel_135556_comb};
  assign p1_add_136311_comb = {{1{p1_sel_135557_comb[15]}}, p1_sel_135557_comb} + {{1{p1_smul_135558_comb[15]}}, p1_smul_135558_comb};
  assign p1_add_136312_comb = {{1{p1_sel_135559_comb[15]}}, p1_sel_135559_comb} + {{1{p1_smul_135560_comb[15]}}, p1_smul_135560_comb};
  assign p1_add_136313_comb = {{1{p1_smul_135561_comb[15]}}, p1_smul_135561_comb} + {{1{p1_smul_135562_comb[15]}}, p1_smul_135562_comb};
  assign p1_add_136314_comb = {{1{p1_smul_135563_comb[15]}}, p1_smul_135563_comb} + {{1{p1_smul_135564_comb[15]}}, p1_smul_135564_comb};
  assign p1_add_136315_comb = {{1{p1_smul_135565_comb[15]}}, p1_smul_135565_comb} + {{1{p1_smul_135566_comb[15]}}, p1_smul_135566_comb};
  assign p1_add_136316_comb = {{1{p1_smul_135567_comb[15]}}, p1_smul_135567_comb} + {{1{p1_smul_135568_comb[15]}}, p1_smul_135568_comb};
  assign p1_add_136317_comb = {{1{p1_smul_135569_comb[15]}}, p1_smul_135569_comb} + {{1{p1_smul_135570_comb[15]}}, p1_smul_135570_comb};
  assign p1_add_136318_comb = {{1{p1_smul_135571_comb[15]}}, p1_smul_135571_comb} + {{1{p1_smul_135572_comb[15]}}, p1_smul_135572_comb};
  assign p1_add_136319_comb = {{1{p1_smul_135573_comb[15]}}, p1_smul_135573_comb} + {{1{p1_smul_135574_comb[15]}}, p1_smul_135574_comb};
  assign p1_add_136320_comb = {{1{p1_smul_135575_comb[15]}}, p1_smul_135575_comb} + {{1{p1_smul_135576_comb[15]}}, p1_smul_135576_comb};
  assign p1_add_136321_comb = {{1{p1_sel_135577_comb[15]}}, p1_sel_135577_comb} + {{1{p1_smul_135578_comb[15]}}, p1_smul_135578_comb};
  assign p1_add_136322_comb = {{1{p1_sel_135579_comb[15]}}, p1_sel_135579_comb} + {{1{p1_smul_135580_comb[15]}}, p1_smul_135580_comb};
  assign p1_add_136323_comb = {{1{p1_smul_135581_comb[15]}}, p1_smul_135581_comb} + {{1{p1_sel_135582_comb[15]}}, p1_sel_135582_comb};
  assign p1_add_136324_comb = {{1{p1_smul_135583_comb[15]}}, p1_smul_135583_comb} + {{1{p1_sel_135584_comb[15]}}, p1_sel_135584_comb};
  assign p1_add_136325_comb = {{1{p1_sel_135585_comb[15]}}, p1_sel_135585_comb} + {{1{p1_smul_135586_comb[15]}}, p1_smul_135586_comb};
  assign p1_add_136326_comb = {{1{p1_sel_135587_comb[15]}}, p1_sel_135587_comb} + {{1{p1_smul_135588_comb[15]}}, p1_smul_135588_comb};
  assign p1_add_136327_comb = {{1{p1_smul_135589_comb[15]}}, p1_smul_135589_comb} + {{1{p1_sel_135590_comb[15]}}, p1_sel_135590_comb};
  assign p1_add_136328_comb = {{1{p1_smul_135591_comb[15]}}, p1_smul_135591_comb} + {{1{p1_sel_135592_comb[15]}}, p1_sel_135592_comb};
  assign p1_add_136329_comb = {{1{p1_sel_135593_comb[15]}}, p1_sel_135593_comb} + {{1{p1_sel_135594_comb[15]}}, p1_sel_135594_comb};
  assign p1_add_136330_comb = {{1{p1_sel_135595_comb[15]}}, p1_sel_135595_comb} + {{1{p1_sel_135596_comb[15]}}, p1_sel_135596_comb};
  assign p1_add_136331_comb = {{1{p1_sel_135597_comb[15]}}, p1_sel_135597_comb} + {{1{p1_sel_135598_comb[15]}}, p1_sel_135598_comb};
  assign p1_add_136332_comb = {{1{p1_sel_135599_comb[15]}}, p1_sel_135599_comb} + {{1{p1_sel_135600_comb[15]}}, p1_sel_135600_comb};
  assign p1_add_136333_comb = {{1{p1_sel_135601_comb[15]}}, p1_sel_135601_comb} + {{1{p1_sel_135602_comb[15]}}, p1_sel_135602_comb};
  assign p1_add_136334_comb = {{1{p1_sel_135603_comb[15]}}, p1_sel_135603_comb} + {{1{p1_sel_135604_comb[15]}}, p1_sel_135604_comb};
  assign p1_add_136335_comb = {{1{p1_sel_135605_comb[15]}}, p1_sel_135605_comb} + {{1{p1_sel_135606_comb[15]}}, p1_sel_135606_comb};
  assign p1_add_136336_comb = {{1{p1_sel_135607_comb[15]}}, p1_sel_135607_comb} + {{1{p1_sel_135608_comb[15]}}, p1_sel_135608_comb};
  assign p1_add_136337_comb = {{1{p1_sel_135609_comb[15]}}, p1_sel_135609_comb} + {{1{p1_sel_135610_comb[15]}}, p1_sel_135610_comb};
  assign p1_add_136338_comb = {{1{p1_smul_135611_comb[15]}}, p1_smul_135611_comb} + {{1{p1_smul_135612_comb[15]}}, p1_smul_135612_comb};
  assign p1_add_136339_comb = {{1{p1_smul_135613_comb[15]}}, p1_smul_135613_comb} + {{1{p1_smul_135614_comb[15]}}, p1_smul_135614_comb};
  assign p1_add_136340_comb = {{1{p1_sel_135615_comb[15]}}, p1_sel_135615_comb} + {{1{p1_sel_135616_comb[15]}}, p1_sel_135616_comb};
  assign p1_add_136341_comb = {{1{p1_sel_135617_comb[15]}}, p1_sel_135617_comb} + {{1{p1_sel_135618_comb[15]}}, p1_sel_135618_comb};
  assign p1_add_136342_comb = {{1{p1_smul_135619_comb[15]}}, p1_smul_135619_comb} + {{1{p1_smul_135620_comb[15]}}, p1_smul_135620_comb};
  assign p1_add_136343_comb = {{1{p1_smul_135621_comb[15]}}, p1_smul_135621_comb} + {{1{p1_smul_135622_comb[15]}}, p1_smul_135622_comb};
  assign p1_add_136344_comb = {{1{p1_sel_135623_comb[15]}}, p1_sel_135623_comb} + {{1{p1_sel_135624_comb[15]}}, p1_sel_135624_comb};
  assign p1_sum__995_comb = p1_sum__993_comb + p1_sum__994_comb;
  assign p1_sum__967_comb = p1_sum__965_comb + p1_sum__966_comb;
  assign p1_sum__932_comb = p1_sum__930_comb + p1_sum__931_comb;
  assign p1_sum__890_comb = p1_sum__888_comb + p1_sum__889_comb;
  assign p1_sum__1784_comb = {{8{p1_add_136113_comb[16]}}, p1_add_136113_comb};
  assign p1_sum__1785_comb = {{8{p1_add_136114_comb[16]}}, p1_add_136114_comb};
  assign p1_sum__1786_comb = {{8{p1_add_136115_comb[16]}}, p1_add_136115_comb};
  assign p1_sum__1787_comb = {{8{p1_add_136116_comb[16]}}, p1_add_136116_comb};
  assign p1_sum__1768_comb = {{8{p1_add_136117_comb[16]}}, p1_add_136117_comb};
  assign p1_sum__1769_comb = {{8{p1_add_136118_comb[16]}}, p1_add_136118_comb};
  assign p1_sum__1770_comb = {{8{p1_add_136119_comb[16]}}, p1_add_136119_comb};
  assign p1_sum__1771_comb = {{8{p1_add_136120_comb[16]}}, p1_add_136120_comb};
  assign p1_sum__1748_comb = {{8{p1_add_136121_comb[16]}}, p1_add_136121_comb};
  assign p1_sum__1749_comb = {{8{p1_add_136122_comb[16]}}, p1_add_136122_comb};
  assign p1_sum__1750_comb = {{8{p1_add_136123_comb[16]}}, p1_add_136123_comb};
  assign p1_sum__1751_comb = {{8{p1_add_136124_comb[16]}}, p1_add_136124_comb};
  assign p1_sum__1724_comb = {{8{p1_add_136125_comb[16]}}, p1_add_136125_comb};
  assign p1_sum__1725_comb = {{8{p1_add_136126_comb[16]}}, p1_add_136126_comb};
  assign p1_sum__1726_comb = {{8{p1_add_136127_comb[16]}}, p1_add_136127_comb};
  assign p1_sum__1727_comb = {{8{p1_add_136128_comb[16]}}, p1_add_136128_comb};
  assign p1_sum__1772_comb = {{8{p1_add_136129_comb[16]}}, p1_add_136129_comb};
  assign p1_sum__1773_comb = {{8{p1_add_136130_comb[16]}}, p1_add_136130_comb};
  assign p1_sum__1774_comb = {{8{p1_add_136131_comb[16]}}, p1_add_136131_comb};
  assign p1_sum__1775_comb = {{8{p1_add_136132_comb[16]}}, p1_add_136132_comb};
  assign p1_sum__1752_comb = {{8{p1_add_136133_comb[16]}}, p1_add_136133_comb};
  assign p1_sum__1753_comb = {{8{p1_add_136134_comb[16]}}, p1_add_136134_comb};
  assign p1_sum__1754_comb = {{8{p1_add_136135_comb[16]}}, p1_add_136135_comb};
  assign p1_sum__1755_comb = {{8{p1_add_136136_comb[16]}}, p1_add_136136_comb};
  assign p1_sum__1728_comb = {{8{p1_add_136137_comb[16]}}, p1_add_136137_comb};
  assign p1_sum__1729_comb = {{8{p1_add_136138_comb[16]}}, p1_add_136138_comb};
  assign p1_sum__1730_comb = {{8{p1_add_136139_comb[16]}}, p1_add_136139_comb};
  assign p1_sum__1731_comb = {{8{p1_add_136140_comb[16]}}, p1_add_136140_comb};
  assign p1_sum__1700_comb = {{8{p1_add_136141_comb[16]}}, p1_add_136141_comb};
  assign p1_sum__1701_comb = {{8{p1_add_136142_comb[16]}}, p1_add_136142_comb};
  assign p1_sum__1702_comb = {{8{p1_add_136143_comb[16]}}, p1_add_136143_comb};
  assign p1_sum__1703_comb = {{8{p1_add_136144_comb[16]}}, p1_add_136144_comb};
  assign p1_sum__1756_comb = {{8{p1_add_136145_comb[16]}}, p1_add_136145_comb};
  assign p1_sum__1757_comb = {{8{p1_add_136146_comb[16]}}, p1_add_136146_comb};
  assign p1_sum__1758_comb = {{8{p1_add_136147_comb[16]}}, p1_add_136147_comb};
  assign p1_sum__1759_comb = {{8{p1_add_136148_comb[16]}}, p1_add_136148_comb};
  assign p1_sum__1732_comb = {{8{p1_add_136149_comb[16]}}, p1_add_136149_comb};
  assign p1_sum__1733_comb = {{8{p1_add_136150_comb[16]}}, p1_add_136150_comb};
  assign p1_sum__1734_comb = {{8{p1_add_136151_comb[16]}}, p1_add_136151_comb};
  assign p1_sum__1735_comb = {{8{p1_add_136152_comb[16]}}, p1_add_136152_comb};
  assign p1_sum__1704_comb = {{8{p1_add_136153_comb[16]}}, p1_add_136153_comb};
  assign p1_sum__1705_comb = {{8{p1_add_136154_comb[16]}}, p1_add_136154_comb};
  assign p1_sum__1706_comb = {{8{p1_add_136155_comb[16]}}, p1_add_136155_comb};
  assign p1_sum__1707_comb = {{8{p1_add_136156_comb[16]}}, p1_add_136156_comb};
  assign p1_sum__1676_comb = {{8{p1_add_136157_comb[16]}}, p1_add_136157_comb};
  assign p1_sum__1677_comb = {{8{p1_add_136158_comb[16]}}, p1_add_136158_comb};
  assign p1_sum__1678_comb = {{8{p1_add_136159_comb[16]}}, p1_add_136159_comb};
  assign p1_sum__1679_comb = {{8{p1_add_136160_comb[16]}}, p1_add_136160_comb};
  assign p1_sum__1736_comb = {{8{p1_add_136161_comb[16]}}, p1_add_136161_comb};
  assign p1_sum__1737_comb = {{8{p1_add_136162_comb[16]}}, p1_add_136162_comb};
  assign p1_sum__1738_comb = {{8{p1_add_136163_comb[16]}}, p1_add_136163_comb};
  assign p1_sum__1739_comb = {{8{p1_add_136164_comb[16]}}, p1_add_136164_comb};
  assign p1_sum__1708_comb = {{8{p1_add_136165_comb[16]}}, p1_add_136165_comb};
  assign p1_sum__1709_comb = {{8{p1_add_136166_comb[16]}}, p1_add_136166_comb};
  assign p1_sum__1710_comb = {{8{p1_add_136167_comb[16]}}, p1_add_136167_comb};
  assign p1_sum__1711_comb = {{8{p1_add_136168_comb[16]}}, p1_add_136168_comb};
  assign p1_sum__1680_comb = {{8{p1_add_136169_comb[16]}}, p1_add_136169_comb};
  assign p1_sum__1681_comb = {{8{p1_add_136170_comb[16]}}, p1_add_136170_comb};
  assign p1_sum__1682_comb = {{8{p1_add_136171_comb[16]}}, p1_add_136171_comb};
  assign p1_sum__1683_comb = {{8{p1_add_136172_comb[16]}}, p1_add_136172_comb};
  assign p1_sum__1652_comb = {{8{p1_add_136173_comb[16]}}, p1_add_136173_comb};
  assign p1_sum__1653_comb = {{8{p1_add_136174_comb[16]}}, p1_add_136174_comb};
  assign p1_sum__1654_comb = {{8{p1_add_136175_comb[16]}}, p1_add_136175_comb};
  assign p1_sum__1655_comb = {{8{p1_add_136176_comb[16]}}, p1_add_136176_comb};
  assign p1_sum__1712_comb = {{8{p1_add_136177_comb[16]}}, p1_add_136177_comb};
  assign p1_sum__1713_comb = {{8{p1_add_136178_comb[16]}}, p1_add_136178_comb};
  assign p1_sum__1714_comb = {{8{p1_add_136179_comb[16]}}, p1_add_136179_comb};
  assign p1_sum__1715_comb = {{8{p1_add_136180_comb[16]}}, p1_add_136180_comb};
  assign p1_sum__1684_comb = {{8{p1_add_136181_comb[16]}}, p1_add_136181_comb};
  assign p1_sum__1685_comb = {{8{p1_add_136182_comb[16]}}, p1_add_136182_comb};
  assign p1_sum__1686_comb = {{8{p1_add_136183_comb[16]}}, p1_add_136183_comb};
  assign p1_sum__1687_comb = {{8{p1_add_136184_comb[16]}}, p1_add_136184_comb};
  assign p1_sum__1656_comb = {{8{p1_add_136185_comb[16]}}, p1_add_136185_comb};
  assign p1_sum__1657_comb = {{8{p1_add_136186_comb[16]}}, p1_add_136186_comb};
  assign p1_sum__1658_comb = {{8{p1_add_136187_comb[16]}}, p1_add_136187_comb};
  assign p1_sum__1659_comb = {{8{p1_add_136188_comb[16]}}, p1_add_136188_comb};
  assign p1_sum__1632_comb = {{8{p1_add_136189_comb[16]}}, p1_add_136189_comb};
  assign p1_sum__1633_comb = {{8{p1_add_136190_comb[16]}}, p1_add_136190_comb};
  assign p1_sum__1634_comb = {{8{p1_add_136191_comb[16]}}, p1_add_136191_comb};
  assign p1_sum__1635_comb = {{8{p1_add_136192_comb[16]}}, p1_add_136192_comb};
  assign p1_sum__1688_comb = {{8{p1_add_136193_comb[16]}}, p1_add_136193_comb};
  assign p1_sum__1689_comb = {{8{p1_add_136194_comb[16]}}, p1_add_136194_comb};
  assign p1_sum__1690_comb = {{8{p1_add_136195_comb[16]}}, p1_add_136195_comb};
  assign p1_sum__1691_comb = {{8{p1_add_136196_comb[16]}}, p1_add_136196_comb};
  assign p1_sum__1660_comb = {{8{p1_add_136197_comb[16]}}, p1_add_136197_comb};
  assign p1_sum__1661_comb = {{8{p1_add_136198_comb[16]}}, p1_add_136198_comb};
  assign p1_sum__1662_comb = {{8{p1_add_136199_comb[16]}}, p1_add_136199_comb};
  assign p1_sum__1663_comb = {{8{p1_add_136200_comb[16]}}, p1_add_136200_comb};
  assign p1_sum__1636_comb = {{8{p1_add_136201_comb[16]}}, p1_add_136201_comb};
  assign p1_sum__1637_comb = {{8{p1_add_136202_comb[16]}}, p1_add_136202_comb};
  assign p1_sum__1638_comb = {{8{p1_add_136203_comb[16]}}, p1_add_136203_comb};
  assign p1_sum__1639_comb = {{8{p1_add_136204_comb[16]}}, p1_add_136204_comb};
  assign p1_sum__1616_comb = {{8{p1_add_136205_comb[16]}}, p1_add_136205_comb};
  assign p1_sum__1617_comb = {{8{p1_add_136206_comb[16]}}, p1_add_136206_comb};
  assign p1_sum__1618_comb = {{8{p1_add_136207_comb[16]}}, p1_add_136207_comb};
  assign p1_sum__1619_comb = {{8{p1_add_136208_comb[16]}}, p1_add_136208_comb};
  assign p1_sum__1664_comb = {{8{p1_add_136209_comb[16]}}, p1_add_136209_comb};
  assign p1_sum__1665_comb = {{8{p1_add_136210_comb[16]}}, p1_add_136210_comb};
  assign p1_sum__1666_comb = {{8{p1_add_136211_comb[16]}}, p1_add_136211_comb};
  assign p1_sum__1667_comb = {{8{p1_add_136212_comb[16]}}, p1_add_136212_comb};
  assign p1_sum__1640_comb = {{8{p1_add_136213_comb[16]}}, p1_add_136213_comb};
  assign p1_sum__1641_comb = {{8{p1_add_136214_comb[16]}}, p1_add_136214_comb};
  assign p1_sum__1642_comb = {{8{p1_add_136215_comb[16]}}, p1_add_136215_comb};
  assign p1_sum__1643_comb = {{8{p1_add_136216_comb[16]}}, p1_add_136216_comb};
  assign p1_sum__1620_comb = {{8{p1_add_136217_comb[16]}}, p1_add_136217_comb};
  assign p1_sum__1621_comb = {{8{p1_add_136218_comb[16]}}, p1_add_136218_comb};
  assign p1_sum__1622_comb = {{8{p1_add_136219_comb[16]}}, p1_add_136219_comb};
  assign p1_sum__1623_comb = {{8{p1_add_136220_comb[16]}}, p1_add_136220_comb};
  assign p1_sum__1604_comb = {{8{p1_add_136221_comb[16]}}, p1_add_136221_comb};
  assign p1_sum__1605_comb = {{8{p1_add_136222_comb[16]}}, p1_add_136222_comb};
  assign p1_sum__1606_comb = {{8{p1_add_136223_comb[16]}}, p1_add_136223_comb};
  assign p1_sum__1607_comb = {{8{p1_add_136224_comb[16]}}, p1_add_136224_comb};
  assign p1_sum__1023_comb = p1_sum__1021_comb + p1_sum__1022_comb;
  assign p1_sum__785_comb = p1_sum__783_comb + p1_sum__784_comb;
  assign p1_sum__1804_comb = {{8{p1_add_136229_comb[16]}}, p1_add_136229_comb};
  assign p1_sum__1805_comb = {{8{p1_add_136230_comb[16]}}, p1_add_136230_comb};
  assign p1_sum__1806_comb = {{8{p1_add_136231_comb[16]}}, p1_add_136231_comb};
  assign p1_sum__1807_comb = {{8{p1_add_136232_comb[16]}}, p1_add_136232_comb};
  assign p1_sum__1668_comb = {{8{p1_add_136233_comb[16]}}, p1_add_136233_comb};
  assign p1_sum__1669_comb = {{8{p1_add_136234_comb[16]}}, p1_add_136234_comb};
  assign p1_sum__1670_comb = {{8{p1_add_136235_comb[16]}}, p1_add_136235_comb};
  assign p1_sum__1671_comb = {{8{p1_add_136236_comb[16]}}, p1_add_136236_comb};
  assign p1_sum__1800_comb = {{8{p1_add_136237_comb[16]}}, p1_add_136237_comb};
  assign p1_sum__1801_comb = {{8{p1_add_136238_comb[16]}}, p1_add_136238_comb};
  assign p1_sum__1802_comb = {{8{p1_add_136239_comb[16]}}, p1_add_136239_comb};
  assign p1_sum__1803_comb = {{8{p1_add_136240_comb[16]}}, p1_add_136240_comb};
  assign p1_sum__1644_comb = {{8{p1_add_136241_comb[16]}}, p1_add_136241_comb};
  assign p1_sum__1645_comb = {{8{p1_add_136242_comb[16]}}, p1_add_136242_comb};
  assign p1_sum__1646_comb = {{8{p1_add_136243_comb[16]}}, p1_add_136243_comb};
  assign p1_sum__1647_comb = {{8{p1_add_136244_comb[16]}}, p1_add_136244_comb};
  assign p1_sum__1792_comb = {{8{p1_add_136245_comb[16]}}, p1_add_136245_comb};
  assign p1_sum__1793_comb = {{8{p1_add_136246_comb[16]}}, p1_add_136246_comb};
  assign p1_sum__1794_comb = {{8{p1_add_136247_comb[16]}}, p1_add_136247_comb};
  assign p1_sum__1795_comb = {{8{p1_add_136248_comb[16]}}, p1_add_136248_comb};
  assign p1_sum__1624_comb = {{8{p1_add_136249_comb[16]}}, p1_add_136249_comb};
  assign p1_sum__1625_comb = {{8{p1_add_136250_comb[16]}}, p1_add_136250_comb};
  assign p1_sum__1626_comb = {{8{p1_add_136251_comb[16]}}, p1_add_136251_comb};
  assign p1_sum__1627_comb = {{8{p1_add_136252_comb[16]}}, p1_add_136252_comb};
  assign p1_sum__1780_comb = {{8{p1_add_136253_comb[16]}}, p1_add_136253_comb};
  assign p1_sum__1781_comb = {{8{p1_add_136254_comb[16]}}, p1_add_136254_comb};
  assign p1_sum__1782_comb = {{8{p1_add_136255_comb[16]}}, p1_add_136255_comb};
  assign p1_sum__1783_comb = {{8{p1_add_136256_comb[16]}}, p1_add_136256_comb};
  assign p1_sum__1608_comb = {{8{p1_add_136257_comb[16]}}, p1_add_136257_comb};
  assign p1_sum__1609_comb = {{8{p1_add_136258_comb[16]}}, p1_add_136258_comb};
  assign p1_sum__1610_comb = {{8{p1_add_136259_comb[16]}}, p1_add_136259_comb};
  assign p1_sum__1611_comb = {{8{p1_add_136260_comb[16]}}, p1_add_136260_comb};
  assign p1_sum__1764_comb = {{8{p1_add_136261_comb[16]}}, p1_add_136261_comb};
  assign p1_sum__1765_comb = {{8{p1_add_136262_comb[16]}}, p1_add_136262_comb};
  assign p1_sum__1766_comb = {{8{p1_add_136263_comb[16]}}, p1_add_136263_comb};
  assign p1_sum__1767_comb = {{8{p1_add_136264_comb[16]}}, p1_add_136264_comb};
  assign p1_sum__1596_comb = {{8{p1_add_136265_comb[16]}}, p1_add_136265_comb};
  assign p1_sum__1597_comb = {{8{p1_add_136266_comb[16]}}, p1_add_136266_comb};
  assign p1_sum__1598_comb = {{8{p1_add_136267_comb[16]}}, p1_add_136267_comb};
  assign p1_sum__1599_comb = {{8{p1_add_136268_comb[16]}}, p1_add_136268_comb};
  assign p1_sum__1744_comb = {{8{p1_add_136269_comb[16]}}, p1_add_136269_comb};
  assign p1_sum__1745_comb = {{8{p1_add_136270_comb[16]}}, p1_add_136270_comb};
  assign p1_sum__1746_comb = {{8{p1_add_136271_comb[16]}}, p1_add_136271_comb};
  assign p1_sum__1747_comb = {{8{p1_add_136272_comb[16]}}, p1_add_136272_comb};
  assign p1_sum__1588_comb = {{8{p1_add_136273_comb[16]}}, p1_add_136273_comb};
  assign p1_sum__1589_comb = {{8{p1_add_136274_comb[16]}}, p1_add_136274_comb};
  assign p1_sum__1590_comb = {{8{p1_add_136275_comb[16]}}, p1_add_136275_comb};
  assign p1_sum__1591_comb = {{8{p1_add_136276_comb[16]}}, p1_add_136276_comb};
  assign p1_sum__1720_comb = {{8{p1_add_136277_comb[16]}}, p1_add_136277_comb};
  assign p1_sum__1721_comb = {{8{p1_add_136278_comb[16]}}, p1_add_136278_comb};
  assign p1_sum__1722_comb = {{8{p1_add_136279_comb[16]}}, p1_add_136279_comb};
  assign p1_sum__1723_comb = {{8{p1_add_136280_comb[16]}}, p1_add_136280_comb};
  assign p1_sum__1584_comb = {{8{p1_add_136281_comb[16]}}, p1_add_136281_comb};
  assign p1_sum__1585_comb = {{8{p1_add_136282_comb[16]}}, p1_add_136282_comb};
  assign p1_sum__1586_comb = {{8{p1_add_136283_comb[16]}}, p1_add_136283_comb};
  assign p1_sum__1587_comb = {{8{p1_add_136284_comb[16]}}, p1_add_136284_comb};
  assign p1_sum__1016_comb = p1_sum__1014_comb + p1_sum__1015_comb;
  assign p1_sum__841_comb = p1_sum__839_comb + p1_sum__840_comb;
  assign p1_sum__1796_comb = {{8{p1_add_136289_comb[16]}}, p1_add_136289_comb};
  assign p1_sum__1797_comb = {{8{p1_add_136290_comb[16]}}, p1_add_136290_comb};
  assign p1_sum__1798_comb = {{8{p1_add_136291_comb[16]}}, p1_add_136291_comb};
  assign p1_sum__1799_comb = {{8{p1_add_136292_comb[16]}}, p1_add_136292_comb};
  assign p1_sum__1696_comb = {{8{p1_add_136293_comb[16]}}, p1_add_136293_comb};
  assign p1_sum__1697_comb = {{8{p1_add_136294_comb[16]}}, p1_add_136294_comb};
  assign p1_sum__1698_comb = {{8{p1_add_136295_comb[16]}}, p1_add_136295_comb};
  assign p1_sum__1699_comb = {{8{p1_add_136296_comb[16]}}, p1_add_136296_comb};
  assign p1_sum__1788_comb = {{8{p1_add_136297_comb[16]}}, p1_add_136297_comb};
  assign p1_sum__1789_comb = {{8{p1_add_136298_comb[16]}}, p1_add_136298_comb};
  assign p1_sum__1790_comb = {{8{p1_add_136299_comb[16]}}, p1_add_136299_comb};
  assign p1_sum__1791_comb = {{8{p1_add_136300_comb[16]}}, p1_add_136300_comb};
  assign p1_sum__1672_comb = {{8{p1_add_136301_comb[16]}}, p1_add_136301_comb};
  assign p1_sum__1673_comb = {{8{p1_add_136302_comb[16]}}, p1_add_136302_comb};
  assign p1_sum__1674_comb = {{8{p1_add_136303_comb[16]}}, p1_add_136303_comb};
  assign p1_sum__1675_comb = {{8{p1_add_136304_comb[16]}}, p1_add_136304_comb};
  assign p1_sum__1776_comb = {{8{p1_add_136305_comb[16]}}, p1_add_136305_comb};
  assign p1_sum__1777_comb = {{8{p1_add_136306_comb[16]}}, p1_add_136306_comb};
  assign p1_sum__1778_comb = {{8{p1_add_136307_comb[16]}}, p1_add_136307_comb};
  assign p1_sum__1779_comb = {{8{p1_add_136308_comb[16]}}, p1_add_136308_comb};
  assign p1_sum__1648_comb = {{8{p1_add_136309_comb[16]}}, p1_add_136309_comb};
  assign p1_sum__1649_comb = {{8{p1_add_136310_comb[16]}}, p1_add_136310_comb};
  assign p1_sum__1650_comb = {{8{p1_add_136311_comb[16]}}, p1_add_136311_comb};
  assign p1_sum__1651_comb = {{8{p1_add_136312_comb[16]}}, p1_add_136312_comb};
  assign p1_sum__1760_comb = {{8{p1_add_136313_comb[16]}}, p1_add_136313_comb};
  assign p1_sum__1761_comb = {{8{p1_add_136314_comb[16]}}, p1_add_136314_comb};
  assign p1_sum__1762_comb = {{8{p1_add_136315_comb[16]}}, p1_add_136315_comb};
  assign p1_sum__1763_comb = {{8{p1_add_136316_comb[16]}}, p1_add_136316_comb};
  assign p1_sum__1628_comb = {{8{p1_add_136317_comb[16]}}, p1_add_136317_comb};
  assign p1_sum__1629_comb = {{8{p1_add_136318_comb[16]}}, p1_add_136318_comb};
  assign p1_sum__1630_comb = {{8{p1_add_136319_comb[16]}}, p1_add_136319_comb};
  assign p1_sum__1631_comb = {{8{p1_add_136320_comb[16]}}, p1_add_136320_comb};
  assign p1_sum__1740_comb = {{8{p1_add_136321_comb[16]}}, p1_add_136321_comb};
  assign p1_sum__1741_comb = {{8{p1_add_136322_comb[16]}}, p1_add_136322_comb};
  assign p1_sum__1742_comb = {{8{p1_add_136323_comb[16]}}, p1_add_136323_comb};
  assign p1_sum__1743_comb = {{8{p1_add_136324_comb[16]}}, p1_add_136324_comb};
  assign p1_sum__1612_comb = {{8{p1_add_136325_comb[16]}}, p1_add_136325_comb};
  assign p1_sum__1613_comb = {{8{p1_add_136326_comb[16]}}, p1_add_136326_comb};
  assign p1_sum__1614_comb = {{8{p1_add_136327_comb[16]}}, p1_add_136327_comb};
  assign p1_sum__1615_comb = {{8{p1_add_136328_comb[16]}}, p1_add_136328_comb};
  assign p1_sum__1716_comb = {{8{p1_add_136329_comb[16]}}, p1_add_136329_comb};
  assign p1_sum__1717_comb = {{8{p1_add_136330_comb[16]}}, p1_add_136330_comb};
  assign p1_sum__1718_comb = {{8{p1_add_136331_comb[16]}}, p1_add_136331_comb};
  assign p1_sum__1719_comb = {{8{p1_add_136332_comb[16]}}, p1_add_136332_comb};
  assign p1_sum__1600_comb = {{8{p1_add_136333_comb[16]}}, p1_add_136333_comb};
  assign p1_sum__1601_comb = {{8{p1_add_136334_comb[16]}}, p1_add_136334_comb};
  assign p1_sum__1602_comb = {{8{p1_add_136335_comb[16]}}, p1_add_136335_comb};
  assign p1_sum__1603_comb = {{8{p1_add_136336_comb[16]}}, p1_add_136336_comb};
  assign p1_sum__1692_comb = {{8{p1_add_136337_comb[16]}}, p1_add_136337_comb};
  assign p1_sum__1693_comb = {{8{p1_add_136338_comb[16]}}, p1_add_136338_comb};
  assign p1_sum__1694_comb = {{8{p1_add_136339_comb[16]}}, p1_add_136339_comb};
  assign p1_sum__1695_comb = {{8{p1_add_136340_comb[16]}}, p1_add_136340_comb};
  assign p1_sum__1592_comb = {{8{p1_add_136341_comb[16]}}, p1_add_136341_comb};
  assign p1_sum__1593_comb = {{8{p1_add_136342_comb[16]}}, p1_add_136342_comb};
  assign p1_sum__1594_comb = {{8{p1_add_136343_comb[16]}}, p1_add_136343_comb};
  assign p1_sum__1595_comb = {{8{p1_add_136344_comb[16]}}, p1_add_136344_comb};
  assign p1_umul_136585_comb = umul32b_32b_x_7b(p1_sum__995_comb, 7'h5b);
  assign p1_umul_136586_comb = umul32b_32b_x_7b(p1_sum__967_comb, 7'h5b);
  assign p1_umul_136587_comb = umul32b_32b_x_7b(p1_sum__932_comb, 7'h5b);
  assign p1_umul_136588_comb = umul32b_32b_x_7b(p1_sum__890_comb, 7'h5b);
  assign p1_sum__1348_comb = p1_sum__1784_comb + p1_sum__1785_comb;
  assign p1_sum__1349_comb = p1_sum__1786_comb + p1_sum__1787_comb;
  assign p1_sum__1340_comb = p1_sum__1768_comb + p1_sum__1769_comb;
  assign p1_sum__1341_comb = p1_sum__1770_comb + p1_sum__1771_comb;
  assign p1_sum__1330_comb = p1_sum__1748_comb + p1_sum__1749_comb;
  assign p1_sum__1331_comb = p1_sum__1750_comb + p1_sum__1751_comb;
  assign p1_sum__1318_comb = p1_sum__1724_comb + p1_sum__1725_comb;
  assign p1_sum__1319_comb = p1_sum__1726_comb + p1_sum__1727_comb;
  assign p1_sum__1342_comb = p1_sum__1772_comb + p1_sum__1773_comb;
  assign p1_sum__1343_comb = p1_sum__1774_comb + p1_sum__1775_comb;
  assign p1_sum__1332_comb = p1_sum__1752_comb + p1_sum__1753_comb;
  assign p1_sum__1333_comb = p1_sum__1754_comb + p1_sum__1755_comb;
  assign p1_sum__1320_comb = p1_sum__1728_comb + p1_sum__1729_comb;
  assign p1_sum__1321_comb = p1_sum__1730_comb + p1_sum__1731_comb;
  assign p1_sum__1306_comb = p1_sum__1700_comb + p1_sum__1701_comb;
  assign p1_sum__1307_comb = p1_sum__1702_comb + p1_sum__1703_comb;
  assign p1_sum__1334_comb = p1_sum__1756_comb + p1_sum__1757_comb;
  assign p1_sum__1335_comb = p1_sum__1758_comb + p1_sum__1759_comb;
  assign p1_sum__1322_comb = p1_sum__1732_comb + p1_sum__1733_comb;
  assign p1_sum__1323_comb = p1_sum__1734_comb + p1_sum__1735_comb;
  assign p1_sum__1308_comb = p1_sum__1704_comb + p1_sum__1705_comb;
  assign p1_sum__1309_comb = p1_sum__1706_comb + p1_sum__1707_comb;
  assign p1_sum__1294_comb = p1_sum__1676_comb + p1_sum__1677_comb;
  assign p1_sum__1295_comb = p1_sum__1678_comb + p1_sum__1679_comb;
  assign p1_sum__1324_comb = p1_sum__1736_comb + p1_sum__1737_comb;
  assign p1_sum__1325_comb = p1_sum__1738_comb + p1_sum__1739_comb;
  assign p1_sum__1310_comb = p1_sum__1708_comb + p1_sum__1709_comb;
  assign p1_sum__1311_comb = p1_sum__1710_comb + p1_sum__1711_comb;
  assign p1_sum__1296_comb = p1_sum__1680_comb + p1_sum__1681_comb;
  assign p1_sum__1297_comb = p1_sum__1682_comb + p1_sum__1683_comb;
  assign p1_sum__1282_comb = p1_sum__1652_comb + p1_sum__1653_comb;
  assign p1_sum__1283_comb = p1_sum__1654_comb + p1_sum__1655_comb;
  assign p1_sum__1312_comb = p1_sum__1712_comb + p1_sum__1713_comb;
  assign p1_sum__1313_comb = p1_sum__1714_comb + p1_sum__1715_comb;
  assign p1_sum__1298_comb = p1_sum__1684_comb + p1_sum__1685_comb;
  assign p1_sum__1299_comb = p1_sum__1686_comb + p1_sum__1687_comb;
  assign p1_sum__1284_comb = p1_sum__1656_comb + p1_sum__1657_comb;
  assign p1_sum__1285_comb = p1_sum__1658_comb + p1_sum__1659_comb;
  assign p1_sum__1272_comb = p1_sum__1632_comb + p1_sum__1633_comb;
  assign p1_sum__1273_comb = p1_sum__1634_comb + p1_sum__1635_comb;
  assign p1_sum__1300_comb = p1_sum__1688_comb + p1_sum__1689_comb;
  assign p1_sum__1301_comb = p1_sum__1690_comb + p1_sum__1691_comb;
  assign p1_sum__1286_comb = p1_sum__1660_comb + p1_sum__1661_comb;
  assign p1_sum__1287_comb = p1_sum__1662_comb + p1_sum__1663_comb;
  assign p1_sum__1274_comb = p1_sum__1636_comb + p1_sum__1637_comb;
  assign p1_sum__1275_comb = p1_sum__1638_comb + p1_sum__1639_comb;
  assign p1_sum__1264_comb = p1_sum__1616_comb + p1_sum__1617_comb;
  assign p1_sum__1265_comb = p1_sum__1618_comb + p1_sum__1619_comb;
  assign p1_sum__1288_comb = p1_sum__1664_comb + p1_sum__1665_comb;
  assign p1_sum__1289_comb = p1_sum__1666_comb + p1_sum__1667_comb;
  assign p1_sum__1276_comb = p1_sum__1640_comb + p1_sum__1641_comb;
  assign p1_sum__1277_comb = p1_sum__1642_comb + p1_sum__1643_comb;
  assign p1_sum__1266_comb = p1_sum__1620_comb + p1_sum__1621_comb;
  assign p1_sum__1267_comb = p1_sum__1622_comb + p1_sum__1623_comb;
  assign p1_sum__1258_comb = p1_sum__1604_comb + p1_sum__1605_comb;
  assign p1_sum__1259_comb = p1_sum__1606_comb + p1_sum__1607_comb;
  assign p1_umul_136645_comb = umul32b_32b_x_7b(p1_sum__1023_comb, 7'h5b);
  assign p1_umul_136646_comb = umul32b_32b_x_7b(p1_sum__785_comb, 7'h5b);
  assign p1_sum__1358_comb = p1_sum__1804_comb + p1_sum__1805_comb;
  assign p1_sum__1359_comb = p1_sum__1806_comb + p1_sum__1807_comb;
  assign p1_sum__1290_comb = p1_sum__1668_comb + p1_sum__1669_comb;
  assign p1_sum__1291_comb = p1_sum__1670_comb + p1_sum__1671_comb;
  assign p1_sum__1356_comb = p1_sum__1800_comb + p1_sum__1801_comb;
  assign p1_sum__1357_comb = p1_sum__1802_comb + p1_sum__1803_comb;
  assign p1_sum__1278_comb = p1_sum__1644_comb + p1_sum__1645_comb;
  assign p1_sum__1279_comb = p1_sum__1646_comb + p1_sum__1647_comb;
  assign p1_sum__1352_comb = p1_sum__1792_comb + p1_sum__1793_comb;
  assign p1_sum__1353_comb = p1_sum__1794_comb + p1_sum__1795_comb;
  assign p1_sum__1268_comb = p1_sum__1624_comb + p1_sum__1625_comb;
  assign p1_sum__1269_comb = p1_sum__1626_comb + p1_sum__1627_comb;
  assign p1_sum__1346_comb = p1_sum__1780_comb + p1_sum__1781_comb;
  assign p1_sum__1347_comb = p1_sum__1782_comb + p1_sum__1783_comb;
  assign p1_sum__1260_comb = p1_sum__1608_comb + p1_sum__1609_comb;
  assign p1_sum__1261_comb = p1_sum__1610_comb + p1_sum__1611_comb;
  assign p1_sum__1338_comb = p1_sum__1764_comb + p1_sum__1765_comb;
  assign p1_sum__1339_comb = p1_sum__1766_comb + p1_sum__1767_comb;
  assign p1_sum__1254_comb = p1_sum__1596_comb + p1_sum__1597_comb;
  assign p1_sum__1255_comb = p1_sum__1598_comb + p1_sum__1599_comb;
  assign p1_sum__1328_comb = p1_sum__1744_comb + p1_sum__1745_comb;
  assign p1_sum__1329_comb = p1_sum__1746_comb + p1_sum__1747_comb;
  assign p1_sum__1250_comb = p1_sum__1588_comb + p1_sum__1589_comb;
  assign p1_sum__1251_comb = p1_sum__1590_comb + p1_sum__1591_comb;
  assign p1_sum__1316_comb = p1_sum__1720_comb + p1_sum__1721_comb;
  assign p1_sum__1317_comb = p1_sum__1722_comb + p1_sum__1723_comb;
  assign p1_sum__1248_comb = p1_sum__1584_comb + p1_sum__1585_comb;
  assign p1_sum__1249_comb = p1_sum__1586_comb + p1_sum__1587_comb;
  assign p1_umul_136675_comb = umul32b_32b_x_7b(p1_sum__1016_comb, 7'h5b);
  assign p1_umul_136676_comb = umul32b_32b_x_7b(p1_sum__841_comb, 7'h5b);
  assign p1_sum__1354_comb = p1_sum__1796_comb + p1_sum__1797_comb;
  assign p1_sum__1355_comb = p1_sum__1798_comb + p1_sum__1799_comb;
  assign p1_sum__1304_comb = p1_sum__1696_comb + p1_sum__1697_comb;
  assign p1_sum__1305_comb = p1_sum__1698_comb + p1_sum__1699_comb;
  assign p1_sum__1350_comb = p1_sum__1788_comb + p1_sum__1789_comb;
  assign p1_sum__1351_comb = p1_sum__1790_comb + p1_sum__1791_comb;
  assign p1_sum__1292_comb = p1_sum__1672_comb + p1_sum__1673_comb;
  assign p1_sum__1293_comb = p1_sum__1674_comb + p1_sum__1675_comb;
  assign p1_sum__1344_comb = p1_sum__1776_comb + p1_sum__1777_comb;
  assign p1_sum__1345_comb = p1_sum__1778_comb + p1_sum__1779_comb;
  assign p1_sum__1280_comb = p1_sum__1648_comb + p1_sum__1649_comb;
  assign p1_sum__1281_comb = p1_sum__1650_comb + p1_sum__1651_comb;
  assign p1_sum__1336_comb = p1_sum__1760_comb + p1_sum__1761_comb;
  assign p1_sum__1337_comb = p1_sum__1762_comb + p1_sum__1763_comb;
  assign p1_sum__1270_comb = p1_sum__1628_comb + p1_sum__1629_comb;
  assign p1_sum__1271_comb = p1_sum__1630_comb + p1_sum__1631_comb;
  assign p1_sum__1326_comb = p1_sum__1740_comb + p1_sum__1741_comb;
  assign p1_sum__1327_comb = p1_sum__1742_comb + p1_sum__1743_comb;
  assign p1_sum__1262_comb = p1_sum__1612_comb + p1_sum__1613_comb;
  assign p1_sum__1263_comb = p1_sum__1614_comb + p1_sum__1615_comb;
  assign p1_sum__1314_comb = p1_sum__1716_comb + p1_sum__1717_comb;
  assign p1_sum__1315_comb = p1_sum__1718_comb + p1_sum__1719_comb;
  assign p1_sum__1256_comb = p1_sum__1600_comb + p1_sum__1601_comb;
  assign p1_sum__1257_comb = p1_sum__1602_comb + p1_sum__1603_comb;
  assign p1_sum__1302_comb = p1_sum__1692_comb + p1_sum__1693_comb;
  assign p1_sum__1303_comb = p1_sum__1694_comb + p1_sum__1695_comb;
  assign p1_sum__1252_comb = p1_sum__1592_comb + p1_sum__1593_comb;
  assign p1_sum__1253_comb = p1_sum__1594_comb + p1_sum__1595_comb;
  assign p1_sum__1130_comb = p1_sum__1348_comb + p1_sum__1349_comb;
  assign p1_sum__1126_comb = p1_sum__1340_comb + p1_sum__1341_comb;
  assign p1_sum__1121_comb = p1_sum__1330_comb + p1_sum__1331_comb;
  assign p1_sum__1115_comb = p1_sum__1318_comb + p1_sum__1319_comb;
  assign p1_sum__1127_comb = p1_sum__1342_comb + p1_sum__1343_comb;
  assign p1_sum__1122_comb = p1_sum__1332_comb + p1_sum__1333_comb;
  assign p1_sum__1116_comb = p1_sum__1320_comb + p1_sum__1321_comb;
  assign p1_sum__1109_comb = p1_sum__1306_comb + p1_sum__1307_comb;
  assign p1_sum__1123_comb = p1_sum__1334_comb + p1_sum__1335_comb;
  assign p1_sum__1117_comb = p1_sum__1322_comb + p1_sum__1323_comb;
  assign p1_sum__1110_comb = p1_sum__1308_comb + p1_sum__1309_comb;
  assign p1_sum__1103_comb = p1_sum__1294_comb + p1_sum__1295_comb;
  assign p1_sum__1118_comb = p1_sum__1324_comb + p1_sum__1325_comb;
  assign p1_sum__1111_comb = p1_sum__1310_comb + p1_sum__1311_comb;
  assign p1_sum__1104_comb = p1_sum__1296_comb + p1_sum__1297_comb;
  assign p1_sum__1097_comb = p1_sum__1282_comb + p1_sum__1283_comb;
  assign p1_sum__1112_comb = p1_sum__1312_comb + p1_sum__1313_comb;
  assign p1_sum__1105_comb = p1_sum__1298_comb + p1_sum__1299_comb;
  assign p1_sum__1098_comb = p1_sum__1284_comb + p1_sum__1285_comb;
  assign p1_sum__1092_comb = p1_sum__1272_comb + p1_sum__1273_comb;
  assign p1_sum__1106_comb = p1_sum__1300_comb + p1_sum__1301_comb;
  assign p1_sum__1099_comb = p1_sum__1286_comb + p1_sum__1287_comb;
  assign p1_sum__1093_comb = p1_sum__1274_comb + p1_sum__1275_comb;
  assign p1_sum__1088_comb = p1_sum__1264_comb + p1_sum__1265_comb;
  assign p1_sum__1100_comb = p1_sum__1288_comb + p1_sum__1289_comb;
  assign p1_sum__1094_comb = p1_sum__1276_comb + p1_sum__1277_comb;
  assign p1_sum__1089_comb = p1_sum__1266_comb + p1_sum__1267_comb;
  assign p1_sum__1085_comb = p1_sum__1258_comb + p1_sum__1259_comb;
  assign p1_sum__1135_comb = p1_sum__1358_comb + p1_sum__1359_comb;
  assign p1_sum__1101_comb = p1_sum__1290_comb + p1_sum__1291_comb;
  assign p1_sum__1134_comb = p1_sum__1356_comb + p1_sum__1357_comb;
  assign p1_sum__1095_comb = p1_sum__1278_comb + p1_sum__1279_comb;
  assign p1_sum__1132_comb = p1_sum__1352_comb + p1_sum__1353_comb;
  assign p1_sum__1090_comb = p1_sum__1268_comb + p1_sum__1269_comb;
  assign p1_sum__1129_comb = p1_sum__1346_comb + p1_sum__1347_comb;
  assign p1_sum__1086_comb = p1_sum__1260_comb + p1_sum__1261_comb;
  assign p1_sum__1125_comb = p1_sum__1338_comb + p1_sum__1339_comb;
  assign p1_sum__1083_comb = p1_sum__1254_comb + p1_sum__1255_comb;
  assign p1_sum__1120_comb = p1_sum__1328_comb + p1_sum__1329_comb;
  assign p1_sum__1081_comb = p1_sum__1250_comb + p1_sum__1251_comb;
  assign p1_sum__1114_comb = p1_sum__1316_comb + p1_sum__1317_comb;
  assign p1_sum__1080_comb = p1_sum__1248_comb + p1_sum__1249_comb;
  assign p1_sum__1133_comb = p1_sum__1354_comb + p1_sum__1355_comb;
  assign p1_sum__1108_comb = p1_sum__1304_comb + p1_sum__1305_comb;
  assign p1_sum__1131_comb = p1_sum__1350_comb + p1_sum__1351_comb;
  assign p1_sum__1102_comb = p1_sum__1292_comb + p1_sum__1293_comb;
  assign p1_sum__1128_comb = p1_sum__1344_comb + p1_sum__1345_comb;
  assign p1_sum__1096_comb = p1_sum__1280_comb + p1_sum__1281_comb;
  assign p1_sum__1124_comb = p1_sum__1336_comb + p1_sum__1337_comb;
  assign p1_sum__1091_comb = p1_sum__1270_comb + p1_sum__1271_comb;
  assign p1_sum__1119_comb = p1_sum__1326_comb + p1_sum__1327_comb;
  assign p1_sum__1087_comb = p1_sum__1262_comb + p1_sum__1263_comb;
  assign p1_sum__1113_comb = p1_sum__1314_comb + p1_sum__1315_comb;
  assign p1_sum__1084_comb = p1_sum__1256_comb + p1_sum__1257_comb;
  assign p1_sum__1107_comb = p1_sum__1302_comb + p1_sum__1303_comb;
  assign p1_sum__1082_comb = p1_sum__1252_comb + p1_sum__1253_comb;
  assign p1_add_136833_comb = p1_umul_136585_comb[31:7] + 25'h000_0001;
  assign p1_add_136834_comb = p1_umul_136586_comb[31:7] + 25'h000_0001;
  assign p1_add_136835_comb = p1_umul_136587_comb[31:7] + 25'h000_0001;
  assign p1_add_136836_comb = p1_umul_136588_comb[31:7] + 25'h000_0001;
  assign p1_add_136837_comb = p1_sum__1130_comb + 25'h000_0001;
  assign p1_add_136838_comb = p1_sum__1126_comb + 25'h000_0001;
  assign p1_add_136839_comb = p1_sum__1121_comb + 25'h000_0001;
  assign p1_add_136840_comb = p1_sum__1115_comb + 25'h000_0001;
  assign p1_add_136841_comb = p1_sum__1127_comb + 25'h000_0001;
  assign p1_add_136842_comb = p1_sum__1122_comb + 25'h000_0001;
  assign p1_add_136843_comb = p1_sum__1116_comb + 25'h000_0001;
  assign p1_add_136844_comb = p1_sum__1109_comb + 25'h000_0001;
  assign p1_add_136845_comb = p1_sum__1123_comb + 25'h000_0001;
  assign p1_add_136846_comb = p1_sum__1117_comb + 25'h000_0001;
  assign p1_add_136847_comb = p1_sum__1110_comb + 25'h000_0001;
  assign p1_add_136848_comb = p1_sum__1103_comb + 25'h000_0001;
  assign p1_add_136849_comb = p1_sum__1118_comb + 25'h000_0001;
  assign p1_add_136850_comb = p1_sum__1111_comb + 25'h000_0001;
  assign p1_add_136851_comb = p1_sum__1104_comb + 25'h000_0001;
  assign p1_add_136852_comb = p1_sum__1097_comb + 25'h000_0001;
  assign p1_add_136853_comb = p1_sum__1112_comb + 25'h000_0001;
  assign p1_add_136854_comb = p1_sum__1105_comb + 25'h000_0001;
  assign p1_add_136855_comb = p1_sum__1098_comb + 25'h000_0001;
  assign p1_add_136856_comb = p1_sum__1092_comb + 25'h000_0001;
  assign p1_add_136857_comb = p1_sum__1106_comb + 25'h000_0001;
  assign p1_add_136858_comb = p1_sum__1099_comb + 25'h000_0001;
  assign p1_add_136859_comb = p1_sum__1093_comb + 25'h000_0001;
  assign p1_add_136860_comb = p1_sum__1088_comb + 25'h000_0001;
  assign p1_add_136861_comb = p1_sum__1100_comb + 25'h000_0001;
  assign p1_add_136862_comb = p1_sum__1094_comb + 25'h000_0001;
  assign p1_add_136863_comb = p1_sum__1089_comb + 25'h000_0001;
  assign p1_add_136864_comb = p1_sum__1085_comb + 25'h000_0001;
  assign p1_add_136865_comb = p1_umul_136645_comb[31:7] + 25'h000_0001;
  assign p1_add_136866_comb = p1_umul_136646_comb[31:7] + 25'h000_0001;
  assign p1_add_136867_comb = p1_sum__1135_comb + 25'h000_0001;
  assign p1_add_136868_comb = p1_sum__1101_comb + 25'h000_0001;
  assign p1_add_136869_comb = p1_sum__1134_comb + 25'h000_0001;
  assign p1_add_136870_comb = p1_sum__1095_comb + 25'h000_0001;
  assign p1_add_136871_comb = p1_sum__1132_comb + 25'h000_0001;
  assign p1_add_136872_comb = p1_sum__1090_comb + 25'h000_0001;
  assign p1_add_136873_comb = p1_sum__1129_comb + 25'h000_0001;
  assign p1_add_136874_comb = p1_sum__1086_comb + 25'h000_0001;
  assign p1_add_136875_comb = p1_sum__1125_comb + 25'h000_0001;
  assign p1_add_136876_comb = p1_sum__1083_comb + 25'h000_0001;
  assign p1_add_136877_comb = p1_sum__1120_comb + 25'h000_0001;
  assign p1_add_136878_comb = p1_sum__1081_comb + 25'h000_0001;
  assign p1_add_136879_comb = p1_sum__1114_comb + 25'h000_0001;
  assign p1_add_136880_comb = p1_sum__1080_comb + 25'h000_0001;
  assign p1_add_136881_comb = p1_umul_136675_comb[31:7] + 25'h000_0001;
  assign p1_add_136882_comb = p1_umul_136676_comb[31:7] + 25'h000_0001;
  assign p1_add_136883_comb = p1_sum__1133_comb + 25'h000_0001;
  assign p1_add_136884_comb = p1_sum__1108_comb + 25'h000_0001;
  assign p1_add_136885_comb = p1_sum__1131_comb + 25'h000_0001;
  assign p1_add_136886_comb = p1_sum__1102_comb + 25'h000_0001;
  assign p1_add_136887_comb = p1_sum__1128_comb + 25'h000_0001;
  assign p1_add_136888_comb = p1_sum__1096_comb + 25'h000_0001;
  assign p1_add_136889_comb = p1_sum__1124_comb + 25'h000_0001;
  assign p1_add_136890_comb = p1_sum__1091_comb + 25'h000_0001;
  assign p1_add_136891_comb = p1_sum__1119_comb + 25'h000_0001;
  assign p1_add_136892_comb = p1_sum__1087_comb + 25'h000_0001;
  assign p1_add_136893_comb = p1_sum__1113_comb + 25'h000_0001;
  assign p1_add_136894_comb = p1_sum__1084_comb + 25'h000_0001;
  assign p1_add_136895_comb = p1_sum__1107_comb + 25'h000_0001;
  assign p1_add_136896_comb = p1_sum__1082_comb + 25'h000_0001;
  assign p1_clipped__256_comb = $signed(p1_add_136833_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136833_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136833_comb[16:8]);
  assign p1_clipped__257_comb = $signed(p1_add_136834_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136834_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136834_comb[16:8]);
  assign p1_clipped__258_comb = $signed(p1_add_136835_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136835_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136835_comb[16:8]);
  assign p1_clipped__259_comb = $signed(p1_add_136836_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136836_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136836_comb[16:8]);
  assign p1_clipped__260_comb = $signed(p1_add_136837_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136837_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136837_comb[16:8]);
  assign p1_clipped__261_comb = $signed(p1_add_136838_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136838_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136838_comb[16:8]);
  assign p1_clipped__262_comb = $signed(p1_add_136839_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136839_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136839_comb[16:8]);
  assign p1_clipped__263_comb = $signed(p1_add_136840_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136840_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136840_comb[16:8]);
  assign p1_clipped__264_comb = $signed(p1_add_136841_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136841_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136841_comb[16:8]);
  assign p1_clipped__265_comb = $signed(p1_add_136842_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136842_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136842_comb[16:8]);
  assign p1_clipped__266_comb = $signed(p1_add_136843_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136843_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136843_comb[16:8]);
  assign p1_clipped__267_comb = $signed(p1_add_136844_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136844_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136844_comb[16:8]);
  assign p1_clipped__268_comb = $signed(p1_add_136845_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136845_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136845_comb[16:8]);
  assign p1_clipped__269_comb = $signed(p1_add_136846_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136846_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136846_comb[16:8]);
  assign p1_clipped__270_comb = $signed(p1_add_136847_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136847_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136847_comb[16:8]);
  assign p1_clipped__271_comb = $signed(p1_add_136848_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136848_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136848_comb[16:8]);
  assign p1_clipped__272_comb = $signed(p1_add_136849_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136849_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136849_comb[16:8]);
  assign p1_clipped__273_comb = $signed(p1_add_136850_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136850_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136850_comb[16:8]);
  assign p1_clipped__274_comb = $signed(p1_add_136851_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136851_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136851_comb[16:8]);
  assign p1_clipped__275_comb = $signed(p1_add_136852_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136852_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136852_comb[16:8]);
  assign p1_clipped__276_comb = $signed(p1_add_136853_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136853_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136853_comb[16:8]);
  assign p1_clipped__277_comb = $signed(p1_add_136854_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136854_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136854_comb[16:8]);
  assign p1_clipped__278_comb = $signed(p1_add_136855_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136855_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136855_comb[16:8]);
  assign p1_clipped__279_comb = $signed(p1_add_136856_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136856_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136856_comb[16:8]);
  assign p1_clipped__280_comb = $signed(p1_add_136857_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136857_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136857_comb[16:8]);
  assign p1_clipped__281_comb = $signed(p1_add_136858_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136858_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136858_comb[16:8]);
  assign p1_clipped__282_comb = $signed(p1_add_136859_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136859_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136859_comb[16:8]);
  assign p1_clipped__283_comb = $signed(p1_add_136860_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136860_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136860_comb[16:8]);
  assign p1_clipped__284_comb = $signed(p1_add_136861_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136861_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136861_comb[16:8]);
  assign p1_clipped__285_comb = $signed(p1_add_136862_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136862_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136862_comb[16:8]);
  assign p1_clipped__286_comb = $signed(p1_add_136863_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136863_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136863_comb[16:8]);
  assign p1_clipped__287_comb = $signed(p1_add_136864_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136864_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136864_comb[16:8]);
  assign p1_clipped__288_comb = $signed(p1_add_136865_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136865_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136865_comb[16:8]);
  assign p1_clipped__291_comb = $signed(p1_add_136866_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136866_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136866_comb[16:8]);
  assign p1_clipped__292_comb = $signed(p1_add_136867_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136867_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136867_comb[16:8]);
  assign p1_clipped__295_comb = $signed(p1_add_136868_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136868_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136868_comb[16:8]);
  assign p1_clipped__296_comb = $signed(p1_add_136869_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136869_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136869_comb[16:8]);
  assign p1_clipped__299_comb = $signed(p1_add_136870_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136870_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136870_comb[16:8]);
  assign p1_clipped__300_comb = $signed(p1_add_136871_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136871_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136871_comb[16:8]);
  assign p1_clipped__303_comb = $signed(p1_add_136872_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136872_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136872_comb[16:8]);
  assign p1_clipped__304_comb = $signed(p1_add_136873_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136873_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136873_comb[16:8]);
  assign p1_clipped__307_comb = $signed(p1_add_136874_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136874_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136874_comb[16:8]);
  assign p1_clipped__308_comb = $signed(p1_add_136875_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136875_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136875_comb[16:8]);
  assign p1_clipped__311_comb = $signed(p1_add_136876_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136876_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136876_comb[16:8]);
  assign p1_clipped__312_comb = $signed(p1_add_136877_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136877_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136877_comb[16:8]);
  assign p1_clipped__315_comb = $signed(p1_add_136878_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136878_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136878_comb[16:8]);
  assign p1_clipped__316_comb = $signed(p1_add_136879_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136879_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136879_comb[16:8]);
  assign p1_clipped__319_comb = $signed(p1_add_136880_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136880_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136880_comb[16:8]);
  assign p1_clipped__289_comb = $signed(p1_add_136881_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136881_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136881_comb[16:8]);
  assign p1_clipped__290_comb = $signed(p1_add_136882_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136882_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136882_comb[16:8]);
  assign p1_clipped__293_comb = $signed(p1_add_136883_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136883_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136883_comb[16:8]);
  assign p1_clipped__294_comb = $signed(p1_add_136884_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136884_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136884_comb[16:8]);
  assign p1_clipped__297_comb = $signed(p1_add_136885_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136885_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136885_comb[16:8]);
  assign p1_clipped__298_comb = $signed(p1_add_136886_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136886_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136886_comb[16:8]);
  assign p1_clipped__301_comb = $signed(p1_add_136887_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136887_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136887_comb[16:8]);
  assign p1_clipped__302_comb = $signed(p1_add_136888_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136888_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136888_comb[16:8]);
  assign p1_clipped__305_comb = $signed(p1_add_136889_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136889_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136889_comb[16:8]);
  assign p1_clipped__306_comb = $signed(p1_add_136890_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136890_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136890_comb[16:8]);
  assign p1_clipped__309_comb = $signed(p1_add_136891_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136891_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136891_comb[16:8]);
  assign p1_clipped__310_comb = $signed(p1_add_136892_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136892_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136892_comb[16:8]);
  assign p1_clipped__313_comb = $signed(p1_add_136893_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136893_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136893_comb[16:8]);
  assign p1_clipped__314_comb = $signed(p1_add_136894_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136894_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136894_comb[16:8]);
  assign p1_clipped__317_comb = $signed(p1_add_136895_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136895_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136895_comb[16:8]);
  assign p1_clipped__318_comb = $signed(p1_add_136896_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_136896_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_136896_comb[16:8]);
  assign p1_add_137665_comb = {{1{p1_clipped__256_comb[8]}}, p1_clipped__256_comb} + 10'h001;
  assign p1_add_137666_comb = {{1{p1_clipped__257_comb[8]}}, p1_clipped__257_comb} + 10'h001;
  assign p1_add_137667_comb = {{1{p1_clipped__258_comb[8]}}, p1_clipped__258_comb} + 10'h001;
  assign p1_add_137668_comb = {{1{p1_clipped__259_comb[8]}}, p1_clipped__259_comb} + 10'h001;
  assign p1_add_137669_comb = {{1{p1_clipped__260_comb[8]}}, p1_clipped__260_comb} + 10'h001;
  assign p1_add_137670_comb = {{1{p1_clipped__261_comb[8]}}, p1_clipped__261_comb} + 10'h001;
  assign p1_add_137671_comb = {{1{p1_clipped__262_comb[8]}}, p1_clipped__262_comb} + 10'h001;
  assign p1_add_137672_comb = {{1{p1_clipped__263_comb[8]}}, p1_clipped__263_comb} + 10'h001;
  assign p1_add_137673_comb = {{1{p1_clipped__264_comb[8]}}, p1_clipped__264_comb} + 10'h001;
  assign p1_add_137674_comb = {{1{p1_clipped__265_comb[8]}}, p1_clipped__265_comb} + 10'h001;
  assign p1_add_137675_comb = {{1{p1_clipped__266_comb[8]}}, p1_clipped__266_comb} + 10'h001;
  assign p1_add_137676_comb = {{1{p1_clipped__267_comb[8]}}, p1_clipped__267_comb} + 10'h001;
  assign p1_add_137677_comb = {{1{p1_clipped__268_comb[8]}}, p1_clipped__268_comb} + 10'h001;
  assign p1_add_137678_comb = {{1{p1_clipped__269_comb[8]}}, p1_clipped__269_comb} + 10'h001;
  assign p1_add_137679_comb = {{1{p1_clipped__270_comb[8]}}, p1_clipped__270_comb} + 10'h001;
  assign p1_add_137680_comb = {{1{p1_clipped__271_comb[8]}}, p1_clipped__271_comb} + 10'h001;
  assign p1_add_137681_comb = {{1{p1_clipped__272_comb[8]}}, p1_clipped__272_comb} + 10'h001;
  assign p1_add_137682_comb = {{1{p1_clipped__273_comb[8]}}, p1_clipped__273_comb} + 10'h001;
  assign p1_add_137683_comb = {{1{p1_clipped__274_comb[8]}}, p1_clipped__274_comb} + 10'h001;
  assign p1_add_137684_comb = {{1{p1_clipped__275_comb[8]}}, p1_clipped__275_comb} + 10'h001;
  assign p1_add_137685_comb = {{1{p1_clipped__276_comb[8]}}, p1_clipped__276_comb} + 10'h001;
  assign p1_add_137686_comb = {{1{p1_clipped__277_comb[8]}}, p1_clipped__277_comb} + 10'h001;
  assign p1_add_137687_comb = {{1{p1_clipped__278_comb[8]}}, p1_clipped__278_comb} + 10'h001;
  assign p1_add_137688_comb = {{1{p1_clipped__279_comb[8]}}, p1_clipped__279_comb} + 10'h001;
  assign p1_add_137689_comb = {{1{p1_clipped__280_comb[8]}}, p1_clipped__280_comb} + 10'h001;
  assign p1_add_137690_comb = {{1{p1_clipped__281_comb[8]}}, p1_clipped__281_comb} + 10'h001;
  assign p1_add_137691_comb = {{1{p1_clipped__282_comb[8]}}, p1_clipped__282_comb} + 10'h001;
  assign p1_add_137692_comb = {{1{p1_clipped__283_comb[8]}}, p1_clipped__283_comb} + 10'h001;
  assign p1_add_137693_comb = {{1{p1_clipped__284_comb[8]}}, p1_clipped__284_comb} + 10'h001;
  assign p1_add_137694_comb = {{1{p1_clipped__285_comb[8]}}, p1_clipped__285_comb} + 10'h001;
  assign p1_add_137695_comb = {{1{p1_clipped__286_comb[8]}}, p1_clipped__286_comb} + 10'h001;
  assign p1_add_137696_comb = {{1{p1_clipped__287_comb[8]}}, p1_clipped__287_comb} + 10'h001;
  assign p1_add_137697_comb = {{1{p1_clipped__288_comb[8]}}, p1_clipped__288_comb} + 10'h001;
  assign p1_add_137698_comb = {{1{p1_clipped__291_comb[8]}}, p1_clipped__291_comb} + 10'h001;
  assign p1_add_137699_comb = {{1{p1_clipped__292_comb[8]}}, p1_clipped__292_comb} + 10'h001;
  assign p1_add_137700_comb = {{1{p1_clipped__295_comb[8]}}, p1_clipped__295_comb} + 10'h001;
  assign p1_add_137701_comb = {{1{p1_clipped__296_comb[8]}}, p1_clipped__296_comb} + 10'h001;
  assign p1_add_137702_comb = {{1{p1_clipped__299_comb[8]}}, p1_clipped__299_comb} + 10'h001;
  assign p1_add_137703_comb = {{1{p1_clipped__300_comb[8]}}, p1_clipped__300_comb} + 10'h001;
  assign p1_add_137704_comb = {{1{p1_clipped__303_comb[8]}}, p1_clipped__303_comb} + 10'h001;
  assign p1_add_137705_comb = {{1{p1_clipped__304_comb[8]}}, p1_clipped__304_comb} + 10'h001;
  assign p1_add_137706_comb = {{1{p1_clipped__307_comb[8]}}, p1_clipped__307_comb} + 10'h001;
  assign p1_add_137707_comb = {{1{p1_clipped__308_comb[8]}}, p1_clipped__308_comb} + 10'h001;
  assign p1_add_137708_comb = {{1{p1_clipped__311_comb[8]}}, p1_clipped__311_comb} + 10'h001;
  assign p1_add_137709_comb = {{1{p1_clipped__312_comb[8]}}, p1_clipped__312_comb} + 10'h001;
  assign p1_add_137710_comb = {{1{p1_clipped__315_comb[8]}}, p1_clipped__315_comb} + 10'h001;
  assign p1_add_137711_comb = {{1{p1_clipped__316_comb[8]}}, p1_clipped__316_comb} + 10'h001;
  assign p1_add_137712_comb = {{1{p1_clipped__319_comb[8]}}, p1_clipped__319_comb} + 10'h001;
  assign p1_add_137713_comb = {{1{p1_clipped__289_comb[8]}}, p1_clipped__289_comb} + 10'h001;
  assign p1_add_137714_comb = {{1{p1_clipped__290_comb[8]}}, p1_clipped__290_comb} + 10'h001;
  assign p1_add_137715_comb = {{1{p1_clipped__293_comb[8]}}, p1_clipped__293_comb} + 10'h001;
  assign p1_add_137716_comb = {{1{p1_clipped__294_comb[8]}}, p1_clipped__294_comb} + 10'h001;
  assign p1_add_137717_comb = {{1{p1_clipped__297_comb[8]}}, p1_clipped__297_comb} + 10'h001;
  assign p1_add_137718_comb = {{1{p1_clipped__298_comb[8]}}, p1_clipped__298_comb} + 10'h001;
  assign p1_add_137719_comb = {{1{p1_clipped__301_comb[8]}}, p1_clipped__301_comb} + 10'h001;
  assign p1_add_137720_comb = {{1{p1_clipped__302_comb[8]}}, p1_clipped__302_comb} + 10'h001;
  assign p1_add_137721_comb = {{1{p1_clipped__305_comb[8]}}, p1_clipped__305_comb} + 10'h001;
  assign p1_add_137722_comb = {{1{p1_clipped__306_comb[8]}}, p1_clipped__306_comb} + 10'h001;
  assign p1_add_137723_comb = {{1{p1_clipped__309_comb[8]}}, p1_clipped__309_comb} + 10'h001;
  assign p1_add_137724_comb = {{1{p1_clipped__310_comb[8]}}, p1_clipped__310_comb} + 10'h001;
  assign p1_add_137725_comb = {{1{p1_clipped__313_comb[8]}}, p1_clipped__313_comb} + 10'h001;
  assign p1_add_137726_comb = {{1{p1_clipped__314_comb[8]}}, p1_clipped__314_comb} + 10'h001;
  assign p1_add_137727_comb = {{1{p1_clipped__317_comb[8]}}, p1_clipped__317_comb} + 10'h001;
  assign p1_add_137728_comb = {{1{p1_clipped__318_comb[8]}}, p1_clipped__318_comb} + 10'h001;
  assign p1_bit_slice_137729_comb = p1_add_137665_comb[9:8];
  assign p1_bit_slice_137730_comb = p1_add_137666_comb[9:8];
  assign p1_bit_slice_137731_comb = p1_add_137667_comb[9:8];
  assign p1_bit_slice_137732_comb = p1_add_137668_comb[9:8];
  assign p1_bit_slice_137733_comb = p1_add_137669_comb[9:8];
  assign p1_bit_slice_137734_comb = p1_add_137670_comb[9:8];
  assign p1_bit_slice_137735_comb = p1_add_137671_comb[9:8];
  assign p1_bit_slice_137736_comb = p1_add_137672_comb[9:8];
  assign p1_bit_slice_137737_comb = p1_add_137673_comb[9:8];
  assign p1_bit_slice_137738_comb = p1_add_137674_comb[9:8];
  assign p1_bit_slice_137739_comb = p1_add_137675_comb[9:8];
  assign p1_bit_slice_137740_comb = p1_add_137676_comb[9:8];
  assign p1_bit_slice_137741_comb = p1_add_137677_comb[9:8];
  assign p1_bit_slice_137742_comb = p1_add_137678_comb[9:8];
  assign p1_bit_slice_137743_comb = p1_add_137679_comb[9:8];
  assign p1_bit_slice_137744_comb = p1_add_137680_comb[9:8];
  assign p1_bit_slice_137745_comb = p1_add_137681_comb[9:8];
  assign p1_bit_slice_137746_comb = p1_add_137682_comb[9:8];
  assign p1_bit_slice_137747_comb = p1_add_137683_comb[9:8];
  assign p1_bit_slice_137748_comb = p1_add_137684_comb[9:8];
  assign p1_bit_slice_137749_comb = p1_add_137685_comb[9:8];
  assign p1_bit_slice_137750_comb = p1_add_137686_comb[9:8];
  assign p1_bit_slice_137751_comb = p1_add_137687_comb[9:8];
  assign p1_bit_slice_137752_comb = p1_add_137688_comb[9:8];
  assign p1_bit_slice_137753_comb = p1_add_137689_comb[9:8];
  assign p1_bit_slice_137754_comb = p1_add_137690_comb[9:8];
  assign p1_bit_slice_137755_comb = p1_add_137691_comb[9:8];
  assign p1_bit_slice_137756_comb = p1_add_137692_comb[9:8];
  assign p1_bit_slice_137757_comb = p1_add_137693_comb[9:8];
  assign p1_bit_slice_137758_comb = p1_add_137694_comb[9:8];
  assign p1_bit_slice_137759_comb = p1_add_137695_comb[9:8];
  assign p1_bit_slice_137760_comb = p1_add_137696_comb[9:8];
  assign p1_bit_slice_137761_comb = p1_add_137697_comb[9:8];
  assign p1_bit_slice_137762_comb = p1_add_137698_comb[9:8];
  assign p1_bit_slice_137763_comb = p1_add_137699_comb[9:8];
  assign p1_bit_slice_137764_comb = p1_add_137700_comb[9:8];
  assign p1_bit_slice_137765_comb = p1_add_137701_comb[9:8];
  assign p1_bit_slice_137766_comb = p1_add_137702_comb[9:8];
  assign p1_bit_slice_137767_comb = p1_add_137703_comb[9:8];
  assign p1_bit_slice_137768_comb = p1_add_137704_comb[9:8];
  assign p1_bit_slice_137769_comb = p1_add_137705_comb[9:8];
  assign p1_bit_slice_137770_comb = p1_add_137706_comb[9:8];
  assign p1_bit_slice_137771_comb = p1_add_137707_comb[9:8];
  assign p1_bit_slice_137772_comb = p1_add_137708_comb[9:8];
  assign p1_bit_slice_137773_comb = p1_add_137709_comb[9:8];
  assign p1_bit_slice_137774_comb = p1_add_137710_comb[9:8];
  assign p1_bit_slice_137775_comb = p1_add_137711_comb[9:8];
  assign p1_bit_slice_137776_comb = p1_add_137712_comb[9:8];
  assign p1_bit_slice_137777_comb = p1_add_137713_comb[9:8];
  assign p1_bit_slice_137778_comb = p1_add_137714_comb[9:8];
  assign p1_bit_slice_137779_comb = p1_add_137715_comb[9:8];
  assign p1_bit_slice_137780_comb = p1_add_137716_comb[9:8];
  assign p1_bit_slice_137781_comb = p1_add_137717_comb[9:8];
  assign p1_bit_slice_137782_comb = p1_add_137718_comb[9:8];
  assign p1_bit_slice_137783_comb = p1_add_137719_comb[9:8];
  assign p1_bit_slice_137784_comb = p1_add_137720_comb[9:8];
  assign p1_bit_slice_137785_comb = p1_add_137721_comb[9:8];
  assign p1_bit_slice_137786_comb = p1_add_137722_comb[9:8];
  assign p1_bit_slice_137787_comb = p1_add_137723_comb[9:8];
  assign p1_bit_slice_137788_comb = p1_add_137724_comb[9:8];
  assign p1_bit_slice_137789_comb = p1_add_137725_comb[9:8];
  assign p1_bit_slice_137790_comb = p1_add_137726_comb[9:8];
  assign p1_bit_slice_137791_comb = p1_add_137727_comb[9:8];
  assign p1_bit_slice_137792_comb = p1_add_137728_comb[9:8];
  assign p1_add_137921_comb = {{1{p1_bit_slice_137729_comb[1]}}, p1_bit_slice_137729_comb} + 3'h1;
  assign p1_add_137922_comb = {{1{p1_bit_slice_137730_comb[1]}}, p1_bit_slice_137730_comb} + 3'h1;
  assign p1_add_137923_comb = {{1{p1_bit_slice_137731_comb[1]}}, p1_bit_slice_137731_comb} + 3'h1;
  assign p1_add_137924_comb = {{1{p1_bit_slice_137732_comb[1]}}, p1_bit_slice_137732_comb} + 3'h1;
  assign p1_add_137925_comb = {{1{p1_bit_slice_137733_comb[1]}}, p1_bit_slice_137733_comb} + 3'h1;
  assign p1_add_137926_comb = {{1{p1_bit_slice_137734_comb[1]}}, p1_bit_slice_137734_comb} + 3'h1;
  assign p1_add_137927_comb = {{1{p1_bit_slice_137735_comb[1]}}, p1_bit_slice_137735_comb} + 3'h1;
  assign p1_add_137928_comb = {{1{p1_bit_slice_137736_comb[1]}}, p1_bit_slice_137736_comb} + 3'h1;
  assign p1_add_137929_comb = {{1{p1_bit_slice_137737_comb[1]}}, p1_bit_slice_137737_comb} + 3'h1;
  assign p1_add_137930_comb = {{1{p1_bit_slice_137738_comb[1]}}, p1_bit_slice_137738_comb} + 3'h1;
  assign p1_add_137931_comb = {{1{p1_bit_slice_137739_comb[1]}}, p1_bit_slice_137739_comb} + 3'h1;
  assign p1_add_137932_comb = {{1{p1_bit_slice_137740_comb[1]}}, p1_bit_slice_137740_comb} + 3'h1;
  assign p1_add_137933_comb = {{1{p1_bit_slice_137741_comb[1]}}, p1_bit_slice_137741_comb} + 3'h1;
  assign p1_add_137934_comb = {{1{p1_bit_slice_137742_comb[1]}}, p1_bit_slice_137742_comb} + 3'h1;
  assign p1_add_137935_comb = {{1{p1_bit_slice_137743_comb[1]}}, p1_bit_slice_137743_comb} + 3'h1;
  assign p1_add_137936_comb = {{1{p1_bit_slice_137744_comb[1]}}, p1_bit_slice_137744_comb} + 3'h1;
  assign p1_add_137937_comb = {{1{p1_bit_slice_137745_comb[1]}}, p1_bit_slice_137745_comb} + 3'h1;
  assign p1_add_137938_comb = {{1{p1_bit_slice_137746_comb[1]}}, p1_bit_slice_137746_comb} + 3'h1;
  assign p1_add_137939_comb = {{1{p1_bit_slice_137747_comb[1]}}, p1_bit_slice_137747_comb} + 3'h1;
  assign p1_add_137940_comb = {{1{p1_bit_slice_137748_comb[1]}}, p1_bit_slice_137748_comb} + 3'h1;
  assign p1_add_137941_comb = {{1{p1_bit_slice_137749_comb[1]}}, p1_bit_slice_137749_comb} + 3'h1;
  assign p1_add_137942_comb = {{1{p1_bit_slice_137750_comb[1]}}, p1_bit_slice_137750_comb} + 3'h1;
  assign p1_add_137943_comb = {{1{p1_bit_slice_137751_comb[1]}}, p1_bit_slice_137751_comb} + 3'h1;
  assign p1_add_137944_comb = {{1{p1_bit_slice_137752_comb[1]}}, p1_bit_slice_137752_comb} + 3'h1;
  assign p1_add_137945_comb = {{1{p1_bit_slice_137753_comb[1]}}, p1_bit_slice_137753_comb} + 3'h1;
  assign p1_add_137946_comb = {{1{p1_bit_slice_137754_comb[1]}}, p1_bit_slice_137754_comb} + 3'h1;
  assign p1_add_137947_comb = {{1{p1_bit_slice_137755_comb[1]}}, p1_bit_slice_137755_comb} + 3'h1;
  assign p1_add_137948_comb = {{1{p1_bit_slice_137756_comb[1]}}, p1_bit_slice_137756_comb} + 3'h1;
  assign p1_add_137949_comb = {{1{p1_bit_slice_137757_comb[1]}}, p1_bit_slice_137757_comb} + 3'h1;
  assign p1_add_137950_comb = {{1{p1_bit_slice_137758_comb[1]}}, p1_bit_slice_137758_comb} + 3'h1;
  assign p1_add_137951_comb = {{1{p1_bit_slice_137759_comb[1]}}, p1_bit_slice_137759_comb} + 3'h1;
  assign p1_add_137952_comb = {{1{p1_bit_slice_137760_comb[1]}}, p1_bit_slice_137760_comb} + 3'h1;
  assign p1_add_137953_comb = {{1{p1_bit_slice_137761_comb[1]}}, p1_bit_slice_137761_comb} + 3'h1;
  assign p1_add_137954_comb = {{1{p1_bit_slice_137762_comb[1]}}, p1_bit_slice_137762_comb} + 3'h1;
  assign p1_add_137955_comb = {{1{p1_bit_slice_137763_comb[1]}}, p1_bit_slice_137763_comb} + 3'h1;
  assign p1_add_137956_comb = {{1{p1_bit_slice_137764_comb[1]}}, p1_bit_slice_137764_comb} + 3'h1;
  assign p1_add_137957_comb = {{1{p1_bit_slice_137765_comb[1]}}, p1_bit_slice_137765_comb} + 3'h1;
  assign p1_add_137958_comb = {{1{p1_bit_slice_137766_comb[1]}}, p1_bit_slice_137766_comb} + 3'h1;
  assign p1_add_137959_comb = {{1{p1_bit_slice_137767_comb[1]}}, p1_bit_slice_137767_comb} + 3'h1;
  assign p1_add_137960_comb = {{1{p1_bit_slice_137768_comb[1]}}, p1_bit_slice_137768_comb} + 3'h1;
  assign p1_add_137961_comb = {{1{p1_bit_slice_137769_comb[1]}}, p1_bit_slice_137769_comb} + 3'h1;
  assign p1_add_137962_comb = {{1{p1_bit_slice_137770_comb[1]}}, p1_bit_slice_137770_comb} + 3'h1;
  assign p1_add_137963_comb = {{1{p1_bit_slice_137771_comb[1]}}, p1_bit_slice_137771_comb} + 3'h1;
  assign p1_add_137964_comb = {{1{p1_bit_slice_137772_comb[1]}}, p1_bit_slice_137772_comb} + 3'h1;
  assign p1_add_137965_comb = {{1{p1_bit_slice_137773_comb[1]}}, p1_bit_slice_137773_comb} + 3'h1;
  assign p1_add_137966_comb = {{1{p1_bit_slice_137774_comb[1]}}, p1_bit_slice_137774_comb} + 3'h1;
  assign p1_add_137967_comb = {{1{p1_bit_slice_137775_comb[1]}}, p1_bit_slice_137775_comb} + 3'h1;
  assign p1_add_137968_comb = {{1{p1_bit_slice_137776_comb[1]}}, p1_bit_slice_137776_comb} + 3'h1;
  assign p1_add_137969_comb = {{1{p1_bit_slice_137777_comb[1]}}, p1_bit_slice_137777_comb} + 3'h1;
  assign p1_add_137970_comb = {{1{p1_bit_slice_137778_comb[1]}}, p1_bit_slice_137778_comb} + 3'h1;
  assign p1_add_137971_comb = {{1{p1_bit_slice_137779_comb[1]}}, p1_bit_slice_137779_comb} + 3'h1;
  assign p1_add_137972_comb = {{1{p1_bit_slice_137780_comb[1]}}, p1_bit_slice_137780_comb} + 3'h1;
  assign p1_add_137973_comb = {{1{p1_bit_slice_137781_comb[1]}}, p1_bit_slice_137781_comb} + 3'h1;
  assign p1_add_137974_comb = {{1{p1_bit_slice_137782_comb[1]}}, p1_bit_slice_137782_comb} + 3'h1;
  assign p1_add_137975_comb = {{1{p1_bit_slice_137783_comb[1]}}, p1_bit_slice_137783_comb} + 3'h1;
  assign p1_add_137976_comb = {{1{p1_bit_slice_137784_comb[1]}}, p1_bit_slice_137784_comb} + 3'h1;
  assign p1_add_137977_comb = {{1{p1_bit_slice_137785_comb[1]}}, p1_bit_slice_137785_comb} + 3'h1;
  assign p1_add_137978_comb = {{1{p1_bit_slice_137786_comb[1]}}, p1_bit_slice_137786_comb} + 3'h1;
  assign p1_add_137979_comb = {{1{p1_bit_slice_137787_comb[1]}}, p1_bit_slice_137787_comb} + 3'h1;
  assign p1_add_137980_comb = {{1{p1_bit_slice_137788_comb[1]}}, p1_bit_slice_137788_comb} + 3'h1;
  assign p1_add_137981_comb = {{1{p1_bit_slice_137789_comb[1]}}, p1_bit_slice_137789_comb} + 3'h1;
  assign p1_add_137982_comb = {{1{p1_bit_slice_137790_comb[1]}}, p1_bit_slice_137790_comb} + 3'h1;
  assign p1_add_137983_comb = {{1{p1_bit_slice_137791_comb[1]}}, p1_bit_slice_137791_comb} + 3'h1;
  assign p1_add_137984_comb = {{1{p1_bit_slice_137792_comb[1]}}, p1_bit_slice_137792_comb} + 3'h1;
  assign p1_clipped__40_comb = p1_add_137921_comb[1] ? 8'hff : {p1_add_137921_comb[0], p1_add_137665_comb[7:1]};
  assign p1_clipped__56_comb = p1_add_137922_comb[1] ? 8'hff : {p1_add_137922_comb[0], p1_add_137666_comb[7:1]};
  assign p1_clipped__72_comb = p1_add_137923_comb[1] ? 8'hff : {p1_add_137923_comb[0], p1_add_137667_comb[7:1]};
  assign p1_clipped__88_comb = p1_add_137924_comb[1] ? 8'hff : {p1_add_137924_comb[0], p1_add_137668_comb[7:1]};
  assign p1_clipped__41_comb = p1_add_137925_comb[1] ? 8'hff : {p1_add_137925_comb[0], p1_add_137669_comb[7:1]};
  assign p1_clipped__57_comb = p1_add_137926_comb[1] ? 8'hff : {p1_add_137926_comb[0], p1_add_137670_comb[7:1]};
  assign p1_clipped__73_comb = p1_add_137927_comb[1] ? 8'hff : {p1_add_137927_comb[0], p1_add_137671_comb[7:1]};
  assign p1_clipped__89_comb = p1_add_137928_comb[1] ? 8'hff : {p1_add_137928_comb[0], p1_add_137672_comb[7:1]};
  assign p1_clipped__42_comb = p1_add_137929_comb[1] ? 8'hff : {p1_add_137929_comb[0], p1_add_137673_comb[7:1]};
  assign p1_clipped__58_comb = p1_add_137930_comb[1] ? 8'hff : {p1_add_137930_comb[0], p1_add_137674_comb[7:1]};
  assign p1_clipped__74_comb = p1_add_137931_comb[1] ? 8'hff : {p1_add_137931_comb[0], p1_add_137675_comb[7:1]};
  assign p1_clipped__90_comb = p1_add_137932_comb[1] ? 8'hff : {p1_add_137932_comb[0], p1_add_137676_comb[7:1]};
  assign p1_clipped__43_comb = p1_add_137933_comb[1] ? 8'hff : {p1_add_137933_comb[0], p1_add_137677_comb[7:1]};
  assign p1_clipped__59_comb = p1_add_137934_comb[1] ? 8'hff : {p1_add_137934_comb[0], p1_add_137678_comb[7:1]};
  assign p1_clipped__75_comb = p1_add_137935_comb[1] ? 8'hff : {p1_add_137935_comb[0], p1_add_137679_comb[7:1]};
  assign p1_clipped__91_comb = p1_add_137936_comb[1] ? 8'hff : {p1_add_137936_comb[0], p1_add_137680_comb[7:1]};
  assign p1_clipped__44_comb = p1_add_137937_comb[1] ? 8'hff : {p1_add_137937_comb[0], p1_add_137681_comb[7:1]};
  assign p1_clipped__60_comb = p1_add_137938_comb[1] ? 8'hff : {p1_add_137938_comb[0], p1_add_137682_comb[7:1]};
  assign p1_clipped__76_comb = p1_add_137939_comb[1] ? 8'hff : {p1_add_137939_comb[0], p1_add_137683_comb[7:1]};
  assign p1_clipped__92_comb = p1_add_137940_comb[1] ? 8'hff : {p1_add_137940_comb[0], p1_add_137684_comb[7:1]};
  assign p1_clipped__45_comb = p1_add_137941_comb[1] ? 8'hff : {p1_add_137941_comb[0], p1_add_137685_comb[7:1]};
  assign p1_clipped__61_comb = p1_add_137942_comb[1] ? 8'hff : {p1_add_137942_comb[0], p1_add_137686_comb[7:1]};
  assign p1_clipped__77_comb = p1_add_137943_comb[1] ? 8'hff : {p1_add_137943_comb[0], p1_add_137687_comb[7:1]};
  assign p1_clipped__93_comb = p1_add_137944_comb[1] ? 8'hff : {p1_add_137944_comb[0], p1_add_137688_comb[7:1]};
  assign p1_clipped__46_comb = p1_add_137945_comb[1] ? 8'hff : {p1_add_137945_comb[0], p1_add_137689_comb[7:1]};
  assign p1_clipped__62_comb = p1_add_137946_comb[1] ? 8'hff : {p1_add_137946_comb[0], p1_add_137690_comb[7:1]};
  assign p1_clipped__78_comb = p1_add_137947_comb[1] ? 8'hff : {p1_add_137947_comb[0], p1_add_137691_comb[7:1]};
  assign p1_clipped__94_comb = p1_add_137948_comb[1] ? 8'hff : {p1_add_137948_comb[0], p1_add_137692_comb[7:1]};
  assign p1_clipped__47_comb = p1_add_137949_comb[1] ? 8'hff : {p1_add_137949_comb[0], p1_add_137693_comb[7:1]};
  assign p1_clipped__63_comb = p1_add_137950_comb[1] ? 8'hff : {p1_add_137950_comb[0], p1_add_137694_comb[7:1]};
  assign p1_clipped__79_comb = p1_add_137951_comb[1] ? 8'hff : {p1_add_137951_comb[0], p1_add_137695_comb[7:1]};
  assign p1_clipped__95_comb = p1_add_137952_comb[1] ? 8'hff : {p1_add_137952_comb[0], p1_add_137696_comb[7:1]};
  assign p1_clipped__8_comb = p1_add_137953_comb[1] ? 8'hff : {p1_add_137953_comb[0], p1_add_137697_comb[7:1]};
  assign p1_clipped__120_comb = p1_add_137954_comb[1] ? 8'hff : {p1_add_137954_comb[0], p1_add_137698_comb[7:1]};
  assign p1_clipped__9_comb = p1_add_137955_comb[1] ? 8'hff : {p1_add_137955_comb[0], p1_add_137699_comb[7:1]};
  assign p1_clipped__121_comb = p1_add_137956_comb[1] ? 8'hff : {p1_add_137956_comb[0], p1_add_137700_comb[7:1]};
  assign p1_clipped__10_comb = p1_add_137957_comb[1] ? 8'hff : {p1_add_137957_comb[0], p1_add_137701_comb[7:1]};
  assign p1_clipped__122_comb = p1_add_137958_comb[1] ? 8'hff : {p1_add_137958_comb[0], p1_add_137702_comb[7:1]};
  assign p1_clipped__11_comb = p1_add_137959_comb[1] ? 8'hff : {p1_add_137959_comb[0], p1_add_137703_comb[7:1]};
  assign p1_clipped__123_comb = p1_add_137960_comb[1] ? 8'hff : {p1_add_137960_comb[0], p1_add_137704_comb[7:1]};
  assign p1_clipped__12_comb = p1_add_137961_comb[1] ? 8'hff : {p1_add_137961_comb[0], p1_add_137705_comb[7:1]};
  assign p1_clipped__124_comb = p1_add_137962_comb[1] ? 8'hff : {p1_add_137962_comb[0], p1_add_137706_comb[7:1]};
  assign p1_clipped__13_comb = p1_add_137963_comb[1] ? 8'hff : {p1_add_137963_comb[0], p1_add_137707_comb[7:1]};
  assign p1_clipped__125_comb = p1_add_137964_comb[1] ? 8'hff : {p1_add_137964_comb[0], p1_add_137708_comb[7:1]};
  assign p1_clipped__14_comb = p1_add_137965_comb[1] ? 8'hff : {p1_add_137965_comb[0], p1_add_137709_comb[7:1]};
  assign p1_clipped__126_comb = p1_add_137966_comb[1] ? 8'hff : {p1_add_137966_comb[0], p1_add_137710_comb[7:1]};
  assign p1_clipped__15_comb = p1_add_137967_comb[1] ? 8'hff : {p1_add_137967_comb[0], p1_add_137711_comb[7:1]};
  assign p1_clipped__127_comb = p1_add_137968_comb[1] ? 8'hff : {p1_add_137968_comb[0], p1_add_137712_comb[7:1]};
  assign p1_clipped__24_comb = p1_add_137969_comb[1] ? 8'hff : {p1_add_137969_comb[0], p1_add_137713_comb[7:1]};
  assign p1_clipped__104_comb = p1_add_137970_comb[1] ? 8'hff : {p1_add_137970_comb[0], p1_add_137714_comb[7:1]};
  assign p1_clipped__25_comb = p1_add_137971_comb[1] ? 8'hff : {p1_add_137971_comb[0], p1_add_137715_comb[7:1]};
  assign p1_clipped__105_comb = p1_add_137972_comb[1] ? 8'hff : {p1_add_137972_comb[0], p1_add_137716_comb[7:1]};
  assign p1_clipped__26_comb = p1_add_137973_comb[1] ? 8'hff : {p1_add_137973_comb[0], p1_add_137717_comb[7:1]};
  assign p1_clipped__106_comb = p1_add_137974_comb[1] ? 8'hff : {p1_add_137974_comb[0], p1_add_137718_comb[7:1]};
  assign p1_clipped__27_comb = p1_add_137975_comb[1] ? 8'hff : {p1_add_137975_comb[0], p1_add_137719_comb[7:1]};
  assign p1_clipped__107_comb = p1_add_137976_comb[1] ? 8'hff : {p1_add_137976_comb[0], p1_add_137720_comb[7:1]};
  assign p1_clipped__28_comb = p1_add_137977_comb[1] ? 8'hff : {p1_add_137977_comb[0], p1_add_137721_comb[7:1]};
  assign p1_clipped__108_comb = p1_add_137978_comb[1] ? 8'hff : {p1_add_137978_comb[0], p1_add_137722_comb[7:1]};
  assign p1_clipped__29_comb = p1_add_137979_comb[1] ? 8'hff : {p1_add_137979_comb[0], p1_add_137723_comb[7:1]};
  assign p1_clipped__109_comb = p1_add_137980_comb[1] ? 8'hff : {p1_add_137980_comb[0], p1_add_137724_comb[7:1]};
  assign p1_clipped__30_comb = p1_add_137981_comb[1] ? 8'hff : {p1_add_137981_comb[0], p1_add_137725_comb[7:1]};
  assign p1_clipped__110_comb = p1_add_137982_comb[1] ? 8'hff : {p1_add_137982_comb[0], p1_add_137726_comb[7:1]};
  assign p1_clipped__31_comb = p1_add_137983_comb[1] ? 8'hff : {p1_add_137983_comb[0], p1_add_137727_comb[7:1]};
  assign p1_clipped__111_comb = p1_add_137984_comb[1] ? 8'hff : {p1_add_137984_comb[0], p1_add_137728_comb[7:1]};
  assign p1_shifted__66_squeezed_comb = {~p1_clipped__40_comb[7], p1_clipped__40_comb[6:0]};
  assign p1_shifted__67_squeezed_comb = {~p1_clipped__56_comb[7], p1_clipped__56_comb[6:0]};
  assign p1_shifted__68_squeezed_comb = {~p1_clipped__72_comb[7], p1_clipped__72_comb[6:0]};
  assign p1_shifted__69_squeezed_comb = {~p1_clipped__88_comb[7], p1_clipped__88_comb[6:0]};
  assign p1_shifted__74_squeezed_comb = {~p1_clipped__41_comb[7], p1_clipped__41_comb[6:0]};
  assign p1_shifted__75_squeezed_comb = {~p1_clipped__57_comb[7], p1_clipped__57_comb[6:0]};
  assign p1_shifted__76_squeezed_comb = {~p1_clipped__73_comb[7], p1_clipped__73_comb[6:0]};
  assign p1_shifted__77_squeezed_comb = {~p1_clipped__89_comb[7], p1_clipped__89_comb[6:0]};
  assign p1_shifted__82_squeezed_comb = {~p1_clipped__42_comb[7], p1_clipped__42_comb[6:0]};
  assign p1_shifted__83_squeezed_comb = {~p1_clipped__58_comb[7], p1_clipped__58_comb[6:0]};
  assign p1_shifted__84_squeezed_comb = {~p1_clipped__74_comb[7], p1_clipped__74_comb[6:0]};
  assign p1_shifted__85_squeezed_comb = {~p1_clipped__90_comb[7], p1_clipped__90_comb[6:0]};
  assign p1_shifted__90_squeezed_comb = {~p1_clipped__43_comb[7], p1_clipped__43_comb[6:0]};
  assign p1_shifted__91_squeezed_comb = {~p1_clipped__59_comb[7], p1_clipped__59_comb[6:0]};
  assign p1_shifted__92_squeezed_comb = {~p1_clipped__75_comb[7], p1_clipped__75_comb[6:0]};
  assign p1_shifted__93_squeezed_comb = {~p1_clipped__91_comb[7], p1_clipped__91_comb[6:0]};
  assign p1_shifted__98_squeezed_comb = {~p1_clipped__44_comb[7], p1_clipped__44_comb[6:0]};
  assign p1_shifted__99_squeezed_comb = {~p1_clipped__60_comb[7], p1_clipped__60_comb[6:0]};
  assign p1_shifted__100_squeezed_comb = {~p1_clipped__76_comb[7], p1_clipped__76_comb[6:0]};
  assign p1_shifted__101_squeezed_comb = {~p1_clipped__92_comb[7], p1_clipped__92_comb[6:0]};
  assign p1_shifted__106_squeezed_comb = {~p1_clipped__45_comb[7], p1_clipped__45_comb[6:0]};
  assign p1_shifted__107_squeezed_comb = {~p1_clipped__61_comb[7], p1_clipped__61_comb[6:0]};
  assign p1_shifted__108_squeezed_comb = {~p1_clipped__77_comb[7], p1_clipped__77_comb[6:0]};
  assign p1_shifted__109_squeezed_comb = {~p1_clipped__93_comb[7], p1_clipped__93_comb[6:0]};
  assign p1_shifted__114_squeezed_comb = {~p1_clipped__46_comb[7], p1_clipped__46_comb[6:0]};
  assign p1_shifted__115_squeezed_comb = {~p1_clipped__62_comb[7], p1_clipped__62_comb[6:0]};
  assign p1_shifted__116_squeezed_comb = {~p1_clipped__78_comb[7], p1_clipped__78_comb[6:0]};
  assign p1_shifted__117_squeezed_comb = {~p1_clipped__94_comb[7], p1_clipped__94_comb[6:0]};
  assign p1_shifted__122_squeezed_comb = {~p1_clipped__47_comb[7], p1_clipped__47_comb[6:0]};
  assign p1_shifted__123_squeezed_comb = {~p1_clipped__63_comb[7], p1_clipped__63_comb[6:0]};
  assign p1_shifted__124_squeezed_comb = {~p1_clipped__79_comb[7], p1_clipped__79_comb[6:0]};
  assign p1_shifted__125_squeezed_comb = {~p1_clipped__95_comb[7], p1_clipped__95_comb[6:0]};
  assign p1_shifted__64_squeezed_comb = {~p1_clipped__8_comb[7], p1_clipped__8_comb[6:0]};
  assign p1_shifted__71_squeezed_comb = {~p1_clipped__120_comb[7], p1_clipped__120_comb[6:0]};
  assign p1_shifted__72_squeezed_comb = {~p1_clipped__9_comb[7], p1_clipped__9_comb[6:0]};
  assign p1_shifted__79_squeezed_comb = {~p1_clipped__121_comb[7], p1_clipped__121_comb[6:0]};
  assign p1_shifted__80_squeezed_comb = {~p1_clipped__10_comb[7], p1_clipped__10_comb[6:0]};
  assign p1_shifted__87_squeezed_comb = {~p1_clipped__122_comb[7], p1_clipped__122_comb[6:0]};
  assign p1_shifted__88_squeezed_comb = {~p1_clipped__11_comb[7], p1_clipped__11_comb[6:0]};
  assign p1_shifted__95_squeezed_comb = {~p1_clipped__123_comb[7], p1_clipped__123_comb[6:0]};
  assign p1_shifted__96_squeezed_comb = {~p1_clipped__12_comb[7], p1_clipped__12_comb[6:0]};
  assign p1_shifted__103_squeezed_comb = {~p1_clipped__124_comb[7], p1_clipped__124_comb[6:0]};
  assign p1_shifted__104_squeezed_comb = {~p1_clipped__13_comb[7], p1_clipped__13_comb[6:0]};
  assign p1_shifted__111_squeezed_comb = {~p1_clipped__125_comb[7], p1_clipped__125_comb[6:0]};
  assign p1_shifted__112_squeezed_comb = {~p1_clipped__14_comb[7], p1_clipped__14_comb[6:0]};
  assign p1_shifted__119_squeezed_comb = {~p1_clipped__126_comb[7], p1_clipped__126_comb[6:0]};
  assign p1_shifted__120_squeezed_comb = {~p1_clipped__15_comb[7], p1_clipped__15_comb[6:0]};
  assign p1_shifted__127_squeezed_comb = {~p1_clipped__127_comb[7], p1_clipped__127_comb[6:0]};
  assign p1_shifted__65_squeezed_comb = {~p1_clipped__24_comb[7], p1_clipped__24_comb[6:0]};
  assign p1_shifted__70_squeezed_comb = {~p1_clipped__104_comb[7], p1_clipped__104_comb[6:0]};
  assign p1_shifted__73_squeezed_comb = {~p1_clipped__25_comb[7], p1_clipped__25_comb[6:0]};
  assign p1_shifted__78_squeezed_comb = {~p1_clipped__105_comb[7], p1_clipped__105_comb[6:0]};
  assign p1_shifted__81_squeezed_comb = {~p1_clipped__26_comb[7], p1_clipped__26_comb[6:0]};
  assign p1_shifted__86_squeezed_comb = {~p1_clipped__106_comb[7], p1_clipped__106_comb[6:0]};
  assign p1_shifted__89_squeezed_comb = {~p1_clipped__27_comb[7], p1_clipped__27_comb[6:0]};
  assign p1_shifted__94_squeezed_comb = {~p1_clipped__107_comb[7], p1_clipped__107_comb[6:0]};
  assign p1_shifted__97_squeezed_comb = {~p1_clipped__28_comb[7], p1_clipped__28_comb[6:0]};
  assign p1_shifted__102_squeezed_comb = {~p1_clipped__108_comb[7], p1_clipped__108_comb[6:0]};
  assign p1_shifted__105_squeezed_comb = {~p1_clipped__29_comb[7], p1_clipped__29_comb[6:0]};
  assign p1_shifted__110_squeezed_comb = {~p1_clipped__109_comb[7], p1_clipped__109_comb[6:0]};
  assign p1_shifted__113_squeezed_comb = {~p1_clipped__30_comb[7], p1_clipped__30_comb[6:0]};
  assign p1_shifted__118_squeezed_comb = {~p1_clipped__110_comb[7], p1_clipped__110_comb[6:0]};
  assign p1_shifted__121_squeezed_comb = {~p1_clipped__31_comb[7], p1_clipped__31_comb[6:0]};
  assign p1_shifted__126_squeezed_comb = {~p1_clipped__111_comb[7], p1_clipped__111_comb[6:0]};
  assign p1_smul_58226_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__66_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___128_comb = 9'h000;
  assign p1_smul_58228_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__67_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___129_comb = 9'h000;
  assign p1_smul_58230_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__68_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___130_comb = 9'h000;
  assign p1_smul_58232_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__69_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___131_comb = 9'h000;
  assign p1_smul_58242_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__74_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___132_comb = 9'h000;
  assign p1_smul_58244_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__75_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___133_comb = 9'h000;
  assign p1_smul_58246_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__76_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___134_comb = 9'h000;
  assign p1_smul_58248_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__77_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___135_comb = 9'h000;
  assign p1_smul_58258_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__82_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___136_comb = 9'h000;
  assign p1_smul_58260_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__83_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___137_comb = 9'h000;
  assign p1_smul_58262_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__84_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___138_comb = 9'h000;
  assign p1_smul_58264_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__85_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___139_comb = 9'h000;
  assign p1_smul_58274_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__90_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___140_comb = 9'h000;
  assign p1_smul_58276_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__91_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___141_comb = 9'h000;
  assign p1_smul_58278_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__92_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___142_comb = 9'h000;
  assign p1_smul_58280_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__93_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___143_comb = 9'h000;
  assign p1_smul_58290_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__98_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___144_comb = 9'h000;
  assign p1_smul_58292_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__99_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___145_comb = 9'h000;
  assign p1_smul_58294_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__100_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___146_comb = 9'h000;
  assign p1_smul_58296_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__101_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___147_comb = 9'h000;
  assign p1_smul_58306_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__106_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___148_comb = 9'h000;
  assign p1_smul_58308_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__107_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___149_comb = 9'h000;
  assign p1_smul_58310_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__108_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___150_comb = 9'h000;
  assign p1_smul_58312_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__109_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___151_comb = 9'h000;
  assign p1_smul_58322_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__114_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___152_comb = 9'h000;
  assign p1_smul_58324_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__115_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___153_comb = 9'h000;
  assign p1_smul_58326_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__116_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___154_comb = 9'h000;
  assign p1_smul_58328_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__117_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___155_comb = 9'h000;
  assign p1_smul_58338_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__122_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___156_comb = 9'h000;
  assign p1_smul_58340_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__123_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___157_comb = 9'h000;
  assign p1_smul_58342_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__124_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___158_comb = 9'h000;
  assign p1_smul_58344_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__125_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___159_comb = 9'h000;
  assign p1_smul_58350_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__64_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___64_comb = 10'h000;
  assign p1_smul_58356_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__67_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___65_comb = 10'h000;
  assign p1_smul_58358_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__68_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___66_comb = 10'h000;
  assign p1_smul_58364_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__71_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___67_comb = 10'h000;
  assign p1_smul_58366_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__72_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___68_comb = 10'h000;
  assign p1_smul_58372_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__75_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___69_comb = 10'h000;
  assign p1_smul_58374_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__76_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___70_comb = 10'h000;
  assign p1_smul_58380_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__79_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___71_comb = 10'h000;
  assign p1_smul_58382_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__80_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___72_comb = 10'h000;
  assign p1_smul_58388_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__83_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___73_comb = 10'h000;
  assign p1_smul_58390_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__84_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___74_comb = 10'h000;
  assign p1_smul_58396_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__87_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___75_comb = 10'h000;
  assign p1_smul_58398_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__88_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___76_comb = 10'h000;
  assign p1_smul_58404_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__91_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___77_comb = 10'h000;
  assign p1_smul_58406_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__92_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___78_comb = 10'h000;
  assign p1_smul_58412_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__95_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___79_comb = 10'h000;
  assign p1_smul_58414_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__96_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___80_comb = 10'h000;
  assign p1_smul_58420_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__99_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___81_comb = 10'h000;
  assign p1_smul_58422_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__100_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___82_comb = 10'h000;
  assign p1_smul_58428_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__103_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___83_comb = 10'h000;
  assign p1_smul_58430_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__104_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___84_comb = 10'h000;
  assign p1_smul_58436_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__107_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___85_comb = 10'h000;
  assign p1_smul_58438_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__108_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___86_comb = 10'h000;
  assign p1_smul_58444_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__111_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___87_comb = 10'h000;
  assign p1_smul_58446_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__112_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___88_comb = 10'h000;
  assign p1_smul_58452_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__115_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___89_comb = 10'h000;
  assign p1_smul_58454_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__116_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___90_comb = 10'h000;
  assign p1_smul_58460_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__119_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___91_comb = 10'h000;
  assign p1_smul_58462_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__120_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___92_comb = 10'h000;
  assign p1_smul_58468_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__123_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___93_comb = 10'h000;
  assign p1_smul_58470_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__124_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___94_comb = 10'h000;
  assign p1_smul_58476_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__127_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___95_comb = 10'h000;
  assign p1_smul_58480_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__65_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___160_comb = 9'h000;
  assign p1_smul_58484_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__67_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___161_comb = 9'h000;
  assign p1_smul_58486_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__68_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___162_comb = 9'h000;
  assign p1_smul_58490_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__70_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___163_comb = 9'h000;
  assign p1_smul_58496_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__73_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___164_comb = 9'h000;
  assign p1_smul_58500_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__75_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___165_comb = 9'h000;
  assign p1_smul_58502_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__76_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___166_comb = 9'h000;
  assign p1_smul_58506_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__78_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___167_comb = 9'h000;
  assign p1_smul_58512_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__81_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___168_comb = 9'h000;
  assign p1_smul_58516_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__83_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___169_comb = 9'h000;
  assign p1_smul_58518_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__84_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___170_comb = 9'h000;
  assign p1_smul_58522_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__86_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___171_comb = 9'h000;
  assign p1_smul_58528_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__89_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___172_comb = 9'h000;
  assign p1_smul_58532_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__91_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___173_comb = 9'h000;
  assign p1_smul_58534_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__92_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___174_comb = 9'h000;
  assign p1_smul_58538_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__94_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___175_comb = 9'h000;
  assign p1_smul_58544_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__97_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___176_comb = 9'h000;
  assign p1_smul_58548_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__99_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___177_comb = 9'h000;
  assign p1_smul_58550_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__100_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___178_comb = 9'h000;
  assign p1_smul_58554_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__102_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___179_comb = 9'h000;
  assign p1_smul_58560_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__105_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___180_comb = 9'h000;
  assign p1_smul_58564_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__107_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___181_comb = 9'h000;
  assign p1_smul_58566_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__108_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___182_comb = 9'h000;
  assign p1_smul_58570_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__110_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___183_comb = 9'h000;
  assign p1_smul_58576_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__113_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___184_comb = 9'h000;
  assign p1_smul_58580_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__115_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___185_comb = 9'h000;
  assign p1_smul_58582_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__116_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___186_comb = 9'h000;
  assign p1_smul_58586_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__118_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___187_comb = 9'h000;
  assign p1_smul_58592_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__121_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___188_comb = 9'h000;
  assign p1_smul_58596_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__123_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___189_comb = 9'h000;
  assign p1_smul_58598_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__124_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___190_comb = 9'h000;
  assign p1_smul_58602_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__126_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___191_comb = 9'h000;
  assign p1_smul_58734_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__64_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___192_comb = 9'h000;
  assign p1_smul_58738_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__66_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___193_comb = 9'h000;
  assign p1_smul_58744_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__69_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___194_comb = 9'h000;
  assign p1_smul_58748_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__71_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___195_comb = 9'h000;
  assign p1_smul_58750_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__72_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___196_comb = 9'h000;
  assign p1_smul_58754_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__74_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___197_comb = 9'h000;
  assign p1_smul_58760_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__77_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___198_comb = 9'h000;
  assign p1_smul_58764_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__79_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___199_comb = 9'h000;
  assign p1_smul_58766_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__80_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___200_comb = 9'h000;
  assign p1_smul_58770_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__82_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___201_comb = 9'h000;
  assign p1_smul_58776_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__85_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___202_comb = 9'h000;
  assign p1_smul_58780_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__87_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___203_comb = 9'h000;
  assign p1_smul_58782_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__88_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___204_comb = 9'h000;
  assign p1_smul_58786_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__90_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___205_comb = 9'h000;
  assign p1_smul_58792_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__93_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___206_comb = 9'h000;
  assign p1_smul_58796_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__95_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___207_comb = 9'h000;
  assign p1_smul_58798_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__96_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___208_comb = 9'h000;
  assign p1_smul_58802_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__98_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___209_comb = 9'h000;
  assign p1_smul_58808_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__101_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___210_comb = 9'h000;
  assign p1_smul_58812_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__103_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___211_comb = 9'h000;
  assign p1_smul_58814_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__104_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___212_comb = 9'h000;
  assign p1_smul_58818_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__106_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___213_comb = 9'h000;
  assign p1_smul_58824_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__109_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___214_comb = 9'h000;
  assign p1_smul_58828_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__111_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___215_comb = 9'h000;
  assign p1_smul_58830_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__112_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___216_comb = 9'h000;
  assign p1_smul_58834_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__114_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___217_comb = 9'h000;
  assign p1_smul_58840_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__117_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___218_comb = 9'h000;
  assign p1_smul_58844_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__119_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___219_comb = 9'h000;
  assign p1_smul_58846_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__120_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___220_comb = 9'h000;
  assign p1_smul_58850_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__122_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___221_comb = 9'h000;
  assign p1_smul_58856_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__125_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___222_comb = 9'h000;
  assign p1_smul_58860_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__127_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___223_comb = 9'h000;
  assign p1_smul_58864_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__65_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___96_comb = 10'h000;
  assign p1_smul_58868_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__67_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___97_comb = 10'h000;
  assign p1_smul_58870_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__68_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___98_comb = 10'h000;
  assign p1_smul_58874_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__70_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___99_comb = 10'h000;
  assign p1_smul_58880_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__73_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___100_comb = 10'h000;
  assign p1_smul_58884_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__75_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___101_comb = 10'h000;
  assign p1_smul_58886_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__76_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___102_comb = 10'h000;
  assign p1_smul_58890_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__78_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___103_comb = 10'h000;
  assign p1_smul_58896_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__81_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___104_comb = 10'h000;
  assign p1_smul_58900_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__83_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___105_comb = 10'h000;
  assign p1_smul_58902_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__84_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___106_comb = 10'h000;
  assign p1_smul_58906_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__86_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___107_comb = 10'h000;
  assign p1_smul_58912_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__89_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___108_comb = 10'h000;
  assign p1_smul_58916_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__91_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___109_comb = 10'h000;
  assign p1_smul_58918_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__92_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___110_comb = 10'h000;
  assign p1_smul_58922_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__94_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___111_comb = 10'h000;
  assign p1_smul_58928_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__97_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___112_comb = 10'h000;
  assign p1_smul_58932_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__99_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___113_comb = 10'h000;
  assign p1_smul_58934_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__100_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___114_comb = 10'h000;
  assign p1_smul_58938_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__102_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___115_comb = 10'h000;
  assign p1_smul_58944_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__105_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___116_comb = 10'h000;
  assign p1_smul_58948_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__107_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___117_comb = 10'h000;
  assign p1_smul_58950_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__108_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___118_comb = 10'h000;
  assign p1_smul_58954_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__110_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___119_comb = 10'h000;
  assign p1_smul_58960_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__113_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___120_comb = 10'h000;
  assign p1_smul_58964_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__115_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___121_comb = 10'h000;
  assign p1_smul_58966_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__116_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___122_comb = 10'h000;
  assign p1_smul_58970_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__118_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___123_comb = 10'h000;
  assign p1_smul_58976_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__121_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___124_comb = 10'h000;
  assign p1_smul_58980_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__123_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___125_comb = 10'h000;
  assign p1_smul_58982_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__124_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___126_comb = 10'h000;
  assign p1_smul_58986_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__126_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___127_comb = 10'h000;
  assign p1_smul_58990_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__64_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___224_comb = 9'h000;
  assign p1_smul_58992_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__65_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___225_comb = 9'h000;
  assign p1_smul_59002_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__70_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___226_comb = 9'h000;
  assign p1_smul_59004_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__71_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___227_comb = 9'h000;
  assign p1_smul_59006_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__72_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___228_comb = 9'h000;
  assign p1_smul_59008_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__73_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___229_comb = 9'h000;
  assign p1_smul_59018_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__78_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___230_comb = 9'h000;
  assign p1_smul_59020_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__79_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___231_comb = 9'h000;
  assign p1_smul_59022_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__80_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___232_comb = 9'h000;
  assign p1_smul_59024_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__81_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___233_comb = 9'h000;
  assign p1_smul_59034_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__86_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___234_comb = 9'h000;
  assign p1_smul_59036_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__87_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___235_comb = 9'h000;
  assign p1_smul_59038_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__88_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___236_comb = 9'h000;
  assign p1_smul_59040_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__89_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___237_comb = 9'h000;
  assign p1_smul_59050_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__94_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___238_comb = 9'h000;
  assign p1_smul_59052_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__95_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___239_comb = 9'h000;
  assign p1_smul_59054_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__96_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___240_comb = 9'h000;
  assign p1_smul_59056_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__97_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___241_comb = 9'h000;
  assign p1_smul_59066_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__102_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___242_comb = 9'h000;
  assign p1_smul_59068_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__103_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___243_comb = 9'h000;
  assign p1_smul_59070_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__104_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___244_comb = 9'h000;
  assign p1_smul_59072_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__105_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___245_comb = 9'h000;
  assign p1_smul_59082_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__110_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___246_comb = 9'h000;
  assign p1_smul_59084_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__111_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___247_comb = 9'h000;
  assign p1_smul_59086_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__112_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___248_comb = 9'h000;
  assign p1_smul_59088_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__113_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___249_comb = 9'h000;
  assign p1_smul_59098_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__118_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___250_comb = 9'h000;
  assign p1_smul_59100_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__119_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___251_comb = 9'h000;
  assign p1_smul_59102_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__120_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___252_comb = 9'h000;
  assign p1_smul_59104_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__121_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___253_comb = 9'h000;
  assign p1_smul_59114_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__126_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___254_comb = 9'h000;
  assign p1_smul_59116_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__127_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___255_comb = 9'h000;
  assign p1_smul_57326_TrailingBits___192_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___193_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___194_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___195_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___196_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___197_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___198_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___199_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___200_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___201_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___202_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___203_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___204_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___205_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___206_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___207_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___208_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___209_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___210_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___211_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___212_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___213_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___214_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___215_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___216_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___217_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___218_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___219_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___220_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___221_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___222_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___223_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___224_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___225_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___226_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___227_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___228_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___229_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___230_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___231_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___232_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___233_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___234_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___235_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___236_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___237_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___238_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___239_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___240_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___241_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___242_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___243_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___244_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___245_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___246_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___247_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___248_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___249_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___250_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___251_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___252_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___253_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___254_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___255_comb = 8'h00;
  assign p1_concat_139457_comb = {p1_smul_58226_NarrowedMult__comb, p1_smul_57330_TrailingBits___128_comb};
  assign p1_concat_139458_comb = {p1_smul_58228_NarrowedMult__comb, p1_smul_57330_TrailingBits___129_comb};
  assign p1_concat_139459_comb = {p1_smul_58230_NarrowedMult__comb, p1_smul_57330_TrailingBits___130_comb};
  assign p1_concat_139460_comb = {p1_smul_58232_NarrowedMult__comb, p1_smul_57330_TrailingBits___131_comb};
  assign p1_concat_139461_comb = {p1_smul_58242_NarrowedMult__comb, p1_smul_57330_TrailingBits___132_comb};
  assign p1_concat_139462_comb = {p1_smul_58244_NarrowedMult__comb, p1_smul_57330_TrailingBits___133_comb};
  assign p1_concat_139463_comb = {p1_smul_58246_NarrowedMult__comb, p1_smul_57330_TrailingBits___134_comb};
  assign p1_concat_139464_comb = {p1_smul_58248_NarrowedMult__comb, p1_smul_57330_TrailingBits___135_comb};
  assign p1_concat_139465_comb = {p1_smul_58258_NarrowedMult__comb, p1_smul_57330_TrailingBits___136_comb};
  assign p1_concat_139466_comb = {p1_smul_58260_NarrowedMult__comb, p1_smul_57330_TrailingBits___137_comb};
  assign p1_concat_139467_comb = {p1_smul_58262_NarrowedMult__comb, p1_smul_57330_TrailingBits___138_comb};
  assign p1_concat_139468_comb = {p1_smul_58264_NarrowedMult__comb, p1_smul_57330_TrailingBits___139_comb};
  assign p1_concat_139469_comb = {p1_smul_58274_NarrowedMult__comb, p1_smul_57330_TrailingBits___140_comb};
  assign p1_concat_139470_comb = {p1_smul_58276_NarrowedMult__comb, p1_smul_57330_TrailingBits___141_comb};
  assign p1_concat_139471_comb = {p1_smul_58278_NarrowedMult__comb, p1_smul_57330_TrailingBits___142_comb};
  assign p1_concat_139472_comb = {p1_smul_58280_NarrowedMult__comb, p1_smul_57330_TrailingBits___143_comb};
  assign p1_concat_139473_comb = {p1_smul_58290_NarrowedMult__comb, p1_smul_57330_TrailingBits___144_comb};
  assign p1_concat_139474_comb = {p1_smul_58292_NarrowedMult__comb, p1_smul_57330_TrailingBits___145_comb};
  assign p1_concat_139475_comb = {p1_smul_58294_NarrowedMult__comb, p1_smul_57330_TrailingBits___146_comb};
  assign p1_concat_139476_comb = {p1_smul_58296_NarrowedMult__comb, p1_smul_57330_TrailingBits___147_comb};
  assign p1_concat_139477_comb = {p1_smul_58306_NarrowedMult__comb, p1_smul_57330_TrailingBits___148_comb};
  assign p1_concat_139478_comb = {p1_smul_58308_NarrowedMult__comb, p1_smul_57330_TrailingBits___149_comb};
  assign p1_concat_139479_comb = {p1_smul_58310_NarrowedMult__comb, p1_smul_57330_TrailingBits___150_comb};
  assign p1_concat_139480_comb = {p1_smul_58312_NarrowedMult__comb, p1_smul_57330_TrailingBits___151_comb};
  assign p1_concat_139481_comb = {p1_smul_58322_NarrowedMult__comb, p1_smul_57330_TrailingBits___152_comb};
  assign p1_concat_139482_comb = {p1_smul_58324_NarrowedMult__comb, p1_smul_57330_TrailingBits___153_comb};
  assign p1_concat_139483_comb = {p1_smul_58326_NarrowedMult__comb, p1_smul_57330_TrailingBits___154_comb};
  assign p1_concat_139484_comb = {p1_smul_58328_NarrowedMult__comb, p1_smul_57330_TrailingBits___155_comb};
  assign p1_concat_139485_comb = {p1_smul_58338_NarrowedMult__comb, p1_smul_57330_TrailingBits___156_comb};
  assign p1_concat_139486_comb = {p1_smul_58340_NarrowedMult__comb, p1_smul_57330_TrailingBits___157_comb};
  assign p1_concat_139487_comb = {p1_smul_58342_NarrowedMult__comb, p1_smul_57330_TrailingBits___158_comb};
  assign p1_concat_139488_comb = {p1_smul_58344_NarrowedMult__comb, p1_smul_57330_TrailingBits___159_comb};
  assign p1_concat_139489_comb = {p1_smul_58350_NarrowedMult__comb, p1_smul_57454_TrailingBits___64_comb};
  assign p1_concat_139490_comb = {p1_smul_58356_NarrowedMult__comb, p1_smul_57454_TrailingBits___65_comb};
  assign p1_concat_139491_comb = {p1_smul_58358_NarrowedMult__comb, p1_smul_57454_TrailingBits___66_comb};
  assign p1_concat_139492_comb = {p1_smul_58364_NarrowedMult__comb, p1_smul_57454_TrailingBits___67_comb};
  assign p1_concat_139493_comb = {p1_smul_58366_NarrowedMult__comb, p1_smul_57454_TrailingBits___68_comb};
  assign p1_concat_139494_comb = {p1_smul_58372_NarrowedMult__comb, p1_smul_57454_TrailingBits___69_comb};
  assign p1_concat_139495_comb = {p1_smul_58374_NarrowedMult__comb, p1_smul_57454_TrailingBits___70_comb};
  assign p1_concat_139496_comb = {p1_smul_58380_NarrowedMult__comb, p1_smul_57454_TrailingBits___71_comb};
  assign p1_concat_139497_comb = {p1_smul_58382_NarrowedMult__comb, p1_smul_57454_TrailingBits___72_comb};
  assign p1_concat_139498_comb = {p1_smul_58388_NarrowedMult__comb, p1_smul_57454_TrailingBits___73_comb};
  assign p1_concat_139499_comb = {p1_smul_58390_NarrowedMult__comb, p1_smul_57454_TrailingBits___74_comb};
  assign p1_concat_139500_comb = {p1_smul_58396_NarrowedMult__comb, p1_smul_57454_TrailingBits___75_comb};
  assign p1_concat_139501_comb = {p1_smul_58398_NarrowedMult__comb, p1_smul_57454_TrailingBits___76_comb};
  assign p1_concat_139502_comb = {p1_smul_58404_NarrowedMult__comb, p1_smul_57454_TrailingBits___77_comb};
  assign p1_concat_139503_comb = {p1_smul_58406_NarrowedMult__comb, p1_smul_57454_TrailingBits___78_comb};
  assign p1_concat_139504_comb = {p1_smul_58412_NarrowedMult__comb, p1_smul_57454_TrailingBits___79_comb};
  assign p1_concat_139505_comb = {p1_smul_58414_NarrowedMult__comb, p1_smul_57454_TrailingBits___80_comb};
  assign p1_concat_139506_comb = {p1_smul_58420_NarrowedMult__comb, p1_smul_57454_TrailingBits___81_comb};
  assign p1_concat_139507_comb = {p1_smul_58422_NarrowedMult__comb, p1_smul_57454_TrailingBits___82_comb};
  assign p1_concat_139508_comb = {p1_smul_58428_NarrowedMult__comb, p1_smul_57454_TrailingBits___83_comb};
  assign p1_concat_139509_comb = {p1_smul_58430_NarrowedMult__comb, p1_smul_57454_TrailingBits___84_comb};
  assign p1_concat_139510_comb = {p1_smul_58436_NarrowedMult__comb, p1_smul_57454_TrailingBits___85_comb};
  assign p1_concat_139511_comb = {p1_smul_58438_NarrowedMult__comb, p1_smul_57454_TrailingBits___86_comb};
  assign p1_concat_139512_comb = {p1_smul_58444_NarrowedMult__comb, p1_smul_57454_TrailingBits___87_comb};
  assign p1_concat_139513_comb = {p1_smul_58446_NarrowedMult__comb, p1_smul_57454_TrailingBits___88_comb};
  assign p1_concat_139514_comb = {p1_smul_58452_NarrowedMult__comb, p1_smul_57454_TrailingBits___89_comb};
  assign p1_concat_139515_comb = {p1_smul_58454_NarrowedMult__comb, p1_smul_57454_TrailingBits___90_comb};
  assign p1_concat_139516_comb = {p1_smul_58460_NarrowedMult__comb, p1_smul_57454_TrailingBits___91_comb};
  assign p1_concat_139517_comb = {p1_smul_58462_NarrowedMult__comb, p1_smul_57454_TrailingBits___92_comb};
  assign p1_concat_139518_comb = {p1_smul_58468_NarrowedMult__comb, p1_smul_57454_TrailingBits___93_comb};
  assign p1_concat_139519_comb = {p1_smul_58470_NarrowedMult__comb, p1_smul_57454_TrailingBits___94_comb};
  assign p1_concat_139520_comb = {p1_smul_58476_NarrowedMult__comb, p1_smul_57454_TrailingBits___95_comb};
  assign p1_concat_139521_comb = {p1_smul_58480_NarrowedMult__comb, p1_smul_57330_TrailingBits___160_comb};
  assign p1_concat_139522_comb = {p1_smul_58484_NarrowedMult__comb, p1_smul_57330_TrailingBits___161_comb};
  assign p1_concat_139523_comb = {p1_smul_58486_NarrowedMult__comb, p1_smul_57330_TrailingBits___162_comb};
  assign p1_concat_139524_comb = {p1_smul_58490_NarrowedMult__comb, p1_smul_57330_TrailingBits___163_comb};
  assign p1_concat_139525_comb = {p1_smul_58496_NarrowedMult__comb, p1_smul_57330_TrailingBits___164_comb};
  assign p1_concat_139526_comb = {p1_smul_58500_NarrowedMult__comb, p1_smul_57330_TrailingBits___165_comb};
  assign p1_concat_139527_comb = {p1_smul_58502_NarrowedMult__comb, p1_smul_57330_TrailingBits___166_comb};
  assign p1_concat_139528_comb = {p1_smul_58506_NarrowedMult__comb, p1_smul_57330_TrailingBits___167_comb};
  assign p1_concat_139529_comb = {p1_smul_58512_NarrowedMult__comb, p1_smul_57330_TrailingBits___168_comb};
  assign p1_concat_139530_comb = {p1_smul_58516_NarrowedMult__comb, p1_smul_57330_TrailingBits___169_comb};
  assign p1_concat_139531_comb = {p1_smul_58518_NarrowedMult__comb, p1_smul_57330_TrailingBits___170_comb};
  assign p1_concat_139532_comb = {p1_smul_58522_NarrowedMult__comb, p1_smul_57330_TrailingBits___171_comb};
  assign p1_concat_139533_comb = {p1_smul_58528_NarrowedMult__comb, p1_smul_57330_TrailingBits___172_comb};
  assign p1_concat_139534_comb = {p1_smul_58532_NarrowedMult__comb, p1_smul_57330_TrailingBits___173_comb};
  assign p1_concat_139535_comb = {p1_smul_58534_NarrowedMult__comb, p1_smul_57330_TrailingBits___174_comb};
  assign p1_concat_139536_comb = {p1_smul_58538_NarrowedMult__comb, p1_smul_57330_TrailingBits___175_comb};
  assign p1_concat_139537_comb = {p1_smul_58544_NarrowedMult__comb, p1_smul_57330_TrailingBits___176_comb};
  assign p1_concat_139538_comb = {p1_smul_58548_NarrowedMult__comb, p1_smul_57330_TrailingBits___177_comb};
  assign p1_concat_139539_comb = {p1_smul_58550_NarrowedMult__comb, p1_smul_57330_TrailingBits___178_comb};
  assign p1_concat_139540_comb = {p1_smul_58554_NarrowedMult__comb, p1_smul_57330_TrailingBits___179_comb};
  assign p1_concat_139541_comb = {p1_smul_58560_NarrowedMult__comb, p1_smul_57330_TrailingBits___180_comb};
  assign p1_concat_139542_comb = {p1_smul_58564_NarrowedMult__comb, p1_smul_57330_TrailingBits___181_comb};
  assign p1_concat_139543_comb = {p1_smul_58566_NarrowedMult__comb, p1_smul_57330_TrailingBits___182_comb};
  assign p1_concat_139544_comb = {p1_smul_58570_NarrowedMult__comb, p1_smul_57330_TrailingBits___183_comb};
  assign p1_concat_139545_comb = {p1_smul_58576_NarrowedMult__comb, p1_smul_57330_TrailingBits___184_comb};
  assign p1_concat_139546_comb = {p1_smul_58580_NarrowedMult__comb, p1_smul_57330_TrailingBits___185_comb};
  assign p1_concat_139547_comb = {p1_smul_58582_NarrowedMult__comb, p1_smul_57330_TrailingBits___186_comb};
  assign p1_concat_139548_comb = {p1_smul_58586_NarrowedMult__comb, p1_smul_57330_TrailingBits___187_comb};
  assign p1_concat_139549_comb = {p1_smul_58592_NarrowedMult__comb, p1_smul_57330_TrailingBits___188_comb};
  assign p1_concat_139550_comb = {p1_smul_58596_NarrowedMult__comb, p1_smul_57330_TrailingBits___189_comb};
  assign p1_concat_139551_comb = {p1_smul_58598_NarrowedMult__comb, p1_smul_57330_TrailingBits___190_comb};
  assign p1_concat_139552_comb = {p1_smul_58602_NarrowedMult__comb, p1_smul_57330_TrailingBits___191_comb};
  assign p1_concat_139553_comb = {p1_smul_58734_NarrowedMult__comb, p1_smul_57330_TrailingBits___192_comb};
  assign p1_concat_139554_comb = {p1_smul_58738_NarrowedMult__comb, p1_smul_57330_TrailingBits___193_comb};
  assign p1_concat_139555_comb = {p1_smul_58744_NarrowedMult__comb, p1_smul_57330_TrailingBits___194_comb};
  assign p1_concat_139556_comb = {p1_smul_58748_NarrowedMult__comb, p1_smul_57330_TrailingBits___195_comb};
  assign p1_concat_139557_comb = {p1_smul_58750_NarrowedMult__comb, p1_smul_57330_TrailingBits___196_comb};
  assign p1_concat_139558_comb = {p1_smul_58754_NarrowedMult__comb, p1_smul_57330_TrailingBits___197_comb};
  assign p1_concat_139559_comb = {p1_smul_58760_NarrowedMult__comb, p1_smul_57330_TrailingBits___198_comb};
  assign p1_concat_139560_comb = {p1_smul_58764_NarrowedMult__comb, p1_smul_57330_TrailingBits___199_comb};
  assign p1_concat_139561_comb = {p1_smul_58766_NarrowedMult__comb, p1_smul_57330_TrailingBits___200_comb};
  assign p1_concat_139562_comb = {p1_smul_58770_NarrowedMult__comb, p1_smul_57330_TrailingBits___201_comb};
  assign p1_concat_139563_comb = {p1_smul_58776_NarrowedMult__comb, p1_smul_57330_TrailingBits___202_comb};
  assign p1_concat_139564_comb = {p1_smul_58780_NarrowedMult__comb, p1_smul_57330_TrailingBits___203_comb};
  assign p1_concat_139565_comb = {p1_smul_58782_NarrowedMult__comb, p1_smul_57330_TrailingBits___204_comb};
  assign p1_concat_139566_comb = {p1_smul_58786_NarrowedMult__comb, p1_smul_57330_TrailingBits___205_comb};
  assign p1_concat_139567_comb = {p1_smul_58792_NarrowedMult__comb, p1_smul_57330_TrailingBits___206_comb};
  assign p1_concat_139568_comb = {p1_smul_58796_NarrowedMult__comb, p1_smul_57330_TrailingBits___207_comb};
  assign p1_concat_139569_comb = {p1_smul_58798_NarrowedMult__comb, p1_smul_57330_TrailingBits___208_comb};
  assign p1_concat_139570_comb = {p1_smul_58802_NarrowedMult__comb, p1_smul_57330_TrailingBits___209_comb};
  assign p1_concat_139571_comb = {p1_smul_58808_NarrowedMult__comb, p1_smul_57330_TrailingBits___210_comb};
  assign p1_concat_139572_comb = {p1_smul_58812_NarrowedMult__comb, p1_smul_57330_TrailingBits___211_comb};
  assign p1_concat_139573_comb = {p1_smul_58814_NarrowedMult__comb, p1_smul_57330_TrailingBits___212_comb};
  assign p1_concat_139574_comb = {p1_smul_58818_NarrowedMult__comb, p1_smul_57330_TrailingBits___213_comb};
  assign p1_concat_139575_comb = {p1_smul_58824_NarrowedMult__comb, p1_smul_57330_TrailingBits___214_comb};
  assign p1_concat_139576_comb = {p1_smul_58828_NarrowedMult__comb, p1_smul_57330_TrailingBits___215_comb};
  assign p1_concat_139577_comb = {p1_smul_58830_NarrowedMult__comb, p1_smul_57330_TrailingBits___216_comb};
  assign p1_concat_139578_comb = {p1_smul_58834_NarrowedMult__comb, p1_smul_57330_TrailingBits___217_comb};
  assign p1_concat_139579_comb = {p1_smul_58840_NarrowedMult__comb, p1_smul_57330_TrailingBits___218_comb};
  assign p1_concat_139580_comb = {p1_smul_58844_NarrowedMult__comb, p1_smul_57330_TrailingBits___219_comb};
  assign p1_concat_139581_comb = {p1_smul_58846_NarrowedMult__comb, p1_smul_57330_TrailingBits___220_comb};
  assign p1_concat_139582_comb = {p1_smul_58850_NarrowedMult__comb, p1_smul_57330_TrailingBits___221_comb};
  assign p1_concat_139583_comb = {p1_smul_58856_NarrowedMult__comb, p1_smul_57330_TrailingBits___222_comb};
  assign p1_concat_139584_comb = {p1_smul_58860_NarrowedMult__comb, p1_smul_57330_TrailingBits___223_comb};
  assign p1_concat_139585_comb = {p1_smul_58864_NarrowedMult__comb, p1_smul_57454_TrailingBits___96_comb};
  assign p1_concat_139586_comb = {p1_smul_58868_NarrowedMult__comb, p1_smul_57454_TrailingBits___97_comb};
  assign p1_concat_139587_comb = {p1_smul_58870_NarrowedMult__comb, p1_smul_57454_TrailingBits___98_comb};
  assign p1_concat_139588_comb = {p1_smul_58874_NarrowedMult__comb, p1_smul_57454_TrailingBits___99_comb};
  assign p1_concat_139589_comb = {p1_smul_58880_NarrowedMult__comb, p1_smul_57454_TrailingBits___100_comb};
  assign p1_concat_139590_comb = {p1_smul_58884_NarrowedMult__comb, p1_smul_57454_TrailingBits___101_comb};
  assign p1_concat_139591_comb = {p1_smul_58886_NarrowedMult__comb, p1_smul_57454_TrailingBits___102_comb};
  assign p1_concat_139592_comb = {p1_smul_58890_NarrowedMult__comb, p1_smul_57454_TrailingBits___103_comb};
  assign p1_concat_139593_comb = {p1_smul_58896_NarrowedMult__comb, p1_smul_57454_TrailingBits___104_comb};
  assign p1_concat_139594_comb = {p1_smul_58900_NarrowedMult__comb, p1_smul_57454_TrailingBits___105_comb};
  assign p1_concat_139595_comb = {p1_smul_58902_NarrowedMult__comb, p1_smul_57454_TrailingBits___106_comb};
  assign p1_concat_139596_comb = {p1_smul_58906_NarrowedMult__comb, p1_smul_57454_TrailingBits___107_comb};
  assign p1_concat_139597_comb = {p1_smul_58912_NarrowedMult__comb, p1_smul_57454_TrailingBits___108_comb};
  assign p1_concat_139598_comb = {p1_smul_58916_NarrowedMult__comb, p1_smul_57454_TrailingBits___109_comb};
  assign p1_concat_139599_comb = {p1_smul_58918_NarrowedMult__comb, p1_smul_57454_TrailingBits___110_comb};
  assign p1_concat_139600_comb = {p1_smul_58922_NarrowedMult__comb, p1_smul_57454_TrailingBits___111_comb};
  assign p1_concat_139601_comb = {p1_smul_58928_NarrowedMult__comb, p1_smul_57454_TrailingBits___112_comb};
  assign p1_concat_139602_comb = {p1_smul_58932_NarrowedMult__comb, p1_smul_57454_TrailingBits___113_comb};
  assign p1_concat_139603_comb = {p1_smul_58934_NarrowedMult__comb, p1_smul_57454_TrailingBits___114_comb};
  assign p1_concat_139604_comb = {p1_smul_58938_NarrowedMult__comb, p1_smul_57454_TrailingBits___115_comb};
  assign p1_concat_139605_comb = {p1_smul_58944_NarrowedMult__comb, p1_smul_57454_TrailingBits___116_comb};
  assign p1_concat_139606_comb = {p1_smul_58948_NarrowedMult__comb, p1_smul_57454_TrailingBits___117_comb};
  assign p1_concat_139607_comb = {p1_smul_58950_NarrowedMult__comb, p1_smul_57454_TrailingBits___118_comb};
  assign p1_concat_139608_comb = {p1_smul_58954_NarrowedMult__comb, p1_smul_57454_TrailingBits___119_comb};
  assign p1_concat_139609_comb = {p1_smul_58960_NarrowedMult__comb, p1_smul_57454_TrailingBits___120_comb};
  assign p1_concat_139610_comb = {p1_smul_58964_NarrowedMult__comb, p1_smul_57454_TrailingBits___121_comb};
  assign p1_concat_139611_comb = {p1_smul_58966_NarrowedMult__comb, p1_smul_57454_TrailingBits___122_comb};
  assign p1_concat_139612_comb = {p1_smul_58970_NarrowedMult__comb, p1_smul_57454_TrailingBits___123_comb};
  assign p1_concat_139613_comb = {p1_smul_58976_NarrowedMult__comb, p1_smul_57454_TrailingBits___124_comb};
  assign p1_concat_139614_comb = {p1_smul_58980_NarrowedMult__comb, p1_smul_57454_TrailingBits___125_comb};
  assign p1_concat_139615_comb = {p1_smul_58982_NarrowedMult__comb, p1_smul_57454_TrailingBits___126_comb};
  assign p1_concat_139616_comb = {p1_smul_58986_NarrowedMult__comb, p1_smul_57454_TrailingBits___127_comb};
  assign p1_concat_139617_comb = {p1_smul_58990_NarrowedMult__comb, p1_smul_57330_TrailingBits___224_comb};
  assign p1_concat_139618_comb = {p1_smul_58992_NarrowedMult__comb, p1_smul_57330_TrailingBits___225_comb};
  assign p1_concat_139619_comb = {p1_smul_59002_NarrowedMult__comb, p1_smul_57330_TrailingBits___226_comb};
  assign p1_concat_139620_comb = {p1_smul_59004_NarrowedMult__comb, p1_smul_57330_TrailingBits___227_comb};
  assign p1_concat_139621_comb = {p1_smul_59006_NarrowedMult__comb, p1_smul_57330_TrailingBits___228_comb};
  assign p1_concat_139622_comb = {p1_smul_59008_NarrowedMult__comb, p1_smul_57330_TrailingBits___229_comb};
  assign p1_concat_139623_comb = {p1_smul_59018_NarrowedMult__comb, p1_smul_57330_TrailingBits___230_comb};
  assign p1_concat_139624_comb = {p1_smul_59020_NarrowedMult__comb, p1_smul_57330_TrailingBits___231_comb};
  assign p1_concat_139625_comb = {p1_smul_59022_NarrowedMult__comb, p1_smul_57330_TrailingBits___232_comb};
  assign p1_concat_139626_comb = {p1_smul_59024_NarrowedMult__comb, p1_smul_57330_TrailingBits___233_comb};
  assign p1_concat_139627_comb = {p1_smul_59034_NarrowedMult__comb, p1_smul_57330_TrailingBits___234_comb};
  assign p1_concat_139628_comb = {p1_smul_59036_NarrowedMult__comb, p1_smul_57330_TrailingBits___235_comb};
  assign p1_concat_139629_comb = {p1_smul_59038_NarrowedMult__comb, p1_smul_57330_TrailingBits___236_comb};
  assign p1_concat_139630_comb = {p1_smul_59040_NarrowedMult__comb, p1_smul_57330_TrailingBits___237_comb};
  assign p1_concat_139631_comb = {p1_smul_59050_NarrowedMult__comb, p1_smul_57330_TrailingBits___238_comb};
  assign p1_concat_139632_comb = {p1_smul_59052_NarrowedMult__comb, p1_smul_57330_TrailingBits___239_comb};
  assign p1_concat_139633_comb = {p1_smul_59054_NarrowedMult__comb, p1_smul_57330_TrailingBits___240_comb};
  assign p1_concat_139634_comb = {p1_smul_59056_NarrowedMult__comb, p1_smul_57330_TrailingBits___241_comb};
  assign p1_concat_139635_comb = {p1_smul_59066_NarrowedMult__comb, p1_smul_57330_TrailingBits___242_comb};
  assign p1_concat_139636_comb = {p1_smul_59068_NarrowedMult__comb, p1_smul_57330_TrailingBits___243_comb};
  assign p1_concat_139637_comb = {p1_smul_59070_NarrowedMult__comb, p1_smul_57330_TrailingBits___244_comb};
  assign p1_concat_139638_comb = {p1_smul_59072_NarrowedMult__comb, p1_smul_57330_TrailingBits___245_comb};
  assign p1_concat_139639_comb = {p1_smul_59082_NarrowedMult__comb, p1_smul_57330_TrailingBits___246_comb};
  assign p1_concat_139640_comb = {p1_smul_59084_NarrowedMult__comb, p1_smul_57330_TrailingBits___247_comb};
  assign p1_concat_139641_comb = {p1_smul_59086_NarrowedMult__comb, p1_smul_57330_TrailingBits___248_comb};
  assign p1_concat_139642_comb = {p1_smul_59088_NarrowedMult__comb, p1_smul_57330_TrailingBits___249_comb};
  assign p1_concat_139643_comb = {p1_smul_59098_NarrowedMult__comb, p1_smul_57330_TrailingBits___250_comb};
  assign p1_concat_139644_comb = {p1_smul_59100_NarrowedMult__comb, p1_smul_57330_TrailingBits___251_comb};
  assign p1_concat_139645_comb = {p1_smul_59102_NarrowedMult__comb, p1_smul_57330_TrailingBits___252_comb};
  assign p1_concat_139646_comb = {p1_smul_59104_NarrowedMult__comb, p1_smul_57330_TrailingBits___253_comb};
  assign p1_concat_139647_comb = {p1_smul_59114_NarrowedMult__comb, p1_smul_57330_TrailingBits___254_comb};
  assign p1_concat_139648_comb = {p1_smul_59116_NarrowedMult__comb, p1_smul_57330_TrailingBits___255_comb};
  assign p1_shifted__64_comb = {~p1_clipped__8_comb[7], p1_clipped__8_comb[6:0], p1_smul_57326_TrailingBits___192_comb};
  assign p1_smul_57326_TrailingBits___64_comb = 8'h00;
  assign p1_shifted__65_comb = {~p1_clipped__24_comb[7], p1_clipped__24_comb[6:0], p1_smul_57326_TrailingBits___193_comb};
  assign p1_smul_57326_TrailingBits___65_comb = 8'h00;
  assign p1_shifted__66_comb = {~p1_clipped__40_comb[7], p1_clipped__40_comb[6:0], p1_smul_57326_TrailingBits___194_comb};
  assign p1_smul_57326_TrailingBits___66_comb = 8'h00;
  assign p1_shifted__67_comb = {~p1_clipped__56_comb[7], p1_clipped__56_comb[6:0], p1_smul_57326_TrailingBits___195_comb};
  assign p1_smul_57326_TrailingBits___67_comb = 8'h00;
  assign p1_shifted__68_comb = {~p1_clipped__72_comb[7], p1_clipped__72_comb[6:0], p1_smul_57326_TrailingBits___196_comb};
  assign p1_smul_57326_TrailingBits___68_comb = 8'h00;
  assign p1_shifted__69_comb = {~p1_clipped__88_comb[7], p1_clipped__88_comb[6:0], p1_smul_57326_TrailingBits___197_comb};
  assign p1_smul_57326_TrailingBits___69_comb = 8'h00;
  assign p1_shifted__70_comb = {~p1_clipped__104_comb[7], p1_clipped__104_comb[6:0], p1_smul_57326_TrailingBits___198_comb};
  assign p1_smul_57326_TrailingBits___70_comb = 8'h00;
  assign p1_shifted__71_comb = {~p1_clipped__120_comb[7], p1_clipped__120_comb[6:0], p1_smul_57326_TrailingBits___199_comb};
  assign p1_smul_57326_TrailingBits___71_comb = 8'h00;
  assign p1_shifted__72_comb = {~p1_clipped__9_comb[7], p1_clipped__9_comb[6:0], p1_smul_57326_TrailingBits___200_comb};
  assign p1_smul_57326_TrailingBits___72_comb = 8'h00;
  assign p1_shifted__73_comb = {~p1_clipped__25_comb[7], p1_clipped__25_comb[6:0], p1_smul_57326_TrailingBits___201_comb};
  assign p1_smul_57326_TrailingBits___73_comb = 8'h00;
  assign p1_shifted__74_comb = {~p1_clipped__41_comb[7], p1_clipped__41_comb[6:0], p1_smul_57326_TrailingBits___202_comb};
  assign p1_smul_57326_TrailingBits___74_comb = 8'h00;
  assign p1_shifted__75_comb = {~p1_clipped__57_comb[7], p1_clipped__57_comb[6:0], p1_smul_57326_TrailingBits___203_comb};
  assign p1_smul_57326_TrailingBits___75_comb = 8'h00;
  assign p1_shifted__76_comb = {~p1_clipped__73_comb[7], p1_clipped__73_comb[6:0], p1_smul_57326_TrailingBits___204_comb};
  assign p1_smul_57326_TrailingBits___76_comb = 8'h00;
  assign p1_shifted__77_comb = {~p1_clipped__89_comb[7], p1_clipped__89_comb[6:0], p1_smul_57326_TrailingBits___205_comb};
  assign p1_smul_57326_TrailingBits___77_comb = 8'h00;
  assign p1_shifted__78_comb = {~p1_clipped__105_comb[7], p1_clipped__105_comb[6:0], p1_smul_57326_TrailingBits___206_comb};
  assign p1_smul_57326_TrailingBits___78_comb = 8'h00;
  assign p1_shifted__79_comb = {~p1_clipped__121_comb[7], p1_clipped__121_comb[6:0], p1_smul_57326_TrailingBits___207_comb};
  assign p1_smul_57326_TrailingBits___79_comb = 8'h00;
  assign p1_shifted__80_comb = {~p1_clipped__10_comb[7], p1_clipped__10_comb[6:0], p1_smul_57326_TrailingBits___208_comb};
  assign p1_smul_57326_TrailingBits___80_comb = 8'h00;
  assign p1_shifted__81_comb = {~p1_clipped__26_comb[7], p1_clipped__26_comb[6:0], p1_smul_57326_TrailingBits___209_comb};
  assign p1_smul_57326_TrailingBits___81_comb = 8'h00;
  assign p1_shifted__82_comb = {~p1_clipped__42_comb[7], p1_clipped__42_comb[6:0], p1_smul_57326_TrailingBits___210_comb};
  assign p1_smul_57326_TrailingBits___82_comb = 8'h00;
  assign p1_shifted__83_comb = {~p1_clipped__58_comb[7], p1_clipped__58_comb[6:0], p1_smul_57326_TrailingBits___211_comb};
  assign p1_smul_57326_TrailingBits___83_comb = 8'h00;
  assign p1_shifted__84_comb = {~p1_clipped__74_comb[7], p1_clipped__74_comb[6:0], p1_smul_57326_TrailingBits___212_comb};
  assign p1_smul_57326_TrailingBits___84_comb = 8'h00;
  assign p1_shifted__85_comb = {~p1_clipped__90_comb[7], p1_clipped__90_comb[6:0], p1_smul_57326_TrailingBits___213_comb};
  assign p1_smul_57326_TrailingBits___85_comb = 8'h00;
  assign p1_shifted__86_comb = {~p1_clipped__106_comb[7], p1_clipped__106_comb[6:0], p1_smul_57326_TrailingBits___214_comb};
  assign p1_smul_57326_TrailingBits___86_comb = 8'h00;
  assign p1_shifted__87_comb = {~p1_clipped__122_comb[7], p1_clipped__122_comb[6:0], p1_smul_57326_TrailingBits___215_comb};
  assign p1_smul_57326_TrailingBits___87_comb = 8'h00;
  assign p1_shifted__88_comb = {~p1_clipped__11_comb[7], p1_clipped__11_comb[6:0], p1_smul_57326_TrailingBits___216_comb};
  assign p1_smul_57326_TrailingBits___88_comb = 8'h00;
  assign p1_shifted__89_comb = {~p1_clipped__27_comb[7], p1_clipped__27_comb[6:0], p1_smul_57326_TrailingBits___217_comb};
  assign p1_smul_57326_TrailingBits___89_comb = 8'h00;
  assign p1_shifted__90_comb = {~p1_clipped__43_comb[7], p1_clipped__43_comb[6:0], p1_smul_57326_TrailingBits___218_comb};
  assign p1_smul_57326_TrailingBits___90_comb = 8'h00;
  assign p1_shifted__91_comb = {~p1_clipped__59_comb[7], p1_clipped__59_comb[6:0], p1_smul_57326_TrailingBits___219_comb};
  assign p1_smul_57326_TrailingBits___91_comb = 8'h00;
  assign p1_shifted__92_comb = {~p1_clipped__75_comb[7], p1_clipped__75_comb[6:0], p1_smul_57326_TrailingBits___220_comb};
  assign p1_smul_57326_TrailingBits___92_comb = 8'h00;
  assign p1_shifted__93_comb = {~p1_clipped__91_comb[7], p1_clipped__91_comb[6:0], p1_smul_57326_TrailingBits___221_comb};
  assign p1_smul_57326_TrailingBits___93_comb = 8'h00;
  assign p1_shifted__94_comb = {~p1_clipped__107_comb[7], p1_clipped__107_comb[6:0], p1_smul_57326_TrailingBits___222_comb};
  assign p1_smul_57326_TrailingBits___94_comb = 8'h00;
  assign p1_shifted__95_comb = {~p1_clipped__123_comb[7], p1_clipped__123_comb[6:0], p1_smul_57326_TrailingBits___223_comb};
  assign p1_smul_57326_TrailingBits___95_comb = 8'h00;
  assign p1_shifted__96_comb = {~p1_clipped__12_comb[7], p1_clipped__12_comb[6:0], p1_smul_57326_TrailingBits___224_comb};
  assign p1_smul_57326_TrailingBits___96_comb = 8'h00;
  assign p1_shifted__97_comb = {~p1_clipped__28_comb[7], p1_clipped__28_comb[6:0], p1_smul_57326_TrailingBits___225_comb};
  assign p1_smul_57326_TrailingBits___97_comb = 8'h00;
  assign p1_shifted__98_comb = {~p1_clipped__44_comb[7], p1_clipped__44_comb[6:0], p1_smul_57326_TrailingBits___226_comb};
  assign p1_smul_57326_TrailingBits___98_comb = 8'h00;
  assign p1_shifted__99_comb = {~p1_clipped__60_comb[7], p1_clipped__60_comb[6:0], p1_smul_57326_TrailingBits___227_comb};
  assign p1_smul_57326_TrailingBits___99_comb = 8'h00;
  assign p1_shifted__100_comb = {~p1_clipped__76_comb[7], p1_clipped__76_comb[6:0], p1_smul_57326_TrailingBits___228_comb};
  assign p1_smul_57326_TrailingBits___100_comb = 8'h00;
  assign p1_shifted__101_comb = {~p1_clipped__92_comb[7], p1_clipped__92_comb[6:0], p1_smul_57326_TrailingBits___229_comb};
  assign p1_smul_57326_TrailingBits___101_comb = 8'h00;
  assign p1_shifted__102_comb = {~p1_clipped__108_comb[7], p1_clipped__108_comb[6:0], p1_smul_57326_TrailingBits___230_comb};
  assign p1_smul_57326_TrailingBits___102_comb = 8'h00;
  assign p1_shifted__103_comb = {~p1_clipped__124_comb[7], p1_clipped__124_comb[6:0], p1_smul_57326_TrailingBits___231_comb};
  assign p1_smul_57326_TrailingBits___103_comb = 8'h00;
  assign p1_shifted__104_comb = {~p1_clipped__13_comb[7], p1_clipped__13_comb[6:0], p1_smul_57326_TrailingBits___232_comb};
  assign p1_smul_57326_TrailingBits___104_comb = 8'h00;
  assign p1_shifted__105_comb = {~p1_clipped__29_comb[7], p1_clipped__29_comb[6:0], p1_smul_57326_TrailingBits___233_comb};
  assign p1_smul_57326_TrailingBits___105_comb = 8'h00;
  assign p1_shifted__106_comb = {~p1_clipped__45_comb[7], p1_clipped__45_comb[6:0], p1_smul_57326_TrailingBits___234_comb};
  assign p1_smul_57326_TrailingBits___106_comb = 8'h00;
  assign p1_shifted__107_comb = {~p1_clipped__61_comb[7], p1_clipped__61_comb[6:0], p1_smul_57326_TrailingBits___235_comb};
  assign p1_smul_57326_TrailingBits___107_comb = 8'h00;
  assign p1_shifted__108_comb = {~p1_clipped__77_comb[7], p1_clipped__77_comb[6:0], p1_smul_57326_TrailingBits___236_comb};
  assign p1_smul_57326_TrailingBits___108_comb = 8'h00;
  assign p1_shifted__109_comb = {~p1_clipped__93_comb[7], p1_clipped__93_comb[6:0], p1_smul_57326_TrailingBits___237_comb};
  assign p1_smul_57326_TrailingBits___109_comb = 8'h00;
  assign p1_shifted__110_comb = {~p1_clipped__109_comb[7], p1_clipped__109_comb[6:0], p1_smul_57326_TrailingBits___238_comb};
  assign p1_smul_57326_TrailingBits___110_comb = 8'h00;
  assign p1_shifted__111_comb = {~p1_clipped__125_comb[7], p1_clipped__125_comb[6:0], p1_smul_57326_TrailingBits___239_comb};
  assign p1_smul_57326_TrailingBits___111_comb = 8'h00;
  assign p1_shifted__112_comb = {~p1_clipped__14_comb[7], p1_clipped__14_comb[6:0], p1_smul_57326_TrailingBits___240_comb};
  assign p1_smul_57326_TrailingBits___112_comb = 8'h00;
  assign p1_shifted__113_comb = {~p1_clipped__30_comb[7], p1_clipped__30_comb[6:0], p1_smul_57326_TrailingBits___241_comb};
  assign p1_smul_57326_TrailingBits___113_comb = 8'h00;
  assign p1_shifted__114_comb = {~p1_clipped__46_comb[7], p1_clipped__46_comb[6:0], p1_smul_57326_TrailingBits___242_comb};
  assign p1_smul_57326_TrailingBits___114_comb = 8'h00;
  assign p1_shifted__115_comb = {~p1_clipped__62_comb[7], p1_clipped__62_comb[6:0], p1_smul_57326_TrailingBits___243_comb};
  assign p1_smul_57326_TrailingBits___115_comb = 8'h00;
  assign p1_shifted__116_comb = {~p1_clipped__78_comb[7], p1_clipped__78_comb[6:0], p1_smul_57326_TrailingBits___244_comb};
  assign p1_smul_57326_TrailingBits___116_comb = 8'h00;
  assign p1_shifted__117_comb = {~p1_clipped__94_comb[7], p1_clipped__94_comb[6:0], p1_smul_57326_TrailingBits___245_comb};
  assign p1_smul_57326_TrailingBits___117_comb = 8'h00;
  assign p1_shifted__118_comb = {~p1_clipped__110_comb[7], p1_clipped__110_comb[6:0], p1_smul_57326_TrailingBits___246_comb};
  assign p1_smul_57326_TrailingBits___118_comb = 8'h00;
  assign p1_shifted__119_comb = {~p1_clipped__126_comb[7], p1_clipped__126_comb[6:0], p1_smul_57326_TrailingBits___247_comb};
  assign p1_smul_57326_TrailingBits___119_comb = 8'h00;
  assign p1_shifted__120_comb = {~p1_clipped__15_comb[7], p1_clipped__15_comb[6:0], p1_smul_57326_TrailingBits___248_comb};
  assign p1_smul_57326_TrailingBits___120_comb = 8'h00;
  assign p1_shifted__121_comb = {~p1_clipped__31_comb[7], p1_clipped__31_comb[6:0], p1_smul_57326_TrailingBits___249_comb};
  assign p1_smul_57326_TrailingBits___121_comb = 8'h00;
  assign p1_shifted__122_comb = {~p1_clipped__47_comb[7], p1_clipped__47_comb[6:0], p1_smul_57326_TrailingBits___250_comb};
  assign p1_smul_57326_TrailingBits___122_comb = 8'h00;
  assign p1_shifted__123_comb = {~p1_clipped__63_comb[7], p1_clipped__63_comb[6:0], p1_smul_57326_TrailingBits___251_comb};
  assign p1_smul_57326_TrailingBits___123_comb = 8'h00;
  assign p1_shifted__124_comb = {~p1_clipped__79_comb[7], p1_clipped__79_comb[6:0], p1_smul_57326_TrailingBits___252_comb};
  assign p1_smul_57326_TrailingBits___124_comb = 8'h00;
  assign p1_shifted__125_comb = {~p1_clipped__95_comb[7], p1_clipped__95_comb[6:0], p1_smul_57326_TrailingBits___253_comb};
  assign p1_smul_57326_TrailingBits___125_comb = 8'h00;
  assign p1_shifted__126_comb = {~p1_clipped__111_comb[7], p1_clipped__111_comb[6:0], p1_smul_57326_TrailingBits___254_comb};
  assign p1_smul_57326_TrailingBits___126_comb = 8'h00;
  assign p1_shifted__127_comb = {~p1_clipped__127_comb[7], p1_clipped__127_comb[6:0], p1_smul_57326_TrailingBits___255_comb};
  assign p1_smul_57326_TrailingBits___127_comb = 8'h00;
  assign p1_prod__519_comb = {{7{p1_concat_139457_comb[24]}}, p1_concat_139457_comb};
  assign p1_prod__523_comb = {{9{p1_concat_139458_comb[22]}}, p1_concat_139458_comb};
  assign p1_prod__528_comb = {{9{p1_concat_139459_comb[22]}}, p1_concat_139459_comb};
  assign p1_prod__534_comb = {{7{p1_concat_139460_comb[24]}}, p1_concat_139460_comb};
  assign p1_prod__583_comb = {{7{p1_concat_139461_comb[24]}}, p1_concat_139461_comb};
  assign p1_prod__587_comb = {{9{p1_concat_139462_comb[22]}}, p1_concat_139462_comb};
  assign p1_prod__592_comb = {{9{p1_concat_139463_comb[22]}}, p1_concat_139463_comb};
  assign p1_prod__598_comb = {{7{p1_concat_139464_comb[24]}}, p1_concat_139464_comb};
  assign p1_prod__647_comb = {{7{p1_concat_139465_comb[24]}}, p1_concat_139465_comb};
  assign p1_prod__651_comb = {{9{p1_concat_139466_comb[22]}}, p1_concat_139466_comb};
  assign p1_prod__656_comb = {{9{p1_concat_139467_comb[22]}}, p1_concat_139467_comb};
  assign p1_prod__662_comb = {{7{p1_concat_139468_comb[24]}}, p1_concat_139468_comb};
  assign p1_prod__711_comb = {{7{p1_concat_139469_comb[24]}}, p1_concat_139469_comb};
  assign p1_prod__715_comb = {{9{p1_concat_139470_comb[22]}}, p1_concat_139470_comb};
  assign p1_prod__720_comb = {{9{p1_concat_139471_comb[22]}}, p1_concat_139471_comb};
  assign p1_prod__726_comb = {{7{p1_concat_139472_comb[24]}}, p1_concat_139472_comb};
  assign p1_prod__775_comb = {{7{p1_concat_139473_comb[24]}}, p1_concat_139473_comb};
  assign p1_prod__779_comb = {{9{p1_concat_139474_comb[22]}}, p1_concat_139474_comb};
  assign p1_prod__784_comb = {{9{p1_concat_139475_comb[22]}}, p1_concat_139475_comb};
  assign p1_prod__790_comb = {{7{p1_concat_139476_comb[24]}}, p1_concat_139476_comb};
  assign p1_prod__839_comb = {{7{p1_concat_139477_comb[24]}}, p1_concat_139477_comb};
  assign p1_prod__843_comb = {{9{p1_concat_139478_comb[22]}}, p1_concat_139478_comb};
  assign p1_prod__848_comb = {{9{p1_concat_139479_comb[22]}}, p1_concat_139479_comb};
  assign p1_prod__854_comb = {{7{p1_concat_139480_comb[24]}}, p1_concat_139480_comb};
  assign p1_prod__903_comb = {{7{p1_concat_139481_comb[24]}}, p1_concat_139481_comb};
  assign p1_prod__907_comb = {{9{p1_concat_139482_comb[22]}}, p1_concat_139482_comb};
  assign p1_prod__912_comb = {{9{p1_concat_139483_comb[22]}}, p1_concat_139483_comb};
  assign p1_prod__918_comb = {{7{p1_concat_139484_comb[24]}}, p1_concat_139484_comb};
  assign p1_prod__967_comb = {{7{p1_concat_139485_comb[24]}}, p1_concat_139485_comb};
  assign p1_prod__971_comb = {{9{p1_concat_139486_comb[22]}}, p1_concat_139486_comb};
  assign p1_prod__976_comb = {{9{p1_concat_139487_comb[22]}}, p1_concat_139487_comb};
  assign p1_prod__982_comb = {{7{p1_concat_139488_comb[24]}}, p1_concat_139488_comb};
  assign p1_prod__517_comb = {{7{p1_concat_139489_comb[24]}}, p1_concat_139489_comb};
  assign p1_prod__529_comb = {{7{p1_concat_139490_comb[24]}}, p1_concat_139490_comb};
  assign p1_prod__535_comb = {{7{p1_concat_139491_comb[24]}}, p1_concat_139491_comb};
  assign p1_prod__555_comb = {{7{p1_concat_139492_comb[24]}}, p1_concat_139492_comb};
  assign p1_prod__581_comb = {{7{p1_concat_139493_comb[24]}}, p1_concat_139493_comb};
  assign p1_prod__593_comb = {{7{p1_concat_139494_comb[24]}}, p1_concat_139494_comb};
  assign p1_prod__599_comb = {{7{p1_concat_139495_comb[24]}}, p1_concat_139495_comb};
  assign p1_prod__619_comb = {{7{p1_concat_139496_comb[24]}}, p1_concat_139496_comb};
  assign p1_prod__645_comb = {{7{p1_concat_139497_comb[24]}}, p1_concat_139497_comb};
  assign p1_prod__657_comb = {{7{p1_concat_139498_comb[24]}}, p1_concat_139498_comb};
  assign p1_prod__663_comb = {{7{p1_concat_139499_comb[24]}}, p1_concat_139499_comb};
  assign p1_prod__683_comb = {{7{p1_concat_139500_comb[24]}}, p1_concat_139500_comb};
  assign p1_prod__709_comb = {{7{p1_concat_139501_comb[24]}}, p1_concat_139501_comb};
  assign p1_prod__721_comb = {{7{p1_concat_139502_comb[24]}}, p1_concat_139502_comb};
  assign p1_prod__727_comb = {{7{p1_concat_139503_comb[24]}}, p1_concat_139503_comb};
  assign p1_prod__747_comb = {{7{p1_concat_139504_comb[24]}}, p1_concat_139504_comb};
  assign p1_prod__773_comb = {{7{p1_concat_139505_comb[24]}}, p1_concat_139505_comb};
  assign p1_prod__785_comb = {{7{p1_concat_139506_comb[24]}}, p1_concat_139506_comb};
  assign p1_prod__791_comb = {{7{p1_concat_139507_comb[24]}}, p1_concat_139507_comb};
  assign p1_prod__811_comb = {{7{p1_concat_139508_comb[24]}}, p1_concat_139508_comb};
  assign p1_prod__837_comb = {{7{p1_concat_139509_comb[24]}}, p1_concat_139509_comb};
  assign p1_prod__849_comb = {{7{p1_concat_139510_comb[24]}}, p1_concat_139510_comb};
  assign p1_prod__855_comb = {{7{p1_concat_139511_comb[24]}}, p1_concat_139511_comb};
  assign p1_prod__875_comb = {{7{p1_concat_139512_comb[24]}}, p1_concat_139512_comb};
  assign p1_prod__901_comb = {{7{p1_concat_139513_comb[24]}}, p1_concat_139513_comb};
  assign p1_prod__913_comb = {{7{p1_concat_139514_comb[24]}}, p1_concat_139514_comb};
  assign p1_prod__919_comb = {{7{p1_concat_139515_comb[24]}}, p1_concat_139515_comb};
  assign p1_prod__939_comb = {{7{p1_concat_139516_comb[24]}}, p1_concat_139516_comb};
  assign p1_prod__965_comb = {{7{p1_concat_139517_comb[24]}}, p1_concat_139517_comb};
  assign p1_prod__977_comb = {{7{p1_concat_139518_comb[24]}}, p1_concat_139518_comb};
  assign p1_prod__983_comb = {{7{p1_concat_139519_comb[24]}}, p1_concat_139519_comb};
  assign p1_prod__1003_comb = {{7{p1_concat_139520_comb[24]}}, p1_concat_139520_comb};
  assign p1_prod__525_comb = {{9{p1_concat_139521_comb[22]}}, p1_concat_139521_comb};
  assign p1_prod__536_comb = {{7{p1_concat_139522_comb[24]}}, p1_concat_139522_comb};
  assign p1_prod__543_comb = {{7{p1_concat_139523_comb[24]}}, p1_concat_139523_comb};
  assign p1_prod__556_comb = {{9{p1_concat_139524_comb[22]}}, p1_concat_139524_comb};
  assign p1_prod__589_comb = {{9{p1_concat_139525_comb[22]}}, p1_concat_139525_comb};
  assign p1_prod__600_comb = {{7{p1_concat_139526_comb[24]}}, p1_concat_139526_comb};
  assign p1_prod__607_comb = {{7{p1_concat_139527_comb[24]}}, p1_concat_139527_comb};
  assign p1_prod__620_comb = {{9{p1_concat_139528_comb[22]}}, p1_concat_139528_comb};
  assign p1_prod__653_comb = {{9{p1_concat_139529_comb[22]}}, p1_concat_139529_comb};
  assign p1_prod__664_comb = {{7{p1_concat_139530_comb[24]}}, p1_concat_139530_comb};
  assign p1_prod__671_comb = {{7{p1_concat_139531_comb[24]}}, p1_concat_139531_comb};
  assign p1_prod__684_comb = {{9{p1_concat_139532_comb[22]}}, p1_concat_139532_comb};
  assign p1_prod__717_comb = {{9{p1_concat_139533_comb[22]}}, p1_concat_139533_comb};
  assign p1_prod__728_comb = {{7{p1_concat_139534_comb[24]}}, p1_concat_139534_comb};
  assign p1_prod__735_comb = {{7{p1_concat_139535_comb[24]}}, p1_concat_139535_comb};
  assign p1_prod__748_comb = {{9{p1_concat_139536_comb[22]}}, p1_concat_139536_comb};
  assign p1_prod__781_comb = {{9{p1_concat_139537_comb[22]}}, p1_concat_139537_comb};
  assign p1_prod__792_comb = {{7{p1_concat_139538_comb[24]}}, p1_concat_139538_comb};
  assign p1_prod__799_comb = {{7{p1_concat_139539_comb[24]}}, p1_concat_139539_comb};
  assign p1_prod__812_comb = {{9{p1_concat_139540_comb[22]}}, p1_concat_139540_comb};
  assign p1_prod__845_comb = {{9{p1_concat_139541_comb[22]}}, p1_concat_139541_comb};
  assign p1_prod__856_comb = {{7{p1_concat_139542_comb[24]}}, p1_concat_139542_comb};
  assign p1_prod__863_comb = {{7{p1_concat_139543_comb[24]}}, p1_concat_139543_comb};
  assign p1_prod__876_comb = {{9{p1_concat_139544_comb[22]}}, p1_concat_139544_comb};
  assign p1_prod__909_comb = {{9{p1_concat_139545_comb[22]}}, p1_concat_139545_comb};
  assign p1_prod__920_comb = {{7{p1_concat_139546_comb[24]}}, p1_concat_139546_comb};
  assign p1_prod__927_comb = {{7{p1_concat_139547_comb[24]}}, p1_concat_139547_comb};
  assign p1_prod__940_comb = {{9{p1_concat_139548_comb[22]}}, p1_concat_139548_comb};
  assign p1_prod__973_comb = {{9{p1_concat_139549_comb[22]}}, p1_concat_139549_comb};
  assign p1_prod__984_comb = {{7{p1_concat_139550_comb[24]}}, p1_concat_139550_comb};
  assign p1_prod__991_comb = {{7{p1_concat_139551_comb[24]}}, p1_concat_139551_comb};
  assign p1_prod__1004_comb = {{9{p1_concat_139552_comb[22]}}, p1_concat_139552_comb};
  assign p1_prod__532_comb = {{7{p1_concat_139553_comb[24]}}, p1_concat_139553_comb};
  assign p1_prod__545_comb = {{9{p1_concat_139554_comb[22]}}, p1_concat_139554_comb};
  assign p1_prod__563_comb = {{9{p1_concat_139555_comb[22]}}, p1_concat_139555_comb};
  assign p1_prod__570_comb = {{7{p1_concat_139556_comb[24]}}, p1_concat_139556_comb};
  assign p1_prod__596_comb = {{7{p1_concat_139557_comb[24]}}, p1_concat_139557_comb};
  assign p1_prod__609_comb = {{9{p1_concat_139558_comb[22]}}, p1_concat_139558_comb};
  assign p1_prod__627_comb = {{9{p1_concat_139559_comb[22]}}, p1_concat_139559_comb};
  assign p1_prod__634_comb = {{7{p1_concat_139560_comb[24]}}, p1_concat_139560_comb};
  assign p1_prod__660_comb = {{7{p1_concat_139561_comb[24]}}, p1_concat_139561_comb};
  assign p1_prod__673_comb = {{9{p1_concat_139562_comb[22]}}, p1_concat_139562_comb};
  assign p1_prod__691_comb = {{9{p1_concat_139563_comb[22]}}, p1_concat_139563_comb};
  assign p1_prod__698_comb = {{7{p1_concat_139564_comb[24]}}, p1_concat_139564_comb};
  assign p1_prod__724_comb = {{7{p1_concat_139565_comb[24]}}, p1_concat_139565_comb};
  assign p1_prod__737_comb = {{9{p1_concat_139566_comb[22]}}, p1_concat_139566_comb};
  assign p1_prod__755_comb = {{9{p1_concat_139567_comb[22]}}, p1_concat_139567_comb};
  assign p1_prod__762_comb = {{7{p1_concat_139568_comb[24]}}, p1_concat_139568_comb};
  assign p1_prod__788_comb = {{7{p1_concat_139569_comb[24]}}, p1_concat_139569_comb};
  assign p1_prod__801_comb = {{9{p1_concat_139570_comb[22]}}, p1_concat_139570_comb};
  assign p1_prod__819_comb = {{9{p1_concat_139571_comb[22]}}, p1_concat_139571_comb};
  assign p1_prod__826_comb = {{7{p1_concat_139572_comb[24]}}, p1_concat_139572_comb};
  assign p1_prod__852_comb = {{7{p1_concat_139573_comb[24]}}, p1_concat_139573_comb};
  assign p1_prod__865_comb = {{9{p1_concat_139574_comb[22]}}, p1_concat_139574_comb};
  assign p1_prod__883_comb = {{9{p1_concat_139575_comb[22]}}, p1_concat_139575_comb};
  assign p1_prod__890_comb = {{7{p1_concat_139576_comb[24]}}, p1_concat_139576_comb};
  assign p1_prod__916_comb = {{7{p1_concat_139577_comb[24]}}, p1_concat_139577_comb};
  assign p1_prod__929_comb = {{9{p1_concat_139578_comb[22]}}, p1_concat_139578_comb};
  assign p1_prod__947_comb = {{9{p1_concat_139579_comb[22]}}, p1_concat_139579_comb};
  assign p1_prod__954_comb = {{7{p1_concat_139580_comb[24]}}, p1_concat_139580_comb};
  assign p1_prod__980_comb = {{7{p1_concat_139581_comb[24]}}, p1_concat_139581_comb};
  assign p1_prod__993_comb = {{9{p1_concat_139582_comb[22]}}, p1_concat_139582_comb};
  assign p1_prod__1011_comb = {{9{p1_concat_139583_comb[22]}}, p1_concat_139583_comb};
  assign p1_prod__1018_comb = {{7{p1_concat_139584_comb[24]}}, p1_concat_139584_comb};
  assign p1_prod__546_comb = {{7{p1_concat_139585_comb[24]}}, p1_concat_139585_comb};
  assign p1_prod__559_comb = {{7{p1_concat_139586_comb[24]}}, p1_concat_139586_comb};
  assign p1_prod__564_comb = {{7{p1_concat_139587_comb[24]}}, p1_concat_139587_comb};
  assign p1_prod__571_comb = {{7{p1_concat_139588_comb[24]}}, p1_concat_139588_comb};
  assign p1_prod__610_comb = {{7{p1_concat_139589_comb[24]}}, p1_concat_139589_comb};
  assign p1_prod__623_comb = {{7{p1_concat_139590_comb[24]}}, p1_concat_139590_comb};
  assign p1_prod__628_comb = {{7{p1_concat_139591_comb[24]}}, p1_concat_139591_comb};
  assign p1_prod__635_comb = {{7{p1_concat_139592_comb[24]}}, p1_concat_139592_comb};
  assign p1_prod__674_comb = {{7{p1_concat_139593_comb[24]}}, p1_concat_139593_comb};
  assign p1_prod__687_comb = {{7{p1_concat_139594_comb[24]}}, p1_concat_139594_comb};
  assign p1_prod__692_comb = {{7{p1_concat_139595_comb[24]}}, p1_concat_139595_comb};
  assign p1_prod__699_comb = {{7{p1_concat_139596_comb[24]}}, p1_concat_139596_comb};
  assign p1_prod__738_comb = {{7{p1_concat_139597_comb[24]}}, p1_concat_139597_comb};
  assign p1_prod__751_comb = {{7{p1_concat_139598_comb[24]}}, p1_concat_139598_comb};
  assign p1_prod__756_comb = {{7{p1_concat_139599_comb[24]}}, p1_concat_139599_comb};
  assign p1_prod__763_comb = {{7{p1_concat_139600_comb[24]}}, p1_concat_139600_comb};
  assign p1_prod__802_comb = {{7{p1_concat_139601_comb[24]}}, p1_concat_139601_comb};
  assign p1_prod__815_comb = {{7{p1_concat_139602_comb[24]}}, p1_concat_139602_comb};
  assign p1_prod__820_comb = {{7{p1_concat_139603_comb[24]}}, p1_concat_139603_comb};
  assign p1_prod__827_comb = {{7{p1_concat_139604_comb[24]}}, p1_concat_139604_comb};
  assign p1_prod__866_comb = {{7{p1_concat_139605_comb[24]}}, p1_concat_139605_comb};
  assign p1_prod__879_comb = {{7{p1_concat_139606_comb[24]}}, p1_concat_139606_comb};
  assign p1_prod__884_comb = {{7{p1_concat_139607_comb[24]}}, p1_concat_139607_comb};
  assign p1_prod__891_comb = {{7{p1_concat_139608_comb[24]}}, p1_concat_139608_comb};
  assign p1_prod__930_comb = {{7{p1_concat_139609_comb[24]}}, p1_concat_139609_comb};
  assign p1_prod__943_comb = {{7{p1_concat_139610_comb[24]}}, p1_concat_139610_comb};
  assign p1_prod__948_comb = {{7{p1_concat_139611_comb[24]}}, p1_concat_139611_comb};
  assign p1_prod__955_comb = {{7{p1_concat_139612_comb[24]}}, p1_concat_139612_comb};
  assign p1_prod__994_comb = {{7{p1_concat_139613_comb[24]}}, p1_concat_139613_comb};
  assign p1_prod__1007_comb = {{7{p1_concat_139614_comb[24]}}, p1_concat_139614_comb};
  assign p1_prod__1012_comb = {{7{p1_concat_139615_comb[24]}}, p1_concat_139615_comb};
  assign p1_prod__1019_comb = {{7{p1_concat_139616_comb[24]}}, p1_concat_139616_comb};
  assign p1_prod__547_comb = {{9{p1_concat_139617_comb[22]}}, p1_concat_139617_comb};
  assign p1_prod__554_comb = {{7{p1_concat_139618_comb[24]}}, p1_concat_139618_comb};
  assign p1_prod__574_comb = {{7{p1_concat_139619_comb[24]}}, p1_concat_139619_comb};
  assign p1_prod__575_comb = {{9{p1_concat_139620_comb[22]}}, p1_concat_139620_comb};
  assign p1_prod__611_comb = {{9{p1_concat_139621_comb[22]}}, p1_concat_139621_comb};
  assign p1_prod__618_comb = {{7{p1_concat_139622_comb[24]}}, p1_concat_139622_comb};
  assign p1_prod__638_comb = {{7{p1_concat_139623_comb[24]}}, p1_concat_139623_comb};
  assign p1_prod__639_comb = {{9{p1_concat_139624_comb[22]}}, p1_concat_139624_comb};
  assign p1_prod__675_comb = {{9{p1_concat_139625_comb[22]}}, p1_concat_139625_comb};
  assign p1_prod__682_comb = {{7{p1_concat_139626_comb[24]}}, p1_concat_139626_comb};
  assign p1_prod__702_comb = {{7{p1_concat_139627_comb[24]}}, p1_concat_139627_comb};
  assign p1_prod__703_comb = {{9{p1_concat_139628_comb[22]}}, p1_concat_139628_comb};
  assign p1_prod__739_comb = {{9{p1_concat_139629_comb[22]}}, p1_concat_139629_comb};
  assign p1_prod__746_comb = {{7{p1_concat_139630_comb[24]}}, p1_concat_139630_comb};
  assign p1_prod__766_comb = {{7{p1_concat_139631_comb[24]}}, p1_concat_139631_comb};
  assign p1_prod__767_comb = {{9{p1_concat_139632_comb[22]}}, p1_concat_139632_comb};
  assign p1_prod__803_comb = {{9{p1_concat_139633_comb[22]}}, p1_concat_139633_comb};
  assign p1_prod__810_comb = {{7{p1_concat_139634_comb[24]}}, p1_concat_139634_comb};
  assign p1_prod__830_comb = {{7{p1_concat_139635_comb[24]}}, p1_concat_139635_comb};
  assign p1_prod__831_comb = {{9{p1_concat_139636_comb[22]}}, p1_concat_139636_comb};
  assign p1_prod__867_comb = {{9{p1_concat_139637_comb[22]}}, p1_concat_139637_comb};
  assign p1_prod__874_comb = {{7{p1_concat_139638_comb[24]}}, p1_concat_139638_comb};
  assign p1_prod__894_comb = {{7{p1_concat_139639_comb[24]}}, p1_concat_139639_comb};
  assign p1_prod__895_comb = {{9{p1_concat_139640_comb[22]}}, p1_concat_139640_comb};
  assign p1_prod__931_comb = {{9{p1_concat_139641_comb[22]}}, p1_concat_139641_comb};
  assign p1_prod__938_comb = {{7{p1_concat_139642_comb[24]}}, p1_concat_139642_comb};
  assign p1_prod__958_comb = {{7{p1_concat_139643_comb[24]}}, p1_concat_139643_comb};
  assign p1_prod__959_comb = {{9{p1_concat_139644_comb[22]}}, p1_concat_139644_comb};
  assign p1_prod__995_comb = {{9{p1_concat_139645_comb[22]}}, p1_concat_139645_comb};
  assign p1_prod__1002_comb = {{7{p1_concat_139646_comb[24]}}, p1_concat_139646_comb};
  assign p1_prod__1022_comb = {{7{p1_concat_139647_comb[24]}}, p1_concat_139647_comb};
  assign p1_prod__1023_comb = {{9{p1_concat_139648_comb[22]}}, p1_concat_139648_comb};
  assign p1_or_140545_comb = p1_prod__519_comb | 32'h0000_0080;
  assign p1_or_140546_comb = p1_prod__523_comb | 32'h0000_0080;
  assign p1_or_140547_comb = p1_prod__528_comb | 32'h0000_0080;
  assign p1_or_140548_comb = p1_prod__534_comb | 32'h0000_0080;
  assign p1_or_140549_comb = p1_prod__583_comb | 32'h0000_0080;
  assign p1_or_140550_comb = p1_prod__587_comb | 32'h0000_0080;
  assign p1_or_140551_comb = p1_prod__592_comb | 32'h0000_0080;
  assign p1_or_140552_comb = p1_prod__598_comb | 32'h0000_0080;
  assign p1_or_140553_comb = p1_prod__647_comb | 32'h0000_0080;
  assign p1_or_140554_comb = p1_prod__651_comb | 32'h0000_0080;
  assign p1_or_140555_comb = p1_prod__656_comb | 32'h0000_0080;
  assign p1_or_140556_comb = p1_prod__662_comb | 32'h0000_0080;
  assign p1_or_140557_comb = p1_prod__711_comb | 32'h0000_0080;
  assign p1_or_140558_comb = p1_prod__715_comb | 32'h0000_0080;
  assign p1_or_140559_comb = p1_prod__720_comb | 32'h0000_0080;
  assign p1_or_140560_comb = p1_prod__726_comb | 32'h0000_0080;
  assign p1_or_140561_comb = p1_prod__775_comb | 32'h0000_0080;
  assign p1_or_140562_comb = p1_prod__779_comb | 32'h0000_0080;
  assign p1_or_140563_comb = p1_prod__784_comb | 32'h0000_0080;
  assign p1_or_140564_comb = p1_prod__790_comb | 32'h0000_0080;
  assign p1_or_140565_comb = p1_prod__839_comb | 32'h0000_0080;
  assign p1_or_140566_comb = p1_prod__843_comb | 32'h0000_0080;
  assign p1_or_140567_comb = p1_prod__848_comb | 32'h0000_0080;
  assign p1_or_140568_comb = p1_prod__854_comb | 32'h0000_0080;
  assign p1_or_140569_comb = p1_prod__903_comb | 32'h0000_0080;
  assign p1_or_140570_comb = p1_prod__907_comb | 32'h0000_0080;
  assign p1_or_140571_comb = p1_prod__912_comb | 32'h0000_0080;
  assign p1_or_140572_comb = p1_prod__918_comb | 32'h0000_0080;
  assign p1_or_140573_comb = p1_prod__967_comb | 32'h0000_0080;
  assign p1_or_140574_comb = p1_prod__971_comb | 32'h0000_0080;
  assign p1_or_140575_comb = p1_prod__976_comb | 32'h0000_0080;
  assign p1_or_140576_comb = p1_prod__982_comb | 32'h0000_0080;
  assign p1_or_140577_comb = p1_prod__517_comb | 32'h0000_0080;
  assign p1_smul_58352_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__65_squeezed_comb, 7'h31);
  assign p1_smul_58354_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__66_squeezed_comb, 7'h4f);
  assign p1_or_140582_comb = p1_prod__529_comb | 32'h0000_0080;
  assign p1_or_140583_comb = p1_prod__535_comb | 32'h0000_0080;
  assign p1_smul_58360_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__69_squeezed_comb, 7'h4f);
  assign p1_smul_58362_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__70_squeezed_comb, 7'h31);
  assign p1_or_140588_comb = p1_prod__555_comb | 32'h0000_0080;
  assign p1_or_140589_comb = p1_prod__581_comb | 32'h0000_0080;
  assign p1_smul_58368_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__73_squeezed_comb, 7'h31);
  assign p1_smul_58370_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__74_squeezed_comb, 7'h4f);
  assign p1_or_140594_comb = p1_prod__593_comb | 32'h0000_0080;
  assign p1_or_140595_comb = p1_prod__599_comb | 32'h0000_0080;
  assign p1_smul_58376_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__77_squeezed_comb, 7'h4f);
  assign p1_smul_58378_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__78_squeezed_comb, 7'h31);
  assign p1_or_140600_comb = p1_prod__619_comb | 32'h0000_0080;
  assign p1_or_140601_comb = p1_prod__645_comb | 32'h0000_0080;
  assign p1_smul_58384_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__81_squeezed_comb, 7'h31);
  assign p1_smul_58386_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__82_squeezed_comb, 7'h4f);
  assign p1_or_140606_comb = p1_prod__657_comb | 32'h0000_0080;
  assign p1_or_140607_comb = p1_prod__663_comb | 32'h0000_0080;
  assign p1_smul_58392_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__85_squeezed_comb, 7'h4f);
  assign p1_smul_58394_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__86_squeezed_comb, 7'h31);
  assign p1_or_140612_comb = p1_prod__683_comb | 32'h0000_0080;
  assign p1_or_140613_comb = p1_prod__709_comb | 32'h0000_0080;
  assign p1_smul_58400_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__89_squeezed_comb, 7'h31);
  assign p1_smul_58402_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__90_squeezed_comb, 7'h4f);
  assign p1_or_140618_comb = p1_prod__721_comb | 32'h0000_0080;
  assign p1_or_140619_comb = p1_prod__727_comb | 32'h0000_0080;
  assign p1_smul_58408_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__93_squeezed_comb, 7'h4f);
  assign p1_smul_58410_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__94_squeezed_comb, 7'h31);
  assign p1_or_140624_comb = p1_prod__747_comb | 32'h0000_0080;
  assign p1_or_140625_comb = p1_prod__773_comb | 32'h0000_0080;
  assign p1_smul_58416_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__97_squeezed_comb, 7'h31);
  assign p1_smul_58418_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__98_squeezed_comb, 7'h4f);
  assign p1_or_140630_comb = p1_prod__785_comb | 32'h0000_0080;
  assign p1_or_140631_comb = p1_prod__791_comb | 32'h0000_0080;
  assign p1_smul_58424_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__101_squeezed_comb, 7'h4f);
  assign p1_smul_58426_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__102_squeezed_comb, 7'h31);
  assign p1_or_140636_comb = p1_prod__811_comb | 32'h0000_0080;
  assign p1_or_140637_comb = p1_prod__837_comb | 32'h0000_0080;
  assign p1_smul_58432_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__105_squeezed_comb, 7'h31);
  assign p1_smul_58434_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__106_squeezed_comb, 7'h4f);
  assign p1_or_140642_comb = p1_prod__849_comb | 32'h0000_0080;
  assign p1_or_140643_comb = p1_prod__855_comb | 32'h0000_0080;
  assign p1_smul_58440_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__109_squeezed_comb, 7'h4f);
  assign p1_smul_58442_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__110_squeezed_comb, 7'h31);
  assign p1_or_140648_comb = p1_prod__875_comb | 32'h0000_0080;
  assign p1_or_140649_comb = p1_prod__901_comb | 32'h0000_0080;
  assign p1_smul_58448_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__113_squeezed_comb, 7'h31);
  assign p1_smul_58450_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__114_squeezed_comb, 7'h4f);
  assign p1_or_140654_comb = p1_prod__913_comb | 32'h0000_0080;
  assign p1_or_140655_comb = p1_prod__919_comb | 32'h0000_0080;
  assign p1_smul_58456_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__117_squeezed_comb, 7'h4f);
  assign p1_smul_58458_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__118_squeezed_comb, 7'h31);
  assign p1_or_140660_comb = p1_prod__939_comb | 32'h0000_0080;
  assign p1_or_140661_comb = p1_prod__965_comb | 32'h0000_0080;
  assign p1_smul_58464_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__121_squeezed_comb, 7'h31);
  assign p1_smul_58466_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__122_squeezed_comb, 7'h4f);
  assign p1_or_140666_comb = p1_prod__977_comb | 32'h0000_0080;
  assign p1_or_140667_comb = p1_prod__983_comb | 32'h0000_0080;
  assign p1_smul_58472_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__125_squeezed_comb, 7'h4f);
  assign p1_smul_58474_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__126_squeezed_comb, 7'h31);
  assign p1_or_140672_comb = p1_prod__1003_comb | 32'h0000_0080;
  assign p1_or_140673_comb = p1_prod__525_comb | 32'h0000_0080;
  assign p1_or_140674_comb = p1_prod__536_comb | 32'h0000_0080;
  assign p1_or_140675_comb = p1_prod__543_comb | 32'h0000_0080;
  assign p1_or_140676_comb = p1_prod__556_comb | 32'h0000_0080;
  assign p1_or_140677_comb = p1_prod__589_comb | 32'h0000_0080;
  assign p1_or_140678_comb = p1_prod__600_comb | 32'h0000_0080;
  assign p1_or_140679_comb = p1_prod__607_comb | 32'h0000_0080;
  assign p1_or_140680_comb = p1_prod__620_comb | 32'h0000_0080;
  assign p1_or_140681_comb = p1_prod__653_comb | 32'h0000_0080;
  assign p1_or_140682_comb = p1_prod__664_comb | 32'h0000_0080;
  assign p1_or_140683_comb = p1_prod__671_comb | 32'h0000_0080;
  assign p1_or_140684_comb = p1_prod__684_comb | 32'h0000_0080;
  assign p1_or_140685_comb = p1_prod__717_comb | 32'h0000_0080;
  assign p1_or_140686_comb = p1_prod__728_comb | 32'h0000_0080;
  assign p1_or_140687_comb = p1_prod__735_comb | 32'h0000_0080;
  assign p1_or_140688_comb = p1_prod__748_comb | 32'h0000_0080;
  assign p1_or_140689_comb = p1_prod__781_comb | 32'h0000_0080;
  assign p1_or_140690_comb = p1_prod__792_comb | 32'h0000_0080;
  assign p1_or_140691_comb = p1_prod__799_comb | 32'h0000_0080;
  assign p1_or_140692_comb = p1_prod__812_comb | 32'h0000_0080;
  assign p1_or_140693_comb = p1_prod__845_comb | 32'h0000_0080;
  assign p1_or_140694_comb = p1_prod__856_comb | 32'h0000_0080;
  assign p1_or_140695_comb = p1_prod__863_comb | 32'h0000_0080;
  assign p1_or_140696_comb = p1_prod__876_comb | 32'h0000_0080;
  assign p1_or_140697_comb = p1_prod__909_comb | 32'h0000_0080;
  assign p1_or_140698_comb = p1_prod__920_comb | 32'h0000_0080;
  assign p1_or_140699_comb = p1_prod__927_comb | 32'h0000_0080;
  assign p1_or_140700_comb = p1_prod__940_comb | 32'h0000_0080;
  assign p1_or_140701_comb = p1_prod__973_comb | 32'h0000_0080;
  assign p1_or_140702_comb = p1_prod__984_comb | 32'h0000_0080;
  assign p1_or_140703_comb = p1_prod__991_comb | 32'h0000_0080;
  assign p1_or_140704_comb = p1_prod__1004_comb | 32'h0000_0080;
  assign p1_or_140705_comb = p1_prod__532_comb | 32'h0000_0080;
  assign p1_or_140706_comb = p1_prod__545_comb | 32'h0000_0080;
  assign p1_or_140707_comb = p1_prod__563_comb | 32'h0000_0080;
  assign p1_or_140708_comb = p1_prod__570_comb | 32'h0000_0080;
  assign p1_or_140709_comb = p1_prod__596_comb | 32'h0000_0080;
  assign p1_or_140710_comb = p1_prod__609_comb | 32'h0000_0080;
  assign p1_or_140711_comb = p1_prod__627_comb | 32'h0000_0080;
  assign p1_or_140712_comb = p1_prod__634_comb | 32'h0000_0080;
  assign p1_or_140713_comb = p1_prod__660_comb | 32'h0000_0080;
  assign p1_or_140714_comb = p1_prod__673_comb | 32'h0000_0080;
  assign p1_or_140715_comb = p1_prod__691_comb | 32'h0000_0080;
  assign p1_or_140716_comb = p1_prod__698_comb | 32'h0000_0080;
  assign p1_or_140717_comb = p1_prod__724_comb | 32'h0000_0080;
  assign p1_or_140718_comb = p1_prod__737_comb | 32'h0000_0080;
  assign p1_or_140719_comb = p1_prod__755_comb | 32'h0000_0080;
  assign p1_or_140720_comb = p1_prod__762_comb | 32'h0000_0080;
  assign p1_or_140721_comb = p1_prod__788_comb | 32'h0000_0080;
  assign p1_or_140722_comb = p1_prod__801_comb | 32'h0000_0080;
  assign p1_or_140723_comb = p1_prod__819_comb | 32'h0000_0080;
  assign p1_or_140724_comb = p1_prod__826_comb | 32'h0000_0080;
  assign p1_or_140725_comb = p1_prod__852_comb | 32'h0000_0080;
  assign p1_or_140726_comb = p1_prod__865_comb | 32'h0000_0080;
  assign p1_or_140727_comb = p1_prod__883_comb | 32'h0000_0080;
  assign p1_or_140728_comb = p1_prod__890_comb | 32'h0000_0080;
  assign p1_or_140729_comb = p1_prod__916_comb | 32'h0000_0080;
  assign p1_or_140730_comb = p1_prod__929_comb | 32'h0000_0080;
  assign p1_or_140731_comb = p1_prod__947_comb | 32'h0000_0080;
  assign p1_or_140732_comb = p1_prod__954_comb | 32'h0000_0080;
  assign p1_or_140733_comb = p1_prod__980_comb | 32'h0000_0080;
  assign p1_or_140734_comb = p1_prod__993_comb | 32'h0000_0080;
  assign p1_or_140735_comb = p1_prod__1011_comb | 32'h0000_0080;
  assign p1_or_140736_comb = p1_prod__1018_comb | 32'h0000_0080;
  assign p1_smul_58862_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__64_squeezed_comb, 7'h31);
  assign p1_or_140739_comb = p1_prod__546_comb | 32'h0000_0080;
  assign p1_smul_58866_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__66_squeezed_comb, 7'h31);
  assign p1_or_140742_comb = p1_prod__559_comb | 32'h0000_0080;
  assign p1_or_140743_comb = p1_prod__564_comb | 32'h0000_0080;
  assign p1_smul_58872_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__69_squeezed_comb, 7'h31);
  assign p1_or_140746_comb = p1_prod__571_comb | 32'h0000_0080;
  assign p1_smul_58876_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__71_squeezed_comb, 7'h31);
  assign p1_smul_58878_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__72_squeezed_comb, 7'h31);
  assign p1_or_140751_comb = p1_prod__610_comb | 32'h0000_0080;
  assign p1_smul_58882_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__74_squeezed_comb, 7'h31);
  assign p1_or_140754_comb = p1_prod__623_comb | 32'h0000_0080;
  assign p1_or_140755_comb = p1_prod__628_comb | 32'h0000_0080;
  assign p1_smul_58888_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__77_squeezed_comb, 7'h31);
  assign p1_or_140758_comb = p1_prod__635_comb | 32'h0000_0080;
  assign p1_smul_58892_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__79_squeezed_comb, 7'h31);
  assign p1_smul_58894_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__80_squeezed_comb, 7'h31);
  assign p1_or_140763_comb = p1_prod__674_comb | 32'h0000_0080;
  assign p1_smul_58898_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__82_squeezed_comb, 7'h31);
  assign p1_or_140766_comb = p1_prod__687_comb | 32'h0000_0080;
  assign p1_or_140767_comb = p1_prod__692_comb | 32'h0000_0080;
  assign p1_smul_58904_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__85_squeezed_comb, 7'h31);
  assign p1_or_140770_comb = p1_prod__699_comb | 32'h0000_0080;
  assign p1_smul_58908_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__87_squeezed_comb, 7'h31);
  assign p1_smul_58910_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__88_squeezed_comb, 7'h31);
  assign p1_or_140775_comb = p1_prod__738_comb | 32'h0000_0080;
  assign p1_smul_58914_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__90_squeezed_comb, 7'h31);
  assign p1_or_140778_comb = p1_prod__751_comb | 32'h0000_0080;
  assign p1_or_140779_comb = p1_prod__756_comb | 32'h0000_0080;
  assign p1_smul_58920_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__93_squeezed_comb, 7'h31);
  assign p1_or_140782_comb = p1_prod__763_comb | 32'h0000_0080;
  assign p1_smul_58924_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__95_squeezed_comb, 7'h31);
  assign p1_smul_58926_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__96_squeezed_comb, 7'h31);
  assign p1_or_140787_comb = p1_prod__802_comb | 32'h0000_0080;
  assign p1_smul_58930_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__98_squeezed_comb, 7'h31);
  assign p1_or_140790_comb = p1_prod__815_comb | 32'h0000_0080;
  assign p1_or_140791_comb = p1_prod__820_comb | 32'h0000_0080;
  assign p1_smul_58936_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__101_squeezed_comb, 7'h31);
  assign p1_or_140794_comb = p1_prod__827_comb | 32'h0000_0080;
  assign p1_smul_58940_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__103_squeezed_comb, 7'h31);
  assign p1_smul_58942_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__104_squeezed_comb, 7'h31);
  assign p1_or_140799_comb = p1_prod__866_comb | 32'h0000_0080;
  assign p1_smul_58946_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__106_squeezed_comb, 7'h31);
  assign p1_or_140802_comb = p1_prod__879_comb | 32'h0000_0080;
  assign p1_or_140803_comb = p1_prod__884_comb | 32'h0000_0080;
  assign p1_smul_58952_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__109_squeezed_comb, 7'h31);
  assign p1_or_140806_comb = p1_prod__891_comb | 32'h0000_0080;
  assign p1_smul_58956_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__111_squeezed_comb, 7'h31);
  assign p1_smul_58958_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__112_squeezed_comb, 7'h31);
  assign p1_or_140811_comb = p1_prod__930_comb | 32'h0000_0080;
  assign p1_smul_58962_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__114_squeezed_comb, 7'h31);
  assign p1_or_140814_comb = p1_prod__943_comb | 32'h0000_0080;
  assign p1_or_140815_comb = p1_prod__948_comb | 32'h0000_0080;
  assign p1_smul_58968_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__117_squeezed_comb, 7'h31);
  assign p1_or_140818_comb = p1_prod__955_comb | 32'h0000_0080;
  assign p1_smul_58972_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__119_squeezed_comb, 7'h31);
  assign p1_smul_58974_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__120_squeezed_comb, 7'h31);
  assign p1_or_140823_comb = p1_prod__994_comb | 32'h0000_0080;
  assign p1_smul_58978_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__122_squeezed_comb, 7'h31);
  assign p1_or_140826_comb = p1_prod__1007_comb | 32'h0000_0080;
  assign p1_or_140827_comb = p1_prod__1012_comb | 32'h0000_0080;
  assign p1_smul_58984_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__125_squeezed_comb, 7'h31);
  assign p1_or_140830_comb = p1_prod__1019_comb | 32'h0000_0080;
  assign p1_smul_58988_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__127_squeezed_comb, 7'h31);
  assign p1_or_140833_comb = p1_prod__547_comb | 32'h0000_0080;
  assign p1_or_140834_comb = p1_prod__554_comb | 32'h0000_0080;
  assign p1_or_140835_comb = p1_prod__574_comb | 32'h0000_0080;
  assign p1_or_140836_comb = p1_prod__575_comb | 32'h0000_0080;
  assign p1_or_140837_comb = p1_prod__611_comb | 32'h0000_0080;
  assign p1_or_140838_comb = p1_prod__618_comb | 32'h0000_0080;
  assign p1_or_140839_comb = p1_prod__638_comb | 32'h0000_0080;
  assign p1_or_140840_comb = p1_prod__639_comb | 32'h0000_0080;
  assign p1_or_140841_comb = p1_prod__675_comb | 32'h0000_0080;
  assign p1_or_140842_comb = p1_prod__682_comb | 32'h0000_0080;
  assign p1_or_140843_comb = p1_prod__702_comb | 32'h0000_0080;
  assign p1_or_140844_comb = p1_prod__703_comb | 32'h0000_0080;
  assign p1_or_140845_comb = p1_prod__739_comb | 32'h0000_0080;
  assign p1_or_140846_comb = p1_prod__746_comb | 32'h0000_0080;
  assign p1_or_140847_comb = p1_prod__766_comb | 32'h0000_0080;
  assign p1_or_140848_comb = p1_prod__767_comb | 32'h0000_0080;
  assign p1_or_140849_comb = p1_prod__803_comb | 32'h0000_0080;
  assign p1_or_140850_comb = p1_prod__810_comb | 32'h0000_0080;
  assign p1_or_140851_comb = p1_prod__830_comb | 32'h0000_0080;
  assign p1_or_140852_comb = p1_prod__831_comb | 32'h0000_0080;
  assign p1_or_140853_comb = p1_prod__867_comb | 32'h0000_0080;
  assign p1_or_140854_comb = p1_prod__874_comb | 32'h0000_0080;
  assign p1_or_140855_comb = p1_prod__894_comb | 32'h0000_0080;
  assign p1_or_140856_comb = p1_prod__895_comb | 32'h0000_0080;
  assign p1_or_140857_comb = p1_prod__931_comb | 32'h0000_0080;
  assign p1_or_140858_comb = p1_prod__938_comb | 32'h0000_0080;
  assign p1_or_140859_comb = p1_prod__958_comb | 32'h0000_0080;
  assign p1_or_140860_comb = p1_prod__959_comb | 32'h0000_0080;
  assign p1_or_140861_comb = p1_prod__995_comb | 32'h0000_0080;
  assign p1_or_140862_comb = p1_prod__1002_comb | 32'h0000_0080;
  assign p1_or_140863_comb = p1_prod__1022_comb | 32'h0000_0080;
  assign p1_or_140864_comb = p1_prod__1023_comb | 32'h0000_0080;
  assign p1_sel_140865_comb = $signed(p1_shifted__64_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__64_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__64_squeezed_comb, p1_smul_57326_TrailingBits___64_comb};
  assign p1_sel_140866_comb = $signed(p1_shifted__65_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__65_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__65_squeezed_comb, p1_smul_57326_TrailingBits___65_comb};
  assign p1_sel_140867_comb = $signed(p1_shifted__66_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__66_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__66_squeezed_comb, p1_smul_57326_TrailingBits___66_comb};
  assign p1_sel_140868_comb = $signed(p1_shifted__67_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__67_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__67_squeezed_comb, p1_smul_57326_TrailingBits___67_comb};
  assign p1_sel_140869_comb = $signed(p1_shifted__68_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__68_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__68_squeezed_comb, p1_smul_57326_TrailingBits___68_comb};
  assign p1_sel_140870_comb = $signed(p1_shifted__69_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__69_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__69_squeezed_comb, p1_smul_57326_TrailingBits___69_comb};
  assign p1_sel_140871_comb = $signed(p1_shifted__70_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__70_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__70_squeezed_comb, p1_smul_57326_TrailingBits___70_comb};
  assign p1_sel_140872_comb = $signed(p1_shifted__71_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__71_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__71_squeezed_comb, p1_smul_57326_TrailingBits___71_comb};
  assign p1_sel_140873_comb = $signed(p1_shifted__72_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__72_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__72_squeezed_comb, p1_smul_57326_TrailingBits___72_comb};
  assign p1_sel_140874_comb = $signed(p1_shifted__73_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__73_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__73_squeezed_comb, p1_smul_57326_TrailingBits___73_comb};
  assign p1_sel_140875_comb = $signed(p1_shifted__74_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__74_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__74_squeezed_comb, p1_smul_57326_TrailingBits___74_comb};
  assign p1_sel_140876_comb = $signed(p1_shifted__75_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__75_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__75_squeezed_comb, p1_smul_57326_TrailingBits___75_comb};
  assign p1_sel_140877_comb = $signed(p1_shifted__76_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__76_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__76_squeezed_comb, p1_smul_57326_TrailingBits___76_comb};
  assign p1_sel_140878_comb = $signed(p1_shifted__77_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__77_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__77_squeezed_comb, p1_smul_57326_TrailingBits___77_comb};
  assign p1_sel_140879_comb = $signed(p1_shifted__78_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__78_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__78_squeezed_comb, p1_smul_57326_TrailingBits___78_comb};
  assign p1_sel_140880_comb = $signed(p1_shifted__79_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__79_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__79_squeezed_comb, p1_smul_57326_TrailingBits___79_comb};
  assign p1_sel_140881_comb = $signed(p1_shifted__80_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__80_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__80_squeezed_comb, p1_smul_57326_TrailingBits___80_comb};
  assign p1_sel_140882_comb = $signed(p1_shifted__81_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__81_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__81_squeezed_comb, p1_smul_57326_TrailingBits___81_comb};
  assign p1_sel_140883_comb = $signed(p1_shifted__82_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__82_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__82_squeezed_comb, p1_smul_57326_TrailingBits___82_comb};
  assign p1_sel_140884_comb = $signed(p1_shifted__83_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__83_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__83_squeezed_comb, p1_smul_57326_TrailingBits___83_comb};
  assign p1_sel_140885_comb = $signed(p1_shifted__84_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__84_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__84_squeezed_comb, p1_smul_57326_TrailingBits___84_comb};
  assign p1_sel_140886_comb = $signed(p1_shifted__85_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__85_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__85_squeezed_comb, p1_smul_57326_TrailingBits___85_comb};
  assign p1_sel_140887_comb = $signed(p1_shifted__86_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__86_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__86_squeezed_comb, p1_smul_57326_TrailingBits___86_comb};
  assign p1_sel_140888_comb = $signed(p1_shifted__87_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__87_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__87_squeezed_comb, p1_smul_57326_TrailingBits___87_comb};
  assign p1_sel_140889_comb = $signed(p1_shifted__88_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__88_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__88_squeezed_comb, p1_smul_57326_TrailingBits___88_comb};
  assign p1_sel_140890_comb = $signed(p1_shifted__89_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__89_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__89_squeezed_comb, p1_smul_57326_TrailingBits___89_comb};
  assign p1_sel_140891_comb = $signed(p1_shifted__90_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__90_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__90_squeezed_comb, p1_smul_57326_TrailingBits___90_comb};
  assign p1_sel_140892_comb = $signed(p1_shifted__91_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__91_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__91_squeezed_comb, p1_smul_57326_TrailingBits___91_comb};
  assign p1_sel_140893_comb = $signed(p1_shifted__92_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__92_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__92_squeezed_comb, p1_smul_57326_TrailingBits___92_comb};
  assign p1_sel_140894_comb = $signed(p1_shifted__93_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__93_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__93_squeezed_comb, p1_smul_57326_TrailingBits___93_comb};
  assign p1_sel_140895_comb = $signed(p1_shifted__94_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__94_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__94_squeezed_comb, p1_smul_57326_TrailingBits___94_comb};
  assign p1_sel_140896_comb = $signed(p1_shifted__95_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__95_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__95_squeezed_comb, p1_smul_57326_TrailingBits___95_comb};
  assign p1_sel_140897_comb = $signed(p1_shifted__96_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__96_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__96_squeezed_comb, p1_smul_57326_TrailingBits___96_comb};
  assign p1_sel_140898_comb = $signed(p1_shifted__97_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__97_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__97_squeezed_comb, p1_smul_57326_TrailingBits___97_comb};
  assign p1_sel_140899_comb = $signed(p1_shifted__98_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__98_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__98_squeezed_comb, p1_smul_57326_TrailingBits___98_comb};
  assign p1_sel_140900_comb = $signed(p1_shifted__99_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__99_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__99_squeezed_comb, p1_smul_57326_TrailingBits___99_comb};
  assign p1_sel_140901_comb = $signed(p1_shifted__100_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__100_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__100_squeezed_comb, p1_smul_57326_TrailingBits___100_comb};
  assign p1_sel_140902_comb = $signed(p1_shifted__101_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__101_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__101_squeezed_comb, p1_smul_57326_TrailingBits___101_comb};
  assign p1_sel_140903_comb = $signed(p1_shifted__102_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__102_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__102_squeezed_comb, p1_smul_57326_TrailingBits___102_comb};
  assign p1_sel_140904_comb = $signed(p1_shifted__103_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__103_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__103_squeezed_comb, p1_smul_57326_TrailingBits___103_comb};
  assign p1_sel_140905_comb = $signed(p1_shifted__104_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__104_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__104_squeezed_comb, p1_smul_57326_TrailingBits___104_comb};
  assign p1_sel_140906_comb = $signed(p1_shifted__105_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__105_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__105_squeezed_comb, p1_smul_57326_TrailingBits___105_comb};
  assign p1_sel_140907_comb = $signed(p1_shifted__106_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__106_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__106_squeezed_comb, p1_smul_57326_TrailingBits___106_comb};
  assign p1_sel_140908_comb = $signed(p1_shifted__107_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__107_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__107_squeezed_comb, p1_smul_57326_TrailingBits___107_comb};
  assign p1_sel_140909_comb = $signed(p1_shifted__108_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__108_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__108_squeezed_comb, p1_smul_57326_TrailingBits___108_comb};
  assign p1_sel_140910_comb = $signed(p1_shifted__109_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__109_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__109_squeezed_comb, p1_smul_57326_TrailingBits___109_comb};
  assign p1_sel_140911_comb = $signed(p1_shifted__110_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__110_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__110_squeezed_comb, p1_smul_57326_TrailingBits___110_comb};
  assign p1_sel_140912_comb = $signed(p1_shifted__111_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__111_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__111_squeezed_comb, p1_smul_57326_TrailingBits___111_comb};
  assign p1_sel_140913_comb = $signed(p1_shifted__112_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__112_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__112_squeezed_comb, p1_smul_57326_TrailingBits___112_comb};
  assign p1_sel_140914_comb = $signed(p1_shifted__113_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__113_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__113_squeezed_comb, p1_smul_57326_TrailingBits___113_comb};
  assign p1_sel_140915_comb = $signed(p1_shifted__114_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__114_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__114_squeezed_comb, p1_smul_57326_TrailingBits___114_comb};
  assign p1_sel_140916_comb = $signed(p1_shifted__115_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__115_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__115_squeezed_comb, p1_smul_57326_TrailingBits___115_comb};
  assign p1_sel_140917_comb = $signed(p1_shifted__116_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__116_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__116_squeezed_comb, p1_smul_57326_TrailingBits___116_comb};
  assign p1_sel_140918_comb = $signed(p1_shifted__117_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__117_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__117_squeezed_comb, p1_smul_57326_TrailingBits___117_comb};
  assign p1_sel_140919_comb = $signed(p1_shifted__118_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__118_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__118_squeezed_comb, p1_smul_57326_TrailingBits___118_comb};
  assign p1_sel_140920_comb = $signed(p1_shifted__119_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__119_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__119_squeezed_comb, p1_smul_57326_TrailingBits___119_comb};
  assign p1_sel_140921_comb = $signed(p1_shifted__120_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__120_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__120_squeezed_comb, p1_smul_57326_TrailingBits___120_comb};
  assign p1_sel_140922_comb = $signed(p1_shifted__121_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__121_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__121_squeezed_comb, p1_smul_57326_TrailingBits___121_comb};
  assign p1_sel_140923_comb = $signed(p1_shifted__122_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__122_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__122_squeezed_comb, p1_smul_57326_TrailingBits___122_comb};
  assign p1_sel_140924_comb = $signed(p1_shifted__123_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__123_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__123_squeezed_comb, p1_smul_57326_TrailingBits___123_comb};
  assign p1_sel_140925_comb = $signed(p1_shifted__124_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__124_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__124_squeezed_comb, p1_smul_57326_TrailingBits___124_comb};
  assign p1_sel_140926_comb = $signed(p1_shifted__125_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__125_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__125_squeezed_comb, p1_smul_57326_TrailingBits___125_comb};
  assign p1_sel_140927_comb = $signed(p1_shifted__126_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__126_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__126_squeezed_comb, p1_smul_57326_TrailingBits___126_comb};
  assign p1_sel_140928_comb = $signed(p1_shifted__127_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__127_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__127_squeezed_comb, p1_smul_57326_TrailingBits___127_comb};
  assign p1_concat_141061_comb = {p1_smul_58352_NarrowedMult__comb, 1'h0};
  assign p1_concat_141063_comb = {p1_smul_58354_NarrowedMult__comb, 1'h0};
  assign p1_concat_141073_comb = {p1_smul_58360_NarrowedMult__comb, 1'h0};
  assign p1_concat_141075_comb = {p1_smul_58362_NarrowedMult__comb, 1'h0};
  assign p1_concat_141085_comb = {p1_smul_58368_NarrowedMult__comb, 1'h0};
  assign p1_concat_141087_comb = {p1_smul_58370_NarrowedMult__comb, 1'h0};
  assign p1_concat_141097_comb = {p1_smul_58376_NarrowedMult__comb, 1'h0};
  assign p1_concat_141099_comb = {p1_smul_58378_NarrowedMult__comb, 1'h0};
  assign p1_concat_141109_comb = {p1_smul_58384_NarrowedMult__comb, 1'h0};
  assign p1_concat_141111_comb = {p1_smul_58386_NarrowedMult__comb, 1'h0};
  assign p1_concat_141121_comb = {p1_smul_58392_NarrowedMult__comb, 1'h0};
  assign p1_concat_141123_comb = {p1_smul_58394_NarrowedMult__comb, 1'h0};
  assign p1_concat_141133_comb = {p1_smul_58400_NarrowedMult__comb, 1'h0};
  assign p1_concat_141135_comb = {p1_smul_58402_NarrowedMult__comb, 1'h0};
  assign p1_concat_141145_comb = {p1_smul_58408_NarrowedMult__comb, 1'h0};
  assign p1_concat_141147_comb = {p1_smul_58410_NarrowedMult__comb, 1'h0};
  assign p1_concat_141157_comb = {p1_smul_58416_NarrowedMult__comb, 1'h0};
  assign p1_concat_141159_comb = {p1_smul_58418_NarrowedMult__comb, 1'h0};
  assign p1_concat_141169_comb = {p1_smul_58424_NarrowedMult__comb, 1'h0};
  assign p1_concat_141171_comb = {p1_smul_58426_NarrowedMult__comb, 1'h0};
  assign p1_concat_141181_comb = {p1_smul_58432_NarrowedMult__comb, 1'h0};
  assign p1_concat_141183_comb = {p1_smul_58434_NarrowedMult__comb, 1'h0};
  assign p1_concat_141193_comb = {p1_smul_58440_NarrowedMult__comb, 1'h0};
  assign p1_concat_141195_comb = {p1_smul_58442_NarrowedMult__comb, 1'h0};
  assign p1_concat_141205_comb = {p1_smul_58448_NarrowedMult__comb, 1'h0};
  assign p1_concat_141207_comb = {p1_smul_58450_NarrowedMult__comb, 1'h0};
  assign p1_concat_141217_comb = {p1_smul_58456_NarrowedMult__comb, 1'h0};
  assign p1_concat_141219_comb = {p1_smul_58458_NarrowedMult__comb, 1'h0};
  assign p1_concat_141229_comb = {p1_smul_58464_NarrowedMult__comb, 1'h0};
  assign p1_concat_141231_comb = {p1_smul_58466_NarrowedMult__comb, 1'h0};
  assign p1_concat_141241_comb = {p1_smul_58472_NarrowedMult__comb, 1'h0};
  assign p1_concat_141243_comb = {p1_smul_58474_NarrowedMult__comb, 1'h0};
  assign p1_concat_141505_comb = {p1_smul_58862_NarrowedMult__comb, 1'h0};
  assign p1_concat_141511_comb = {p1_smul_58866_NarrowedMult__comb, 1'h0};
  assign p1_concat_141521_comb = {p1_smul_58872_NarrowedMult__comb, 1'h0};
  assign p1_concat_141527_comb = {p1_smul_58876_NarrowedMult__comb, 1'h0};
  assign p1_concat_141529_comb = {p1_smul_58878_NarrowedMult__comb, 1'h0};
  assign p1_concat_141535_comb = {p1_smul_58882_NarrowedMult__comb, 1'h0};
  assign p1_concat_141545_comb = {p1_smul_58888_NarrowedMult__comb, 1'h0};
  assign p1_concat_141551_comb = {p1_smul_58892_NarrowedMult__comb, 1'h0};
  assign p1_concat_141553_comb = {p1_smul_58894_NarrowedMult__comb, 1'h0};
  assign p1_concat_141559_comb = {p1_smul_58898_NarrowedMult__comb, 1'h0};
  assign p1_concat_141569_comb = {p1_smul_58904_NarrowedMult__comb, 1'h0};
  assign p1_concat_141575_comb = {p1_smul_58908_NarrowedMult__comb, 1'h0};
  assign p1_concat_141577_comb = {p1_smul_58910_NarrowedMult__comb, 1'h0};
  assign p1_concat_141583_comb = {p1_smul_58914_NarrowedMult__comb, 1'h0};
  assign p1_concat_141593_comb = {p1_smul_58920_NarrowedMult__comb, 1'h0};
  assign p1_concat_141599_comb = {p1_smul_58924_NarrowedMult__comb, 1'h0};
  assign p1_concat_141601_comb = {p1_smul_58926_NarrowedMult__comb, 1'h0};
  assign p1_concat_141607_comb = {p1_smul_58930_NarrowedMult__comb, 1'h0};
  assign p1_concat_141617_comb = {p1_smul_58936_NarrowedMult__comb, 1'h0};
  assign p1_concat_141623_comb = {p1_smul_58940_NarrowedMult__comb, 1'h0};
  assign p1_concat_141625_comb = {p1_smul_58942_NarrowedMult__comb, 1'h0};
  assign p1_concat_141631_comb = {p1_smul_58946_NarrowedMult__comb, 1'h0};
  assign p1_concat_141641_comb = {p1_smul_58952_NarrowedMult__comb, 1'h0};
  assign p1_concat_141647_comb = {p1_smul_58956_NarrowedMult__comb, 1'h0};
  assign p1_concat_141649_comb = {p1_smul_58958_NarrowedMult__comb, 1'h0};
  assign p1_concat_141655_comb = {p1_smul_58962_NarrowedMult__comb, 1'h0};
  assign p1_concat_141665_comb = {p1_smul_58968_NarrowedMult__comb, 1'h0};
  assign p1_concat_141671_comb = {p1_smul_58972_NarrowedMult__comb, 1'h0};
  assign p1_concat_141673_comb = {p1_smul_58974_NarrowedMult__comb, 1'h0};
  assign p1_concat_141679_comb = {p1_smul_58978_NarrowedMult__comb, 1'h0};
  assign p1_concat_141689_comb = {p1_smul_58984_NarrowedMult__comb, 1'h0};
  assign p1_concat_141695_comb = {p1_smul_58988_NarrowedMult__comb, 1'h0};
  assign p1_add_142785_comb = {{1{p1_sel_140865_comb[15]}}, p1_sel_140865_comb} + {{1{p1_sel_140866_comb[15]}}, p1_sel_140866_comb};
  assign p1_add_142786_comb = {{1{p1_sel_140867_comb[15]}}, p1_sel_140867_comb} + {{1{p1_sel_140868_comb[15]}}, p1_sel_140868_comb};
  assign p1_add_142787_comb = {{1{p1_sel_140869_comb[15]}}, p1_sel_140869_comb} + {{1{p1_sel_140870_comb[15]}}, p1_sel_140870_comb};
  assign p1_add_142788_comb = {{1{p1_sel_140871_comb[15]}}, p1_sel_140871_comb} + {{1{p1_sel_140872_comb[15]}}, p1_sel_140872_comb};
  assign p1_add_142789_comb = {{1{p1_sel_140873_comb[15]}}, p1_sel_140873_comb} + {{1{p1_sel_140874_comb[15]}}, p1_sel_140874_comb};
  assign p1_add_142790_comb = {{1{p1_sel_140875_comb[15]}}, p1_sel_140875_comb} + {{1{p1_sel_140876_comb[15]}}, p1_sel_140876_comb};
  assign p1_add_142791_comb = {{1{p1_sel_140877_comb[15]}}, p1_sel_140877_comb} + {{1{p1_sel_140878_comb[15]}}, p1_sel_140878_comb};
  assign p1_add_142792_comb = {{1{p1_sel_140879_comb[15]}}, p1_sel_140879_comb} + {{1{p1_sel_140880_comb[15]}}, p1_sel_140880_comb};
  assign p1_add_142793_comb = {{1{p1_sel_140881_comb[15]}}, p1_sel_140881_comb} + {{1{p1_sel_140882_comb[15]}}, p1_sel_140882_comb};
  assign p1_add_142794_comb = {{1{p1_sel_140883_comb[15]}}, p1_sel_140883_comb} + {{1{p1_sel_140884_comb[15]}}, p1_sel_140884_comb};
  assign p1_add_142795_comb = {{1{p1_sel_140885_comb[15]}}, p1_sel_140885_comb} + {{1{p1_sel_140886_comb[15]}}, p1_sel_140886_comb};
  assign p1_add_142796_comb = {{1{p1_sel_140887_comb[15]}}, p1_sel_140887_comb} + {{1{p1_sel_140888_comb[15]}}, p1_sel_140888_comb};
  assign p1_add_142797_comb = {{1{p1_sel_140889_comb[15]}}, p1_sel_140889_comb} + {{1{p1_sel_140890_comb[15]}}, p1_sel_140890_comb};
  assign p1_add_142798_comb = {{1{p1_sel_140891_comb[15]}}, p1_sel_140891_comb} + {{1{p1_sel_140892_comb[15]}}, p1_sel_140892_comb};
  assign p1_add_142799_comb = {{1{p1_sel_140893_comb[15]}}, p1_sel_140893_comb} + {{1{p1_sel_140894_comb[15]}}, p1_sel_140894_comb};
  assign p1_add_142800_comb = {{1{p1_sel_140895_comb[15]}}, p1_sel_140895_comb} + {{1{p1_sel_140896_comb[15]}}, p1_sel_140896_comb};
  assign p1_add_142801_comb = {{1{p1_sel_140897_comb[15]}}, p1_sel_140897_comb} + {{1{p1_sel_140898_comb[15]}}, p1_sel_140898_comb};
  assign p1_add_142802_comb = {{1{p1_sel_140899_comb[15]}}, p1_sel_140899_comb} + {{1{p1_sel_140900_comb[15]}}, p1_sel_140900_comb};
  assign p1_add_142803_comb = {{1{p1_sel_140901_comb[15]}}, p1_sel_140901_comb} + {{1{p1_sel_140902_comb[15]}}, p1_sel_140902_comb};
  assign p1_add_142804_comb = {{1{p1_sel_140903_comb[15]}}, p1_sel_140903_comb} + {{1{p1_sel_140904_comb[15]}}, p1_sel_140904_comb};
  assign p1_add_142805_comb = {{1{p1_sel_140905_comb[15]}}, p1_sel_140905_comb} + {{1{p1_sel_140906_comb[15]}}, p1_sel_140906_comb};
  assign p1_add_142806_comb = {{1{p1_sel_140907_comb[15]}}, p1_sel_140907_comb} + {{1{p1_sel_140908_comb[15]}}, p1_sel_140908_comb};
  assign p1_add_142807_comb = {{1{p1_sel_140909_comb[15]}}, p1_sel_140909_comb} + {{1{p1_sel_140910_comb[15]}}, p1_sel_140910_comb};
  assign p1_add_142808_comb = {{1{p1_sel_140911_comb[15]}}, p1_sel_140911_comb} + {{1{p1_sel_140912_comb[15]}}, p1_sel_140912_comb};
  assign p1_add_142809_comb = {{1{p1_sel_140913_comb[15]}}, p1_sel_140913_comb} + {{1{p1_sel_140914_comb[15]}}, p1_sel_140914_comb};
  assign p1_add_142810_comb = {{1{p1_sel_140915_comb[15]}}, p1_sel_140915_comb} + {{1{p1_sel_140916_comb[15]}}, p1_sel_140916_comb};
  assign p1_add_142811_comb = {{1{p1_sel_140917_comb[15]}}, p1_sel_140917_comb} + {{1{p1_sel_140918_comb[15]}}, p1_sel_140918_comb};
  assign p1_add_142812_comb = {{1{p1_sel_140919_comb[15]}}, p1_sel_140919_comb} + {{1{p1_sel_140920_comb[15]}}, p1_sel_140920_comb};
  assign p1_add_142813_comb = {{1{p1_sel_140921_comb[15]}}, p1_sel_140921_comb} + {{1{p1_sel_140922_comb[15]}}, p1_sel_140922_comb};
  assign p1_add_142814_comb = {{1{p1_sel_140923_comb[15]}}, p1_sel_140923_comb} + {{1{p1_sel_140924_comb[15]}}, p1_sel_140924_comb};
  assign p1_add_142815_comb = {{1{p1_sel_140925_comb[15]}}, p1_sel_140925_comb} + {{1{p1_sel_140926_comb[15]}}, p1_sel_140926_comb};
  assign p1_add_142816_comb = {{1{p1_sel_140927_comb[15]}}, p1_sel_140927_comb} + {{1{p1_sel_140928_comb[15]}}, p1_sel_140928_comb};
  assign p1_smul_142817_comb = smul16b_8b_x_9b(p1_shifted__64_squeezed_comb, 9'h0fb);
  assign p1_smul_142818_comb = smul16b_8b_x_9b(p1_shifted__65_squeezed_comb, 9'h0d5);
  assign p1_sel_142819_comb = $signed(p1_or_140545_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140545_comb[23:9], 1'h0};
  assign p1_sel_142820_comb = $signed(p1_or_140546_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140546_comb[23:9], 1'h0};
  assign p1_sel_142821_comb = $signed(p1_or_140547_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140547_comb[23:9], 1'h0};
  assign p1_sel_142822_comb = $signed(p1_or_140548_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140548_comb[23:9], 1'h0};
  assign p1_smul_142823_comb = smul16b_8b_x_9b(p1_shifted__70_squeezed_comb, 9'h12b);
  assign p1_smul_142824_comb = smul16b_8b_x_9b(p1_shifted__71_squeezed_comb, 9'h105);
  assign p1_smul_142825_comb = smul16b_8b_x_9b(p1_shifted__72_squeezed_comb, 9'h0fb);
  assign p1_smul_142826_comb = smul16b_8b_x_9b(p1_shifted__73_squeezed_comb, 9'h0d5);
  assign p1_sel_142827_comb = $signed(p1_or_140549_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140549_comb[23:9], 1'h0};
  assign p1_sel_142828_comb = $signed(p1_or_140550_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140550_comb[23:9], 1'h0};
  assign p1_sel_142829_comb = $signed(p1_or_140551_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140551_comb[23:9], 1'h0};
  assign p1_sel_142830_comb = $signed(p1_or_140552_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140552_comb[23:9], 1'h0};
  assign p1_smul_142831_comb = smul16b_8b_x_9b(p1_shifted__78_squeezed_comb, 9'h12b);
  assign p1_smul_142832_comb = smul16b_8b_x_9b(p1_shifted__79_squeezed_comb, 9'h105);
  assign p1_smul_142833_comb = smul16b_8b_x_9b(p1_shifted__80_squeezed_comb, 9'h0fb);
  assign p1_smul_142834_comb = smul16b_8b_x_9b(p1_shifted__81_squeezed_comb, 9'h0d5);
  assign p1_sel_142835_comb = $signed(p1_or_140553_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140553_comb[23:9], 1'h0};
  assign p1_sel_142836_comb = $signed(p1_or_140554_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140554_comb[23:9], 1'h0};
  assign p1_sel_142837_comb = $signed(p1_or_140555_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140555_comb[23:9], 1'h0};
  assign p1_sel_142838_comb = $signed(p1_or_140556_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140556_comb[23:9], 1'h0};
  assign p1_smul_142839_comb = smul16b_8b_x_9b(p1_shifted__86_squeezed_comb, 9'h12b);
  assign p1_smul_142840_comb = smul16b_8b_x_9b(p1_shifted__87_squeezed_comb, 9'h105);
  assign p1_smul_142841_comb = smul16b_8b_x_9b(p1_shifted__88_squeezed_comb, 9'h0fb);
  assign p1_smul_142842_comb = smul16b_8b_x_9b(p1_shifted__89_squeezed_comb, 9'h0d5);
  assign p1_sel_142843_comb = $signed(p1_or_140557_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140557_comb[23:9], 1'h0};
  assign p1_sel_142844_comb = $signed(p1_or_140558_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140558_comb[23:9], 1'h0};
  assign p1_sel_142845_comb = $signed(p1_or_140559_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140559_comb[23:9], 1'h0};
  assign p1_sel_142846_comb = $signed(p1_or_140560_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140560_comb[23:9], 1'h0};
  assign p1_smul_142847_comb = smul16b_8b_x_9b(p1_shifted__94_squeezed_comb, 9'h12b);
  assign p1_smul_142848_comb = smul16b_8b_x_9b(p1_shifted__95_squeezed_comb, 9'h105);
  assign p1_smul_142849_comb = smul16b_8b_x_9b(p1_shifted__96_squeezed_comb, 9'h0fb);
  assign p1_smul_142850_comb = smul16b_8b_x_9b(p1_shifted__97_squeezed_comb, 9'h0d5);
  assign p1_sel_142851_comb = $signed(p1_or_140561_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140561_comb[23:9], 1'h0};
  assign p1_sel_142852_comb = $signed(p1_or_140562_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140562_comb[23:9], 1'h0};
  assign p1_sel_142853_comb = $signed(p1_or_140563_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140563_comb[23:9], 1'h0};
  assign p1_sel_142854_comb = $signed(p1_or_140564_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140564_comb[23:9], 1'h0};
  assign p1_smul_142855_comb = smul16b_8b_x_9b(p1_shifted__102_squeezed_comb, 9'h12b);
  assign p1_smul_142856_comb = smul16b_8b_x_9b(p1_shifted__103_squeezed_comb, 9'h105);
  assign p1_smul_142857_comb = smul16b_8b_x_9b(p1_shifted__104_squeezed_comb, 9'h0fb);
  assign p1_smul_142858_comb = smul16b_8b_x_9b(p1_shifted__105_squeezed_comb, 9'h0d5);
  assign p1_sel_142859_comb = $signed(p1_or_140565_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140565_comb[23:9], 1'h0};
  assign p1_sel_142860_comb = $signed(p1_or_140566_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140566_comb[23:9], 1'h0};
  assign p1_sel_142861_comb = $signed(p1_or_140567_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140567_comb[23:9], 1'h0};
  assign p1_sel_142862_comb = $signed(p1_or_140568_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140568_comb[23:9], 1'h0};
  assign p1_smul_142863_comb = smul16b_8b_x_9b(p1_shifted__110_squeezed_comb, 9'h12b);
  assign p1_smul_142864_comb = smul16b_8b_x_9b(p1_shifted__111_squeezed_comb, 9'h105);
  assign p1_smul_142865_comb = smul16b_8b_x_9b(p1_shifted__112_squeezed_comb, 9'h0fb);
  assign p1_smul_142866_comb = smul16b_8b_x_9b(p1_shifted__113_squeezed_comb, 9'h0d5);
  assign p1_sel_142867_comb = $signed(p1_or_140569_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140569_comb[23:9], 1'h0};
  assign p1_sel_142868_comb = $signed(p1_or_140570_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140570_comb[23:9], 1'h0};
  assign p1_sel_142869_comb = $signed(p1_or_140571_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140571_comb[23:9], 1'h0};
  assign p1_sel_142870_comb = $signed(p1_or_140572_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140572_comb[23:9], 1'h0};
  assign p1_smul_142871_comb = smul16b_8b_x_9b(p1_shifted__118_squeezed_comb, 9'h12b);
  assign p1_smul_142872_comb = smul16b_8b_x_9b(p1_shifted__119_squeezed_comb, 9'h105);
  assign p1_smul_142873_comb = smul16b_8b_x_9b(p1_shifted__120_squeezed_comb, 9'h0fb);
  assign p1_smul_142874_comb = smul16b_8b_x_9b(p1_shifted__121_squeezed_comb, 9'h0d5);
  assign p1_sel_142875_comb = $signed(p1_or_140573_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140573_comb[23:9], 1'h0};
  assign p1_sel_142876_comb = $signed(p1_or_140574_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140574_comb[23:9], 1'h0};
  assign p1_sel_142877_comb = $signed(p1_or_140575_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140575_comb[23:9], 1'h0};
  assign p1_sel_142878_comb = $signed(p1_or_140576_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140576_comb[23:9], 1'h0};
  assign p1_smul_142879_comb = smul16b_8b_x_9b(p1_shifted__126_squeezed_comb, 9'h12b);
  assign p1_smul_142880_comb = smul16b_8b_x_9b(p1_shifted__127_squeezed_comb, 9'h105);
  assign p1_sel_142881_comb = $signed(p1_or_140577_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140577_comb[23:10], 2'h0};
  assign p1_sel_142882_comb = $signed(p1_concat_141061_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141061_comb;
  assign p1_sel_142883_comb = $signed(p1_concat_141063_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141063_comb;
  assign p1_sel_142884_comb = $signed(p1_or_140582_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140582_comb[23:10], 2'h0};
  assign p1_sel_142885_comb = $signed(p1_or_140583_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140583_comb[23:10], 2'h0};
  assign p1_sel_142886_comb = $signed(p1_concat_141073_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141073_comb;
  assign p1_sel_142887_comb = $signed(p1_concat_141075_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141075_comb;
  assign p1_sel_142888_comb = $signed(p1_or_140588_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140588_comb[23:10], 2'h0};
  assign p1_sel_142889_comb = $signed(p1_or_140589_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140589_comb[23:10], 2'h0};
  assign p1_sel_142890_comb = $signed(p1_concat_141085_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141085_comb;
  assign p1_sel_142891_comb = $signed(p1_concat_141087_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141087_comb;
  assign p1_sel_142892_comb = $signed(p1_or_140594_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140594_comb[23:10], 2'h0};
  assign p1_sel_142893_comb = $signed(p1_or_140595_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140595_comb[23:10], 2'h0};
  assign p1_sel_142894_comb = $signed(p1_concat_141097_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141097_comb;
  assign p1_sel_142895_comb = $signed(p1_concat_141099_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141099_comb;
  assign p1_sel_142896_comb = $signed(p1_or_140600_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140600_comb[23:10], 2'h0};
  assign p1_sel_142897_comb = $signed(p1_or_140601_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140601_comb[23:10], 2'h0};
  assign p1_sel_142898_comb = $signed(p1_concat_141109_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141109_comb;
  assign p1_sel_142899_comb = $signed(p1_concat_141111_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141111_comb;
  assign p1_sel_142900_comb = $signed(p1_or_140606_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140606_comb[23:10], 2'h0};
  assign p1_sel_142901_comb = $signed(p1_or_140607_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140607_comb[23:10], 2'h0};
  assign p1_sel_142902_comb = $signed(p1_concat_141121_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141121_comb;
  assign p1_sel_142903_comb = $signed(p1_concat_141123_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141123_comb;
  assign p1_sel_142904_comb = $signed(p1_or_140612_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140612_comb[23:10], 2'h0};
  assign p1_sel_142905_comb = $signed(p1_or_140613_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140613_comb[23:10], 2'h0};
  assign p1_sel_142906_comb = $signed(p1_concat_141133_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141133_comb;
  assign p1_sel_142907_comb = $signed(p1_concat_141135_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141135_comb;
  assign p1_sel_142908_comb = $signed(p1_or_140618_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140618_comb[23:10], 2'h0};
  assign p1_sel_142909_comb = $signed(p1_or_140619_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140619_comb[23:10], 2'h0};
  assign p1_sel_142910_comb = $signed(p1_concat_141145_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141145_comb;
  assign p1_sel_142911_comb = $signed(p1_concat_141147_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141147_comb;
  assign p1_sel_142912_comb = $signed(p1_or_140624_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140624_comb[23:10], 2'h0};
  assign p1_sel_142913_comb = $signed(p1_or_140625_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140625_comb[23:10], 2'h0};
  assign p1_sel_142914_comb = $signed(p1_concat_141157_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141157_comb;
  assign p1_sel_142915_comb = $signed(p1_concat_141159_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141159_comb;
  assign p1_sel_142916_comb = $signed(p1_or_140630_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140630_comb[23:10], 2'h0};
  assign p1_sel_142917_comb = $signed(p1_or_140631_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140631_comb[23:10], 2'h0};
  assign p1_sel_142918_comb = $signed(p1_concat_141169_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141169_comb;
  assign p1_sel_142919_comb = $signed(p1_concat_141171_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141171_comb;
  assign p1_sel_142920_comb = $signed(p1_or_140636_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140636_comb[23:10], 2'h0};
  assign p1_sel_142921_comb = $signed(p1_or_140637_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140637_comb[23:10], 2'h0};
  assign p1_sel_142922_comb = $signed(p1_concat_141181_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141181_comb;
  assign p1_sel_142923_comb = $signed(p1_concat_141183_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141183_comb;
  assign p1_sel_142924_comb = $signed(p1_or_140642_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140642_comb[23:10], 2'h0};
  assign p1_sel_142925_comb = $signed(p1_or_140643_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140643_comb[23:10], 2'h0};
  assign p1_sel_142926_comb = $signed(p1_concat_141193_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141193_comb;
  assign p1_sel_142927_comb = $signed(p1_concat_141195_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141195_comb;
  assign p1_sel_142928_comb = $signed(p1_or_140648_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140648_comb[23:10], 2'h0};
  assign p1_sel_142929_comb = $signed(p1_or_140649_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140649_comb[23:10], 2'h0};
  assign p1_sel_142930_comb = $signed(p1_concat_141205_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141205_comb;
  assign p1_sel_142931_comb = $signed(p1_concat_141207_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141207_comb;
  assign p1_sel_142932_comb = $signed(p1_or_140654_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140654_comb[23:10], 2'h0};
  assign p1_sel_142933_comb = $signed(p1_or_140655_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140655_comb[23:10], 2'h0};
  assign p1_sel_142934_comb = $signed(p1_concat_141217_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141217_comb;
  assign p1_sel_142935_comb = $signed(p1_concat_141219_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141219_comb;
  assign p1_sel_142936_comb = $signed(p1_or_140660_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140660_comb[23:10], 2'h0};
  assign p1_sel_142937_comb = $signed(p1_or_140661_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140661_comb[23:10], 2'h0};
  assign p1_sel_142938_comb = $signed(p1_concat_141229_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141229_comb;
  assign p1_sel_142939_comb = $signed(p1_concat_141231_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141231_comb;
  assign p1_sel_142940_comb = $signed(p1_or_140666_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140666_comb[23:10], 2'h0};
  assign p1_sel_142941_comb = $signed(p1_or_140667_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140667_comb[23:10], 2'h0};
  assign p1_sel_142942_comb = $signed(p1_concat_141241_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141241_comb;
  assign p1_sel_142943_comb = $signed(p1_concat_141243_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141243_comb;
  assign p1_sel_142944_comb = $signed(p1_or_140672_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140672_comb[23:10], 2'h0};
  assign p1_smul_142945_comb = smul16b_8b_x_9b(p1_shifted__64_squeezed_comb, 9'h0d5);
  assign p1_sel_142946_comb = $signed(p1_or_140673_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140673_comb[23:9], 1'h0};
  assign p1_smul_142947_comb = smul16b_8b_x_9b(p1_shifted__66_squeezed_comb, 9'h105);
  assign p1_sel_142948_comb = $signed(p1_or_140674_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140674_comb[23:9], 1'h0};
  assign p1_sel_142949_comb = $signed(p1_or_140675_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140675_comb[23:9], 1'h0};
  assign p1_smul_142950_comb = smul16b_8b_x_9b(p1_shifted__69_squeezed_comb, 9'h0fb);
  assign p1_sel_142951_comb = $signed(p1_or_140676_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140676_comb[23:9], 1'h0};
  assign p1_smul_142952_comb = smul16b_8b_x_9b(p1_shifted__71_squeezed_comb, 9'h12b);
  assign p1_smul_142953_comb = smul16b_8b_x_9b(p1_shifted__72_squeezed_comb, 9'h0d5);
  assign p1_sel_142954_comb = $signed(p1_or_140677_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140677_comb[23:9], 1'h0};
  assign p1_smul_142955_comb = smul16b_8b_x_9b(p1_shifted__74_squeezed_comb, 9'h105);
  assign p1_sel_142956_comb = $signed(p1_or_140678_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140678_comb[23:9], 1'h0};
  assign p1_sel_142957_comb = $signed(p1_or_140679_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140679_comb[23:9], 1'h0};
  assign p1_smul_142958_comb = smul16b_8b_x_9b(p1_shifted__77_squeezed_comb, 9'h0fb);
  assign p1_sel_142959_comb = $signed(p1_or_140680_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140680_comb[23:9], 1'h0};
  assign p1_smul_142960_comb = smul16b_8b_x_9b(p1_shifted__79_squeezed_comb, 9'h12b);
  assign p1_smul_142961_comb = smul16b_8b_x_9b(p1_shifted__80_squeezed_comb, 9'h0d5);
  assign p1_sel_142962_comb = $signed(p1_or_140681_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140681_comb[23:9], 1'h0};
  assign p1_smul_142963_comb = smul16b_8b_x_9b(p1_shifted__82_squeezed_comb, 9'h105);
  assign p1_sel_142964_comb = $signed(p1_or_140682_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140682_comb[23:9], 1'h0};
  assign p1_sel_142965_comb = $signed(p1_or_140683_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140683_comb[23:9], 1'h0};
  assign p1_smul_142966_comb = smul16b_8b_x_9b(p1_shifted__85_squeezed_comb, 9'h0fb);
  assign p1_sel_142967_comb = $signed(p1_or_140684_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140684_comb[23:9], 1'h0};
  assign p1_smul_142968_comb = smul16b_8b_x_9b(p1_shifted__87_squeezed_comb, 9'h12b);
  assign p1_smul_142969_comb = smul16b_8b_x_9b(p1_shifted__88_squeezed_comb, 9'h0d5);
  assign p1_sel_142970_comb = $signed(p1_or_140685_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140685_comb[23:9], 1'h0};
  assign p1_smul_142971_comb = smul16b_8b_x_9b(p1_shifted__90_squeezed_comb, 9'h105);
  assign p1_sel_142972_comb = $signed(p1_or_140686_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140686_comb[23:9], 1'h0};
  assign p1_sel_142973_comb = $signed(p1_or_140687_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140687_comb[23:9], 1'h0};
  assign p1_smul_142974_comb = smul16b_8b_x_9b(p1_shifted__93_squeezed_comb, 9'h0fb);
  assign p1_sel_142975_comb = $signed(p1_or_140688_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140688_comb[23:9], 1'h0};
  assign p1_smul_142976_comb = smul16b_8b_x_9b(p1_shifted__95_squeezed_comb, 9'h12b);
  assign p1_smul_142977_comb = smul16b_8b_x_9b(p1_shifted__96_squeezed_comb, 9'h0d5);
  assign p1_sel_142978_comb = $signed(p1_or_140689_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140689_comb[23:9], 1'h0};
  assign p1_smul_142979_comb = smul16b_8b_x_9b(p1_shifted__98_squeezed_comb, 9'h105);
  assign p1_sel_142980_comb = $signed(p1_or_140690_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140690_comb[23:9], 1'h0};
  assign p1_sel_142981_comb = $signed(p1_or_140691_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140691_comb[23:9], 1'h0};
  assign p1_smul_142982_comb = smul16b_8b_x_9b(p1_shifted__101_squeezed_comb, 9'h0fb);
  assign p1_sel_142983_comb = $signed(p1_or_140692_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140692_comb[23:9], 1'h0};
  assign p1_smul_142984_comb = smul16b_8b_x_9b(p1_shifted__103_squeezed_comb, 9'h12b);
  assign p1_smul_142985_comb = smul16b_8b_x_9b(p1_shifted__104_squeezed_comb, 9'h0d5);
  assign p1_sel_142986_comb = $signed(p1_or_140693_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140693_comb[23:9], 1'h0};
  assign p1_smul_142987_comb = smul16b_8b_x_9b(p1_shifted__106_squeezed_comb, 9'h105);
  assign p1_sel_142988_comb = $signed(p1_or_140694_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140694_comb[23:9], 1'h0};
  assign p1_sel_142989_comb = $signed(p1_or_140695_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140695_comb[23:9], 1'h0};
  assign p1_smul_142990_comb = smul16b_8b_x_9b(p1_shifted__109_squeezed_comb, 9'h0fb);
  assign p1_sel_142991_comb = $signed(p1_or_140696_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140696_comb[23:9], 1'h0};
  assign p1_smul_142992_comb = smul16b_8b_x_9b(p1_shifted__111_squeezed_comb, 9'h12b);
  assign p1_smul_142993_comb = smul16b_8b_x_9b(p1_shifted__112_squeezed_comb, 9'h0d5);
  assign p1_sel_142994_comb = $signed(p1_or_140697_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140697_comb[23:9], 1'h0};
  assign p1_smul_142995_comb = smul16b_8b_x_9b(p1_shifted__114_squeezed_comb, 9'h105);
  assign p1_sel_142996_comb = $signed(p1_or_140698_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140698_comb[23:9], 1'h0};
  assign p1_sel_142997_comb = $signed(p1_or_140699_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140699_comb[23:9], 1'h0};
  assign p1_smul_142998_comb = smul16b_8b_x_9b(p1_shifted__117_squeezed_comb, 9'h0fb);
  assign p1_sel_142999_comb = $signed(p1_or_140700_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140700_comb[23:9], 1'h0};
  assign p1_smul_143000_comb = smul16b_8b_x_9b(p1_shifted__119_squeezed_comb, 9'h12b);
  assign p1_smul_143001_comb = smul16b_8b_x_9b(p1_shifted__120_squeezed_comb, 9'h0d5);
  assign p1_sel_143002_comb = $signed(p1_or_140701_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140701_comb[23:9], 1'h0};
  assign p1_smul_143003_comb = smul16b_8b_x_9b(p1_shifted__122_squeezed_comb, 9'h105);
  assign p1_sel_143004_comb = $signed(p1_or_140702_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140702_comb[23:9], 1'h0};
  assign p1_sel_143005_comb = $signed(p1_or_140703_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140703_comb[23:9], 1'h0};
  assign p1_smul_143006_comb = smul16b_8b_x_9b(p1_shifted__125_squeezed_comb, 9'h0fb);
  assign p1_sel_143007_comb = $signed(p1_or_140704_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140704_comb[23:9], 1'h0};
  assign p1_smul_143008_comb = smul16b_8b_x_9b(p1_shifted__127_squeezed_comb, 9'h12b);
  assign p1_smul_143009_comb = smul16b_8b_x_9b(p1_shifted__64_squeezed_comb, 9'h0b5);
  assign p1_smul_143010_comb = smul16b_8b_x_9b(p1_shifted__65_squeezed_comb, 9'h14b);
  assign p1_smul_143011_comb = smul16b_8b_x_9b(p1_shifted__66_squeezed_comb, 9'h14b);
  assign p1_smul_143012_comb = smul16b_8b_x_9b(p1_shifted__67_squeezed_comb, 9'h0b5);
  assign p1_smul_143013_comb = smul16b_8b_x_9b(p1_shifted__68_squeezed_comb, 9'h0b5);
  assign p1_smul_143014_comb = smul16b_8b_x_9b(p1_shifted__69_squeezed_comb, 9'h14b);
  assign p1_smul_143015_comb = smul16b_8b_x_9b(p1_shifted__70_squeezed_comb, 9'h14b);
  assign p1_smul_143016_comb = smul16b_8b_x_9b(p1_shifted__71_squeezed_comb, 9'h0b5);
  assign p1_smul_143017_comb = smul16b_8b_x_9b(p1_shifted__72_squeezed_comb, 9'h0b5);
  assign p1_smul_143018_comb = smul16b_8b_x_9b(p1_shifted__73_squeezed_comb, 9'h14b);
  assign p1_smul_143019_comb = smul16b_8b_x_9b(p1_shifted__74_squeezed_comb, 9'h14b);
  assign p1_smul_143020_comb = smul16b_8b_x_9b(p1_shifted__75_squeezed_comb, 9'h0b5);
  assign p1_smul_143021_comb = smul16b_8b_x_9b(p1_shifted__76_squeezed_comb, 9'h0b5);
  assign p1_smul_143022_comb = smul16b_8b_x_9b(p1_shifted__77_squeezed_comb, 9'h14b);
  assign p1_smul_143023_comb = smul16b_8b_x_9b(p1_shifted__78_squeezed_comb, 9'h14b);
  assign p1_smul_143024_comb = smul16b_8b_x_9b(p1_shifted__79_squeezed_comb, 9'h0b5);
  assign p1_smul_143025_comb = smul16b_8b_x_9b(p1_shifted__80_squeezed_comb, 9'h0b5);
  assign p1_smul_143026_comb = smul16b_8b_x_9b(p1_shifted__81_squeezed_comb, 9'h14b);
  assign p1_smul_143027_comb = smul16b_8b_x_9b(p1_shifted__82_squeezed_comb, 9'h14b);
  assign p1_smul_143028_comb = smul16b_8b_x_9b(p1_shifted__83_squeezed_comb, 9'h0b5);
  assign p1_smul_143029_comb = smul16b_8b_x_9b(p1_shifted__84_squeezed_comb, 9'h0b5);
  assign p1_smul_143030_comb = smul16b_8b_x_9b(p1_shifted__85_squeezed_comb, 9'h14b);
  assign p1_smul_143031_comb = smul16b_8b_x_9b(p1_shifted__86_squeezed_comb, 9'h14b);
  assign p1_smul_143032_comb = smul16b_8b_x_9b(p1_shifted__87_squeezed_comb, 9'h0b5);
  assign p1_smul_143033_comb = smul16b_8b_x_9b(p1_shifted__88_squeezed_comb, 9'h0b5);
  assign p1_smul_143034_comb = smul16b_8b_x_9b(p1_shifted__89_squeezed_comb, 9'h14b);
  assign p1_smul_143035_comb = smul16b_8b_x_9b(p1_shifted__90_squeezed_comb, 9'h14b);
  assign p1_smul_143036_comb = smul16b_8b_x_9b(p1_shifted__91_squeezed_comb, 9'h0b5);
  assign p1_smul_143037_comb = smul16b_8b_x_9b(p1_shifted__92_squeezed_comb, 9'h0b5);
  assign p1_smul_143038_comb = smul16b_8b_x_9b(p1_shifted__93_squeezed_comb, 9'h14b);
  assign p1_smul_143039_comb = smul16b_8b_x_9b(p1_shifted__94_squeezed_comb, 9'h14b);
  assign p1_smul_143040_comb = smul16b_8b_x_9b(p1_shifted__95_squeezed_comb, 9'h0b5);
  assign p1_smul_143041_comb = smul16b_8b_x_9b(p1_shifted__96_squeezed_comb, 9'h0b5);
  assign p1_smul_143042_comb = smul16b_8b_x_9b(p1_shifted__97_squeezed_comb, 9'h14b);
  assign p1_smul_143043_comb = smul16b_8b_x_9b(p1_shifted__98_squeezed_comb, 9'h14b);
  assign p1_smul_143044_comb = smul16b_8b_x_9b(p1_shifted__99_squeezed_comb, 9'h0b5);
  assign p1_smul_143045_comb = smul16b_8b_x_9b(p1_shifted__100_squeezed_comb, 9'h0b5);
  assign p1_smul_143046_comb = smul16b_8b_x_9b(p1_shifted__101_squeezed_comb, 9'h14b);
  assign p1_smul_143047_comb = smul16b_8b_x_9b(p1_shifted__102_squeezed_comb, 9'h14b);
  assign p1_smul_143048_comb = smul16b_8b_x_9b(p1_shifted__103_squeezed_comb, 9'h0b5);
  assign p1_smul_143049_comb = smul16b_8b_x_9b(p1_shifted__104_squeezed_comb, 9'h0b5);
  assign p1_smul_143050_comb = smul16b_8b_x_9b(p1_shifted__105_squeezed_comb, 9'h14b);
  assign p1_smul_143051_comb = smul16b_8b_x_9b(p1_shifted__106_squeezed_comb, 9'h14b);
  assign p1_smul_143052_comb = smul16b_8b_x_9b(p1_shifted__107_squeezed_comb, 9'h0b5);
  assign p1_smul_143053_comb = smul16b_8b_x_9b(p1_shifted__108_squeezed_comb, 9'h0b5);
  assign p1_smul_143054_comb = smul16b_8b_x_9b(p1_shifted__109_squeezed_comb, 9'h14b);
  assign p1_smul_143055_comb = smul16b_8b_x_9b(p1_shifted__110_squeezed_comb, 9'h14b);
  assign p1_smul_143056_comb = smul16b_8b_x_9b(p1_shifted__111_squeezed_comb, 9'h0b5);
  assign p1_smul_143057_comb = smul16b_8b_x_9b(p1_shifted__112_squeezed_comb, 9'h0b5);
  assign p1_smul_143058_comb = smul16b_8b_x_9b(p1_shifted__113_squeezed_comb, 9'h14b);
  assign p1_smul_143059_comb = smul16b_8b_x_9b(p1_shifted__114_squeezed_comb, 9'h14b);
  assign p1_smul_143060_comb = smul16b_8b_x_9b(p1_shifted__115_squeezed_comb, 9'h0b5);
  assign p1_smul_143061_comb = smul16b_8b_x_9b(p1_shifted__116_squeezed_comb, 9'h0b5);
  assign p1_smul_143062_comb = smul16b_8b_x_9b(p1_shifted__117_squeezed_comb, 9'h14b);
  assign p1_smul_143063_comb = smul16b_8b_x_9b(p1_shifted__118_squeezed_comb, 9'h14b);
  assign p1_smul_143064_comb = smul16b_8b_x_9b(p1_shifted__119_squeezed_comb, 9'h0b5);
  assign p1_smul_143065_comb = smul16b_8b_x_9b(p1_shifted__120_squeezed_comb, 9'h0b5);
  assign p1_smul_143066_comb = smul16b_8b_x_9b(p1_shifted__121_squeezed_comb, 9'h14b);
  assign p1_smul_143067_comb = smul16b_8b_x_9b(p1_shifted__122_squeezed_comb, 9'h14b);
  assign p1_smul_143068_comb = smul16b_8b_x_9b(p1_shifted__123_squeezed_comb, 9'h0b5);
  assign p1_smul_143069_comb = smul16b_8b_x_9b(p1_shifted__124_squeezed_comb, 9'h0b5);
  assign p1_smul_143070_comb = smul16b_8b_x_9b(p1_shifted__125_squeezed_comb, 9'h14b);
  assign p1_smul_143071_comb = smul16b_8b_x_9b(p1_shifted__126_squeezed_comb, 9'h14b);
  assign p1_smul_143072_comb = smul16b_8b_x_9b(p1_shifted__127_squeezed_comb, 9'h0b5);
  assign p1_sel_143073_comb = $signed(p1_or_140705_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140705_comb[23:9], 1'h0};
  assign p1_smul_143074_comb = smul16b_8b_x_9b(p1_shifted__65_squeezed_comb, 9'h105);
  assign p1_sel_143075_comb = $signed(p1_or_140706_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140706_comb[23:9], 1'h0};
  assign p1_smul_143076_comb = smul16b_8b_x_9b(p1_shifted__67_squeezed_comb, 9'h0d5);
  assign p1_smul_143077_comb = smul16b_8b_x_9b(p1_shifted__68_squeezed_comb, 9'h0d5);
  assign p1_sel_143078_comb = $signed(p1_or_140707_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140707_comb[23:9], 1'h0};
  assign p1_smul_143079_comb = smul16b_8b_x_9b(p1_shifted__70_squeezed_comb, 9'h105);
  assign p1_sel_143080_comb = $signed(p1_or_140708_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140708_comb[23:9], 1'h0};
  assign p1_sel_143081_comb = $signed(p1_or_140709_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140709_comb[23:9], 1'h0};
  assign p1_smul_143082_comb = smul16b_8b_x_9b(p1_shifted__73_squeezed_comb, 9'h105);
  assign p1_sel_143083_comb = $signed(p1_or_140710_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140710_comb[23:9], 1'h0};
  assign p1_smul_143084_comb = smul16b_8b_x_9b(p1_shifted__75_squeezed_comb, 9'h0d5);
  assign p1_smul_143085_comb = smul16b_8b_x_9b(p1_shifted__76_squeezed_comb, 9'h0d5);
  assign p1_sel_143086_comb = $signed(p1_or_140711_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140711_comb[23:9], 1'h0};
  assign p1_smul_143087_comb = smul16b_8b_x_9b(p1_shifted__78_squeezed_comb, 9'h105);
  assign p1_sel_143088_comb = $signed(p1_or_140712_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140712_comb[23:9], 1'h0};
  assign p1_sel_143089_comb = $signed(p1_or_140713_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140713_comb[23:9], 1'h0};
  assign p1_smul_143090_comb = smul16b_8b_x_9b(p1_shifted__81_squeezed_comb, 9'h105);
  assign p1_sel_143091_comb = $signed(p1_or_140714_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140714_comb[23:9], 1'h0};
  assign p1_smul_143092_comb = smul16b_8b_x_9b(p1_shifted__83_squeezed_comb, 9'h0d5);
  assign p1_smul_143093_comb = smul16b_8b_x_9b(p1_shifted__84_squeezed_comb, 9'h0d5);
  assign p1_sel_143094_comb = $signed(p1_or_140715_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140715_comb[23:9], 1'h0};
  assign p1_smul_143095_comb = smul16b_8b_x_9b(p1_shifted__86_squeezed_comb, 9'h105);
  assign p1_sel_143096_comb = $signed(p1_or_140716_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140716_comb[23:9], 1'h0};
  assign p1_sel_143097_comb = $signed(p1_or_140717_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140717_comb[23:9], 1'h0};
  assign p1_smul_143098_comb = smul16b_8b_x_9b(p1_shifted__89_squeezed_comb, 9'h105);
  assign p1_sel_143099_comb = $signed(p1_or_140718_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140718_comb[23:9], 1'h0};
  assign p1_smul_143100_comb = smul16b_8b_x_9b(p1_shifted__91_squeezed_comb, 9'h0d5);
  assign p1_smul_143101_comb = smul16b_8b_x_9b(p1_shifted__92_squeezed_comb, 9'h0d5);
  assign p1_sel_143102_comb = $signed(p1_or_140719_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140719_comb[23:9], 1'h0};
  assign p1_smul_143103_comb = smul16b_8b_x_9b(p1_shifted__94_squeezed_comb, 9'h105);
  assign p1_sel_143104_comb = $signed(p1_or_140720_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140720_comb[23:9], 1'h0};
  assign p1_sel_143105_comb = $signed(p1_or_140721_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140721_comb[23:9], 1'h0};
  assign p1_smul_143106_comb = smul16b_8b_x_9b(p1_shifted__97_squeezed_comb, 9'h105);
  assign p1_sel_143107_comb = $signed(p1_or_140722_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140722_comb[23:9], 1'h0};
  assign p1_smul_143108_comb = smul16b_8b_x_9b(p1_shifted__99_squeezed_comb, 9'h0d5);
  assign p1_smul_143109_comb = smul16b_8b_x_9b(p1_shifted__100_squeezed_comb, 9'h0d5);
  assign p1_sel_143110_comb = $signed(p1_or_140723_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140723_comb[23:9], 1'h0};
  assign p1_smul_143111_comb = smul16b_8b_x_9b(p1_shifted__102_squeezed_comb, 9'h105);
  assign p1_sel_143112_comb = $signed(p1_or_140724_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140724_comb[23:9], 1'h0};
  assign p1_sel_143113_comb = $signed(p1_or_140725_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140725_comb[23:9], 1'h0};
  assign p1_smul_143114_comb = smul16b_8b_x_9b(p1_shifted__105_squeezed_comb, 9'h105);
  assign p1_sel_143115_comb = $signed(p1_or_140726_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140726_comb[23:9], 1'h0};
  assign p1_smul_143116_comb = smul16b_8b_x_9b(p1_shifted__107_squeezed_comb, 9'h0d5);
  assign p1_smul_143117_comb = smul16b_8b_x_9b(p1_shifted__108_squeezed_comb, 9'h0d5);
  assign p1_sel_143118_comb = $signed(p1_or_140727_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140727_comb[23:9], 1'h0};
  assign p1_smul_143119_comb = smul16b_8b_x_9b(p1_shifted__110_squeezed_comb, 9'h105);
  assign p1_sel_143120_comb = $signed(p1_or_140728_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140728_comb[23:9], 1'h0};
  assign p1_sel_143121_comb = $signed(p1_or_140729_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140729_comb[23:9], 1'h0};
  assign p1_smul_143122_comb = smul16b_8b_x_9b(p1_shifted__113_squeezed_comb, 9'h105);
  assign p1_sel_143123_comb = $signed(p1_or_140730_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140730_comb[23:9], 1'h0};
  assign p1_smul_143124_comb = smul16b_8b_x_9b(p1_shifted__115_squeezed_comb, 9'h0d5);
  assign p1_smul_143125_comb = smul16b_8b_x_9b(p1_shifted__116_squeezed_comb, 9'h0d5);
  assign p1_sel_143126_comb = $signed(p1_or_140731_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140731_comb[23:9], 1'h0};
  assign p1_smul_143127_comb = smul16b_8b_x_9b(p1_shifted__118_squeezed_comb, 9'h105);
  assign p1_sel_143128_comb = $signed(p1_or_140732_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140732_comb[23:9], 1'h0};
  assign p1_sel_143129_comb = $signed(p1_or_140733_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140733_comb[23:9], 1'h0};
  assign p1_smul_143130_comb = smul16b_8b_x_9b(p1_shifted__121_squeezed_comb, 9'h105);
  assign p1_sel_143131_comb = $signed(p1_or_140734_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140734_comb[23:9], 1'h0};
  assign p1_smul_143132_comb = smul16b_8b_x_9b(p1_shifted__123_squeezed_comb, 9'h0d5);
  assign p1_smul_143133_comb = smul16b_8b_x_9b(p1_shifted__124_squeezed_comb, 9'h0d5);
  assign p1_sel_143134_comb = $signed(p1_or_140735_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140735_comb[23:9], 1'h0};
  assign p1_smul_143135_comb = smul16b_8b_x_9b(p1_shifted__126_squeezed_comb, 9'h105);
  assign p1_sel_143136_comb = $signed(p1_or_140736_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140736_comb[23:9], 1'h0};
  assign p1_sel_143137_comb = $signed(p1_concat_141505_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141505_comb;
  assign p1_sel_143138_comb = $signed(p1_or_140739_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140739_comb[23:10], 2'h0};
  assign p1_sel_143139_comb = $signed(p1_concat_141511_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141511_comb;
  assign p1_sel_143140_comb = $signed(p1_or_140742_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140742_comb[23:10], 2'h0};
  assign p1_sel_143141_comb = $signed(p1_or_140743_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140743_comb[23:10], 2'h0};
  assign p1_sel_143142_comb = $signed(p1_concat_141521_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141521_comb;
  assign p1_sel_143143_comb = $signed(p1_or_140746_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140746_comb[23:10], 2'h0};
  assign p1_sel_143144_comb = $signed(p1_concat_141527_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141527_comb;
  assign p1_sel_143145_comb = $signed(p1_concat_141529_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141529_comb;
  assign p1_sel_143146_comb = $signed(p1_or_140751_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140751_comb[23:10], 2'h0};
  assign p1_sel_143147_comb = $signed(p1_concat_141535_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141535_comb;
  assign p1_sel_143148_comb = $signed(p1_or_140754_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140754_comb[23:10], 2'h0};
  assign p1_sel_143149_comb = $signed(p1_or_140755_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140755_comb[23:10], 2'h0};
  assign p1_sel_143150_comb = $signed(p1_concat_141545_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141545_comb;
  assign p1_sel_143151_comb = $signed(p1_or_140758_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140758_comb[23:10], 2'h0};
  assign p1_sel_143152_comb = $signed(p1_concat_141551_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141551_comb;
  assign p1_sel_143153_comb = $signed(p1_concat_141553_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141553_comb;
  assign p1_sel_143154_comb = $signed(p1_or_140763_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140763_comb[23:10], 2'h0};
  assign p1_sel_143155_comb = $signed(p1_concat_141559_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141559_comb;
  assign p1_sel_143156_comb = $signed(p1_or_140766_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140766_comb[23:10], 2'h0};
  assign p1_sel_143157_comb = $signed(p1_or_140767_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140767_comb[23:10], 2'h0};
  assign p1_sel_143158_comb = $signed(p1_concat_141569_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141569_comb;
  assign p1_sel_143159_comb = $signed(p1_or_140770_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140770_comb[23:10], 2'h0};
  assign p1_sel_143160_comb = $signed(p1_concat_141575_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141575_comb;
  assign p1_sel_143161_comb = $signed(p1_concat_141577_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141577_comb;
  assign p1_sel_143162_comb = $signed(p1_or_140775_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140775_comb[23:10], 2'h0};
  assign p1_sel_143163_comb = $signed(p1_concat_141583_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141583_comb;
  assign p1_sel_143164_comb = $signed(p1_or_140778_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140778_comb[23:10], 2'h0};
  assign p1_sel_143165_comb = $signed(p1_or_140779_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140779_comb[23:10], 2'h0};
  assign p1_sel_143166_comb = $signed(p1_concat_141593_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141593_comb;
  assign p1_sel_143167_comb = $signed(p1_or_140782_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140782_comb[23:10], 2'h0};
  assign p1_sel_143168_comb = $signed(p1_concat_141599_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141599_comb;
  assign p1_sel_143169_comb = $signed(p1_concat_141601_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141601_comb;
  assign p1_sel_143170_comb = $signed(p1_or_140787_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140787_comb[23:10], 2'h0};
  assign p1_sel_143171_comb = $signed(p1_concat_141607_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141607_comb;
  assign p1_sel_143172_comb = $signed(p1_or_140790_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140790_comb[23:10], 2'h0};
  assign p1_sel_143173_comb = $signed(p1_or_140791_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140791_comb[23:10], 2'h0};
  assign p1_sel_143174_comb = $signed(p1_concat_141617_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141617_comb;
  assign p1_sel_143175_comb = $signed(p1_or_140794_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140794_comb[23:10], 2'h0};
  assign p1_sel_143176_comb = $signed(p1_concat_141623_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141623_comb;
  assign p1_sel_143177_comb = $signed(p1_concat_141625_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141625_comb;
  assign p1_sel_143178_comb = $signed(p1_or_140799_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140799_comb[23:10], 2'h0};
  assign p1_sel_143179_comb = $signed(p1_concat_141631_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141631_comb;
  assign p1_sel_143180_comb = $signed(p1_or_140802_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140802_comb[23:10], 2'h0};
  assign p1_sel_143181_comb = $signed(p1_or_140803_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140803_comb[23:10], 2'h0};
  assign p1_sel_143182_comb = $signed(p1_concat_141641_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141641_comb;
  assign p1_sel_143183_comb = $signed(p1_or_140806_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140806_comb[23:10], 2'h0};
  assign p1_sel_143184_comb = $signed(p1_concat_141647_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141647_comb;
  assign p1_sel_143185_comb = $signed(p1_concat_141649_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141649_comb;
  assign p1_sel_143186_comb = $signed(p1_or_140811_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140811_comb[23:10], 2'h0};
  assign p1_sel_143187_comb = $signed(p1_concat_141655_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141655_comb;
  assign p1_sel_143188_comb = $signed(p1_or_140814_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140814_comb[23:10], 2'h0};
  assign p1_sel_143189_comb = $signed(p1_or_140815_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140815_comb[23:10], 2'h0};
  assign p1_sel_143190_comb = $signed(p1_concat_141665_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141665_comb;
  assign p1_sel_143191_comb = $signed(p1_or_140818_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140818_comb[23:10], 2'h0};
  assign p1_sel_143192_comb = $signed(p1_concat_141671_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141671_comb;
  assign p1_sel_143193_comb = $signed(p1_concat_141673_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141673_comb;
  assign p1_sel_143194_comb = $signed(p1_or_140823_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140823_comb[23:10], 2'h0};
  assign p1_sel_143195_comb = $signed(p1_concat_141679_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141679_comb;
  assign p1_sel_143196_comb = $signed(p1_or_140826_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140826_comb[23:10], 2'h0};
  assign p1_sel_143197_comb = $signed(p1_or_140827_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140827_comb[23:10], 2'h0};
  assign p1_sel_143198_comb = $signed(p1_concat_141689_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141689_comb;
  assign p1_sel_143199_comb = $signed(p1_or_140830_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140830_comb[23:10], 2'h0};
  assign p1_sel_143200_comb = $signed(p1_concat_141695_comb) > $signed(16'h7fff) ? 16'h7fff : p1_concat_141695_comb;
  assign p1_sel_143201_comb = $signed(p1_or_140833_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140833_comb[23:9], 1'h0};
  assign p1_sel_143202_comb = $signed(p1_or_140834_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140834_comb[23:9], 1'h0};
  assign p1_smul_143203_comb = smul16b_8b_x_9b(p1_shifted__66_squeezed_comb, 9'h0d5);
  assign p1_smul_143204_comb = smul16b_8b_x_9b(p1_shifted__67_squeezed_comb, 9'h105);
  assign p1_smul_143205_comb = smul16b_8b_x_9b(p1_shifted__68_squeezed_comb, 9'h105);
  assign p1_smul_143206_comb = smul16b_8b_x_9b(p1_shifted__69_squeezed_comb, 9'h0d5);
  assign p1_sel_143207_comb = $signed(p1_or_140835_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140835_comb[23:9], 1'h0};
  assign p1_sel_143208_comb = $signed(p1_or_140836_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140836_comb[23:9], 1'h0};
  assign p1_sel_143209_comb = $signed(p1_or_140837_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140837_comb[23:9], 1'h0};
  assign p1_sel_143210_comb = $signed(p1_or_140838_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140838_comb[23:9], 1'h0};
  assign p1_smul_143211_comb = smul16b_8b_x_9b(p1_shifted__74_squeezed_comb, 9'h0d5);
  assign p1_smul_143212_comb = smul16b_8b_x_9b(p1_shifted__75_squeezed_comb, 9'h105);
  assign p1_smul_143213_comb = smul16b_8b_x_9b(p1_shifted__76_squeezed_comb, 9'h105);
  assign p1_smul_143214_comb = smul16b_8b_x_9b(p1_shifted__77_squeezed_comb, 9'h0d5);
  assign p1_sel_143215_comb = $signed(p1_or_140839_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140839_comb[23:9], 1'h0};
  assign p1_sel_143216_comb = $signed(p1_or_140840_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140840_comb[23:9], 1'h0};
  assign p1_sel_143217_comb = $signed(p1_or_140841_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140841_comb[23:9], 1'h0};
  assign p1_sel_143218_comb = $signed(p1_or_140842_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140842_comb[23:9], 1'h0};
  assign p1_smul_143219_comb = smul16b_8b_x_9b(p1_shifted__82_squeezed_comb, 9'h0d5);
  assign p1_smul_143220_comb = smul16b_8b_x_9b(p1_shifted__83_squeezed_comb, 9'h105);
  assign p1_smul_143221_comb = smul16b_8b_x_9b(p1_shifted__84_squeezed_comb, 9'h105);
  assign p1_smul_143222_comb = smul16b_8b_x_9b(p1_shifted__85_squeezed_comb, 9'h0d5);
  assign p1_sel_143223_comb = $signed(p1_or_140843_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140843_comb[23:9], 1'h0};
  assign p1_sel_143224_comb = $signed(p1_or_140844_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140844_comb[23:9], 1'h0};
  assign p1_sel_143225_comb = $signed(p1_or_140845_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140845_comb[23:9], 1'h0};
  assign p1_sel_143226_comb = $signed(p1_or_140846_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140846_comb[23:9], 1'h0};
  assign p1_smul_143227_comb = smul16b_8b_x_9b(p1_shifted__90_squeezed_comb, 9'h0d5);
  assign p1_smul_143228_comb = smul16b_8b_x_9b(p1_shifted__91_squeezed_comb, 9'h105);
  assign p1_smul_143229_comb = smul16b_8b_x_9b(p1_shifted__92_squeezed_comb, 9'h105);
  assign p1_smul_143230_comb = smul16b_8b_x_9b(p1_shifted__93_squeezed_comb, 9'h0d5);
  assign p1_sel_143231_comb = $signed(p1_or_140847_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140847_comb[23:9], 1'h0};
  assign p1_sel_143232_comb = $signed(p1_or_140848_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140848_comb[23:9], 1'h0};
  assign p1_sel_143233_comb = $signed(p1_or_140849_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140849_comb[23:9], 1'h0};
  assign p1_sel_143234_comb = $signed(p1_or_140850_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140850_comb[23:9], 1'h0};
  assign p1_smul_143235_comb = smul16b_8b_x_9b(p1_shifted__98_squeezed_comb, 9'h0d5);
  assign p1_smul_143236_comb = smul16b_8b_x_9b(p1_shifted__99_squeezed_comb, 9'h105);
  assign p1_smul_143237_comb = smul16b_8b_x_9b(p1_shifted__100_squeezed_comb, 9'h105);
  assign p1_smul_143238_comb = smul16b_8b_x_9b(p1_shifted__101_squeezed_comb, 9'h0d5);
  assign p1_sel_143239_comb = $signed(p1_or_140851_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140851_comb[23:9], 1'h0};
  assign p1_sel_143240_comb = $signed(p1_or_140852_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140852_comb[23:9], 1'h0};
  assign p1_sel_143241_comb = $signed(p1_or_140853_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140853_comb[23:9], 1'h0};
  assign p1_sel_143242_comb = $signed(p1_or_140854_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140854_comb[23:9], 1'h0};
  assign p1_smul_143243_comb = smul16b_8b_x_9b(p1_shifted__106_squeezed_comb, 9'h0d5);
  assign p1_smul_143244_comb = smul16b_8b_x_9b(p1_shifted__107_squeezed_comb, 9'h105);
  assign p1_smul_143245_comb = smul16b_8b_x_9b(p1_shifted__108_squeezed_comb, 9'h105);
  assign p1_smul_143246_comb = smul16b_8b_x_9b(p1_shifted__109_squeezed_comb, 9'h0d5);
  assign p1_sel_143247_comb = $signed(p1_or_140855_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140855_comb[23:9], 1'h0};
  assign p1_sel_143248_comb = $signed(p1_or_140856_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140856_comb[23:9], 1'h0};
  assign p1_sel_143249_comb = $signed(p1_or_140857_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140857_comb[23:9], 1'h0};
  assign p1_sel_143250_comb = $signed(p1_or_140858_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140858_comb[23:9], 1'h0};
  assign p1_smul_143251_comb = smul16b_8b_x_9b(p1_shifted__114_squeezed_comb, 9'h0d5);
  assign p1_smul_143252_comb = smul16b_8b_x_9b(p1_shifted__115_squeezed_comb, 9'h105);
  assign p1_smul_143253_comb = smul16b_8b_x_9b(p1_shifted__116_squeezed_comb, 9'h105);
  assign p1_smul_143254_comb = smul16b_8b_x_9b(p1_shifted__117_squeezed_comb, 9'h0d5);
  assign p1_sel_143255_comb = $signed(p1_or_140859_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140859_comb[23:9], 1'h0};
  assign p1_sel_143256_comb = $signed(p1_or_140860_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140860_comb[23:9], 1'h0};
  assign p1_sel_143257_comb = $signed(p1_or_140861_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140861_comb[23:9], 1'h0};
  assign p1_sel_143258_comb = $signed(p1_or_140862_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140862_comb[23:9], 1'h0};
  assign p1_smul_143259_comb = smul16b_8b_x_9b(p1_shifted__122_squeezed_comb, 9'h0d5);
  assign p1_smul_143260_comb = smul16b_8b_x_9b(p1_shifted__123_squeezed_comb, 9'h105);
  assign p1_smul_143261_comb = smul16b_8b_x_9b(p1_shifted__124_squeezed_comb, 9'h105);
  assign p1_smul_143262_comb = smul16b_8b_x_9b(p1_shifted__125_squeezed_comb, 9'h0d5);
  assign p1_sel_143263_comb = $signed(p1_or_140863_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140863_comb[23:9], 1'h0};
  assign p1_sel_143264_comb = $signed(p1_or_140864_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_140864_comb[23:9], 1'h0};
  assign p1_sum__520_comb = {{15{p1_add_142785_comb[16]}}, p1_add_142785_comb};
  assign p1_sum__521_comb = {{15{p1_add_142786_comb[16]}}, p1_add_142786_comb};
  assign p1_sum__522_comb = {{15{p1_add_142787_comb[16]}}, p1_add_142787_comb};
  assign p1_sum__523_comb = {{15{p1_add_142788_comb[16]}}, p1_add_142788_comb};
  assign p1_sum__464_comb = {{15{p1_add_142789_comb[16]}}, p1_add_142789_comb};
  assign p1_sum__465_comb = {{15{p1_add_142790_comb[16]}}, p1_add_142790_comb};
  assign p1_sum__466_comb = {{15{p1_add_142791_comb[16]}}, p1_add_142791_comb};
  assign p1_sum__467_comb = {{15{p1_add_142792_comb[16]}}, p1_add_142792_comb};
  assign p1_sum__408_comb = {{15{p1_add_142793_comb[16]}}, p1_add_142793_comb};
  assign p1_sum__409_comb = {{15{p1_add_142794_comb[16]}}, p1_add_142794_comb};
  assign p1_sum__410_comb = {{15{p1_add_142795_comb[16]}}, p1_add_142795_comb};
  assign p1_sum__411_comb = {{15{p1_add_142796_comb[16]}}, p1_add_142796_comb};
  assign p1_sum__352_comb = {{15{p1_add_142797_comb[16]}}, p1_add_142797_comb};
  assign p1_sum__353_comb = {{15{p1_add_142798_comb[16]}}, p1_add_142798_comb};
  assign p1_sum__354_comb = {{15{p1_add_142799_comb[16]}}, p1_add_142799_comb};
  assign p1_sum__355_comb = {{15{p1_add_142800_comb[16]}}, p1_add_142800_comb};
  assign p1_sum__296_comb = {{15{p1_add_142801_comb[16]}}, p1_add_142801_comb};
  assign p1_sum__297_comb = {{15{p1_add_142802_comb[16]}}, p1_add_142802_comb};
  assign p1_sum__298_comb = {{15{p1_add_142803_comb[16]}}, p1_add_142803_comb};
  assign p1_sum__299_comb = {{15{p1_add_142804_comb[16]}}, p1_add_142804_comb};
  assign p1_sum__240_comb = {{15{p1_add_142805_comb[16]}}, p1_add_142805_comb};
  assign p1_sum__241_comb = {{15{p1_add_142806_comb[16]}}, p1_add_142806_comb};
  assign p1_sum__242_comb = {{15{p1_add_142807_comb[16]}}, p1_add_142807_comb};
  assign p1_sum__243_comb = {{15{p1_add_142808_comb[16]}}, p1_add_142808_comb};
  assign p1_sum__184_comb = {{15{p1_add_142809_comb[16]}}, p1_add_142809_comb};
  assign p1_sum__185_comb = {{15{p1_add_142810_comb[16]}}, p1_add_142810_comb};
  assign p1_sum__186_comb = {{15{p1_add_142811_comb[16]}}, p1_add_142811_comb};
  assign p1_sum__187_comb = {{15{p1_add_142812_comb[16]}}, p1_add_142812_comb};
  assign p1_sum__128_comb = {{15{p1_add_142813_comb[16]}}, p1_add_142813_comb};
  assign p1_sum__129_comb = {{15{p1_add_142814_comb[16]}}, p1_add_142814_comb};
  assign p1_sum__130_comb = {{15{p1_add_142815_comb[16]}}, p1_add_142815_comb};
  assign p1_sum__131_comb = {{15{p1_add_142816_comb[16]}}, p1_add_142816_comb};
  assign p1_sum__524_comb = p1_sum__520_comb + p1_sum__521_comb;
  assign p1_sum__525_comb = p1_sum__522_comb + p1_sum__523_comb;
  assign p1_sum__468_comb = p1_sum__464_comb + p1_sum__465_comb;
  assign p1_sum__469_comb = p1_sum__466_comb + p1_sum__467_comb;
  assign p1_sum__412_comb = p1_sum__408_comb + p1_sum__409_comb;
  assign p1_sum__413_comb = p1_sum__410_comb + p1_sum__411_comb;
  assign p1_sum__356_comb = p1_sum__352_comb + p1_sum__353_comb;
  assign p1_sum__357_comb = p1_sum__354_comb + p1_sum__355_comb;
  assign p1_sum__300_comb = p1_sum__296_comb + p1_sum__297_comb;
  assign p1_sum__301_comb = p1_sum__298_comb + p1_sum__299_comb;
  assign p1_sum__244_comb = p1_sum__240_comb + p1_sum__241_comb;
  assign p1_sum__245_comb = p1_sum__242_comb + p1_sum__243_comb;
  assign p1_sum__188_comb = p1_sum__184_comb + p1_sum__185_comb;
  assign p1_sum__189_comb = p1_sum__186_comb + p1_sum__187_comb;
  assign p1_sum__132_comb = p1_sum__128_comb + p1_sum__129_comb;
  assign p1_sum__133_comb = p1_sum__130_comb + p1_sum__131_comb;
  assign p1_add_143761_comb = {{1{p1_smul_142817_comb[15]}}, p1_smul_142817_comb} + {{1{p1_smul_142818_comb[15]}}, p1_smul_142818_comb};
  assign p1_add_143762_comb = {{1{p1_sel_142819_comb[15]}}, p1_sel_142819_comb} + {{1{p1_sel_142820_comb[15]}}, p1_sel_142820_comb};
  assign p1_add_143763_comb = {{1{p1_sel_142821_comb[15]}}, p1_sel_142821_comb} + {{1{p1_sel_142822_comb[15]}}, p1_sel_142822_comb};
  assign p1_add_143764_comb = {{1{p1_smul_142823_comb[15]}}, p1_smul_142823_comb} + {{1{p1_smul_142824_comb[15]}}, p1_smul_142824_comb};
  assign p1_add_143765_comb = {{1{p1_smul_142825_comb[15]}}, p1_smul_142825_comb} + {{1{p1_smul_142826_comb[15]}}, p1_smul_142826_comb};
  assign p1_add_143766_comb = {{1{p1_sel_142827_comb[15]}}, p1_sel_142827_comb} + {{1{p1_sel_142828_comb[15]}}, p1_sel_142828_comb};
  assign p1_add_143767_comb = {{1{p1_sel_142829_comb[15]}}, p1_sel_142829_comb} + {{1{p1_sel_142830_comb[15]}}, p1_sel_142830_comb};
  assign p1_add_143768_comb = {{1{p1_smul_142831_comb[15]}}, p1_smul_142831_comb} + {{1{p1_smul_142832_comb[15]}}, p1_smul_142832_comb};
  assign p1_add_143769_comb = {{1{p1_smul_142833_comb[15]}}, p1_smul_142833_comb} + {{1{p1_smul_142834_comb[15]}}, p1_smul_142834_comb};
  assign p1_add_143770_comb = {{1{p1_sel_142835_comb[15]}}, p1_sel_142835_comb} + {{1{p1_sel_142836_comb[15]}}, p1_sel_142836_comb};
  assign p1_add_143771_comb = {{1{p1_sel_142837_comb[15]}}, p1_sel_142837_comb} + {{1{p1_sel_142838_comb[15]}}, p1_sel_142838_comb};
  assign p1_add_143772_comb = {{1{p1_smul_142839_comb[15]}}, p1_smul_142839_comb} + {{1{p1_smul_142840_comb[15]}}, p1_smul_142840_comb};
  assign p1_add_143773_comb = {{1{p1_smul_142841_comb[15]}}, p1_smul_142841_comb} + {{1{p1_smul_142842_comb[15]}}, p1_smul_142842_comb};
  assign p1_add_143774_comb = {{1{p1_sel_142843_comb[15]}}, p1_sel_142843_comb} + {{1{p1_sel_142844_comb[15]}}, p1_sel_142844_comb};
  assign p1_add_143775_comb = {{1{p1_sel_142845_comb[15]}}, p1_sel_142845_comb} + {{1{p1_sel_142846_comb[15]}}, p1_sel_142846_comb};
  assign p1_add_143776_comb = {{1{p1_smul_142847_comb[15]}}, p1_smul_142847_comb} + {{1{p1_smul_142848_comb[15]}}, p1_smul_142848_comb};
  assign p1_add_143777_comb = {{1{p1_smul_142849_comb[15]}}, p1_smul_142849_comb} + {{1{p1_smul_142850_comb[15]}}, p1_smul_142850_comb};
  assign p1_add_143778_comb = {{1{p1_sel_142851_comb[15]}}, p1_sel_142851_comb} + {{1{p1_sel_142852_comb[15]}}, p1_sel_142852_comb};
  assign p1_add_143779_comb = {{1{p1_sel_142853_comb[15]}}, p1_sel_142853_comb} + {{1{p1_sel_142854_comb[15]}}, p1_sel_142854_comb};
  assign p1_add_143780_comb = {{1{p1_smul_142855_comb[15]}}, p1_smul_142855_comb} + {{1{p1_smul_142856_comb[15]}}, p1_smul_142856_comb};
  assign p1_add_143781_comb = {{1{p1_smul_142857_comb[15]}}, p1_smul_142857_comb} + {{1{p1_smul_142858_comb[15]}}, p1_smul_142858_comb};
  assign p1_add_143782_comb = {{1{p1_sel_142859_comb[15]}}, p1_sel_142859_comb} + {{1{p1_sel_142860_comb[15]}}, p1_sel_142860_comb};
  assign p1_add_143783_comb = {{1{p1_sel_142861_comb[15]}}, p1_sel_142861_comb} + {{1{p1_sel_142862_comb[15]}}, p1_sel_142862_comb};
  assign p1_add_143784_comb = {{1{p1_smul_142863_comb[15]}}, p1_smul_142863_comb} + {{1{p1_smul_142864_comb[15]}}, p1_smul_142864_comb};
  assign p1_add_143785_comb = {{1{p1_smul_142865_comb[15]}}, p1_smul_142865_comb} + {{1{p1_smul_142866_comb[15]}}, p1_smul_142866_comb};
  assign p1_add_143786_comb = {{1{p1_sel_142867_comb[15]}}, p1_sel_142867_comb} + {{1{p1_sel_142868_comb[15]}}, p1_sel_142868_comb};
  assign p1_add_143787_comb = {{1{p1_sel_142869_comb[15]}}, p1_sel_142869_comb} + {{1{p1_sel_142870_comb[15]}}, p1_sel_142870_comb};
  assign p1_add_143788_comb = {{1{p1_smul_142871_comb[15]}}, p1_smul_142871_comb} + {{1{p1_smul_142872_comb[15]}}, p1_smul_142872_comb};
  assign p1_add_143789_comb = {{1{p1_smul_142873_comb[15]}}, p1_smul_142873_comb} + {{1{p1_smul_142874_comb[15]}}, p1_smul_142874_comb};
  assign p1_add_143790_comb = {{1{p1_sel_142875_comb[15]}}, p1_sel_142875_comb} + {{1{p1_sel_142876_comb[15]}}, p1_sel_142876_comb};
  assign p1_add_143791_comb = {{1{p1_sel_142877_comb[15]}}, p1_sel_142877_comb} + {{1{p1_sel_142878_comb[15]}}, p1_sel_142878_comb};
  assign p1_add_143792_comb = {{1{p1_smul_142879_comb[15]}}, p1_smul_142879_comb} + {{1{p1_smul_142880_comb[15]}}, p1_smul_142880_comb};
  assign p1_add_143793_comb = {{1{p1_sel_142881_comb[15]}}, p1_sel_142881_comb} + {{1{p1_sel_142882_comb[15]}}, p1_sel_142882_comb};
  assign p1_add_143794_comb = {{1{p1_sel_142883_comb[15]}}, p1_sel_142883_comb} + {{1{p1_sel_142884_comb[15]}}, p1_sel_142884_comb};
  assign p1_add_143795_comb = {{1{p1_sel_142885_comb[15]}}, p1_sel_142885_comb} + {{1{p1_sel_142886_comb[15]}}, p1_sel_142886_comb};
  assign p1_add_143796_comb = {{1{p1_sel_142887_comb[15]}}, p1_sel_142887_comb} + {{1{p1_sel_142888_comb[15]}}, p1_sel_142888_comb};
  assign p1_add_143797_comb = {{1{p1_sel_142889_comb[15]}}, p1_sel_142889_comb} + {{1{p1_sel_142890_comb[15]}}, p1_sel_142890_comb};
  assign p1_add_143798_comb = {{1{p1_sel_142891_comb[15]}}, p1_sel_142891_comb} + {{1{p1_sel_142892_comb[15]}}, p1_sel_142892_comb};
  assign p1_add_143799_comb = {{1{p1_sel_142893_comb[15]}}, p1_sel_142893_comb} + {{1{p1_sel_142894_comb[15]}}, p1_sel_142894_comb};
  assign p1_add_143800_comb = {{1{p1_sel_142895_comb[15]}}, p1_sel_142895_comb} + {{1{p1_sel_142896_comb[15]}}, p1_sel_142896_comb};
  assign p1_add_143801_comb = {{1{p1_sel_142897_comb[15]}}, p1_sel_142897_comb} + {{1{p1_sel_142898_comb[15]}}, p1_sel_142898_comb};
  assign p1_add_143802_comb = {{1{p1_sel_142899_comb[15]}}, p1_sel_142899_comb} + {{1{p1_sel_142900_comb[15]}}, p1_sel_142900_comb};
  assign p1_add_143803_comb = {{1{p1_sel_142901_comb[15]}}, p1_sel_142901_comb} + {{1{p1_sel_142902_comb[15]}}, p1_sel_142902_comb};
  assign p1_add_143804_comb = {{1{p1_sel_142903_comb[15]}}, p1_sel_142903_comb} + {{1{p1_sel_142904_comb[15]}}, p1_sel_142904_comb};
  assign p1_add_143805_comb = {{1{p1_sel_142905_comb[15]}}, p1_sel_142905_comb} + {{1{p1_sel_142906_comb[15]}}, p1_sel_142906_comb};
  assign p1_add_143806_comb = {{1{p1_sel_142907_comb[15]}}, p1_sel_142907_comb} + {{1{p1_sel_142908_comb[15]}}, p1_sel_142908_comb};
  assign p1_add_143807_comb = {{1{p1_sel_142909_comb[15]}}, p1_sel_142909_comb} + {{1{p1_sel_142910_comb[15]}}, p1_sel_142910_comb};
  assign p1_add_143808_comb = {{1{p1_sel_142911_comb[15]}}, p1_sel_142911_comb} + {{1{p1_sel_142912_comb[15]}}, p1_sel_142912_comb};
  assign p1_add_143809_comb = {{1{p1_sel_142913_comb[15]}}, p1_sel_142913_comb} + {{1{p1_sel_142914_comb[15]}}, p1_sel_142914_comb};
  assign p1_add_143810_comb = {{1{p1_sel_142915_comb[15]}}, p1_sel_142915_comb} + {{1{p1_sel_142916_comb[15]}}, p1_sel_142916_comb};
  assign p1_add_143811_comb = {{1{p1_sel_142917_comb[15]}}, p1_sel_142917_comb} + {{1{p1_sel_142918_comb[15]}}, p1_sel_142918_comb};
  assign p1_add_143812_comb = {{1{p1_sel_142919_comb[15]}}, p1_sel_142919_comb} + {{1{p1_sel_142920_comb[15]}}, p1_sel_142920_comb};
  assign p1_add_143813_comb = {{1{p1_sel_142921_comb[15]}}, p1_sel_142921_comb} + {{1{p1_sel_142922_comb[15]}}, p1_sel_142922_comb};
  assign p1_add_143814_comb = {{1{p1_sel_142923_comb[15]}}, p1_sel_142923_comb} + {{1{p1_sel_142924_comb[15]}}, p1_sel_142924_comb};
  assign p1_add_143815_comb = {{1{p1_sel_142925_comb[15]}}, p1_sel_142925_comb} + {{1{p1_sel_142926_comb[15]}}, p1_sel_142926_comb};
  assign p1_add_143816_comb = {{1{p1_sel_142927_comb[15]}}, p1_sel_142927_comb} + {{1{p1_sel_142928_comb[15]}}, p1_sel_142928_comb};
  assign p1_add_143817_comb = {{1{p1_sel_142929_comb[15]}}, p1_sel_142929_comb} + {{1{p1_sel_142930_comb[15]}}, p1_sel_142930_comb};
  assign p1_add_143818_comb = {{1{p1_sel_142931_comb[15]}}, p1_sel_142931_comb} + {{1{p1_sel_142932_comb[15]}}, p1_sel_142932_comb};
  assign p1_add_143819_comb = {{1{p1_sel_142933_comb[15]}}, p1_sel_142933_comb} + {{1{p1_sel_142934_comb[15]}}, p1_sel_142934_comb};
  assign p1_add_143820_comb = {{1{p1_sel_142935_comb[15]}}, p1_sel_142935_comb} + {{1{p1_sel_142936_comb[15]}}, p1_sel_142936_comb};
  assign p1_add_143821_comb = {{1{p1_sel_142937_comb[15]}}, p1_sel_142937_comb} + {{1{p1_sel_142938_comb[15]}}, p1_sel_142938_comb};
  assign p1_add_143822_comb = {{1{p1_sel_142939_comb[15]}}, p1_sel_142939_comb} + {{1{p1_sel_142940_comb[15]}}, p1_sel_142940_comb};
  assign p1_add_143823_comb = {{1{p1_sel_142941_comb[15]}}, p1_sel_142941_comb} + {{1{p1_sel_142942_comb[15]}}, p1_sel_142942_comb};
  assign p1_add_143824_comb = {{1{p1_sel_142943_comb[15]}}, p1_sel_142943_comb} + {{1{p1_sel_142944_comb[15]}}, p1_sel_142944_comb};
  assign p1_add_143825_comb = {{1{p1_smul_142945_comb[15]}}, p1_smul_142945_comb} + {{1{p1_sel_142946_comb[15]}}, p1_sel_142946_comb};
  assign p1_add_143826_comb = {{1{p1_smul_142947_comb[15]}}, p1_smul_142947_comb} + {{1{p1_sel_142948_comb[15]}}, p1_sel_142948_comb};
  assign p1_add_143827_comb = {{1{p1_sel_142949_comb[15]}}, p1_sel_142949_comb} + {{1{p1_smul_142950_comb[15]}}, p1_smul_142950_comb};
  assign p1_add_143828_comb = {{1{p1_sel_142951_comb[15]}}, p1_sel_142951_comb} + {{1{p1_smul_142952_comb[15]}}, p1_smul_142952_comb};
  assign p1_add_143829_comb = {{1{p1_smul_142953_comb[15]}}, p1_smul_142953_comb} + {{1{p1_sel_142954_comb[15]}}, p1_sel_142954_comb};
  assign p1_add_143830_comb = {{1{p1_smul_142955_comb[15]}}, p1_smul_142955_comb} + {{1{p1_sel_142956_comb[15]}}, p1_sel_142956_comb};
  assign p1_add_143831_comb = {{1{p1_sel_142957_comb[15]}}, p1_sel_142957_comb} + {{1{p1_smul_142958_comb[15]}}, p1_smul_142958_comb};
  assign p1_add_143832_comb = {{1{p1_sel_142959_comb[15]}}, p1_sel_142959_comb} + {{1{p1_smul_142960_comb[15]}}, p1_smul_142960_comb};
  assign p1_add_143833_comb = {{1{p1_smul_142961_comb[15]}}, p1_smul_142961_comb} + {{1{p1_sel_142962_comb[15]}}, p1_sel_142962_comb};
  assign p1_add_143834_comb = {{1{p1_smul_142963_comb[15]}}, p1_smul_142963_comb} + {{1{p1_sel_142964_comb[15]}}, p1_sel_142964_comb};
  assign p1_add_143835_comb = {{1{p1_sel_142965_comb[15]}}, p1_sel_142965_comb} + {{1{p1_smul_142966_comb[15]}}, p1_smul_142966_comb};
  assign p1_add_143836_comb = {{1{p1_sel_142967_comb[15]}}, p1_sel_142967_comb} + {{1{p1_smul_142968_comb[15]}}, p1_smul_142968_comb};
  assign p1_add_143837_comb = {{1{p1_smul_142969_comb[15]}}, p1_smul_142969_comb} + {{1{p1_sel_142970_comb[15]}}, p1_sel_142970_comb};
  assign p1_add_143838_comb = {{1{p1_smul_142971_comb[15]}}, p1_smul_142971_comb} + {{1{p1_sel_142972_comb[15]}}, p1_sel_142972_comb};
  assign p1_add_143839_comb = {{1{p1_sel_142973_comb[15]}}, p1_sel_142973_comb} + {{1{p1_smul_142974_comb[15]}}, p1_smul_142974_comb};
  assign p1_add_143840_comb = {{1{p1_sel_142975_comb[15]}}, p1_sel_142975_comb} + {{1{p1_smul_142976_comb[15]}}, p1_smul_142976_comb};
  assign p1_add_143841_comb = {{1{p1_smul_142977_comb[15]}}, p1_smul_142977_comb} + {{1{p1_sel_142978_comb[15]}}, p1_sel_142978_comb};
  assign p1_add_143842_comb = {{1{p1_smul_142979_comb[15]}}, p1_smul_142979_comb} + {{1{p1_sel_142980_comb[15]}}, p1_sel_142980_comb};
  assign p1_add_143843_comb = {{1{p1_sel_142981_comb[15]}}, p1_sel_142981_comb} + {{1{p1_smul_142982_comb[15]}}, p1_smul_142982_comb};
  assign p1_add_143844_comb = {{1{p1_sel_142983_comb[15]}}, p1_sel_142983_comb} + {{1{p1_smul_142984_comb[15]}}, p1_smul_142984_comb};
  assign p1_add_143845_comb = {{1{p1_smul_142985_comb[15]}}, p1_smul_142985_comb} + {{1{p1_sel_142986_comb[15]}}, p1_sel_142986_comb};
  assign p1_add_143846_comb = {{1{p1_smul_142987_comb[15]}}, p1_smul_142987_comb} + {{1{p1_sel_142988_comb[15]}}, p1_sel_142988_comb};
  assign p1_add_143847_comb = {{1{p1_sel_142989_comb[15]}}, p1_sel_142989_comb} + {{1{p1_smul_142990_comb[15]}}, p1_smul_142990_comb};
  assign p1_add_143848_comb = {{1{p1_sel_142991_comb[15]}}, p1_sel_142991_comb} + {{1{p1_smul_142992_comb[15]}}, p1_smul_142992_comb};
  assign p1_add_143849_comb = {{1{p1_smul_142993_comb[15]}}, p1_smul_142993_comb} + {{1{p1_sel_142994_comb[15]}}, p1_sel_142994_comb};
  assign p1_add_143850_comb = {{1{p1_smul_142995_comb[15]}}, p1_smul_142995_comb} + {{1{p1_sel_142996_comb[15]}}, p1_sel_142996_comb};
  assign p1_add_143851_comb = {{1{p1_sel_142997_comb[15]}}, p1_sel_142997_comb} + {{1{p1_smul_142998_comb[15]}}, p1_smul_142998_comb};
  assign p1_add_143852_comb = {{1{p1_sel_142999_comb[15]}}, p1_sel_142999_comb} + {{1{p1_smul_143000_comb[15]}}, p1_smul_143000_comb};
  assign p1_add_143853_comb = {{1{p1_smul_143001_comb[15]}}, p1_smul_143001_comb} + {{1{p1_sel_143002_comb[15]}}, p1_sel_143002_comb};
  assign p1_add_143854_comb = {{1{p1_smul_143003_comb[15]}}, p1_smul_143003_comb} + {{1{p1_sel_143004_comb[15]}}, p1_sel_143004_comb};
  assign p1_add_143855_comb = {{1{p1_sel_143005_comb[15]}}, p1_sel_143005_comb} + {{1{p1_smul_143006_comb[15]}}, p1_smul_143006_comb};
  assign p1_add_143856_comb = {{1{p1_sel_143007_comb[15]}}, p1_sel_143007_comb} + {{1{p1_smul_143008_comb[15]}}, p1_smul_143008_comb};
  assign p1_add_143857_comb = {{1{p1_smul_143009_comb[15]}}, p1_smul_143009_comb} + {{1{p1_smul_143010_comb[15]}}, p1_smul_143010_comb};
  assign p1_add_143858_comb = {{1{p1_smul_143011_comb[15]}}, p1_smul_143011_comb} + {{1{p1_smul_143012_comb[15]}}, p1_smul_143012_comb};
  assign p1_add_143859_comb = {{1{p1_smul_143013_comb[15]}}, p1_smul_143013_comb} + {{1{p1_smul_143014_comb[15]}}, p1_smul_143014_comb};
  assign p1_add_143860_comb = {{1{p1_smul_143015_comb[15]}}, p1_smul_143015_comb} + {{1{p1_smul_143016_comb[15]}}, p1_smul_143016_comb};
  assign p1_add_143861_comb = {{1{p1_smul_143017_comb[15]}}, p1_smul_143017_comb} + {{1{p1_smul_143018_comb[15]}}, p1_smul_143018_comb};
  assign p1_add_143862_comb = {{1{p1_smul_143019_comb[15]}}, p1_smul_143019_comb} + {{1{p1_smul_143020_comb[15]}}, p1_smul_143020_comb};
  assign p1_add_143863_comb = {{1{p1_smul_143021_comb[15]}}, p1_smul_143021_comb} + {{1{p1_smul_143022_comb[15]}}, p1_smul_143022_comb};
  assign p1_add_143864_comb = {{1{p1_smul_143023_comb[15]}}, p1_smul_143023_comb} + {{1{p1_smul_143024_comb[15]}}, p1_smul_143024_comb};
  assign p1_add_143865_comb = {{1{p1_smul_143025_comb[15]}}, p1_smul_143025_comb} + {{1{p1_smul_143026_comb[15]}}, p1_smul_143026_comb};
  assign p1_add_143866_comb = {{1{p1_smul_143027_comb[15]}}, p1_smul_143027_comb} + {{1{p1_smul_143028_comb[15]}}, p1_smul_143028_comb};
  assign p1_add_143867_comb = {{1{p1_smul_143029_comb[15]}}, p1_smul_143029_comb} + {{1{p1_smul_143030_comb[15]}}, p1_smul_143030_comb};
  assign p1_add_143868_comb = {{1{p1_smul_143031_comb[15]}}, p1_smul_143031_comb} + {{1{p1_smul_143032_comb[15]}}, p1_smul_143032_comb};
  assign p1_add_143869_comb = {{1{p1_smul_143033_comb[15]}}, p1_smul_143033_comb} + {{1{p1_smul_143034_comb[15]}}, p1_smul_143034_comb};
  assign p1_add_143870_comb = {{1{p1_smul_143035_comb[15]}}, p1_smul_143035_comb} + {{1{p1_smul_143036_comb[15]}}, p1_smul_143036_comb};
  assign p1_add_143871_comb = {{1{p1_smul_143037_comb[15]}}, p1_smul_143037_comb} + {{1{p1_smul_143038_comb[15]}}, p1_smul_143038_comb};
  assign p1_add_143872_comb = {{1{p1_smul_143039_comb[15]}}, p1_smul_143039_comb} + {{1{p1_smul_143040_comb[15]}}, p1_smul_143040_comb};
  assign p1_add_143873_comb = {{1{p1_smul_143041_comb[15]}}, p1_smul_143041_comb} + {{1{p1_smul_143042_comb[15]}}, p1_smul_143042_comb};
  assign p1_add_143874_comb = {{1{p1_smul_143043_comb[15]}}, p1_smul_143043_comb} + {{1{p1_smul_143044_comb[15]}}, p1_smul_143044_comb};
  assign p1_add_143875_comb = {{1{p1_smul_143045_comb[15]}}, p1_smul_143045_comb} + {{1{p1_smul_143046_comb[15]}}, p1_smul_143046_comb};
  assign p1_add_143876_comb = {{1{p1_smul_143047_comb[15]}}, p1_smul_143047_comb} + {{1{p1_smul_143048_comb[15]}}, p1_smul_143048_comb};
  assign p1_add_143877_comb = {{1{p1_smul_143049_comb[15]}}, p1_smul_143049_comb} + {{1{p1_smul_143050_comb[15]}}, p1_smul_143050_comb};
  assign p1_add_143878_comb = {{1{p1_smul_143051_comb[15]}}, p1_smul_143051_comb} + {{1{p1_smul_143052_comb[15]}}, p1_smul_143052_comb};
  assign p1_add_143879_comb = {{1{p1_smul_143053_comb[15]}}, p1_smul_143053_comb} + {{1{p1_smul_143054_comb[15]}}, p1_smul_143054_comb};
  assign p1_add_143880_comb = {{1{p1_smul_143055_comb[15]}}, p1_smul_143055_comb} + {{1{p1_smul_143056_comb[15]}}, p1_smul_143056_comb};
  assign p1_add_143881_comb = {{1{p1_smul_143057_comb[15]}}, p1_smul_143057_comb} + {{1{p1_smul_143058_comb[15]}}, p1_smul_143058_comb};
  assign p1_add_143882_comb = {{1{p1_smul_143059_comb[15]}}, p1_smul_143059_comb} + {{1{p1_smul_143060_comb[15]}}, p1_smul_143060_comb};
  assign p1_add_143883_comb = {{1{p1_smul_143061_comb[15]}}, p1_smul_143061_comb} + {{1{p1_smul_143062_comb[15]}}, p1_smul_143062_comb};
  assign p1_add_143884_comb = {{1{p1_smul_143063_comb[15]}}, p1_smul_143063_comb} + {{1{p1_smul_143064_comb[15]}}, p1_smul_143064_comb};
  assign p1_add_143885_comb = {{1{p1_smul_143065_comb[15]}}, p1_smul_143065_comb} + {{1{p1_smul_143066_comb[15]}}, p1_smul_143066_comb};
  assign p1_add_143886_comb = {{1{p1_smul_143067_comb[15]}}, p1_smul_143067_comb} + {{1{p1_smul_143068_comb[15]}}, p1_smul_143068_comb};
  assign p1_add_143887_comb = {{1{p1_smul_143069_comb[15]}}, p1_smul_143069_comb} + {{1{p1_smul_143070_comb[15]}}, p1_smul_143070_comb};
  assign p1_add_143888_comb = {{1{p1_smul_143071_comb[15]}}, p1_smul_143071_comb} + {{1{p1_smul_143072_comb[15]}}, p1_smul_143072_comb};
  assign p1_add_143889_comb = {{1{p1_sel_143073_comb[15]}}, p1_sel_143073_comb} + {{1{p1_smul_143074_comb[15]}}, p1_smul_143074_comb};
  assign p1_add_143890_comb = {{1{p1_sel_143075_comb[15]}}, p1_sel_143075_comb} + {{1{p1_smul_143076_comb[15]}}, p1_smul_143076_comb};
  assign p1_add_143891_comb = {{1{p1_smul_143077_comb[15]}}, p1_smul_143077_comb} + {{1{p1_sel_143078_comb[15]}}, p1_sel_143078_comb};
  assign p1_add_143892_comb = {{1{p1_smul_143079_comb[15]}}, p1_smul_143079_comb} + {{1{p1_sel_143080_comb[15]}}, p1_sel_143080_comb};
  assign p1_add_143893_comb = {{1{p1_sel_143081_comb[15]}}, p1_sel_143081_comb} + {{1{p1_smul_143082_comb[15]}}, p1_smul_143082_comb};
  assign p1_add_143894_comb = {{1{p1_sel_143083_comb[15]}}, p1_sel_143083_comb} + {{1{p1_smul_143084_comb[15]}}, p1_smul_143084_comb};
  assign p1_add_143895_comb = {{1{p1_smul_143085_comb[15]}}, p1_smul_143085_comb} + {{1{p1_sel_143086_comb[15]}}, p1_sel_143086_comb};
  assign p1_add_143896_comb = {{1{p1_smul_143087_comb[15]}}, p1_smul_143087_comb} + {{1{p1_sel_143088_comb[15]}}, p1_sel_143088_comb};
  assign p1_add_143897_comb = {{1{p1_sel_143089_comb[15]}}, p1_sel_143089_comb} + {{1{p1_smul_143090_comb[15]}}, p1_smul_143090_comb};
  assign p1_add_143898_comb = {{1{p1_sel_143091_comb[15]}}, p1_sel_143091_comb} + {{1{p1_smul_143092_comb[15]}}, p1_smul_143092_comb};
  assign p1_add_143899_comb = {{1{p1_smul_143093_comb[15]}}, p1_smul_143093_comb} + {{1{p1_sel_143094_comb[15]}}, p1_sel_143094_comb};
  assign p1_add_143900_comb = {{1{p1_smul_143095_comb[15]}}, p1_smul_143095_comb} + {{1{p1_sel_143096_comb[15]}}, p1_sel_143096_comb};
  assign p1_add_143901_comb = {{1{p1_sel_143097_comb[15]}}, p1_sel_143097_comb} + {{1{p1_smul_143098_comb[15]}}, p1_smul_143098_comb};
  assign p1_add_143902_comb = {{1{p1_sel_143099_comb[15]}}, p1_sel_143099_comb} + {{1{p1_smul_143100_comb[15]}}, p1_smul_143100_comb};
  assign p1_add_143903_comb = {{1{p1_smul_143101_comb[15]}}, p1_smul_143101_comb} + {{1{p1_sel_143102_comb[15]}}, p1_sel_143102_comb};
  assign p1_add_143904_comb = {{1{p1_smul_143103_comb[15]}}, p1_smul_143103_comb} + {{1{p1_sel_143104_comb[15]}}, p1_sel_143104_comb};
  assign p1_add_143905_comb = {{1{p1_sel_143105_comb[15]}}, p1_sel_143105_comb} + {{1{p1_smul_143106_comb[15]}}, p1_smul_143106_comb};
  assign p1_add_143906_comb = {{1{p1_sel_143107_comb[15]}}, p1_sel_143107_comb} + {{1{p1_smul_143108_comb[15]}}, p1_smul_143108_comb};
  assign p1_add_143907_comb = {{1{p1_smul_143109_comb[15]}}, p1_smul_143109_comb} + {{1{p1_sel_143110_comb[15]}}, p1_sel_143110_comb};
  assign p1_add_143908_comb = {{1{p1_smul_143111_comb[15]}}, p1_smul_143111_comb} + {{1{p1_sel_143112_comb[15]}}, p1_sel_143112_comb};
  assign p1_add_143909_comb = {{1{p1_sel_143113_comb[15]}}, p1_sel_143113_comb} + {{1{p1_smul_143114_comb[15]}}, p1_smul_143114_comb};
  assign p1_add_143910_comb = {{1{p1_sel_143115_comb[15]}}, p1_sel_143115_comb} + {{1{p1_smul_143116_comb[15]}}, p1_smul_143116_comb};
  assign p1_add_143911_comb = {{1{p1_smul_143117_comb[15]}}, p1_smul_143117_comb} + {{1{p1_sel_143118_comb[15]}}, p1_sel_143118_comb};
  assign p1_add_143912_comb = {{1{p1_smul_143119_comb[15]}}, p1_smul_143119_comb} + {{1{p1_sel_143120_comb[15]}}, p1_sel_143120_comb};
  assign p1_add_143913_comb = {{1{p1_sel_143121_comb[15]}}, p1_sel_143121_comb} + {{1{p1_smul_143122_comb[15]}}, p1_smul_143122_comb};
  assign p1_add_143914_comb = {{1{p1_sel_143123_comb[15]}}, p1_sel_143123_comb} + {{1{p1_smul_143124_comb[15]}}, p1_smul_143124_comb};
  assign p1_add_143915_comb = {{1{p1_smul_143125_comb[15]}}, p1_smul_143125_comb} + {{1{p1_sel_143126_comb[15]}}, p1_sel_143126_comb};
  assign p1_add_143916_comb = {{1{p1_smul_143127_comb[15]}}, p1_smul_143127_comb} + {{1{p1_sel_143128_comb[15]}}, p1_sel_143128_comb};
  assign p1_add_143917_comb = {{1{p1_sel_143129_comb[15]}}, p1_sel_143129_comb} + {{1{p1_smul_143130_comb[15]}}, p1_smul_143130_comb};
  assign p1_add_143918_comb = {{1{p1_sel_143131_comb[15]}}, p1_sel_143131_comb} + {{1{p1_smul_143132_comb[15]}}, p1_smul_143132_comb};
  assign p1_add_143919_comb = {{1{p1_smul_143133_comb[15]}}, p1_smul_143133_comb} + {{1{p1_sel_143134_comb[15]}}, p1_sel_143134_comb};
  assign p1_add_143920_comb = {{1{p1_smul_143135_comb[15]}}, p1_smul_143135_comb} + {{1{p1_sel_143136_comb[15]}}, p1_sel_143136_comb};
  assign p1_add_143921_comb = {{1{p1_sel_143137_comb[15]}}, p1_sel_143137_comb} + {{1{p1_sel_143138_comb[15]}}, p1_sel_143138_comb};
  assign p1_add_143922_comb = {{1{p1_sel_143139_comb[15]}}, p1_sel_143139_comb} + {{1{p1_sel_143140_comb[15]}}, p1_sel_143140_comb};
  assign p1_add_143923_comb = {{1{p1_sel_143141_comb[15]}}, p1_sel_143141_comb} + {{1{p1_sel_143142_comb[15]}}, p1_sel_143142_comb};
  assign p1_add_143924_comb = {{1{p1_sel_143143_comb[15]}}, p1_sel_143143_comb} + {{1{p1_sel_143144_comb[15]}}, p1_sel_143144_comb};
  assign p1_add_143925_comb = {{1{p1_sel_143145_comb[15]}}, p1_sel_143145_comb} + {{1{p1_sel_143146_comb[15]}}, p1_sel_143146_comb};
  assign p1_add_143926_comb = {{1{p1_sel_143147_comb[15]}}, p1_sel_143147_comb} + {{1{p1_sel_143148_comb[15]}}, p1_sel_143148_comb};
  assign p1_add_143927_comb = {{1{p1_sel_143149_comb[15]}}, p1_sel_143149_comb} + {{1{p1_sel_143150_comb[15]}}, p1_sel_143150_comb};
  assign p1_add_143928_comb = {{1{p1_sel_143151_comb[15]}}, p1_sel_143151_comb} + {{1{p1_sel_143152_comb[15]}}, p1_sel_143152_comb};
  assign p1_add_143929_comb = {{1{p1_sel_143153_comb[15]}}, p1_sel_143153_comb} + {{1{p1_sel_143154_comb[15]}}, p1_sel_143154_comb};
  assign p1_add_143930_comb = {{1{p1_sel_143155_comb[15]}}, p1_sel_143155_comb} + {{1{p1_sel_143156_comb[15]}}, p1_sel_143156_comb};
  assign p1_add_143931_comb = {{1{p1_sel_143157_comb[15]}}, p1_sel_143157_comb} + {{1{p1_sel_143158_comb[15]}}, p1_sel_143158_comb};
  assign p1_add_143932_comb = {{1{p1_sel_143159_comb[15]}}, p1_sel_143159_comb} + {{1{p1_sel_143160_comb[15]}}, p1_sel_143160_comb};
  assign p1_add_143933_comb = {{1{p1_sel_143161_comb[15]}}, p1_sel_143161_comb} + {{1{p1_sel_143162_comb[15]}}, p1_sel_143162_comb};
  assign p1_add_143934_comb = {{1{p1_sel_143163_comb[15]}}, p1_sel_143163_comb} + {{1{p1_sel_143164_comb[15]}}, p1_sel_143164_comb};
  assign p1_add_143935_comb = {{1{p1_sel_143165_comb[15]}}, p1_sel_143165_comb} + {{1{p1_sel_143166_comb[15]}}, p1_sel_143166_comb};
  assign p1_add_143936_comb = {{1{p1_sel_143167_comb[15]}}, p1_sel_143167_comb} + {{1{p1_sel_143168_comb[15]}}, p1_sel_143168_comb};
  assign p1_add_143937_comb = {{1{p1_sel_143169_comb[15]}}, p1_sel_143169_comb} + {{1{p1_sel_143170_comb[15]}}, p1_sel_143170_comb};
  assign p1_add_143938_comb = {{1{p1_sel_143171_comb[15]}}, p1_sel_143171_comb} + {{1{p1_sel_143172_comb[15]}}, p1_sel_143172_comb};
  assign p1_add_143939_comb = {{1{p1_sel_143173_comb[15]}}, p1_sel_143173_comb} + {{1{p1_sel_143174_comb[15]}}, p1_sel_143174_comb};
  assign p1_add_143940_comb = {{1{p1_sel_143175_comb[15]}}, p1_sel_143175_comb} + {{1{p1_sel_143176_comb[15]}}, p1_sel_143176_comb};
  assign p1_add_143941_comb = {{1{p1_sel_143177_comb[15]}}, p1_sel_143177_comb} + {{1{p1_sel_143178_comb[15]}}, p1_sel_143178_comb};
  assign p1_add_143942_comb = {{1{p1_sel_143179_comb[15]}}, p1_sel_143179_comb} + {{1{p1_sel_143180_comb[15]}}, p1_sel_143180_comb};
  assign p1_add_143943_comb = {{1{p1_sel_143181_comb[15]}}, p1_sel_143181_comb} + {{1{p1_sel_143182_comb[15]}}, p1_sel_143182_comb};
  assign p1_add_143944_comb = {{1{p1_sel_143183_comb[15]}}, p1_sel_143183_comb} + {{1{p1_sel_143184_comb[15]}}, p1_sel_143184_comb};
  assign p1_add_143945_comb = {{1{p1_sel_143185_comb[15]}}, p1_sel_143185_comb} + {{1{p1_sel_143186_comb[15]}}, p1_sel_143186_comb};
  assign p1_add_143946_comb = {{1{p1_sel_143187_comb[15]}}, p1_sel_143187_comb} + {{1{p1_sel_143188_comb[15]}}, p1_sel_143188_comb};
  assign p1_add_143947_comb = {{1{p1_sel_143189_comb[15]}}, p1_sel_143189_comb} + {{1{p1_sel_143190_comb[15]}}, p1_sel_143190_comb};
  assign p1_add_143948_comb = {{1{p1_sel_143191_comb[15]}}, p1_sel_143191_comb} + {{1{p1_sel_143192_comb[15]}}, p1_sel_143192_comb};
  assign p1_add_143949_comb = {{1{p1_sel_143193_comb[15]}}, p1_sel_143193_comb} + {{1{p1_sel_143194_comb[15]}}, p1_sel_143194_comb};
  assign p1_add_143950_comb = {{1{p1_sel_143195_comb[15]}}, p1_sel_143195_comb} + {{1{p1_sel_143196_comb[15]}}, p1_sel_143196_comb};
  assign p1_add_143951_comb = {{1{p1_sel_143197_comb[15]}}, p1_sel_143197_comb} + {{1{p1_sel_143198_comb[15]}}, p1_sel_143198_comb};
  assign p1_add_143952_comb = {{1{p1_sel_143199_comb[15]}}, p1_sel_143199_comb} + {{1{p1_sel_143200_comb[15]}}, p1_sel_143200_comb};
  assign p1_add_143953_comb = {{1{p1_sel_143201_comb[15]}}, p1_sel_143201_comb} + {{1{p1_sel_143202_comb[15]}}, p1_sel_143202_comb};
  assign p1_add_143954_comb = {{1{p1_smul_143203_comb[15]}}, p1_smul_143203_comb} + {{1{p1_smul_143204_comb[15]}}, p1_smul_143204_comb};
  assign p1_add_143955_comb = {{1{p1_smul_143205_comb[15]}}, p1_smul_143205_comb} + {{1{p1_smul_143206_comb[15]}}, p1_smul_143206_comb};
  assign p1_add_143956_comb = {{1{p1_sel_143207_comb[15]}}, p1_sel_143207_comb} + {{1{p1_sel_143208_comb[15]}}, p1_sel_143208_comb};
  assign p1_add_143957_comb = {{1{p1_sel_143209_comb[15]}}, p1_sel_143209_comb} + {{1{p1_sel_143210_comb[15]}}, p1_sel_143210_comb};
  assign p1_add_143958_comb = {{1{p1_smul_143211_comb[15]}}, p1_smul_143211_comb} + {{1{p1_smul_143212_comb[15]}}, p1_smul_143212_comb};
  assign p1_add_143959_comb = {{1{p1_smul_143213_comb[15]}}, p1_smul_143213_comb} + {{1{p1_smul_143214_comb[15]}}, p1_smul_143214_comb};
  assign p1_add_143960_comb = {{1{p1_sel_143215_comb[15]}}, p1_sel_143215_comb} + {{1{p1_sel_143216_comb[15]}}, p1_sel_143216_comb};
  assign p1_add_143961_comb = {{1{p1_sel_143217_comb[15]}}, p1_sel_143217_comb} + {{1{p1_sel_143218_comb[15]}}, p1_sel_143218_comb};
  assign p1_add_143962_comb = {{1{p1_smul_143219_comb[15]}}, p1_smul_143219_comb} + {{1{p1_smul_143220_comb[15]}}, p1_smul_143220_comb};
  assign p1_add_143963_comb = {{1{p1_smul_143221_comb[15]}}, p1_smul_143221_comb} + {{1{p1_smul_143222_comb[15]}}, p1_smul_143222_comb};
  assign p1_add_143964_comb = {{1{p1_sel_143223_comb[15]}}, p1_sel_143223_comb} + {{1{p1_sel_143224_comb[15]}}, p1_sel_143224_comb};
  assign p1_add_143965_comb = {{1{p1_sel_143225_comb[15]}}, p1_sel_143225_comb} + {{1{p1_sel_143226_comb[15]}}, p1_sel_143226_comb};
  assign p1_add_143966_comb = {{1{p1_smul_143227_comb[15]}}, p1_smul_143227_comb} + {{1{p1_smul_143228_comb[15]}}, p1_smul_143228_comb};
  assign p1_add_143967_comb = {{1{p1_smul_143229_comb[15]}}, p1_smul_143229_comb} + {{1{p1_smul_143230_comb[15]}}, p1_smul_143230_comb};
  assign p1_add_143968_comb = {{1{p1_sel_143231_comb[15]}}, p1_sel_143231_comb} + {{1{p1_sel_143232_comb[15]}}, p1_sel_143232_comb};
  assign p1_add_143969_comb = {{1{p1_sel_143233_comb[15]}}, p1_sel_143233_comb} + {{1{p1_sel_143234_comb[15]}}, p1_sel_143234_comb};
  assign p1_add_143970_comb = {{1{p1_smul_143235_comb[15]}}, p1_smul_143235_comb} + {{1{p1_smul_143236_comb[15]}}, p1_smul_143236_comb};
  assign p1_add_143971_comb = {{1{p1_smul_143237_comb[15]}}, p1_smul_143237_comb} + {{1{p1_smul_143238_comb[15]}}, p1_smul_143238_comb};
  assign p1_add_143972_comb = {{1{p1_sel_143239_comb[15]}}, p1_sel_143239_comb} + {{1{p1_sel_143240_comb[15]}}, p1_sel_143240_comb};
  assign p1_add_143973_comb = {{1{p1_sel_143241_comb[15]}}, p1_sel_143241_comb} + {{1{p1_sel_143242_comb[15]}}, p1_sel_143242_comb};
  assign p1_add_143974_comb = {{1{p1_smul_143243_comb[15]}}, p1_smul_143243_comb} + {{1{p1_smul_143244_comb[15]}}, p1_smul_143244_comb};
  assign p1_add_143975_comb = {{1{p1_smul_143245_comb[15]}}, p1_smul_143245_comb} + {{1{p1_smul_143246_comb[15]}}, p1_smul_143246_comb};
  assign p1_add_143976_comb = {{1{p1_sel_143247_comb[15]}}, p1_sel_143247_comb} + {{1{p1_sel_143248_comb[15]}}, p1_sel_143248_comb};
  assign p1_add_143977_comb = {{1{p1_sel_143249_comb[15]}}, p1_sel_143249_comb} + {{1{p1_sel_143250_comb[15]}}, p1_sel_143250_comb};
  assign p1_add_143978_comb = {{1{p1_smul_143251_comb[15]}}, p1_smul_143251_comb} + {{1{p1_smul_143252_comb[15]}}, p1_smul_143252_comb};
  assign p1_add_143979_comb = {{1{p1_smul_143253_comb[15]}}, p1_smul_143253_comb} + {{1{p1_smul_143254_comb[15]}}, p1_smul_143254_comb};
  assign p1_add_143980_comb = {{1{p1_sel_143255_comb[15]}}, p1_sel_143255_comb} + {{1{p1_sel_143256_comb[15]}}, p1_sel_143256_comb};
  assign p1_add_143981_comb = {{1{p1_sel_143257_comb[15]}}, p1_sel_143257_comb} + {{1{p1_sel_143258_comb[15]}}, p1_sel_143258_comb};
  assign p1_add_143982_comb = {{1{p1_smul_143259_comb[15]}}, p1_smul_143259_comb} + {{1{p1_smul_143260_comb[15]}}, p1_smul_143260_comb};
  assign p1_add_143983_comb = {{1{p1_smul_143261_comb[15]}}, p1_smul_143261_comb} + {{1{p1_smul_143262_comb[15]}}, p1_smul_143262_comb};
  assign p1_add_143984_comb = {{1{p1_sel_143263_comb[15]}}, p1_sel_143263_comb} + {{1{p1_sel_143264_comb[15]}}, p1_sel_143264_comb};
  assign p1_sum__526_comb = p1_sum__524_comb + p1_sum__525_comb;
  assign p1_sum__470_comb = p1_sum__468_comb + p1_sum__469_comb;
  assign p1_sum__414_comb = p1_sum__412_comb + p1_sum__413_comb;
  assign p1_sum__358_comb = p1_sum__356_comb + p1_sum__357_comb;
  assign p1_sum__302_comb = p1_sum__300_comb + p1_sum__301_comb;
  assign p1_sum__246_comb = p1_sum__244_comb + p1_sum__245_comb;
  assign p1_sum__190_comb = p1_sum__188_comb + p1_sum__189_comb;
  assign p1_sum__134_comb = p1_sum__132_comb + p1_sum__133_comb;
  assign p1_sum__1580_comb = {{8{p1_add_143761_comb[16]}}, p1_add_143761_comb};
  assign p1_sum__1581_comb = {{8{p1_add_143762_comb[16]}}, p1_add_143762_comb};
  assign p1_sum__1582_comb = {{8{p1_add_143763_comb[16]}}, p1_add_143763_comb};
  assign p1_sum__1583_comb = {{8{p1_add_143764_comb[16]}}, p1_add_143764_comb};
  assign p1_sum__1552_comb = {{8{p1_add_143765_comb[16]}}, p1_add_143765_comb};
  assign p1_sum__1553_comb = {{8{p1_add_143766_comb[16]}}, p1_add_143766_comb};
  assign p1_sum__1554_comb = {{8{p1_add_143767_comb[16]}}, p1_add_143767_comb};
  assign p1_sum__1555_comb = {{8{p1_add_143768_comb[16]}}, p1_add_143768_comb};
  assign p1_sum__1524_comb = {{8{p1_add_143769_comb[16]}}, p1_add_143769_comb};
  assign p1_sum__1525_comb = {{8{p1_add_143770_comb[16]}}, p1_add_143770_comb};
  assign p1_sum__1526_comb = {{8{p1_add_143771_comb[16]}}, p1_add_143771_comb};
  assign p1_sum__1527_comb = {{8{p1_add_143772_comb[16]}}, p1_add_143772_comb};
  assign p1_sum__1496_comb = {{8{p1_add_143773_comb[16]}}, p1_add_143773_comb};
  assign p1_sum__1497_comb = {{8{p1_add_143774_comb[16]}}, p1_add_143774_comb};
  assign p1_sum__1498_comb = {{8{p1_add_143775_comb[16]}}, p1_add_143775_comb};
  assign p1_sum__1499_comb = {{8{p1_add_143776_comb[16]}}, p1_add_143776_comb};
  assign p1_sum__1468_comb = {{8{p1_add_143777_comb[16]}}, p1_add_143777_comb};
  assign p1_sum__1469_comb = {{8{p1_add_143778_comb[16]}}, p1_add_143778_comb};
  assign p1_sum__1470_comb = {{8{p1_add_143779_comb[16]}}, p1_add_143779_comb};
  assign p1_sum__1471_comb = {{8{p1_add_143780_comb[16]}}, p1_add_143780_comb};
  assign p1_sum__1440_comb = {{8{p1_add_143781_comb[16]}}, p1_add_143781_comb};
  assign p1_sum__1441_comb = {{8{p1_add_143782_comb[16]}}, p1_add_143782_comb};
  assign p1_sum__1442_comb = {{8{p1_add_143783_comb[16]}}, p1_add_143783_comb};
  assign p1_sum__1443_comb = {{8{p1_add_143784_comb[16]}}, p1_add_143784_comb};
  assign p1_sum__1412_comb = {{8{p1_add_143785_comb[16]}}, p1_add_143785_comb};
  assign p1_sum__1413_comb = {{8{p1_add_143786_comb[16]}}, p1_add_143786_comb};
  assign p1_sum__1414_comb = {{8{p1_add_143787_comb[16]}}, p1_add_143787_comb};
  assign p1_sum__1415_comb = {{8{p1_add_143788_comb[16]}}, p1_add_143788_comb};
  assign p1_sum__1384_comb = {{8{p1_add_143789_comb[16]}}, p1_add_143789_comb};
  assign p1_sum__1385_comb = {{8{p1_add_143790_comb[16]}}, p1_add_143790_comb};
  assign p1_sum__1386_comb = {{8{p1_add_143791_comb[16]}}, p1_add_143791_comb};
  assign p1_sum__1387_comb = {{8{p1_add_143792_comb[16]}}, p1_add_143792_comb};
  assign p1_sum__1576_comb = {{8{p1_add_143793_comb[16]}}, p1_add_143793_comb};
  assign p1_sum__1577_comb = {{8{p1_add_143794_comb[16]}}, p1_add_143794_comb};
  assign p1_sum__1578_comb = {{8{p1_add_143795_comb[16]}}, p1_add_143795_comb};
  assign p1_sum__1579_comb = {{8{p1_add_143796_comb[16]}}, p1_add_143796_comb};
  assign p1_sum__1548_comb = {{8{p1_add_143797_comb[16]}}, p1_add_143797_comb};
  assign p1_sum__1549_comb = {{8{p1_add_143798_comb[16]}}, p1_add_143798_comb};
  assign p1_sum__1550_comb = {{8{p1_add_143799_comb[16]}}, p1_add_143799_comb};
  assign p1_sum__1551_comb = {{8{p1_add_143800_comb[16]}}, p1_add_143800_comb};
  assign p1_sum__1520_comb = {{8{p1_add_143801_comb[16]}}, p1_add_143801_comb};
  assign p1_sum__1521_comb = {{8{p1_add_143802_comb[16]}}, p1_add_143802_comb};
  assign p1_sum__1522_comb = {{8{p1_add_143803_comb[16]}}, p1_add_143803_comb};
  assign p1_sum__1523_comb = {{8{p1_add_143804_comb[16]}}, p1_add_143804_comb};
  assign p1_sum__1492_comb = {{8{p1_add_143805_comb[16]}}, p1_add_143805_comb};
  assign p1_sum__1493_comb = {{8{p1_add_143806_comb[16]}}, p1_add_143806_comb};
  assign p1_sum__1494_comb = {{8{p1_add_143807_comb[16]}}, p1_add_143807_comb};
  assign p1_sum__1495_comb = {{8{p1_add_143808_comb[16]}}, p1_add_143808_comb};
  assign p1_sum__1464_comb = {{8{p1_add_143809_comb[16]}}, p1_add_143809_comb};
  assign p1_sum__1465_comb = {{8{p1_add_143810_comb[16]}}, p1_add_143810_comb};
  assign p1_sum__1466_comb = {{8{p1_add_143811_comb[16]}}, p1_add_143811_comb};
  assign p1_sum__1467_comb = {{8{p1_add_143812_comb[16]}}, p1_add_143812_comb};
  assign p1_sum__1436_comb = {{8{p1_add_143813_comb[16]}}, p1_add_143813_comb};
  assign p1_sum__1437_comb = {{8{p1_add_143814_comb[16]}}, p1_add_143814_comb};
  assign p1_sum__1438_comb = {{8{p1_add_143815_comb[16]}}, p1_add_143815_comb};
  assign p1_sum__1439_comb = {{8{p1_add_143816_comb[16]}}, p1_add_143816_comb};
  assign p1_sum__1408_comb = {{8{p1_add_143817_comb[16]}}, p1_add_143817_comb};
  assign p1_sum__1409_comb = {{8{p1_add_143818_comb[16]}}, p1_add_143818_comb};
  assign p1_sum__1410_comb = {{8{p1_add_143819_comb[16]}}, p1_add_143819_comb};
  assign p1_sum__1411_comb = {{8{p1_add_143820_comb[16]}}, p1_add_143820_comb};
  assign p1_sum__1380_comb = {{8{p1_add_143821_comb[16]}}, p1_add_143821_comb};
  assign p1_sum__1381_comb = {{8{p1_add_143822_comb[16]}}, p1_add_143822_comb};
  assign p1_sum__1382_comb = {{8{p1_add_143823_comb[16]}}, p1_add_143823_comb};
  assign p1_sum__1383_comb = {{8{p1_add_143824_comb[16]}}, p1_add_143824_comb};
  assign p1_sum__1572_comb = {{8{p1_add_143825_comb[16]}}, p1_add_143825_comb};
  assign p1_sum__1573_comb = {{8{p1_add_143826_comb[16]}}, p1_add_143826_comb};
  assign p1_sum__1574_comb = {{8{p1_add_143827_comb[16]}}, p1_add_143827_comb};
  assign p1_sum__1575_comb = {{8{p1_add_143828_comb[16]}}, p1_add_143828_comb};
  assign p1_sum__1544_comb = {{8{p1_add_143829_comb[16]}}, p1_add_143829_comb};
  assign p1_sum__1545_comb = {{8{p1_add_143830_comb[16]}}, p1_add_143830_comb};
  assign p1_sum__1546_comb = {{8{p1_add_143831_comb[16]}}, p1_add_143831_comb};
  assign p1_sum__1547_comb = {{8{p1_add_143832_comb[16]}}, p1_add_143832_comb};
  assign p1_sum__1516_comb = {{8{p1_add_143833_comb[16]}}, p1_add_143833_comb};
  assign p1_sum__1517_comb = {{8{p1_add_143834_comb[16]}}, p1_add_143834_comb};
  assign p1_sum__1518_comb = {{8{p1_add_143835_comb[16]}}, p1_add_143835_comb};
  assign p1_sum__1519_comb = {{8{p1_add_143836_comb[16]}}, p1_add_143836_comb};
  assign p1_sum__1488_comb = {{8{p1_add_143837_comb[16]}}, p1_add_143837_comb};
  assign p1_sum__1489_comb = {{8{p1_add_143838_comb[16]}}, p1_add_143838_comb};
  assign p1_sum__1490_comb = {{8{p1_add_143839_comb[16]}}, p1_add_143839_comb};
  assign p1_sum__1491_comb = {{8{p1_add_143840_comb[16]}}, p1_add_143840_comb};
  assign p1_sum__1460_comb = {{8{p1_add_143841_comb[16]}}, p1_add_143841_comb};
  assign p1_sum__1461_comb = {{8{p1_add_143842_comb[16]}}, p1_add_143842_comb};
  assign p1_sum__1462_comb = {{8{p1_add_143843_comb[16]}}, p1_add_143843_comb};
  assign p1_sum__1463_comb = {{8{p1_add_143844_comb[16]}}, p1_add_143844_comb};
  assign p1_sum__1432_comb = {{8{p1_add_143845_comb[16]}}, p1_add_143845_comb};
  assign p1_sum__1433_comb = {{8{p1_add_143846_comb[16]}}, p1_add_143846_comb};
  assign p1_sum__1434_comb = {{8{p1_add_143847_comb[16]}}, p1_add_143847_comb};
  assign p1_sum__1435_comb = {{8{p1_add_143848_comb[16]}}, p1_add_143848_comb};
  assign p1_sum__1404_comb = {{8{p1_add_143849_comb[16]}}, p1_add_143849_comb};
  assign p1_sum__1405_comb = {{8{p1_add_143850_comb[16]}}, p1_add_143850_comb};
  assign p1_sum__1406_comb = {{8{p1_add_143851_comb[16]}}, p1_add_143851_comb};
  assign p1_sum__1407_comb = {{8{p1_add_143852_comb[16]}}, p1_add_143852_comb};
  assign p1_sum__1376_comb = {{8{p1_add_143853_comb[16]}}, p1_add_143853_comb};
  assign p1_sum__1377_comb = {{8{p1_add_143854_comb[16]}}, p1_add_143854_comb};
  assign p1_sum__1378_comb = {{8{p1_add_143855_comb[16]}}, p1_add_143855_comb};
  assign p1_sum__1379_comb = {{8{p1_add_143856_comb[16]}}, p1_add_143856_comb};
  assign p1_sum__1568_comb = {{8{p1_add_143857_comb[16]}}, p1_add_143857_comb};
  assign p1_sum__1569_comb = {{8{p1_add_143858_comb[16]}}, p1_add_143858_comb};
  assign p1_sum__1570_comb = {{8{p1_add_143859_comb[16]}}, p1_add_143859_comb};
  assign p1_sum__1571_comb = {{8{p1_add_143860_comb[16]}}, p1_add_143860_comb};
  assign p1_sum__1540_comb = {{8{p1_add_143861_comb[16]}}, p1_add_143861_comb};
  assign p1_sum__1541_comb = {{8{p1_add_143862_comb[16]}}, p1_add_143862_comb};
  assign p1_sum__1542_comb = {{8{p1_add_143863_comb[16]}}, p1_add_143863_comb};
  assign p1_sum__1543_comb = {{8{p1_add_143864_comb[16]}}, p1_add_143864_comb};
  assign p1_sum__1512_comb = {{8{p1_add_143865_comb[16]}}, p1_add_143865_comb};
  assign p1_sum__1513_comb = {{8{p1_add_143866_comb[16]}}, p1_add_143866_comb};
  assign p1_sum__1514_comb = {{8{p1_add_143867_comb[16]}}, p1_add_143867_comb};
  assign p1_sum__1515_comb = {{8{p1_add_143868_comb[16]}}, p1_add_143868_comb};
  assign p1_sum__1484_comb = {{8{p1_add_143869_comb[16]}}, p1_add_143869_comb};
  assign p1_sum__1485_comb = {{8{p1_add_143870_comb[16]}}, p1_add_143870_comb};
  assign p1_sum__1486_comb = {{8{p1_add_143871_comb[16]}}, p1_add_143871_comb};
  assign p1_sum__1487_comb = {{8{p1_add_143872_comb[16]}}, p1_add_143872_comb};
  assign p1_sum__1456_comb = {{8{p1_add_143873_comb[16]}}, p1_add_143873_comb};
  assign p1_sum__1457_comb = {{8{p1_add_143874_comb[16]}}, p1_add_143874_comb};
  assign p1_sum__1458_comb = {{8{p1_add_143875_comb[16]}}, p1_add_143875_comb};
  assign p1_sum__1459_comb = {{8{p1_add_143876_comb[16]}}, p1_add_143876_comb};
  assign p1_sum__1428_comb = {{8{p1_add_143877_comb[16]}}, p1_add_143877_comb};
  assign p1_sum__1429_comb = {{8{p1_add_143878_comb[16]}}, p1_add_143878_comb};
  assign p1_sum__1430_comb = {{8{p1_add_143879_comb[16]}}, p1_add_143879_comb};
  assign p1_sum__1431_comb = {{8{p1_add_143880_comb[16]}}, p1_add_143880_comb};
  assign p1_sum__1400_comb = {{8{p1_add_143881_comb[16]}}, p1_add_143881_comb};
  assign p1_sum__1401_comb = {{8{p1_add_143882_comb[16]}}, p1_add_143882_comb};
  assign p1_sum__1402_comb = {{8{p1_add_143883_comb[16]}}, p1_add_143883_comb};
  assign p1_sum__1403_comb = {{8{p1_add_143884_comb[16]}}, p1_add_143884_comb};
  assign p1_sum__1372_comb = {{8{p1_add_143885_comb[16]}}, p1_add_143885_comb};
  assign p1_sum__1373_comb = {{8{p1_add_143886_comb[16]}}, p1_add_143886_comb};
  assign p1_sum__1374_comb = {{8{p1_add_143887_comb[16]}}, p1_add_143887_comb};
  assign p1_sum__1375_comb = {{8{p1_add_143888_comb[16]}}, p1_add_143888_comb};
  assign p1_sum__1564_comb = {{8{p1_add_143889_comb[16]}}, p1_add_143889_comb};
  assign p1_sum__1565_comb = {{8{p1_add_143890_comb[16]}}, p1_add_143890_comb};
  assign p1_sum__1566_comb = {{8{p1_add_143891_comb[16]}}, p1_add_143891_comb};
  assign p1_sum__1567_comb = {{8{p1_add_143892_comb[16]}}, p1_add_143892_comb};
  assign p1_sum__1536_comb = {{8{p1_add_143893_comb[16]}}, p1_add_143893_comb};
  assign p1_sum__1537_comb = {{8{p1_add_143894_comb[16]}}, p1_add_143894_comb};
  assign p1_sum__1538_comb = {{8{p1_add_143895_comb[16]}}, p1_add_143895_comb};
  assign p1_sum__1539_comb = {{8{p1_add_143896_comb[16]}}, p1_add_143896_comb};
  assign p1_sum__1508_comb = {{8{p1_add_143897_comb[16]}}, p1_add_143897_comb};
  assign p1_sum__1509_comb = {{8{p1_add_143898_comb[16]}}, p1_add_143898_comb};
  assign p1_sum__1510_comb = {{8{p1_add_143899_comb[16]}}, p1_add_143899_comb};
  assign p1_sum__1511_comb = {{8{p1_add_143900_comb[16]}}, p1_add_143900_comb};
  assign p1_sum__1480_comb = {{8{p1_add_143901_comb[16]}}, p1_add_143901_comb};
  assign p1_sum__1481_comb = {{8{p1_add_143902_comb[16]}}, p1_add_143902_comb};
  assign p1_sum__1482_comb = {{8{p1_add_143903_comb[16]}}, p1_add_143903_comb};
  assign p1_sum__1483_comb = {{8{p1_add_143904_comb[16]}}, p1_add_143904_comb};
  assign p1_sum__1452_comb = {{8{p1_add_143905_comb[16]}}, p1_add_143905_comb};
  assign p1_sum__1453_comb = {{8{p1_add_143906_comb[16]}}, p1_add_143906_comb};
  assign p1_sum__1454_comb = {{8{p1_add_143907_comb[16]}}, p1_add_143907_comb};
  assign p1_sum__1455_comb = {{8{p1_add_143908_comb[16]}}, p1_add_143908_comb};
  assign p1_sum__1424_comb = {{8{p1_add_143909_comb[16]}}, p1_add_143909_comb};
  assign p1_sum__1425_comb = {{8{p1_add_143910_comb[16]}}, p1_add_143910_comb};
  assign p1_sum__1426_comb = {{8{p1_add_143911_comb[16]}}, p1_add_143911_comb};
  assign p1_sum__1427_comb = {{8{p1_add_143912_comb[16]}}, p1_add_143912_comb};
  assign p1_sum__1396_comb = {{8{p1_add_143913_comb[16]}}, p1_add_143913_comb};
  assign p1_sum__1397_comb = {{8{p1_add_143914_comb[16]}}, p1_add_143914_comb};
  assign p1_sum__1398_comb = {{8{p1_add_143915_comb[16]}}, p1_add_143915_comb};
  assign p1_sum__1399_comb = {{8{p1_add_143916_comb[16]}}, p1_add_143916_comb};
  assign p1_sum__1368_comb = {{8{p1_add_143917_comb[16]}}, p1_add_143917_comb};
  assign p1_sum__1369_comb = {{8{p1_add_143918_comb[16]}}, p1_add_143918_comb};
  assign p1_sum__1370_comb = {{8{p1_add_143919_comb[16]}}, p1_add_143919_comb};
  assign p1_sum__1371_comb = {{8{p1_add_143920_comb[16]}}, p1_add_143920_comb};
  assign p1_sum__1560_comb = {{8{p1_add_143921_comb[16]}}, p1_add_143921_comb};
  assign p1_sum__1561_comb = {{8{p1_add_143922_comb[16]}}, p1_add_143922_comb};
  assign p1_sum__1562_comb = {{8{p1_add_143923_comb[16]}}, p1_add_143923_comb};
  assign p1_sum__1563_comb = {{8{p1_add_143924_comb[16]}}, p1_add_143924_comb};
  assign p1_sum__1532_comb = {{8{p1_add_143925_comb[16]}}, p1_add_143925_comb};
  assign p1_sum__1533_comb = {{8{p1_add_143926_comb[16]}}, p1_add_143926_comb};
  assign p1_sum__1534_comb = {{8{p1_add_143927_comb[16]}}, p1_add_143927_comb};
  assign p1_sum__1535_comb = {{8{p1_add_143928_comb[16]}}, p1_add_143928_comb};
  assign p1_sum__1504_comb = {{8{p1_add_143929_comb[16]}}, p1_add_143929_comb};
  assign p1_sum__1505_comb = {{8{p1_add_143930_comb[16]}}, p1_add_143930_comb};
  assign p1_sum__1506_comb = {{8{p1_add_143931_comb[16]}}, p1_add_143931_comb};
  assign p1_sum__1507_comb = {{8{p1_add_143932_comb[16]}}, p1_add_143932_comb};
  assign p1_sum__1476_comb = {{8{p1_add_143933_comb[16]}}, p1_add_143933_comb};
  assign p1_sum__1477_comb = {{8{p1_add_143934_comb[16]}}, p1_add_143934_comb};
  assign p1_sum__1478_comb = {{8{p1_add_143935_comb[16]}}, p1_add_143935_comb};
  assign p1_sum__1479_comb = {{8{p1_add_143936_comb[16]}}, p1_add_143936_comb};
  assign p1_sum__1448_comb = {{8{p1_add_143937_comb[16]}}, p1_add_143937_comb};
  assign p1_sum__1449_comb = {{8{p1_add_143938_comb[16]}}, p1_add_143938_comb};
  assign p1_sum__1450_comb = {{8{p1_add_143939_comb[16]}}, p1_add_143939_comb};
  assign p1_sum__1451_comb = {{8{p1_add_143940_comb[16]}}, p1_add_143940_comb};
  assign p1_sum__1420_comb = {{8{p1_add_143941_comb[16]}}, p1_add_143941_comb};
  assign p1_sum__1421_comb = {{8{p1_add_143942_comb[16]}}, p1_add_143942_comb};
  assign p1_sum__1422_comb = {{8{p1_add_143943_comb[16]}}, p1_add_143943_comb};
  assign p1_sum__1423_comb = {{8{p1_add_143944_comb[16]}}, p1_add_143944_comb};
  assign p1_sum__1392_comb = {{8{p1_add_143945_comb[16]}}, p1_add_143945_comb};
  assign p1_sum__1393_comb = {{8{p1_add_143946_comb[16]}}, p1_add_143946_comb};
  assign p1_sum__1394_comb = {{8{p1_add_143947_comb[16]}}, p1_add_143947_comb};
  assign p1_sum__1395_comb = {{8{p1_add_143948_comb[16]}}, p1_add_143948_comb};
  assign p1_sum__1364_comb = {{8{p1_add_143949_comb[16]}}, p1_add_143949_comb};
  assign p1_sum__1365_comb = {{8{p1_add_143950_comb[16]}}, p1_add_143950_comb};
  assign p1_sum__1366_comb = {{8{p1_add_143951_comb[16]}}, p1_add_143951_comb};
  assign p1_sum__1367_comb = {{8{p1_add_143952_comb[16]}}, p1_add_143952_comb};
  assign p1_sum__1556_comb = {{8{p1_add_143953_comb[16]}}, p1_add_143953_comb};
  assign p1_sum__1557_comb = {{8{p1_add_143954_comb[16]}}, p1_add_143954_comb};
  assign p1_sum__1558_comb = {{8{p1_add_143955_comb[16]}}, p1_add_143955_comb};
  assign p1_sum__1559_comb = {{8{p1_add_143956_comb[16]}}, p1_add_143956_comb};
  assign p1_sum__1528_comb = {{8{p1_add_143957_comb[16]}}, p1_add_143957_comb};
  assign p1_sum__1529_comb = {{8{p1_add_143958_comb[16]}}, p1_add_143958_comb};
  assign p1_sum__1530_comb = {{8{p1_add_143959_comb[16]}}, p1_add_143959_comb};
  assign p1_sum__1531_comb = {{8{p1_add_143960_comb[16]}}, p1_add_143960_comb};
  assign p1_sum__1500_comb = {{8{p1_add_143961_comb[16]}}, p1_add_143961_comb};
  assign p1_sum__1501_comb = {{8{p1_add_143962_comb[16]}}, p1_add_143962_comb};
  assign p1_sum__1502_comb = {{8{p1_add_143963_comb[16]}}, p1_add_143963_comb};
  assign p1_sum__1503_comb = {{8{p1_add_143964_comb[16]}}, p1_add_143964_comb};
  assign p1_sum__1472_comb = {{8{p1_add_143965_comb[16]}}, p1_add_143965_comb};
  assign p1_sum__1473_comb = {{8{p1_add_143966_comb[16]}}, p1_add_143966_comb};
  assign p1_sum__1474_comb = {{8{p1_add_143967_comb[16]}}, p1_add_143967_comb};
  assign p1_sum__1475_comb = {{8{p1_add_143968_comb[16]}}, p1_add_143968_comb};
  assign p1_sum__1444_comb = {{8{p1_add_143969_comb[16]}}, p1_add_143969_comb};
  assign p1_sum__1445_comb = {{8{p1_add_143970_comb[16]}}, p1_add_143970_comb};
  assign p1_sum__1446_comb = {{8{p1_add_143971_comb[16]}}, p1_add_143971_comb};
  assign p1_sum__1447_comb = {{8{p1_add_143972_comb[16]}}, p1_add_143972_comb};
  assign p1_sum__1416_comb = {{8{p1_add_143973_comb[16]}}, p1_add_143973_comb};
  assign p1_sum__1417_comb = {{8{p1_add_143974_comb[16]}}, p1_add_143974_comb};
  assign p1_sum__1418_comb = {{8{p1_add_143975_comb[16]}}, p1_add_143975_comb};
  assign p1_sum__1419_comb = {{8{p1_add_143976_comb[16]}}, p1_add_143976_comb};
  assign p1_sum__1388_comb = {{8{p1_add_143977_comb[16]}}, p1_add_143977_comb};
  assign p1_sum__1389_comb = {{8{p1_add_143978_comb[16]}}, p1_add_143978_comb};
  assign p1_sum__1390_comb = {{8{p1_add_143979_comb[16]}}, p1_add_143979_comb};
  assign p1_sum__1391_comb = {{8{p1_add_143980_comb[16]}}, p1_add_143980_comb};
  assign p1_sum__1360_comb = {{8{p1_add_143981_comb[16]}}, p1_add_143981_comb};
  assign p1_sum__1361_comb = {{8{p1_add_143982_comb[16]}}, p1_add_143982_comb};
  assign p1_sum__1362_comb = {{8{p1_add_143983_comb[16]}}, p1_add_143983_comb};
  assign p1_sum__1363_comb = {{8{p1_add_143984_comb[16]}}, p1_add_143984_comb};
  assign p1_umul_144225_comb = umul32b_32b_x_7b(p1_sum__526_comb, 7'h5b);
  assign p1_umul_144226_comb = umul32b_32b_x_7b(p1_sum__470_comb, 7'h5b);
  assign p1_umul_144227_comb = umul32b_32b_x_7b(p1_sum__414_comb, 7'h5b);
  assign p1_umul_144228_comb = umul32b_32b_x_7b(p1_sum__358_comb, 7'h5b);
  assign p1_umul_144229_comb = umul32b_32b_x_7b(p1_sum__302_comb, 7'h5b);
  assign p1_umul_144230_comb = umul32b_32b_x_7b(p1_sum__246_comb, 7'h5b);
  assign p1_umul_144231_comb = umul32b_32b_x_7b(p1_sum__190_comb, 7'h5b);
  assign p1_umul_144232_comb = umul32b_32b_x_7b(p1_sum__134_comb, 7'h5b);
  assign p1_sum__1246_comb = p1_sum__1580_comb + p1_sum__1581_comb;
  assign p1_sum__1247_comb = p1_sum__1582_comb + p1_sum__1583_comb;
  assign p1_sum__1232_comb = p1_sum__1552_comb + p1_sum__1553_comb;
  assign p1_sum__1233_comb = p1_sum__1554_comb + p1_sum__1555_comb;
  assign p1_sum__1218_comb = p1_sum__1524_comb + p1_sum__1525_comb;
  assign p1_sum__1219_comb = p1_sum__1526_comb + p1_sum__1527_comb;
  assign p1_sum__1204_comb = p1_sum__1496_comb + p1_sum__1497_comb;
  assign p1_sum__1205_comb = p1_sum__1498_comb + p1_sum__1499_comb;
  assign p1_sum__1190_comb = p1_sum__1468_comb + p1_sum__1469_comb;
  assign p1_sum__1191_comb = p1_sum__1470_comb + p1_sum__1471_comb;
  assign p1_sum__1176_comb = p1_sum__1440_comb + p1_sum__1441_comb;
  assign p1_sum__1177_comb = p1_sum__1442_comb + p1_sum__1443_comb;
  assign p1_sum__1162_comb = p1_sum__1412_comb + p1_sum__1413_comb;
  assign p1_sum__1163_comb = p1_sum__1414_comb + p1_sum__1415_comb;
  assign p1_sum__1148_comb = p1_sum__1384_comb + p1_sum__1385_comb;
  assign p1_sum__1149_comb = p1_sum__1386_comb + p1_sum__1387_comb;
  assign p1_sum__1244_comb = p1_sum__1576_comb + p1_sum__1577_comb;
  assign p1_sum__1245_comb = p1_sum__1578_comb + p1_sum__1579_comb;
  assign p1_sum__1230_comb = p1_sum__1548_comb + p1_sum__1549_comb;
  assign p1_sum__1231_comb = p1_sum__1550_comb + p1_sum__1551_comb;
  assign p1_sum__1216_comb = p1_sum__1520_comb + p1_sum__1521_comb;
  assign p1_sum__1217_comb = p1_sum__1522_comb + p1_sum__1523_comb;
  assign p1_sum__1202_comb = p1_sum__1492_comb + p1_sum__1493_comb;
  assign p1_sum__1203_comb = p1_sum__1494_comb + p1_sum__1495_comb;
  assign p1_sum__1188_comb = p1_sum__1464_comb + p1_sum__1465_comb;
  assign p1_sum__1189_comb = p1_sum__1466_comb + p1_sum__1467_comb;
  assign p1_sum__1174_comb = p1_sum__1436_comb + p1_sum__1437_comb;
  assign p1_sum__1175_comb = p1_sum__1438_comb + p1_sum__1439_comb;
  assign p1_sum__1160_comb = p1_sum__1408_comb + p1_sum__1409_comb;
  assign p1_sum__1161_comb = p1_sum__1410_comb + p1_sum__1411_comb;
  assign p1_sum__1146_comb = p1_sum__1380_comb + p1_sum__1381_comb;
  assign p1_sum__1147_comb = p1_sum__1382_comb + p1_sum__1383_comb;
  assign p1_sum__1242_comb = p1_sum__1572_comb + p1_sum__1573_comb;
  assign p1_sum__1243_comb = p1_sum__1574_comb + p1_sum__1575_comb;
  assign p1_sum__1228_comb = p1_sum__1544_comb + p1_sum__1545_comb;
  assign p1_sum__1229_comb = p1_sum__1546_comb + p1_sum__1547_comb;
  assign p1_sum__1214_comb = p1_sum__1516_comb + p1_sum__1517_comb;
  assign p1_sum__1215_comb = p1_sum__1518_comb + p1_sum__1519_comb;
  assign p1_sum__1200_comb = p1_sum__1488_comb + p1_sum__1489_comb;
  assign p1_sum__1201_comb = p1_sum__1490_comb + p1_sum__1491_comb;
  assign p1_sum__1186_comb = p1_sum__1460_comb + p1_sum__1461_comb;
  assign p1_sum__1187_comb = p1_sum__1462_comb + p1_sum__1463_comb;
  assign p1_sum__1172_comb = p1_sum__1432_comb + p1_sum__1433_comb;
  assign p1_sum__1173_comb = p1_sum__1434_comb + p1_sum__1435_comb;
  assign p1_sum__1158_comb = p1_sum__1404_comb + p1_sum__1405_comb;
  assign p1_sum__1159_comb = p1_sum__1406_comb + p1_sum__1407_comb;
  assign p1_sum__1144_comb = p1_sum__1376_comb + p1_sum__1377_comb;
  assign p1_sum__1145_comb = p1_sum__1378_comb + p1_sum__1379_comb;
  assign p1_sum__1240_comb = p1_sum__1568_comb + p1_sum__1569_comb;
  assign p1_sum__1241_comb = p1_sum__1570_comb + p1_sum__1571_comb;
  assign p1_sum__1226_comb = p1_sum__1540_comb + p1_sum__1541_comb;
  assign p1_sum__1227_comb = p1_sum__1542_comb + p1_sum__1543_comb;
  assign p1_sum__1212_comb = p1_sum__1512_comb + p1_sum__1513_comb;
  assign p1_sum__1213_comb = p1_sum__1514_comb + p1_sum__1515_comb;
  assign p1_sum__1198_comb = p1_sum__1484_comb + p1_sum__1485_comb;
  assign p1_sum__1199_comb = p1_sum__1486_comb + p1_sum__1487_comb;
  assign p1_sum__1184_comb = p1_sum__1456_comb + p1_sum__1457_comb;
  assign p1_sum__1185_comb = p1_sum__1458_comb + p1_sum__1459_comb;
  assign p1_sum__1170_comb = p1_sum__1428_comb + p1_sum__1429_comb;
  assign p1_sum__1171_comb = p1_sum__1430_comb + p1_sum__1431_comb;
  assign p1_sum__1156_comb = p1_sum__1400_comb + p1_sum__1401_comb;
  assign p1_sum__1157_comb = p1_sum__1402_comb + p1_sum__1403_comb;
  assign p1_sum__1142_comb = p1_sum__1372_comb + p1_sum__1373_comb;
  assign p1_sum__1143_comb = p1_sum__1374_comb + p1_sum__1375_comb;
  assign p1_sum__1238_comb = p1_sum__1564_comb + p1_sum__1565_comb;
  assign p1_sum__1239_comb = p1_sum__1566_comb + p1_sum__1567_comb;
  assign p1_sum__1224_comb = p1_sum__1536_comb + p1_sum__1537_comb;
  assign p1_sum__1225_comb = p1_sum__1538_comb + p1_sum__1539_comb;
  assign p1_sum__1210_comb = p1_sum__1508_comb + p1_sum__1509_comb;
  assign p1_sum__1211_comb = p1_sum__1510_comb + p1_sum__1511_comb;
  assign p1_sum__1196_comb = p1_sum__1480_comb + p1_sum__1481_comb;
  assign p1_sum__1197_comb = p1_sum__1482_comb + p1_sum__1483_comb;
  assign p1_sum__1182_comb = p1_sum__1452_comb + p1_sum__1453_comb;
  assign p1_sum__1183_comb = p1_sum__1454_comb + p1_sum__1455_comb;
  assign p1_sum__1168_comb = p1_sum__1424_comb + p1_sum__1425_comb;
  assign p1_sum__1169_comb = p1_sum__1426_comb + p1_sum__1427_comb;
  assign p1_sum__1154_comb = p1_sum__1396_comb + p1_sum__1397_comb;
  assign p1_sum__1155_comb = p1_sum__1398_comb + p1_sum__1399_comb;
  assign p1_sum__1140_comb = p1_sum__1368_comb + p1_sum__1369_comb;
  assign p1_sum__1141_comb = p1_sum__1370_comb + p1_sum__1371_comb;
  assign p1_sum__1236_comb = p1_sum__1560_comb + p1_sum__1561_comb;
  assign p1_sum__1237_comb = p1_sum__1562_comb + p1_sum__1563_comb;
  assign p1_sum__1222_comb = p1_sum__1532_comb + p1_sum__1533_comb;
  assign p1_sum__1223_comb = p1_sum__1534_comb + p1_sum__1535_comb;
  assign p1_sum__1208_comb = p1_sum__1504_comb + p1_sum__1505_comb;
  assign p1_sum__1209_comb = p1_sum__1506_comb + p1_sum__1507_comb;
  assign p1_sum__1194_comb = p1_sum__1476_comb + p1_sum__1477_comb;
  assign p1_sum__1195_comb = p1_sum__1478_comb + p1_sum__1479_comb;
  assign p1_sum__1180_comb = p1_sum__1448_comb + p1_sum__1449_comb;
  assign p1_sum__1181_comb = p1_sum__1450_comb + p1_sum__1451_comb;
  assign p1_sum__1166_comb = p1_sum__1420_comb + p1_sum__1421_comb;
  assign p1_sum__1167_comb = p1_sum__1422_comb + p1_sum__1423_comb;
  assign p1_sum__1152_comb = p1_sum__1392_comb + p1_sum__1393_comb;
  assign p1_sum__1153_comb = p1_sum__1394_comb + p1_sum__1395_comb;
  assign p1_sum__1138_comb = p1_sum__1364_comb + p1_sum__1365_comb;
  assign p1_sum__1139_comb = p1_sum__1366_comb + p1_sum__1367_comb;
  assign p1_sum__1234_comb = p1_sum__1556_comb + p1_sum__1557_comb;
  assign p1_sum__1235_comb = p1_sum__1558_comb + p1_sum__1559_comb;
  assign p1_sum__1220_comb = p1_sum__1528_comb + p1_sum__1529_comb;
  assign p1_sum__1221_comb = p1_sum__1530_comb + p1_sum__1531_comb;
  assign p1_sum__1206_comb = p1_sum__1500_comb + p1_sum__1501_comb;
  assign p1_sum__1207_comb = p1_sum__1502_comb + p1_sum__1503_comb;
  assign p1_sum__1192_comb = p1_sum__1472_comb + p1_sum__1473_comb;
  assign p1_sum__1193_comb = p1_sum__1474_comb + p1_sum__1475_comb;
  assign p1_sum__1178_comb = p1_sum__1444_comb + p1_sum__1445_comb;
  assign p1_sum__1179_comb = p1_sum__1446_comb + p1_sum__1447_comb;
  assign p1_sum__1164_comb = p1_sum__1416_comb + p1_sum__1417_comb;
  assign p1_sum__1165_comb = p1_sum__1418_comb + p1_sum__1419_comb;
  assign p1_sum__1150_comb = p1_sum__1388_comb + p1_sum__1389_comb;
  assign p1_sum__1151_comb = p1_sum__1390_comb + p1_sum__1391_comb;
  assign p1_sum__1136_comb = p1_sum__1360_comb + p1_sum__1361_comb;
  assign p1_sum__1137_comb = p1_sum__1362_comb + p1_sum__1363_comb;
  assign p1_sum__1079_comb = p1_sum__1246_comb + p1_sum__1247_comb;
  assign p1_sum__1072_comb = p1_sum__1232_comb + p1_sum__1233_comb;
  assign p1_sum__1065_comb = p1_sum__1218_comb + p1_sum__1219_comb;
  assign p1_sum__1058_comb = p1_sum__1204_comb + p1_sum__1205_comb;
  assign p1_sum__1051_comb = p1_sum__1190_comb + p1_sum__1191_comb;
  assign p1_sum__1044_comb = p1_sum__1176_comb + p1_sum__1177_comb;
  assign p1_sum__1037_comb = p1_sum__1162_comb + p1_sum__1163_comb;
  assign p1_sum__1030_comb = p1_sum__1148_comb + p1_sum__1149_comb;
  assign p1_sum__1078_comb = p1_sum__1244_comb + p1_sum__1245_comb;
  assign p1_sum__1071_comb = p1_sum__1230_comb + p1_sum__1231_comb;
  assign p1_sum__1064_comb = p1_sum__1216_comb + p1_sum__1217_comb;
  assign p1_sum__1057_comb = p1_sum__1202_comb + p1_sum__1203_comb;
  assign p1_sum__1050_comb = p1_sum__1188_comb + p1_sum__1189_comb;
  assign p1_sum__1043_comb = p1_sum__1174_comb + p1_sum__1175_comb;
  assign p1_sum__1036_comb = p1_sum__1160_comb + p1_sum__1161_comb;
  assign p1_sum__1029_comb = p1_sum__1146_comb + p1_sum__1147_comb;
  assign p1_sum__1077_comb = p1_sum__1242_comb + p1_sum__1243_comb;
  assign p1_sum__1070_comb = p1_sum__1228_comb + p1_sum__1229_comb;
  assign p1_sum__1063_comb = p1_sum__1214_comb + p1_sum__1215_comb;
  assign p1_sum__1056_comb = p1_sum__1200_comb + p1_sum__1201_comb;
  assign p1_sum__1049_comb = p1_sum__1186_comb + p1_sum__1187_comb;
  assign p1_sum__1042_comb = p1_sum__1172_comb + p1_sum__1173_comb;
  assign p1_sum__1035_comb = p1_sum__1158_comb + p1_sum__1159_comb;
  assign p1_sum__1028_comb = p1_sum__1144_comb + p1_sum__1145_comb;
  assign p1_sum__1076_comb = p1_sum__1240_comb + p1_sum__1241_comb;
  assign p1_sum__1069_comb = p1_sum__1226_comb + p1_sum__1227_comb;
  assign p1_sum__1062_comb = p1_sum__1212_comb + p1_sum__1213_comb;
  assign p1_sum__1055_comb = p1_sum__1198_comb + p1_sum__1199_comb;
  assign p1_sum__1048_comb = p1_sum__1184_comb + p1_sum__1185_comb;
  assign p1_sum__1041_comb = p1_sum__1170_comb + p1_sum__1171_comb;
  assign p1_sum__1034_comb = p1_sum__1156_comb + p1_sum__1157_comb;
  assign p1_sum__1027_comb = p1_sum__1142_comb + p1_sum__1143_comb;
  assign p1_sum__1075_comb = p1_sum__1238_comb + p1_sum__1239_comb;
  assign p1_sum__1068_comb = p1_sum__1224_comb + p1_sum__1225_comb;
  assign p1_sum__1061_comb = p1_sum__1210_comb + p1_sum__1211_comb;
  assign p1_sum__1054_comb = p1_sum__1196_comb + p1_sum__1197_comb;
  assign p1_sum__1047_comb = p1_sum__1182_comb + p1_sum__1183_comb;
  assign p1_sum__1040_comb = p1_sum__1168_comb + p1_sum__1169_comb;
  assign p1_sum__1033_comb = p1_sum__1154_comb + p1_sum__1155_comb;
  assign p1_sum__1026_comb = p1_sum__1140_comb + p1_sum__1141_comb;
  assign p1_sum__1074_comb = p1_sum__1236_comb + p1_sum__1237_comb;
  assign p1_sum__1067_comb = p1_sum__1222_comb + p1_sum__1223_comb;
  assign p1_sum__1060_comb = p1_sum__1208_comb + p1_sum__1209_comb;
  assign p1_sum__1053_comb = p1_sum__1194_comb + p1_sum__1195_comb;
  assign p1_sum__1046_comb = p1_sum__1180_comb + p1_sum__1181_comb;
  assign p1_sum__1039_comb = p1_sum__1166_comb + p1_sum__1167_comb;
  assign p1_sum__1032_comb = p1_sum__1152_comb + p1_sum__1153_comb;
  assign p1_sum__1025_comb = p1_sum__1138_comb + p1_sum__1139_comb;
  assign p1_sum__1073_comb = p1_sum__1234_comb + p1_sum__1235_comb;
  assign p1_sum__1066_comb = p1_sum__1220_comb + p1_sum__1221_comb;
  assign p1_sum__1059_comb = p1_sum__1206_comb + p1_sum__1207_comb;
  assign p1_sum__1052_comb = p1_sum__1192_comb + p1_sum__1193_comb;
  assign p1_sum__1045_comb = p1_sum__1178_comb + p1_sum__1179_comb;
  assign p1_sum__1038_comb = p1_sum__1164_comb + p1_sum__1165_comb;
  assign p1_sum__1031_comb = p1_sum__1150_comb + p1_sum__1151_comb;
  assign p1_sum__1024_comb = p1_sum__1136_comb + p1_sum__1137_comb;
  assign p1_add_144473_comb = p1_umul_144225_comb[31:7] + 25'h000_0001;
  assign p1_add_144474_comb = p1_umul_144226_comb[31:7] + 25'h000_0001;
  assign p1_add_144475_comb = p1_umul_144227_comb[31:7] + 25'h000_0001;
  assign p1_add_144476_comb = p1_umul_144228_comb[31:7] + 25'h000_0001;
  assign p1_add_144477_comb = p1_umul_144229_comb[31:7] + 25'h000_0001;
  assign p1_add_144478_comb = p1_umul_144230_comb[31:7] + 25'h000_0001;
  assign p1_add_144479_comb = p1_umul_144231_comb[31:7] + 25'h000_0001;
  assign p1_add_144480_comb = p1_umul_144232_comb[31:7] + 25'h000_0001;
  assign p1_add_144481_comb = p1_sum__1079_comb + 25'h000_0001;
  assign p1_add_144482_comb = p1_sum__1072_comb + 25'h000_0001;
  assign p1_add_144483_comb = p1_sum__1065_comb + 25'h000_0001;
  assign p1_add_144484_comb = p1_sum__1058_comb + 25'h000_0001;
  assign p1_add_144485_comb = p1_sum__1051_comb + 25'h000_0001;
  assign p1_add_144486_comb = p1_sum__1044_comb + 25'h000_0001;
  assign p1_add_144487_comb = p1_sum__1037_comb + 25'h000_0001;
  assign p1_add_144488_comb = p1_sum__1030_comb + 25'h000_0001;
  assign p1_add_144489_comb = p1_sum__1078_comb + 25'h000_0001;
  assign p1_add_144490_comb = p1_sum__1071_comb + 25'h000_0001;
  assign p1_add_144491_comb = p1_sum__1064_comb + 25'h000_0001;
  assign p1_add_144492_comb = p1_sum__1057_comb + 25'h000_0001;
  assign p1_add_144493_comb = p1_sum__1050_comb + 25'h000_0001;
  assign p1_add_144494_comb = p1_sum__1043_comb + 25'h000_0001;
  assign p1_add_144495_comb = p1_sum__1036_comb + 25'h000_0001;
  assign p1_add_144496_comb = p1_sum__1029_comb + 25'h000_0001;
  assign p1_add_144497_comb = p1_sum__1077_comb + 25'h000_0001;
  assign p1_add_144498_comb = p1_sum__1070_comb + 25'h000_0001;
  assign p1_add_144499_comb = p1_sum__1063_comb + 25'h000_0001;
  assign p1_add_144500_comb = p1_sum__1056_comb + 25'h000_0001;
  assign p1_add_144501_comb = p1_sum__1049_comb + 25'h000_0001;
  assign p1_add_144502_comb = p1_sum__1042_comb + 25'h000_0001;
  assign p1_add_144503_comb = p1_sum__1035_comb + 25'h000_0001;
  assign p1_add_144504_comb = p1_sum__1028_comb + 25'h000_0001;
  assign p1_add_144505_comb = p1_sum__1076_comb + 25'h000_0001;
  assign p1_add_144506_comb = p1_sum__1069_comb + 25'h000_0001;
  assign p1_add_144507_comb = p1_sum__1062_comb + 25'h000_0001;
  assign p1_add_144508_comb = p1_sum__1055_comb + 25'h000_0001;
  assign p1_add_144509_comb = p1_sum__1048_comb + 25'h000_0001;
  assign p1_add_144510_comb = p1_sum__1041_comb + 25'h000_0001;
  assign p1_add_144511_comb = p1_sum__1034_comb + 25'h000_0001;
  assign p1_add_144512_comb = p1_sum__1027_comb + 25'h000_0001;
  assign p1_add_144513_comb = p1_sum__1075_comb + 25'h000_0001;
  assign p1_add_144514_comb = p1_sum__1068_comb + 25'h000_0001;
  assign p1_add_144515_comb = p1_sum__1061_comb + 25'h000_0001;
  assign p1_add_144516_comb = p1_sum__1054_comb + 25'h000_0001;
  assign p1_add_144517_comb = p1_sum__1047_comb + 25'h000_0001;
  assign p1_add_144518_comb = p1_sum__1040_comb + 25'h000_0001;
  assign p1_add_144519_comb = p1_sum__1033_comb + 25'h000_0001;
  assign p1_add_144520_comb = p1_sum__1026_comb + 25'h000_0001;
  assign p1_add_144521_comb = p1_sum__1074_comb + 25'h000_0001;
  assign p1_add_144522_comb = p1_sum__1067_comb + 25'h000_0001;
  assign p1_add_144523_comb = p1_sum__1060_comb + 25'h000_0001;
  assign p1_add_144524_comb = p1_sum__1053_comb + 25'h000_0001;
  assign p1_add_144525_comb = p1_sum__1046_comb + 25'h000_0001;
  assign p1_add_144526_comb = p1_sum__1039_comb + 25'h000_0001;
  assign p1_add_144527_comb = p1_sum__1032_comb + 25'h000_0001;
  assign p1_add_144528_comb = p1_sum__1025_comb + 25'h000_0001;
  assign p1_add_144529_comb = p1_sum__1073_comb + 25'h000_0001;
  assign p1_add_144530_comb = p1_sum__1066_comb + 25'h000_0001;
  assign p1_add_144531_comb = p1_sum__1059_comb + 25'h000_0001;
  assign p1_add_144532_comb = p1_sum__1052_comb + 25'h000_0001;
  assign p1_add_144533_comb = p1_sum__1045_comb + 25'h000_0001;
  assign p1_add_144534_comb = p1_sum__1038_comb + 25'h000_0001;
  assign p1_add_144535_comb = p1_sum__1031_comb + 25'h000_0001;
  assign p1_add_144536_comb = p1_sum__1024_comb + 25'h000_0001;
  assign p1_clipped__320_comb = $signed(p1_add_144473_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144473_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144473_comb[16:8]);
  assign p1_clipped__321_comb = $signed(p1_add_144474_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144474_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144474_comb[16:8]);
  assign p1_clipped__322_comb = $signed(p1_add_144475_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144475_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144475_comb[16:8]);
  assign p1_clipped__323_comb = $signed(p1_add_144476_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144476_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144476_comb[16:8]);
  assign p1_clipped__324_comb = $signed(p1_add_144477_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144477_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144477_comb[16:8]);
  assign p1_clipped__325_comb = $signed(p1_add_144478_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144478_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144478_comb[16:8]);
  assign p1_clipped__326_comb = $signed(p1_add_144479_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144479_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144479_comb[16:8]);
  assign p1_clipped__327_comb = $signed(p1_add_144480_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144480_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144480_comb[16:8]);
  assign p1_clipped__328_comb = $signed(p1_add_144481_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144481_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144481_comb[16:8]);
  assign p1_clipped__329_comb = $signed(p1_add_144482_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144482_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144482_comb[16:8]);
  assign p1_clipped__330_comb = $signed(p1_add_144483_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144483_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144483_comb[16:8]);
  assign p1_clipped__331_comb = $signed(p1_add_144484_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144484_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144484_comb[16:8]);
  assign p1_clipped__332_comb = $signed(p1_add_144485_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144485_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144485_comb[16:8]);
  assign p1_clipped__333_comb = $signed(p1_add_144486_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144486_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144486_comb[16:8]);
  assign p1_clipped__334_comb = $signed(p1_add_144487_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144487_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144487_comb[16:8]);
  assign p1_clipped__335_comb = $signed(p1_add_144488_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144488_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144488_comb[16:8]);
  assign p1_clipped__336_comb = $signed(p1_add_144489_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144489_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144489_comb[16:8]);
  assign p1_clipped__337_comb = $signed(p1_add_144490_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144490_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144490_comb[16:8]);
  assign p1_clipped__338_comb = $signed(p1_add_144491_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144491_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144491_comb[16:8]);
  assign p1_clipped__339_comb = $signed(p1_add_144492_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144492_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144492_comb[16:8]);
  assign p1_clipped__340_comb = $signed(p1_add_144493_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144493_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144493_comb[16:8]);
  assign p1_clipped__341_comb = $signed(p1_add_144494_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144494_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144494_comb[16:8]);
  assign p1_clipped__342_comb = $signed(p1_add_144495_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144495_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144495_comb[16:8]);
  assign p1_clipped__343_comb = $signed(p1_add_144496_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144496_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144496_comb[16:8]);
  assign p1_clipped__344_comb = $signed(p1_add_144497_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144497_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144497_comb[16:8]);
  assign p1_clipped__345_comb = $signed(p1_add_144498_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144498_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144498_comb[16:8]);
  assign p1_clipped__346_comb = $signed(p1_add_144499_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144499_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144499_comb[16:8]);
  assign p1_clipped__347_comb = $signed(p1_add_144500_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144500_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144500_comb[16:8]);
  assign p1_clipped__348_comb = $signed(p1_add_144501_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144501_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144501_comb[16:8]);
  assign p1_clipped__349_comb = $signed(p1_add_144502_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144502_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144502_comb[16:8]);
  assign p1_clipped__350_comb = $signed(p1_add_144503_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144503_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144503_comb[16:8]);
  assign p1_clipped__351_comb = $signed(p1_add_144504_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144504_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144504_comb[16:8]);
  assign p1_clipped__352_comb = $signed(p1_add_144505_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144505_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144505_comb[16:8]);
  assign p1_clipped__353_comb = $signed(p1_add_144506_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144506_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144506_comb[16:8]);
  assign p1_clipped__354_comb = $signed(p1_add_144507_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144507_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144507_comb[16:8]);
  assign p1_clipped__355_comb = $signed(p1_add_144508_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144508_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144508_comb[16:8]);
  assign p1_clipped__356_comb = $signed(p1_add_144509_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144509_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144509_comb[16:8]);
  assign p1_clipped__357_comb = $signed(p1_add_144510_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144510_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144510_comb[16:8]);
  assign p1_clipped__358_comb = $signed(p1_add_144511_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144511_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144511_comb[16:8]);
  assign p1_clipped__359_comb = $signed(p1_add_144512_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144512_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144512_comb[16:8]);
  assign p1_clipped__360_comb = $signed(p1_add_144513_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144513_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144513_comb[16:8]);
  assign p1_clipped__361_comb = $signed(p1_add_144514_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144514_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144514_comb[16:8]);
  assign p1_clipped__362_comb = $signed(p1_add_144515_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144515_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144515_comb[16:8]);
  assign p1_clipped__363_comb = $signed(p1_add_144516_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144516_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144516_comb[16:8]);
  assign p1_clipped__364_comb = $signed(p1_add_144517_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144517_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144517_comb[16:8]);
  assign p1_clipped__365_comb = $signed(p1_add_144518_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144518_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144518_comb[16:8]);
  assign p1_clipped__366_comb = $signed(p1_add_144519_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144519_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144519_comb[16:8]);
  assign p1_clipped__367_comb = $signed(p1_add_144520_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144520_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144520_comb[16:8]);
  assign p1_clipped__368_comb = $signed(p1_add_144521_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144521_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144521_comb[16:8]);
  assign p1_clipped__369_comb = $signed(p1_add_144522_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144522_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144522_comb[16:8]);
  assign p1_clipped__370_comb = $signed(p1_add_144523_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144523_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144523_comb[16:8]);
  assign p1_clipped__371_comb = $signed(p1_add_144524_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144524_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144524_comb[16:8]);
  assign p1_clipped__372_comb = $signed(p1_add_144525_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144525_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144525_comb[16:8]);
  assign p1_clipped__373_comb = $signed(p1_add_144526_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144526_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144526_comb[16:8]);
  assign p1_clipped__374_comb = $signed(p1_add_144527_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144527_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144527_comb[16:8]);
  assign p1_clipped__375_comb = $signed(p1_add_144528_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144528_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144528_comb[16:8]);
  assign p1_clipped__376_comb = $signed(p1_add_144529_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144529_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144529_comb[16:8]);
  assign p1_clipped__377_comb = $signed(p1_add_144530_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144530_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144530_comb[16:8]);
  assign p1_clipped__378_comb = $signed(p1_add_144531_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144531_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144531_comb[16:8]);
  assign p1_clipped__379_comb = $signed(p1_add_144532_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144532_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144532_comb[16:8]);
  assign p1_clipped__380_comb = $signed(p1_add_144533_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144533_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144533_comb[16:8]);
  assign p1_clipped__381_comb = $signed(p1_add_144534_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144534_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144534_comb[16:8]);
  assign p1_clipped__382_comb = $signed(p1_add_144535_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144535_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144535_comb[16:8]);
  assign p1_clipped__383_comb = $signed(p1_add_144536_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_144536_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_144536_comb[16:8]);
  assign p1_add_145305_comb = {{1{p1_clipped__320_comb[8]}}, p1_clipped__320_comb} + 10'h001;
  assign p1_add_145306_comb = {{1{p1_clipped__321_comb[8]}}, p1_clipped__321_comb} + 10'h001;
  assign p1_add_145307_comb = {{1{p1_clipped__322_comb[8]}}, p1_clipped__322_comb} + 10'h001;
  assign p1_add_145308_comb = {{1{p1_clipped__323_comb[8]}}, p1_clipped__323_comb} + 10'h001;
  assign p1_add_145309_comb = {{1{p1_clipped__324_comb[8]}}, p1_clipped__324_comb} + 10'h001;
  assign p1_add_145310_comb = {{1{p1_clipped__325_comb[8]}}, p1_clipped__325_comb} + 10'h001;
  assign p1_add_145311_comb = {{1{p1_clipped__326_comb[8]}}, p1_clipped__326_comb} + 10'h001;
  assign p1_add_145312_comb = {{1{p1_clipped__327_comb[8]}}, p1_clipped__327_comb} + 10'h001;
  assign p1_add_145313_comb = {{1{p1_clipped__328_comb[8]}}, p1_clipped__328_comb} + 10'h001;
  assign p1_add_145314_comb = {{1{p1_clipped__329_comb[8]}}, p1_clipped__329_comb} + 10'h001;
  assign p1_add_145315_comb = {{1{p1_clipped__330_comb[8]}}, p1_clipped__330_comb} + 10'h001;
  assign p1_add_145316_comb = {{1{p1_clipped__331_comb[8]}}, p1_clipped__331_comb} + 10'h001;
  assign p1_add_145317_comb = {{1{p1_clipped__332_comb[8]}}, p1_clipped__332_comb} + 10'h001;
  assign p1_add_145318_comb = {{1{p1_clipped__333_comb[8]}}, p1_clipped__333_comb} + 10'h001;
  assign p1_add_145319_comb = {{1{p1_clipped__334_comb[8]}}, p1_clipped__334_comb} + 10'h001;
  assign p1_add_145320_comb = {{1{p1_clipped__335_comb[8]}}, p1_clipped__335_comb} + 10'h001;
  assign p1_add_145321_comb = {{1{p1_clipped__336_comb[8]}}, p1_clipped__336_comb} + 10'h001;
  assign p1_add_145322_comb = {{1{p1_clipped__337_comb[8]}}, p1_clipped__337_comb} + 10'h001;
  assign p1_add_145323_comb = {{1{p1_clipped__338_comb[8]}}, p1_clipped__338_comb} + 10'h001;
  assign p1_add_145324_comb = {{1{p1_clipped__339_comb[8]}}, p1_clipped__339_comb} + 10'h001;
  assign p1_add_145325_comb = {{1{p1_clipped__340_comb[8]}}, p1_clipped__340_comb} + 10'h001;
  assign p1_add_145326_comb = {{1{p1_clipped__341_comb[8]}}, p1_clipped__341_comb} + 10'h001;
  assign p1_add_145327_comb = {{1{p1_clipped__342_comb[8]}}, p1_clipped__342_comb} + 10'h001;
  assign p1_add_145328_comb = {{1{p1_clipped__343_comb[8]}}, p1_clipped__343_comb} + 10'h001;
  assign p1_add_145329_comb = {{1{p1_clipped__344_comb[8]}}, p1_clipped__344_comb} + 10'h001;
  assign p1_add_145330_comb = {{1{p1_clipped__345_comb[8]}}, p1_clipped__345_comb} + 10'h001;
  assign p1_add_145331_comb = {{1{p1_clipped__346_comb[8]}}, p1_clipped__346_comb} + 10'h001;
  assign p1_add_145332_comb = {{1{p1_clipped__347_comb[8]}}, p1_clipped__347_comb} + 10'h001;
  assign p1_add_145333_comb = {{1{p1_clipped__348_comb[8]}}, p1_clipped__348_comb} + 10'h001;
  assign p1_add_145334_comb = {{1{p1_clipped__349_comb[8]}}, p1_clipped__349_comb} + 10'h001;
  assign p1_add_145335_comb = {{1{p1_clipped__350_comb[8]}}, p1_clipped__350_comb} + 10'h001;
  assign p1_add_145336_comb = {{1{p1_clipped__351_comb[8]}}, p1_clipped__351_comb} + 10'h001;
  assign p1_add_145337_comb = {{1{p1_clipped__352_comb[8]}}, p1_clipped__352_comb} + 10'h001;
  assign p1_add_145338_comb = {{1{p1_clipped__353_comb[8]}}, p1_clipped__353_comb} + 10'h001;
  assign p1_add_145339_comb = {{1{p1_clipped__354_comb[8]}}, p1_clipped__354_comb} + 10'h001;
  assign p1_add_145340_comb = {{1{p1_clipped__355_comb[8]}}, p1_clipped__355_comb} + 10'h001;
  assign p1_add_145341_comb = {{1{p1_clipped__356_comb[8]}}, p1_clipped__356_comb} + 10'h001;
  assign p1_add_145342_comb = {{1{p1_clipped__357_comb[8]}}, p1_clipped__357_comb} + 10'h001;
  assign p1_add_145343_comb = {{1{p1_clipped__358_comb[8]}}, p1_clipped__358_comb} + 10'h001;
  assign p1_add_145344_comb = {{1{p1_clipped__359_comb[8]}}, p1_clipped__359_comb} + 10'h001;
  assign p1_add_145345_comb = {{1{p1_clipped__360_comb[8]}}, p1_clipped__360_comb} + 10'h001;
  assign p1_add_145346_comb = {{1{p1_clipped__361_comb[8]}}, p1_clipped__361_comb} + 10'h001;
  assign p1_add_145347_comb = {{1{p1_clipped__362_comb[8]}}, p1_clipped__362_comb} + 10'h001;
  assign p1_add_145348_comb = {{1{p1_clipped__363_comb[8]}}, p1_clipped__363_comb} + 10'h001;
  assign p1_add_145349_comb = {{1{p1_clipped__364_comb[8]}}, p1_clipped__364_comb} + 10'h001;
  assign p1_add_145350_comb = {{1{p1_clipped__365_comb[8]}}, p1_clipped__365_comb} + 10'h001;
  assign p1_add_145351_comb = {{1{p1_clipped__366_comb[8]}}, p1_clipped__366_comb} + 10'h001;
  assign p1_add_145352_comb = {{1{p1_clipped__367_comb[8]}}, p1_clipped__367_comb} + 10'h001;
  assign p1_add_145353_comb = {{1{p1_clipped__368_comb[8]}}, p1_clipped__368_comb} + 10'h001;
  assign p1_add_145354_comb = {{1{p1_clipped__369_comb[8]}}, p1_clipped__369_comb} + 10'h001;
  assign p1_add_145355_comb = {{1{p1_clipped__370_comb[8]}}, p1_clipped__370_comb} + 10'h001;
  assign p1_add_145356_comb = {{1{p1_clipped__371_comb[8]}}, p1_clipped__371_comb} + 10'h001;
  assign p1_add_145357_comb = {{1{p1_clipped__372_comb[8]}}, p1_clipped__372_comb} + 10'h001;
  assign p1_add_145358_comb = {{1{p1_clipped__373_comb[8]}}, p1_clipped__373_comb} + 10'h001;
  assign p1_add_145359_comb = {{1{p1_clipped__374_comb[8]}}, p1_clipped__374_comb} + 10'h001;
  assign p1_add_145360_comb = {{1{p1_clipped__375_comb[8]}}, p1_clipped__375_comb} + 10'h001;
  assign p1_add_145361_comb = {{1{p1_clipped__376_comb[8]}}, p1_clipped__376_comb} + 10'h001;
  assign p1_add_145362_comb = {{1{p1_clipped__377_comb[8]}}, p1_clipped__377_comb} + 10'h001;
  assign p1_add_145363_comb = {{1{p1_clipped__378_comb[8]}}, p1_clipped__378_comb} + 10'h001;
  assign p1_add_145364_comb = {{1{p1_clipped__379_comb[8]}}, p1_clipped__379_comb} + 10'h001;
  assign p1_add_145365_comb = {{1{p1_clipped__380_comb[8]}}, p1_clipped__380_comb} + 10'h001;
  assign p1_add_145366_comb = {{1{p1_clipped__381_comb[8]}}, p1_clipped__381_comb} + 10'h001;
  assign p1_add_145367_comb = {{1{p1_clipped__382_comb[8]}}, p1_clipped__382_comb} + 10'h001;
  assign p1_add_145368_comb = {{1{p1_clipped__383_comb[8]}}, p1_clipped__383_comb} + 10'h001;
  assign p1_bit_slice_145369_comb = p1_add_145305_comb[9:8];
  assign p1_bit_slice_145370_comb = p1_add_145306_comb[9:8];
  assign p1_bit_slice_145371_comb = p1_add_145307_comb[9:8];
  assign p1_bit_slice_145372_comb = p1_add_145308_comb[9:8];
  assign p1_bit_slice_145373_comb = p1_add_145309_comb[9:8];
  assign p1_bit_slice_145374_comb = p1_add_145310_comb[9:8];
  assign p1_bit_slice_145375_comb = p1_add_145311_comb[9:8];
  assign p1_bit_slice_145376_comb = p1_add_145312_comb[9:8];
  assign p1_bit_slice_145377_comb = p1_add_145313_comb[9:8];
  assign p1_bit_slice_145378_comb = p1_add_145314_comb[9:8];
  assign p1_bit_slice_145379_comb = p1_add_145315_comb[9:8];
  assign p1_bit_slice_145380_comb = p1_add_145316_comb[9:8];
  assign p1_bit_slice_145381_comb = p1_add_145317_comb[9:8];
  assign p1_bit_slice_145382_comb = p1_add_145318_comb[9:8];
  assign p1_bit_slice_145383_comb = p1_add_145319_comb[9:8];
  assign p1_bit_slice_145384_comb = p1_add_145320_comb[9:8];
  assign p1_bit_slice_145385_comb = p1_add_145321_comb[9:8];
  assign p1_bit_slice_145386_comb = p1_add_145322_comb[9:8];
  assign p1_bit_slice_145387_comb = p1_add_145323_comb[9:8];
  assign p1_bit_slice_145388_comb = p1_add_145324_comb[9:8];
  assign p1_bit_slice_145389_comb = p1_add_145325_comb[9:8];
  assign p1_bit_slice_145390_comb = p1_add_145326_comb[9:8];
  assign p1_bit_slice_145391_comb = p1_add_145327_comb[9:8];
  assign p1_bit_slice_145392_comb = p1_add_145328_comb[9:8];
  assign p1_bit_slice_145393_comb = p1_add_145329_comb[9:8];
  assign p1_bit_slice_145394_comb = p1_add_145330_comb[9:8];
  assign p1_bit_slice_145395_comb = p1_add_145331_comb[9:8];
  assign p1_bit_slice_145396_comb = p1_add_145332_comb[9:8];
  assign p1_bit_slice_145397_comb = p1_add_145333_comb[9:8];
  assign p1_bit_slice_145398_comb = p1_add_145334_comb[9:8];
  assign p1_bit_slice_145399_comb = p1_add_145335_comb[9:8];
  assign p1_bit_slice_145400_comb = p1_add_145336_comb[9:8];
  assign p1_bit_slice_145401_comb = p1_add_145337_comb[9:8];
  assign p1_bit_slice_145402_comb = p1_add_145338_comb[9:8];
  assign p1_bit_slice_145403_comb = p1_add_145339_comb[9:8];
  assign p1_bit_slice_145404_comb = p1_add_145340_comb[9:8];
  assign p1_bit_slice_145405_comb = p1_add_145341_comb[9:8];
  assign p1_bit_slice_145406_comb = p1_add_145342_comb[9:8];
  assign p1_bit_slice_145407_comb = p1_add_145343_comb[9:8];
  assign p1_bit_slice_145408_comb = p1_add_145344_comb[9:8];
  assign p1_bit_slice_145409_comb = p1_add_145345_comb[9:8];
  assign p1_bit_slice_145410_comb = p1_add_145346_comb[9:8];
  assign p1_bit_slice_145411_comb = p1_add_145347_comb[9:8];
  assign p1_bit_slice_145412_comb = p1_add_145348_comb[9:8];
  assign p1_bit_slice_145413_comb = p1_add_145349_comb[9:8];
  assign p1_bit_slice_145414_comb = p1_add_145350_comb[9:8];
  assign p1_bit_slice_145415_comb = p1_add_145351_comb[9:8];
  assign p1_bit_slice_145416_comb = p1_add_145352_comb[9:8];
  assign p1_bit_slice_145417_comb = p1_add_145353_comb[9:8];
  assign p1_bit_slice_145418_comb = p1_add_145354_comb[9:8];
  assign p1_bit_slice_145419_comb = p1_add_145355_comb[9:8];
  assign p1_bit_slice_145420_comb = p1_add_145356_comb[9:8];
  assign p1_bit_slice_145421_comb = p1_add_145357_comb[9:8];
  assign p1_bit_slice_145422_comb = p1_add_145358_comb[9:8];
  assign p1_bit_slice_145423_comb = p1_add_145359_comb[9:8];
  assign p1_bit_slice_145424_comb = p1_add_145360_comb[9:8];
  assign p1_bit_slice_145425_comb = p1_add_145361_comb[9:8];
  assign p1_bit_slice_145426_comb = p1_add_145362_comb[9:8];
  assign p1_bit_slice_145427_comb = p1_add_145363_comb[9:8];
  assign p1_bit_slice_145428_comb = p1_add_145364_comb[9:8];
  assign p1_bit_slice_145429_comb = p1_add_145365_comb[9:8];
  assign p1_bit_slice_145430_comb = p1_add_145366_comb[9:8];
  assign p1_bit_slice_145431_comb = p1_add_145367_comb[9:8];
  assign p1_bit_slice_145432_comb = p1_add_145368_comb[9:8];
  assign p1_add_145561_comb = {{1{p1_bit_slice_145369_comb[1]}}, p1_bit_slice_145369_comb} + 3'h1;
  assign p1_add_145562_comb = {{1{p1_bit_slice_145370_comb[1]}}, p1_bit_slice_145370_comb} + 3'h1;
  assign p1_add_145563_comb = {{1{p1_bit_slice_145371_comb[1]}}, p1_bit_slice_145371_comb} + 3'h1;
  assign p1_add_145564_comb = {{1{p1_bit_slice_145372_comb[1]}}, p1_bit_slice_145372_comb} + 3'h1;
  assign p1_add_145565_comb = {{1{p1_bit_slice_145373_comb[1]}}, p1_bit_slice_145373_comb} + 3'h1;
  assign p1_add_145566_comb = {{1{p1_bit_slice_145374_comb[1]}}, p1_bit_slice_145374_comb} + 3'h1;
  assign p1_add_145567_comb = {{1{p1_bit_slice_145375_comb[1]}}, p1_bit_slice_145375_comb} + 3'h1;
  assign p1_add_145568_comb = {{1{p1_bit_slice_145376_comb[1]}}, p1_bit_slice_145376_comb} + 3'h1;
  assign p1_add_145569_comb = {{1{p1_bit_slice_145377_comb[1]}}, p1_bit_slice_145377_comb} + 3'h1;
  assign p1_add_145570_comb = {{1{p1_bit_slice_145378_comb[1]}}, p1_bit_slice_145378_comb} + 3'h1;
  assign p1_add_145571_comb = {{1{p1_bit_slice_145379_comb[1]}}, p1_bit_slice_145379_comb} + 3'h1;
  assign p1_add_145572_comb = {{1{p1_bit_slice_145380_comb[1]}}, p1_bit_slice_145380_comb} + 3'h1;
  assign p1_add_145573_comb = {{1{p1_bit_slice_145381_comb[1]}}, p1_bit_slice_145381_comb} + 3'h1;
  assign p1_add_145574_comb = {{1{p1_bit_slice_145382_comb[1]}}, p1_bit_slice_145382_comb} + 3'h1;
  assign p1_add_145575_comb = {{1{p1_bit_slice_145383_comb[1]}}, p1_bit_slice_145383_comb} + 3'h1;
  assign p1_add_145576_comb = {{1{p1_bit_slice_145384_comb[1]}}, p1_bit_slice_145384_comb} + 3'h1;
  assign p1_add_145577_comb = {{1{p1_bit_slice_145385_comb[1]}}, p1_bit_slice_145385_comb} + 3'h1;
  assign p1_add_145578_comb = {{1{p1_bit_slice_145386_comb[1]}}, p1_bit_slice_145386_comb} + 3'h1;
  assign p1_add_145579_comb = {{1{p1_bit_slice_145387_comb[1]}}, p1_bit_slice_145387_comb} + 3'h1;
  assign p1_add_145580_comb = {{1{p1_bit_slice_145388_comb[1]}}, p1_bit_slice_145388_comb} + 3'h1;
  assign p1_add_145581_comb = {{1{p1_bit_slice_145389_comb[1]}}, p1_bit_slice_145389_comb} + 3'h1;
  assign p1_add_145582_comb = {{1{p1_bit_slice_145390_comb[1]}}, p1_bit_slice_145390_comb} + 3'h1;
  assign p1_add_145583_comb = {{1{p1_bit_slice_145391_comb[1]}}, p1_bit_slice_145391_comb} + 3'h1;
  assign p1_add_145584_comb = {{1{p1_bit_slice_145392_comb[1]}}, p1_bit_slice_145392_comb} + 3'h1;
  assign p1_add_145585_comb = {{1{p1_bit_slice_145393_comb[1]}}, p1_bit_slice_145393_comb} + 3'h1;
  assign p1_add_145586_comb = {{1{p1_bit_slice_145394_comb[1]}}, p1_bit_slice_145394_comb} + 3'h1;
  assign p1_add_145587_comb = {{1{p1_bit_slice_145395_comb[1]}}, p1_bit_slice_145395_comb} + 3'h1;
  assign p1_add_145588_comb = {{1{p1_bit_slice_145396_comb[1]}}, p1_bit_slice_145396_comb} + 3'h1;
  assign p1_add_145589_comb = {{1{p1_bit_slice_145397_comb[1]}}, p1_bit_slice_145397_comb} + 3'h1;
  assign p1_add_145590_comb = {{1{p1_bit_slice_145398_comb[1]}}, p1_bit_slice_145398_comb} + 3'h1;
  assign p1_add_145591_comb = {{1{p1_bit_slice_145399_comb[1]}}, p1_bit_slice_145399_comb} + 3'h1;
  assign p1_add_145592_comb = {{1{p1_bit_slice_145400_comb[1]}}, p1_bit_slice_145400_comb} + 3'h1;
  assign p1_add_145593_comb = {{1{p1_bit_slice_145401_comb[1]}}, p1_bit_slice_145401_comb} + 3'h1;
  assign p1_add_145594_comb = {{1{p1_bit_slice_145402_comb[1]}}, p1_bit_slice_145402_comb} + 3'h1;
  assign p1_add_145595_comb = {{1{p1_bit_slice_145403_comb[1]}}, p1_bit_slice_145403_comb} + 3'h1;
  assign p1_add_145596_comb = {{1{p1_bit_slice_145404_comb[1]}}, p1_bit_slice_145404_comb} + 3'h1;
  assign p1_add_145597_comb = {{1{p1_bit_slice_145405_comb[1]}}, p1_bit_slice_145405_comb} + 3'h1;
  assign p1_add_145598_comb = {{1{p1_bit_slice_145406_comb[1]}}, p1_bit_slice_145406_comb} + 3'h1;
  assign p1_add_145599_comb = {{1{p1_bit_slice_145407_comb[1]}}, p1_bit_slice_145407_comb} + 3'h1;
  assign p1_add_145600_comb = {{1{p1_bit_slice_145408_comb[1]}}, p1_bit_slice_145408_comb} + 3'h1;
  assign p1_add_145601_comb = {{1{p1_bit_slice_145409_comb[1]}}, p1_bit_slice_145409_comb} + 3'h1;
  assign p1_add_145602_comb = {{1{p1_bit_slice_145410_comb[1]}}, p1_bit_slice_145410_comb} + 3'h1;
  assign p1_add_145603_comb = {{1{p1_bit_slice_145411_comb[1]}}, p1_bit_slice_145411_comb} + 3'h1;
  assign p1_add_145604_comb = {{1{p1_bit_slice_145412_comb[1]}}, p1_bit_slice_145412_comb} + 3'h1;
  assign p1_add_145605_comb = {{1{p1_bit_slice_145413_comb[1]}}, p1_bit_slice_145413_comb} + 3'h1;
  assign p1_add_145606_comb = {{1{p1_bit_slice_145414_comb[1]}}, p1_bit_slice_145414_comb} + 3'h1;
  assign p1_add_145607_comb = {{1{p1_bit_slice_145415_comb[1]}}, p1_bit_slice_145415_comb} + 3'h1;
  assign p1_add_145608_comb = {{1{p1_bit_slice_145416_comb[1]}}, p1_bit_slice_145416_comb} + 3'h1;
  assign p1_add_145609_comb = {{1{p1_bit_slice_145417_comb[1]}}, p1_bit_slice_145417_comb} + 3'h1;
  assign p1_add_145610_comb = {{1{p1_bit_slice_145418_comb[1]}}, p1_bit_slice_145418_comb} + 3'h1;
  assign p1_add_145611_comb = {{1{p1_bit_slice_145419_comb[1]}}, p1_bit_slice_145419_comb} + 3'h1;
  assign p1_add_145612_comb = {{1{p1_bit_slice_145420_comb[1]}}, p1_bit_slice_145420_comb} + 3'h1;
  assign p1_add_145613_comb = {{1{p1_bit_slice_145421_comb[1]}}, p1_bit_slice_145421_comb} + 3'h1;
  assign p1_add_145614_comb = {{1{p1_bit_slice_145422_comb[1]}}, p1_bit_slice_145422_comb} + 3'h1;
  assign p1_add_145615_comb = {{1{p1_bit_slice_145423_comb[1]}}, p1_bit_slice_145423_comb} + 3'h1;
  assign p1_add_145616_comb = {{1{p1_bit_slice_145424_comb[1]}}, p1_bit_slice_145424_comb} + 3'h1;
  assign p1_add_145617_comb = {{1{p1_bit_slice_145425_comb[1]}}, p1_bit_slice_145425_comb} + 3'h1;
  assign p1_add_145618_comb = {{1{p1_bit_slice_145426_comb[1]}}, p1_bit_slice_145426_comb} + 3'h1;
  assign p1_add_145619_comb = {{1{p1_bit_slice_145427_comb[1]}}, p1_bit_slice_145427_comb} + 3'h1;
  assign p1_add_145620_comb = {{1{p1_bit_slice_145428_comb[1]}}, p1_bit_slice_145428_comb} + 3'h1;
  assign p1_add_145621_comb = {{1{p1_bit_slice_145429_comb[1]}}, p1_bit_slice_145429_comb} + 3'h1;
  assign p1_add_145622_comb = {{1{p1_bit_slice_145430_comb[1]}}, p1_bit_slice_145430_comb} + 3'h1;
  assign p1_add_145623_comb = {{1{p1_bit_slice_145431_comb[1]}}, p1_bit_slice_145431_comb} + 3'h1;
  assign p1_add_145624_comb = {{1{p1_bit_slice_145432_comb[1]}}, p1_bit_slice_145432_comb} + 3'h1;
  assign p1_clipped__136_comb = p1_add_145561_comb[1] ? 8'hff : {p1_add_145561_comb[0], p1_add_145305_comb[7:1]};
  assign p1_clipped__152_comb = p1_add_145562_comb[1] ? 8'hff : {p1_add_145562_comb[0], p1_add_145306_comb[7:1]};
  assign p1_clipped__168_comb = p1_add_145563_comb[1] ? 8'hff : {p1_add_145563_comb[0], p1_add_145307_comb[7:1]};
  assign p1_clipped__184_comb = p1_add_145564_comb[1] ? 8'hff : {p1_add_145564_comb[0], p1_add_145308_comb[7:1]};
  assign p1_clipped__200_comb = p1_add_145565_comb[1] ? 8'hff : {p1_add_145565_comb[0], p1_add_145309_comb[7:1]};
  assign p1_clipped__216_comb = p1_add_145566_comb[1] ? 8'hff : {p1_add_145566_comb[0], p1_add_145310_comb[7:1]};
  assign p1_clipped__232_comb = p1_add_145567_comb[1] ? 8'hff : {p1_add_145567_comb[0], p1_add_145311_comb[7:1]};
  assign p1_clipped__248_comb = p1_add_145568_comb[1] ? 8'hff : {p1_add_145568_comb[0], p1_add_145312_comb[7:1]};
  assign p1_clipped__137_comb = p1_add_145569_comb[1] ? 8'hff : {p1_add_145569_comb[0], p1_add_145313_comb[7:1]};
  assign p1_clipped__153_comb = p1_add_145570_comb[1] ? 8'hff : {p1_add_145570_comb[0], p1_add_145314_comb[7:1]};
  assign p1_clipped__169_comb = p1_add_145571_comb[1] ? 8'hff : {p1_add_145571_comb[0], p1_add_145315_comb[7:1]};
  assign p1_clipped__185_comb = p1_add_145572_comb[1] ? 8'hff : {p1_add_145572_comb[0], p1_add_145316_comb[7:1]};
  assign p1_clipped__201_comb = p1_add_145573_comb[1] ? 8'hff : {p1_add_145573_comb[0], p1_add_145317_comb[7:1]};
  assign p1_clipped__217_comb = p1_add_145574_comb[1] ? 8'hff : {p1_add_145574_comb[0], p1_add_145318_comb[7:1]};
  assign p1_clipped__233_comb = p1_add_145575_comb[1] ? 8'hff : {p1_add_145575_comb[0], p1_add_145319_comb[7:1]};
  assign p1_clipped__249_comb = p1_add_145576_comb[1] ? 8'hff : {p1_add_145576_comb[0], p1_add_145320_comb[7:1]};
  assign p1_clipped__138_comb = p1_add_145577_comb[1] ? 8'hff : {p1_add_145577_comb[0], p1_add_145321_comb[7:1]};
  assign p1_clipped__154_comb = p1_add_145578_comb[1] ? 8'hff : {p1_add_145578_comb[0], p1_add_145322_comb[7:1]};
  assign p1_clipped__170_comb = p1_add_145579_comb[1] ? 8'hff : {p1_add_145579_comb[0], p1_add_145323_comb[7:1]};
  assign p1_clipped__186_comb = p1_add_145580_comb[1] ? 8'hff : {p1_add_145580_comb[0], p1_add_145324_comb[7:1]};
  assign p1_clipped__202_comb = p1_add_145581_comb[1] ? 8'hff : {p1_add_145581_comb[0], p1_add_145325_comb[7:1]};
  assign p1_clipped__218_comb = p1_add_145582_comb[1] ? 8'hff : {p1_add_145582_comb[0], p1_add_145326_comb[7:1]};
  assign p1_clipped__234_comb = p1_add_145583_comb[1] ? 8'hff : {p1_add_145583_comb[0], p1_add_145327_comb[7:1]};
  assign p1_clipped__250_comb = p1_add_145584_comb[1] ? 8'hff : {p1_add_145584_comb[0], p1_add_145328_comb[7:1]};
  assign p1_clipped__139_comb = p1_add_145585_comb[1] ? 8'hff : {p1_add_145585_comb[0], p1_add_145329_comb[7:1]};
  assign p1_clipped__155_comb = p1_add_145586_comb[1] ? 8'hff : {p1_add_145586_comb[0], p1_add_145330_comb[7:1]};
  assign p1_clipped__171_comb = p1_add_145587_comb[1] ? 8'hff : {p1_add_145587_comb[0], p1_add_145331_comb[7:1]};
  assign p1_clipped__187_comb = p1_add_145588_comb[1] ? 8'hff : {p1_add_145588_comb[0], p1_add_145332_comb[7:1]};
  assign p1_clipped__203_comb = p1_add_145589_comb[1] ? 8'hff : {p1_add_145589_comb[0], p1_add_145333_comb[7:1]};
  assign p1_clipped__219_comb = p1_add_145590_comb[1] ? 8'hff : {p1_add_145590_comb[0], p1_add_145334_comb[7:1]};
  assign p1_clipped__235_comb = p1_add_145591_comb[1] ? 8'hff : {p1_add_145591_comb[0], p1_add_145335_comb[7:1]};
  assign p1_clipped__251_comb = p1_add_145592_comb[1] ? 8'hff : {p1_add_145592_comb[0], p1_add_145336_comb[7:1]};
  assign p1_clipped__140_comb = p1_add_145593_comb[1] ? 8'hff : {p1_add_145593_comb[0], p1_add_145337_comb[7:1]};
  assign p1_clipped__156_comb = p1_add_145594_comb[1] ? 8'hff : {p1_add_145594_comb[0], p1_add_145338_comb[7:1]};
  assign p1_clipped__172_comb = p1_add_145595_comb[1] ? 8'hff : {p1_add_145595_comb[0], p1_add_145339_comb[7:1]};
  assign p1_clipped__188_comb = p1_add_145596_comb[1] ? 8'hff : {p1_add_145596_comb[0], p1_add_145340_comb[7:1]};
  assign p1_clipped__204_comb = p1_add_145597_comb[1] ? 8'hff : {p1_add_145597_comb[0], p1_add_145341_comb[7:1]};
  assign p1_clipped__220_comb = p1_add_145598_comb[1] ? 8'hff : {p1_add_145598_comb[0], p1_add_145342_comb[7:1]};
  assign p1_clipped__236_comb = p1_add_145599_comb[1] ? 8'hff : {p1_add_145599_comb[0], p1_add_145343_comb[7:1]};
  assign p1_clipped__252_comb = p1_add_145600_comb[1] ? 8'hff : {p1_add_145600_comb[0], p1_add_145344_comb[7:1]};
  assign p1_clipped__141_comb = p1_add_145601_comb[1] ? 8'hff : {p1_add_145601_comb[0], p1_add_145345_comb[7:1]};
  assign p1_clipped__157_comb = p1_add_145602_comb[1] ? 8'hff : {p1_add_145602_comb[0], p1_add_145346_comb[7:1]};
  assign p1_clipped__173_comb = p1_add_145603_comb[1] ? 8'hff : {p1_add_145603_comb[0], p1_add_145347_comb[7:1]};
  assign p1_clipped__189_comb = p1_add_145604_comb[1] ? 8'hff : {p1_add_145604_comb[0], p1_add_145348_comb[7:1]};
  assign p1_clipped__205_comb = p1_add_145605_comb[1] ? 8'hff : {p1_add_145605_comb[0], p1_add_145349_comb[7:1]};
  assign p1_clipped__221_comb = p1_add_145606_comb[1] ? 8'hff : {p1_add_145606_comb[0], p1_add_145350_comb[7:1]};
  assign p1_clipped__237_comb = p1_add_145607_comb[1] ? 8'hff : {p1_add_145607_comb[0], p1_add_145351_comb[7:1]};
  assign p1_clipped__253_comb = p1_add_145608_comb[1] ? 8'hff : {p1_add_145608_comb[0], p1_add_145352_comb[7:1]};
  assign p1_clipped__142_comb = p1_add_145609_comb[1] ? 8'hff : {p1_add_145609_comb[0], p1_add_145353_comb[7:1]};
  assign p1_clipped__158_comb = p1_add_145610_comb[1] ? 8'hff : {p1_add_145610_comb[0], p1_add_145354_comb[7:1]};
  assign p1_clipped__174_comb = p1_add_145611_comb[1] ? 8'hff : {p1_add_145611_comb[0], p1_add_145355_comb[7:1]};
  assign p1_clipped__190_comb = p1_add_145612_comb[1] ? 8'hff : {p1_add_145612_comb[0], p1_add_145356_comb[7:1]};
  assign p1_clipped__206_comb = p1_add_145613_comb[1] ? 8'hff : {p1_add_145613_comb[0], p1_add_145357_comb[7:1]};
  assign p1_clipped__222_comb = p1_add_145614_comb[1] ? 8'hff : {p1_add_145614_comb[0], p1_add_145358_comb[7:1]};
  assign p1_clipped__238_comb = p1_add_145615_comb[1] ? 8'hff : {p1_add_145615_comb[0], p1_add_145359_comb[7:1]};
  assign p1_clipped__254_comb = p1_add_145616_comb[1] ? 8'hff : {p1_add_145616_comb[0], p1_add_145360_comb[7:1]};
  assign p1_clipped__143_comb = p1_add_145617_comb[1] ? 8'hff : {p1_add_145617_comb[0], p1_add_145361_comb[7:1]};
  assign p1_clipped__159_comb = p1_add_145618_comb[1] ? 8'hff : {p1_add_145618_comb[0], p1_add_145362_comb[7:1]};
  assign p1_clipped__175_comb = p1_add_145619_comb[1] ? 8'hff : {p1_add_145619_comb[0], p1_add_145363_comb[7:1]};
  assign p1_clipped__191_comb = p1_add_145620_comb[1] ? 8'hff : {p1_add_145620_comb[0], p1_add_145364_comb[7:1]};
  assign p1_clipped__207_comb = p1_add_145621_comb[1] ? 8'hff : {p1_add_145621_comb[0], p1_add_145365_comb[7:1]};
  assign p1_clipped__223_comb = p1_add_145622_comb[1] ? 8'hff : {p1_add_145622_comb[0], p1_add_145366_comb[7:1]};
  assign p1_clipped__239_comb = p1_add_145623_comb[1] ? 8'hff : {p1_add_145623_comb[0], p1_add_145367_comb[7:1]};
  assign p1_clipped__255_comb = p1_add_145624_comb[1] ? 8'hff : {p1_add_145624_comb[0], p1_add_145368_comb[7:1]};
  assign p1_array_146009_comb[0] = p1_clipped__136_comb;
  assign p1_array_146009_comb[1] = p1_clipped__152_comb;
  assign p1_array_146009_comb[2] = p1_clipped__168_comb;
  assign p1_array_146009_comb[3] = p1_clipped__184_comb;
  assign p1_array_146009_comb[4] = p1_clipped__200_comb;
  assign p1_array_146009_comb[5] = p1_clipped__216_comb;
  assign p1_array_146009_comb[6] = p1_clipped__232_comb;
  assign p1_array_146009_comb[7] = p1_clipped__248_comb;
  assign p1_array_146010_comb[0] = p1_clipped__137_comb;
  assign p1_array_146010_comb[1] = p1_clipped__153_comb;
  assign p1_array_146010_comb[2] = p1_clipped__169_comb;
  assign p1_array_146010_comb[3] = p1_clipped__185_comb;
  assign p1_array_146010_comb[4] = p1_clipped__201_comb;
  assign p1_array_146010_comb[5] = p1_clipped__217_comb;
  assign p1_array_146010_comb[6] = p1_clipped__233_comb;
  assign p1_array_146010_comb[7] = p1_clipped__249_comb;
  assign p1_array_146011_comb[0] = p1_clipped__138_comb;
  assign p1_array_146011_comb[1] = p1_clipped__154_comb;
  assign p1_array_146011_comb[2] = p1_clipped__170_comb;
  assign p1_array_146011_comb[3] = p1_clipped__186_comb;
  assign p1_array_146011_comb[4] = p1_clipped__202_comb;
  assign p1_array_146011_comb[5] = p1_clipped__218_comb;
  assign p1_array_146011_comb[6] = p1_clipped__234_comb;
  assign p1_array_146011_comb[7] = p1_clipped__250_comb;
  assign p1_array_146012_comb[0] = p1_clipped__139_comb;
  assign p1_array_146012_comb[1] = p1_clipped__155_comb;
  assign p1_array_146012_comb[2] = p1_clipped__171_comb;
  assign p1_array_146012_comb[3] = p1_clipped__187_comb;
  assign p1_array_146012_comb[4] = p1_clipped__203_comb;
  assign p1_array_146012_comb[5] = p1_clipped__219_comb;
  assign p1_array_146012_comb[6] = p1_clipped__235_comb;
  assign p1_array_146012_comb[7] = p1_clipped__251_comb;
  assign p1_array_146013_comb[0] = p1_clipped__140_comb;
  assign p1_array_146013_comb[1] = p1_clipped__156_comb;
  assign p1_array_146013_comb[2] = p1_clipped__172_comb;
  assign p1_array_146013_comb[3] = p1_clipped__188_comb;
  assign p1_array_146013_comb[4] = p1_clipped__204_comb;
  assign p1_array_146013_comb[5] = p1_clipped__220_comb;
  assign p1_array_146013_comb[6] = p1_clipped__236_comb;
  assign p1_array_146013_comb[7] = p1_clipped__252_comb;
  assign p1_array_146014_comb[0] = p1_clipped__141_comb;
  assign p1_array_146014_comb[1] = p1_clipped__157_comb;
  assign p1_array_146014_comb[2] = p1_clipped__173_comb;
  assign p1_array_146014_comb[3] = p1_clipped__189_comb;
  assign p1_array_146014_comb[4] = p1_clipped__205_comb;
  assign p1_array_146014_comb[5] = p1_clipped__221_comb;
  assign p1_array_146014_comb[6] = p1_clipped__237_comb;
  assign p1_array_146014_comb[7] = p1_clipped__253_comb;
  assign p1_array_146015_comb[0] = p1_clipped__142_comb;
  assign p1_array_146015_comb[1] = p1_clipped__158_comb;
  assign p1_array_146015_comb[2] = p1_clipped__174_comb;
  assign p1_array_146015_comb[3] = p1_clipped__190_comb;
  assign p1_array_146015_comb[4] = p1_clipped__206_comb;
  assign p1_array_146015_comb[5] = p1_clipped__222_comb;
  assign p1_array_146015_comb[6] = p1_clipped__238_comb;
  assign p1_array_146015_comb[7] = p1_clipped__254_comb;
  assign p1_array_146016_comb[0] = p1_clipped__143_comb;
  assign p1_array_146016_comb[1] = p1_clipped__159_comb;
  assign p1_array_146016_comb[2] = p1_clipped__175_comb;
  assign p1_array_146016_comb[3] = p1_clipped__191_comb;
  assign p1_array_146016_comb[4] = p1_clipped__207_comb;
  assign p1_array_146016_comb[5] = p1_clipped__223_comb;
  assign p1_array_146016_comb[6] = p1_clipped__239_comb;
  assign p1_array_146016_comb[7] = p1_clipped__255_comb;
  assign p1_col_transformed_comb[0][0] = p1_array_146009_comb[0];
  assign p1_col_transformed_comb[0][1] = p1_array_146009_comb[1];
  assign p1_col_transformed_comb[0][2] = p1_array_146009_comb[2];
  assign p1_col_transformed_comb[0][3] = p1_array_146009_comb[3];
  assign p1_col_transformed_comb[0][4] = p1_array_146009_comb[4];
  assign p1_col_transformed_comb[0][5] = p1_array_146009_comb[5];
  assign p1_col_transformed_comb[0][6] = p1_array_146009_comb[6];
  assign p1_col_transformed_comb[0][7] = p1_array_146009_comb[7];
  assign p1_col_transformed_comb[1][0] = p1_array_146010_comb[0];
  assign p1_col_transformed_comb[1][1] = p1_array_146010_comb[1];
  assign p1_col_transformed_comb[1][2] = p1_array_146010_comb[2];
  assign p1_col_transformed_comb[1][3] = p1_array_146010_comb[3];
  assign p1_col_transformed_comb[1][4] = p1_array_146010_comb[4];
  assign p1_col_transformed_comb[1][5] = p1_array_146010_comb[5];
  assign p1_col_transformed_comb[1][6] = p1_array_146010_comb[6];
  assign p1_col_transformed_comb[1][7] = p1_array_146010_comb[7];
  assign p1_col_transformed_comb[2][0] = p1_array_146011_comb[0];
  assign p1_col_transformed_comb[2][1] = p1_array_146011_comb[1];
  assign p1_col_transformed_comb[2][2] = p1_array_146011_comb[2];
  assign p1_col_transformed_comb[2][3] = p1_array_146011_comb[3];
  assign p1_col_transformed_comb[2][4] = p1_array_146011_comb[4];
  assign p1_col_transformed_comb[2][5] = p1_array_146011_comb[5];
  assign p1_col_transformed_comb[2][6] = p1_array_146011_comb[6];
  assign p1_col_transformed_comb[2][7] = p1_array_146011_comb[7];
  assign p1_col_transformed_comb[3][0] = p1_array_146012_comb[0];
  assign p1_col_transformed_comb[3][1] = p1_array_146012_comb[1];
  assign p1_col_transformed_comb[3][2] = p1_array_146012_comb[2];
  assign p1_col_transformed_comb[3][3] = p1_array_146012_comb[3];
  assign p1_col_transformed_comb[3][4] = p1_array_146012_comb[4];
  assign p1_col_transformed_comb[3][5] = p1_array_146012_comb[5];
  assign p1_col_transformed_comb[3][6] = p1_array_146012_comb[6];
  assign p1_col_transformed_comb[3][7] = p1_array_146012_comb[7];
  assign p1_col_transformed_comb[4][0] = p1_array_146013_comb[0];
  assign p1_col_transformed_comb[4][1] = p1_array_146013_comb[1];
  assign p1_col_transformed_comb[4][2] = p1_array_146013_comb[2];
  assign p1_col_transformed_comb[4][3] = p1_array_146013_comb[3];
  assign p1_col_transformed_comb[4][4] = p1_array_146013_comb[4];
  assign p1_col_transformed_comb[4][5] = p1_array_146013_comb[5];
  assign p1_col_transformed_comb[4][6] = p1_array_146013_comb[6];
  assign p1_col_transformed_comb[4][7] = p1_array_146013_comb[7];
  assign p1_col_transformed_comb[5][0] = p1_array_146014_comb[0];
  assign p1_col_transformed_comb[5][1] = p1_array_146014_comb[1];
  assign p1_col_transformed_comb[5][2] = p1_array_146014_comb[2];
  assign p1_col_transformed_comb[5][3] = p1_array_146014_comb[3];
  assign p1_col_transformed_comb[5][4] = p1_array_146014_comb[4];
  assign p1_col_transformed_comb[5][5] = p1_array_146014_comb[5];
  assign p1_col_transformed_comb[5][6] = p1_array_146014_comb[6];
  assign p1_col_transformed_comb[5][7] = p1_array_146014_comb[7];
  assign p1_col_transformed_comb[6][0] = p1_array_146015_comb[0];
  assign p1_col_transformed_comb[6][1] = p1_array_146015_comb[1];
  assign p1_col_transformed_comb[6][2] = p1_array_146015_comb[2];
  assign p1_col_transformed_comb[6][3] = p1_array_146015_comb[3];
  assign p1_col_transformed_comb[6][4] = p1_array_146015_comb[4];
  assign p1_col_transformed_comb[6][5] = p1_array_146015_comb[5];
  assign p1_col_transformed_comb[6][6] = p1_array_146015_comb[6];
  assign p1_col_transformed_comb[6][7] = p1_array_146015_comb[7];
  assign p1_col_transformed_comb[7][0] = p1_array_146016_comb[0];
  assign p1_col_transformed_comb[7][1] = p1_array_146016_comb[1];
  assign p1_col_transformed_comb[7][2] = p1_array_146016_comb[2];
  assign p1_col_transformed_comb[7][3] = p1_array_146016_comb[3];
  assign p1_col_transformed_comb[7][4] = p1_array_146016_comb[4];
  assign p1_col_transformed_comb[7][5] = p1_array_146016_comb[5];
  assign p1_col_transformed_comb[7][6] = p1_array_146016_comb[6];
  assign p1_col_transformed_comb[7][7] = p1_array_146016_comb[7];

  // Registers for pipe stage 1:
  reg [7:0] p1_col_transformed[0:7][0:7];
  always @ (posedge clk) begin
    p1_col_transformed[0][0] <= p1_col_transformed_comb[0][0];
    p1_col_transformed[0][1] <= p1_col_transformed_comb[0][1];
    p1_col_transformed[0][2] <= p1_col_transformed_comb[0][2];
    p1_col_transformed[0][3] <= p1_col_transformed_comb[0][3];
    p1_col_transformed[0][4] <= p1_col_transformed_comb[0][4];
    p1_col_transformed[0][5] <= p1_col_transformed_comb[0][5];
    p1_col_transformed[0][6] <= p1_col_transformed_comb[0][6];
    p1_col_transformed[0][7] <= p1_col_transformed_comb[0][7];
    p1_col_transformed[1][0] <= p1_col_transformed_comb[1][0];
    p1_col_transformed[1][1] <= p1_col_transformed_comb[1][1];
    p1_col_transformed[1][2] <= p1_col_transformed_comb[1][2];
    p1_col_transformed[1][3] <= p1_col_transformed_comb[1][3];
    p1_col_transformed[1][4] <= p1_col_transformed_comb[1][4];
    p1_col_transformed[1][5] <= p1_col_transformed_comb[1][5];
    p1_col_transformed[1][6] <= p1_col_transformed_comb[1][6];
    p1_col_transformed[1][7] <= p1_col_transformed_comb[1][7];
    p1_col_transformed[2][0] <= p1_col_transformed_comb[2][0];
    p1_col_transformed[2][1] <= p1_col_transformed_comb[2][1];
    p1_col_transformed[2][2] <= p1_col_transformed_comb[2][2];
    p1_col_transformed[2][3] <= p1_col_transformed_comb[2][3];
    p1_col_transformed[2][4] <= p1_col_transformed_comb[2][4];
    p1_col_transformed[2][5] <= p1_col_transformed_comb[2][5];
    p1_col_transformed[2][6] <= p1_col_transformed_comb[2][6];
    p1_col_transformed[2][7] <= p1_col_transformed_comb[2][7];
    p1_col_transformed[3][0] <= p1_col_transformed_comb[3][0];
    p1_col_transformed[3][1] <= p1_col_transformed_comb[3][1];
    p1_col_transformed[3][2] <= p1_col_transformed_comb[3][2];
    p1_col_transformed[3][3] <= p1_col_transformed_comb[3][3];
    p1_col_transformed[3][4] <= p1_col_transformed_comb[3][4];
    p1_col_transformed[3][5] <= p1_col_transformed_comb[3][5];
    p1_col_transformed[3][6] <= p1_col_transformed_comb[3][6];
    p1_col_transformed[3][7] <= p1_col_transformed_comb[3][7];
    p1_col_transformed[4][0] <= p1_col_transformed_comb[4][0];
    p1_col_transformed[4][1] <= p1_col_transformed_comb[4][1];
    p1_col_transformed[4][2] <= p1_col_transformed_comb[4][2];
    p1_col_transformed[4][3] <= p1_col_transformed_comb[4][3];
    p1_col_transformed[4][4] <= p1_col_transformed_comb[4][4];
    p1_col_transformed[4][5] <= p1_col_transformed_comb[4][5];
    p1_col_transformed[4][6] <= p1_col_transformed_comb[4][6];
    p1_col_transformed[4][7] <= p1_col_transformed_comb[4][7];
    p1_col_transformed[5][0] <= p1_col_transformed_comb[5][0];
    p1_col_transformed[5][1] <= p1_col_transformed_comb[5][1];
    p1_col_transformed[5][2] <= p1_col_transformed_comb[5][2];
    p1_col_transformed[5][3] <= p1_col_transformed_comb[5][3];
    p1_col_transformed[5][4] <= p1_col_transformed_comb[5][4];
    p1_col_transformed[5][5] <= p1_col_transformed_comb[5][5];
    p1_col_transformed[5][6] <= p1_col_transformed_comb[5][6];
    p1_col_transformed[5][7] <= p1_col_transformed_comb[5][7];
    p1_col_transformed[6][0] <= p1_col_transformed_comb[6][0];
    p1_col_transformed[6][1] <= p1_col_transformed_comb[6][1];
    p1_col_transformed[6][2] <= p1_col_transformed_comb[6][2];
    p1_col_transformed[6][3] <= p1_col_transformed_comb[6][3];
    p1_col_transformed[6][4] <= p1_col_transformed_comb[6][4];
    p1_col_transformed[6][5] <= p1_col_transformed_comb[6][5];
    p1_col_transformed[6][6] <= p1_col_transformed_comb[6][6];
    p1_col_transformed[6][7] <= p1_col_transformed_comb[6][7];
    p1_col_transformed[7][0] <= p1_col_transformed_comb[7][0];
    p1_col_transformed[7][1] <= p1_col_transformed_comb[7][1];
    p1_col_transformed[7][2] <= p1_col_transformed_comb[7][2];
    p1_col_transformed[7][3] <= p1_col_transformed_comb[7][3];
    p1_col_transformed[7][4] <= p1_col_transformed_comb[7][4];
    p1_col_transformed[7][5] <= p1_col_transformed_comb[7][5];
    p1_col_transformed[7][6] <= p1_col_transformed_comb[7][6];
    p1_col_transformed[7][7] <= p1_col_transformed_comb[7][7];
  end
  assign out = {{p1_col_transformed[7][7], p1_col_transformed[7][6], p1_col_transformed[7][5], p1_col_transformed[7][4], p1_col_transformed[7][3], p1_col_transformed[7][2], p1_col_transformed[7][1], p1_col_transformed[7][0]}, {p1_col_transformed[6][7], p1_col_transformed[6][6], p1_col_transformed[6][5], p1_col_transformed[6][4], p1_col_transformed[6][3], p1_col_transformed[6][2], p1_col_transformed[6][1], p1_col_transformed[6][0]}, {p1_col_transformed[5][7], p1_col_transformed[5][6], p1_col_transformed[5][5], p1_col_transformed[5][4], p1_col_transformed[5][3], p1_col_transformed[5][2], p1_col_transformed[5][1], p1_col_transformed[5][0]}, {p1_col_transformed[4][7], p1_col_transformed[4][6], p1_col_transformed[4][5], p1_col_transformed[4][4], p1_col_transformed[4][3], p1_col_transformed[4][2], p1_col_transformed[4][1], p1_col_transformed[4][0]}, {p1_col_transformed[3][7], p1_col_transformed[3][6], p1_col_transformed[3][5], p1_col_transformed[3][4], p1_col_transformed[3][3], p1_col_transformed[3][2], p1_col_transformed[3][1], p1_col_transformed[3][0]}, {p1_col_transformed[2][7], p1_col_transformed[2][6], p1_col_transformed[2][5], p1_col_transformed[2][4], p1_col_transformed[2][3], p1_col_transformed[2][2], p1_col_transformed[2][1], p1_col_transformed[2][0]}, {p1_col_transformed[1][7], p1_col_transformed[1][6], p1_col_transformed[1][5], p1_col_transformed[1][4], p1_col_transformed[1][3], p1_col_transformed[1][2], p1_col_transformed[1][1], p1_col_transformed[1][0]}, {p1_col_transformed[0][7], p1_col_transformed[0][6], p1_col_transformed[0][5], p1_col_transformed[0][4], p1_col_transformed[0][3], p1_col_transformed[0][2], p1_col_transformed[0][1], p1_col_transformed[0][0]}};
endmodule
