module Huffman_ACenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [43:0] out
);
  wire [4:0] literal_9350[0:251];
  assign literal_9350[0] = 5'h02;
  assign literal_9350[1] = 5'h02;
  assign literal_9350[2] = 5'h03;
  assign literal_9350[3] = 5'h04;
  assign literal_9350[4] = 5'h05;
  assign literal_9350[5] = 5'h07;
  assign literal_9350[6] = 5'h08;
  assign literal_9350[7] = 5'h0e;
  assign literal_9350[8] = 5'h10;
  assign literal_9350[9] = 5'h10;
  assign literal_9350[10] = 5'h10;
  assign literal_9350[11] = 5'h00;
  assign literal_9350[12] = 5'h00;
  assign literal_9350[13] = 5'h00;
  assign literal_9350[14] = 5'h00;
  assign literal_9350[15] = 5'h00;
  assign literal_9350[16] = 5'h00;
  assign literal_9350[17] = 5'h03;
  assign literal_9350[18] = 5'h06;
  assign literal_9350[19] = 5'h07;
  assign literal_9350[20] = 5'h09;
  assign literal_9350[21] = 5'h0b;
  assign literal_9350[22] = 5'h0d;
  assign literal_9350[23] = 5'h10;
  assign literal_9350[24] = 5'h10;
  assign literal_9350[25] = 5'h10;
  assign literal_9350[26] = 5'h10;
  assign literal_9350[27] = 5'h00;
  assign literal_9350[28] = 5'h00;
  assign literal_9350[29] = 5'h00;
  assign literal_9350[30] = 5'h00;
  assign literal_9350[31] = 5'h00;
  assign literal_9350[32] = 5'h00;
  assign literal_9350[33] = 5'h05;
  assign literal_9350[34] = 5'h07;
  assign literal_9350[35] = 5'h0a;
  assign literal_9350[36] = 5'h0c;
  assign literal_9350[37] = 5'h0d;
  assign literal_9350[38] = 5'h10;
  assign literal_9350[39] = 5'h10;
  assign literal_9350[40] = 5'h10;
  assign literal_9350[41] = 5'h10;
  assign literal_9350[42] = 5'h10;
  assign literal_9350[43] = 5'h00;
  assign literal_9350[44] = 5'h00;
  assign literal_9350[45] = 5'h00;
  assign literal_9350[46] = 5'h00;
  assign literal_9350[47] = 5'h00;
  assign literal_9350[48] = 5'h00;
  assign literal_9350[49] = 5'h06;
  assign literal_9350[50] = 5'h08;
  assign literal_9350[51] = 5'h0b;
  assign literal_9350[52] = 5'h0c;
  assign literal_9350[53] = 5'h0f;
  assign literal_9350[54] = 5'h10;
  assign literal_9350[55] = 5'h10;
  assign literal_9350[56] = 5'h10;
  assign literal_9350[57] = 5'h10;
  assign literal_9350[58] = 5'h10;
  assign literal_9350[59] = 5'h00;
  assign literal_9350[60] = 5'h00;
  assign literal_9350[61] = 5'h00;
  assign literal_9350[62] = 5'h00;
  assign literal_9350[63] = 5'h00;
  assign literal_9350[64] = 5'h00;
  assign literal_9350[65] = 5'h06;
  assign literal_9350[66] = 5'h0a;
  assign literal_9350[67] = 5'h0c;
  assign literal_9350[68] = 5'h0f;
  assign literal_9350[69] = 5'h10;
  assign literal_9350[70] = 5'h10;
  assign literal_9350[71] = 5'h10;
  assign literal_9350[72] = 5'h10;
  assign literal_9350[73] = 5'h10;
  assign literal_9350[74] = 5'h10;
  assign literal_9350[75] = 5'h00;
  assign literal_9350[76] = 5'h00;
  assign literal_9350[77] = 5'h00;
  assign literal_9350[78] = 5'h00;
  assign literal_9350[79] = 5'h00;
  assign literal_9350[80] = 5'h00;
  assign literal_9350[81] = 5'h07;
  assign literal_9350[82] = 5'h0b;
  assign literal_9350[83] = 5'h0d;
  assign literal_9350[84] = 5'h10;
  assign literal_9350[85] = 5'h10;
  assign literal_9350[86] = 5'h10;
  assign literal_9350[87] = 5'h10;
  assign literal_9350[88] = 5'h10;
  assign literal_9350[89] = 5'h10;
  assign literal_9350[90] = 5'h10;
  assign literal_9350[91] = 5'h00;
  assign literal_9350[92] = 5'h00;
  assign literal_9350[93] = 5'h00;
  assign literal_9350[94] = 5'h00;
  assign literal_9350[95] = 5'h00;
  assign literal_9350[96] = 5'h00;
  assign literal_9350[97] = 5'h07;
  assign literal_9350[98] = 5'h0b;
  assign literal_9350[99] = 5'h0d;
  assign literal_9350[100] = 5'h10;
  assign literal_9350[101] = 5'h10;
  assign literal_9350[102] = 5'h10;
  assign literal_9350[103] = 5'h10;
  assign literal_9350[104] = 5'h10;
  assign literal_9350[105] = 5'h10;
  assign literal_9350[106] = 5'h10;
  assign literal_9350[107] = 5'h00;
  assign literal_9350[108] = 5'h00;
  assign literal_9350[109] = 5'h00;
  assign literal_9350[110] = 5'h00;
  assign literal_9350[111] = 5'h00;
  assign literal_9350[112] = 5'h00;
  assign literal_9350[113] = 5'h08;
  assign literal_9350[114] = 5'h0b;
  assign literal_9350[115] = 5'h0e;
  assign literal_9350[116] = 5'h10;
  assign literal_9350[117] = 5'h10;
  assign literal_9350[118] = 5'h10;
  assign literal_9350[119] = 5'h10;
  assign literal_9350[120] = 5'h10;
  assign literal_9350[121] = 5'h10;
  assign literal_9350[122] = 5'h10;
  assign literal_9350[123] = 5'h00;
  assign literal_9350[124] = 5'h00;
  assign literal_9350[125] = 5'h00;
  assign literal_9350[126] = 5'h00;
  assign literal_9350[127] = 5'h00;
  assign literal_9350[128] = 5'h00;
  assign literal_9350[129] = 5'h08;
  assign literal_9350[130] = 5'h0c;
  assign literal_9350[131] = 5'h10;
  assign literal_9350[132] = 5'h10;
  assign literal_9350[133] = 5'h10;
  assign literal_9350[134] = 5'h10;
  assign literal_9350[135] = 5'h10;
  assign literal_9350[136] = 5'h10;
  assign literal_9350[137] = 5'h10;
  assign literal_9350[138] = 5'h10;
  assign literal_9350[139] = 5'h00;
  assign literal_9350[140] = 5'h00;
  assign literal_9350[141] = 5'h00;
  assign literal_9350[142] = 5'h00;
  assign literal_9350[143] = 5'h00;
  assign literal_9350[144] = 5'h00;
  assign literal_9350[145] = 5'h08;
  assign literal_9350[146] = 5'h0d;
  assign literal_9350[147] = 5'h10;
  assign literal_9350[148] = 5'h10;
  assign literal_9350[149] = 5'h10;
  assign literal_9350[150] = 5'h10;
  assign literal_9350[151] = 5'h10;
  assign literal_9350[152] = 5'h10;
  assign literal_9350[153] = 5'h10;
  assign literal_9350[154] = 5'h10;
  assign literal_9350[155] = 5'h00;
  assign literal_9350[156] = 5'h00;
  assign literal_9350[157] = 5'h00;
  assign literal_9350[158] = 5'h00;
  assign literal_9350[159] = 5'h00;
  assign literal_9350[160] = 5'h00;
  assign literal_9350[161] = 5'h09;
  assign literal_9350[162] = 5'h0d;
  assign literal_9350[163] = 5'h10;
  assign literal_9350[164] = 5'h10;
  assign literal_9350[165] = 5'h10;
  assign literal_9350[166] = 5'h10;
  assign literal_9350[167] = 5'h10;
  assign literal_9350[168] = 5'h10;
  assign literal_9350[169] = 5'h10;
  assign literal_9350[170] = 5'h10;
  assign literal_9350[171] = 5'h00;
  assign literal_9350[172] = 5'h00;
  assign literal_9350[173] = 5'h00;
  assign literal_9350[174] = 5'h00;
  assign literal_9350[175] = 5'h00;
  assign literal_9350[176] = 5'h00;
  assign literal_9350[177] = 5'h09;
  assign literal_9350[178] = 5'h0d;
  assign literal_9350[179] = 5'h10;
  assign literal_9350[180] = 5'h10;
  assign literal_9350[181] = 5'h10;
  assign literal_9350[182] = 5'h10;
  assign literal_9350[183] = 5'h10;
  assign literal_9350[184] = 5'h10;
  assign literal_9350[185] = 5'h10;
  assign literal_9350[186] = 5'h10;
  assign literal_9350[187] = 5'h00;
  assign literal_9350[188] = 5'h00;
  assign literal_9350[189] = 5'h00;
  assign literal_9350[190] = 5'h00;
  assign literal_9350[191] = 5'h00;
  assign literal_9350[192] = 5'h00;
  assign literal_9350[193] = 5'h0a;
  assign literal_9350[194] = 5'h0d;
  assign literal_9350[195] = 5'h10;
  assign literal_9350[196] = 5'h10;
  assign literal_9350[197] = 5'h10;
  assign literal_9350[198] = 5'h10;
  assign literal_9350[199] = 5'h10;
  assign literal_9350[200] = 5'h10;
  assign literal_9350[201] = 5'h10;
  assign literal_9350[202] = 5'h10;
  assign literal_9350[203] = 5'h00;
  assign literal_9350[204] = 5'h00;
  assign literal_9350[205] = 5'h00;
  assign literal_9350[206] = 5'h00;
  assign literal_9350[207] = 5'h00;
  assign literal_9350[208] = 5'h00;
  assign literal_9350[209] = 5'h0a;
  assign literal_9350[210] = 5'h0e;
  assign literal_9350[211] = 5'h10;
  assign literal_9350[212] = 5'h10;
  assign literal_9350[213] = 5'h10;
  assign literal_9350[214] = 5'h10;
  assign literal_9350[215] = 5'h10;
  assign literal_9350[216] = 5'h10;
  assign literal_9350[217] = 5'h10;
  assign literal_9350[218] = 5'h10;
  assign literal_9350[219] = 5'h00;
  assign literal_9350[220] = 5'h00;
  assign literal_9350[221] = 5'h00;
  assign literal_9350[222] = 5'h00;
  assign literal_9350[223] = 5'h00;
  assign literal_9350[224] = 5'h00;
  assign literal_9350[225] = 5'h0a;
  assign literal_9350[226] = 5'h0f;
  assign literal_9350[227] = 5'h10;
  assign literal_9350[228] = 5'h10;
  assign literal_9350[229] = 5'h10;
  assign literal_9350[230] = 5'h10;
  assign literal_9350[231] = 5'h10;
  assign literal_9350[232] = 5'h10;
  assign literal_9350[233] = 5'h10;
  assign literal_9350[234] = 5'h10;
  assign literal_9350[235] = 5'h00;
  assign literal_9350[236] = 5'h00;
  assign literal_9350[237] = 5'h00;
  assign literal_9350[238] = 5'h00;
  assign literal_9350[239] = 5'h00;
  assign literal_9350[240] = 5'h09;
  assign literal_9350[241] = 5'h0b;
  assign literal_9350[242] = 5'h10;
  assign literal_9350[243] = 5'h10;
  assign literal_9350[244] = 5'h10;
  assign literal_9350[245] = 5'h10;
  assign literal_9350[246] = 5'h10;
  assign literal_9350[247] = 5'h10;
  assign literal_9350[248] = 5'h10;
  assign literal_9350[249] = 5'h10;
  assign literal_9350[250] = 5'h10;
  assign literal_9350[251] = 5'h00;
  wire [4:0] literal_9352[0:251];
  assign literal_9352[0] = 5'h04;
  assign literal_9352[1] = 5'h02;
  assign literal_9352[2] = 5'h02;
  assign literal_9352[3] = 5'h03;
  assign literal_9352[4] = 5'h04;
  assign literal_9352[5] = 5'h05;
  assign literal_9352[6] = 5'h07;
  assign literal_9352[7] = 5'h09;
  assign literal_9352[8] = 5'h10;
  assign literal_9352[9] = 5'h10;
  assign literal_9352[10] = 5'h10;
  assign literal_9352[11] = 5'h00;
  assign literal_9352[12] = 5'h00;
  assign literal_9352[13] = 5'h00;
  assign literal_9352[14] = 5'h00;
  assign literal_9352[15] = 5'h00;
  assign literal_9352[16] = 5'h00;
  assign literal_9352[17] = 5'h04;
  assign literal_9352[18] = 5'h05;
  assign literal_9352[19] = 5'h07;
  assign literal_9352[20] = 5'h09;
  assign literal_9352[21] = 5'h0a;
  assign literal_9352[22] = 5'h0b;
  assign literal_9352[23] = 5'h10;
  assign literal_9352[24] = 5'h10;
  assign literal_9352[25] = 5'h10;
  assign literal_9352[26] = 5'h10;
  assign literal_9352[27] = 5'h00;
  assign literal_9352[28] = 5'h00;
  assign literal_9352[29] = 5'h00;
  assign literal_9352[30] = 5'h00;
  assign literal_9352[31] = 5'h00;
  assign literal_9352[32] = 5'h00;
  assign literal_9352[33] = 5'h05;
  assign literal_9352[34] = 5'h08;
  assign literal_9352[35] = 5'h0a;
  assign literal_9352[36] = 5'h0c;
  assign literal_9352[37] = 5'h0e;
  assign literal_9352[38] = 5'h10;
  assign literal_9352[39] = 5'h10;
  assign literal_9352[40] = 5'h10;
  assign literal_9352[41] = 5'h10;
  assign literal_9352[42] = 5'h10;
  assign literal_9352[43] = 5'h00;
  assign literal_9352[44] = 5'h00;
  assign literal_9352[45] = 5'h00;
  assign literal_9352[46] = 5'h00;
  assign literal_9352[47] = 5'h00;
  assign literal_9352[48] = 5'h00;
  assign literal_9352[49] = 5'h06;
  assign literal_9352[50] = 5'h09;
  assign literal_9352[51] = 5'h0b;
  assign literal_9352[52] = 5'h0e;
  assign literal_9352[53] = 5'h10;
  assign literal_9352[54] = 5'h10;
  assign literal_9352[55] = 5'h10;
  assign literal_9352[56] = 5'h10;
  assign literal_9352[57] = 5'h10;
  assign literal_9352[58] = 5'h10;
  assign literal_9352[59] = 5'h00;
  assign literal_9352[60] = 5'h00;
  assign literal_9352[61] = 5'h00;
  assign literal_9352[62] = 5'h00;
  assign literal_9352[63] = 5'h00;
  assign literal_9352[64] = 5'h00;
  assign literal_9352[65] = 5'h06;
  assign literal_9352[66] = 5'h0a;
  assign literal_9352[67] = 5'h0e;
  assign literal_9352[68] = 5'h10;
  assign literal_9352[69] = 5'h10;
  assign literal_9352[70] = 5'h10;
  assign literal_9352[71] = 5'h10;
  assign literal_9352[72] = 5'h10;
  assign literal_9352[73] = 5'h10;
  assign literal_9352[74] = 5'h10;
  assign literal_9352[75] = 5'h00;
  assign literal_9352[76] = 5'h00;
  assign literal_9352[77] = 5'h00;
  assign literal_9352[78] = 5'h00;
  assign literal_9352[79] = 5'h00;
  assign literal_9352[80] = 5'h00;
  assign literal_9352[81] = 5'h07;
  assign literal_9352[82] = 5'h0a;
  assign literal_9352[83] = 5'h0e;
  assign literal_9352[84] = 5'h10;
  assign literal_9352[85] = 5'h10;
  assign literal_9352[86] = 5'h10;
  assign literal_9352[87] = 5'h10;
  assign literal_9352[88] = 5'h10;
  assign literal_9352[89] = 5'h10;
  assign literal_9352[90] = 5'h10;
  assign literal_9352[91] = 5'h00;
  assign literal_9352[92] = 5'h00;
  assign literal_9352[93] = 5'h00;
  assign literal_9352[94] = 5'h00;
  assign literal_9352[95] = 5'h00;
  assign literal_9352[96] = 5'h00;
  assign literal_9352[97] = 5'h07;
  assign literal_9352[98] = 5'h0c;
  assign literal_9352[99] = 5'h0f;
  assign literal_9352[100] = 5'h10;
  assign literal_9352[101] = 5'h10;
  assign literal_9352[102] = 5'h10;
  assign literal_9352[103] = 5'h10;
  assign literal_9352[104] = 5'h10;
  assign literal_9352[105] = 5'h10;
  assign literal_9352[106] = 5'h10;
  assign literal_9352[107] = 5'h00;
  assign literal_9352[108] = 5'h00;
  assign literal_9352[109] = 5'h00;
  assign literal_9352[110] = 5'h00;
  assign literal_9352[111] = 5'h00;
  assign literal_9352[112] = 5'h00;
  assign literal_9352[113] = 5'h08;
  assign literal_9352[114] = 5'h0c;
  assign literal_9352[115] = 5'h10;
  assign literal_9352[116] = 5'h10;
  assign literal_9352[117] = 5'h10;
  assign literal_9352[118] = 5'h10;
  assign literal_9352[119] = 5'h10;
  assign literal_9352[120] = 5'h10;
  assign literal_9352[121] = 5'h10;
  assign literal_9352[122] = 5'h10;
  assign literal_9352[123] = 5'h00;
  assign literal_9352[124] = 5'h00;
  assign literal_9352[125] = 5'h00;
  assign literal_9352[126] = 5'h00;
  assign literal_9352[127] = 5'h00;
  assign literal_9352[128] = 5'h00;
  assign literal_9352[129] = 5'h09;
  assign literal_9352[130] = 5'h0d;
  assign literal_9352[131] = 5'h10;
  assign literal_9352[132] = 5'h10;
  assign literal_9352[133] = 5'h10;
  assign literal_9352[134] = 5'h10;
  assign literal_9352[135] = 5'h10;
  assign literal_9352[136] = 5'h10;
  assign literal_9352[137] = 5'h10;
  assign literal_9352[138] = 5'h10;
  assign literal_9352[139] = 5'h00;
  assign literal_9352[140] = 5'h00;
  assign literal_9352[141] = 5'h00;
  assign literal_9352[142] = 5'h00;
  assign literal_9352[143] = 5'h00;
  assign literal_9352[144] = 5'h00;
  assign literal_9352[145] = 5'h09;
  assign literal_9352[146] = 5'h0e;
  assign literal_9352[147] = 5'h10;
  assign literal_9352[148] = 5'h10;
  assign literal_9352[149] = 5'h10;
  assign literal_9352[150] = 5'h10;
  assign literal_9352[151] = 5'h10;
  assign literal_9352[152] = 5'h10;
  assign literal_9352[153] = 5'h10;
  assign literal_9352[154] = 5'h10;
  assign literal_9352[155] = 5'h00;
  assign literal_9352[156] = 5'h00;
  assign literal_9352[157] = 5'h00;
  assign literal_9352[158] = 5'h00;
  assign literal_9352[159] = 5'h00;
  assign literal_9352[160] = 5'h00;
  assign literal_9352[161] = 5'h09;
  assign literal_9352[162] = 5'h0e;
  assign literal_9352[163] = 5'h10;
  assign literal_9352[164] = 5'h10;
  assign literal_9352[165] = 5'h10;
  assign literal_9352[166] = 5'h10;
  assign literal_9352[167] = 5'h10;
  assign literal_9352[168] = 5'h10;
  assign literal_9352[169] = 5'h10;
  assign literal_9352[170] = 5'h10;
  assign literal_9352[171] = 5'h00;
  assign literal_9352[172] = 5'h00;
  assign literal_9352[173] = 5'h00;
  assign literal_9352[174] = 5'h00;
  assign literal_9352[175] = 5'h00;
  assign literal_9352[176] = 5'h00;
  assign literal_9352[177] = 5'h0a;
  assign literal_9352[178] = 5'h0f;
  assign literal_9352[179] = 5'h10;
  assign literal_9352[180] = 5'h10;
  assign literal_9352[181] = 5'h10;
  assign literal_9352[182] = 5'h10;
  assign literal_9352[183] = 5'h10;
  assign literal_9352[184] = 5'h10;
  assign literal_9352[185] = 5'h10;
  assign literal_9352[186] = 5'h10;
  assign literal_9352[187] = 5'h00;
  assign literal_9352[188] = 5'h00;
  assign literal_9352[189] = 5'h00;
  assign literal_9352[190] = 5'h00;
  assign literal_9352[191] = 5'h00;
  assign literal_9352[192] = 5'h00;
  assign literal_9352[193] = 5'h0a;
  assign literal_9352[194] = 5'h10;
  assign literal_9352[195] = 5'h10;
  assign literal_9352[196] = 5'h10;
  assign literal_9352[197] = 5'h10;
  assign literal_9352[198] = 5'h10;
  assign literal_9352[199] = 5'h10;
  assign literal_9352[200] = 5'h10;
  assign literal_9352[201] = 5'h10;
  assign literal_9352[202] = 5'h10;
  assign literal_9352[203] = 5'h00;
  assign literal_9352[204] = 5'h00;
  assign literal_9352[205] = 5'h00;
  assign literal_9352[206] = 5'h00;
  assign literal_9352[207] = 5'h00;
  assign literal_9352[208] = 5'h00;
  assign literal_9352[209] = 5'h0a;
  assign literal_9352[210] = 5'h10;
  assign literal_9352[211] = 5'h10;
  assign literal_9352[212] = 5'h10;
  assign literal_9352[213] = 5'h10;
  assign literal_9352[214] = 5'h10;
  assign literal_9352[215] = 5'h10;
  assign literal_9352[216] = 5'h10;
  assign literal_9352[217] = 5'h10;
  assign literal_9352[218] = 5'h10;
  assign literal_9352[219] = 5'h00;
  assign literal_9352[220] = 5'h00;
  assign literal_9352[221] = 5'h00;
  assign literal_9352[222] = 5'h00;
  assign literal_9352[223] = 5'h00;
  assign literal_9352[224] = 5'h00;
  assign literal_9352[225] = 5'h0b;
  assign literal_9352[226] = 5'h10;
  assign literal_9352[227] = 5'h10;
  assign literal_9352[228] = 5'h10;
  assign literal_9352[229] = 5'h10;
  assign literal_9352[230] = 5'h10;
  assign literal_9352[231] = 5'h10;
  assign literal_9352[232] = 5'h10;
  assign literal_9352[233] = 5'h10;
  assign literal_9352[234] = 5'h10;
  assign literal_9352[235] = 5'h00;
  assign literal_9352[236] = 5'h00;
  assign literal_9352[237] = 5'h00;
  assign literal_9352[238] = 5'h00;
  assign literal_9352[239] = 5'h00;
  assign literal_9352[240] = 5'h0c;
  assign literal_9352[241] = 5'h0d;
  assign literal_9352[242] = 5'h10;
  assign literal_9352[243] = 5'h10;
  assign literal_9352[244] = 5'h10;
  assign literal_9352[245] = 5'h10;
  assign literal_9352[246] = 5'h10;
  assign literal_9352[247] = 5'h10;
  assign literal_9352[248] = 5'h10;
  assign literal_9352[249] = 5'h10;
  assign literal_9352[250] = 5'h10;
  assign literal_9352[251] = 5'h00;
  wire [15:0] literal_9355[0:251];
  assign literal_9355[0] = 16'h0001;
  assign literal_9355[1] = 16'h0000;
  assign literal_9355[2] = 16'h0004;
  assign literal_9355[3] = 16'h000c;
  assign literal_9355[4] = 16'h001a;
  assign literal_9355[5] = 16'h0076;
  assign literal_9355[6] = 16'h00f6;
  assign literal_9355[7] = 16'h3fe0;
  assign literal_9355[8] = 16'hff96;
  assign literal_9355[9] = 16'hff97;
  assign literal_9355[10] = 16'hff98;
  assign literal_9355[11] = 16'h0000;
  assign literal_9355[12] = 16'h0000;
  assign literal_9355[13] = 16'h0000;
  assign literal_9355[14] = 16'h0000;
  assign literal_9355[15] = 16'h0000;
  assign literal_9355[16] = 16'h0000;
  assign literal_9355[17] = 16'h0005;
  assign literal_9355[18] = 16'h0038;
  assign literal_9355[19] = 16'h0078;
  assign literal_9355[20] = 16'h01f9;
  assign literal_9355[21] = 16'h07f2;
  assign literal_9355[22] = 16'h1fe8;
  assign literal_9355[23] = 16'hff93;
  assign literal_9355[24] = 16'hff99;
  assign literal_9355[25] = 16'hff9a;
  assign literal_9355[26] = 16'hff9e;
  assign literal_9355[27] = 16'h0000;
  assign literal_9355[28] = 16'h0000;
  assign literal_9355[29] = 16'h0000;
  assign literal_9355[30] = 16'h0000;
  assign literal_9355[31] = 16'h0000;
  assign literal_9355[32] = 16'h0000;
  assign literal_9355[33] = 16'h001b;
  assign literal_9355[34] = 16'h007a;
  assign literal_9355[35] = 16'h03f7;
  assign literal_9355[36] = 16'h0ff0;
  assign literal_9355[37] = 16'h1feb;
  assign literal_9355[38] = 16'hff9b;
  assign literal_9355[39] = 16'hff9f;
  assign literal_9355[40] = 16'hffa8;
  assign literal_9355[41] = 16'hffa9;
  assign literal_9355[42] = 16'hfff1;
  assign literal_9355[43] = 16'h0000;
  assign literal_9355[44] = 16'h0000;
  assign literal_9355[45] = 16'h0000;
  assign literal_9355[46] = 16'h0000;
  assign literal_9355[47] = 16'h0000;
  assign literal_9355[48] = 16'h0000;
  assign literal_9355[49] = 16'h0039;
  assign literal_9355[50] = 16'h00fa;
  assign literal_9355[51] = 16'h07f7;
  assign literal_9355[52] = 16'h0ff1;
  assign literal_9355[53] = 16'h7fc6;
  assign literal_9355[54] = 16'hff9c;
  assign literal_9355[55] = 16'hffa3;
  assign literal_9355[56] = 16'hffd7;
  assign literal_9355[57] = 16'hffe4;
  assign literal_9355[58] = 16'hfff2;
  assign literal_9355[59] = 16'h0000;
  assign literal_9355[60] = 16'h0000;
  assign literal_9355[61] = 16'h0000;
  assign literal_9355[62] = 16'h0000;
  assign literal_9355[63] = 16'h0000;
  assign literal_9355[64] = 16'h0000;
  assign literal_9355[65] = 16'h003a;
  assign literal_9355[66] = 16'h03f8;
  assign literal_9355[67] = 16'h0ff2;
  assign literal_9355[68] = 16'h7fc8;
  assign literal_9355[69] = 16'hff9d;
  assign literal_9355[70] = 16'hffbf;
  assign literal_9355[71] = 16'hffcb;
  assign literal_9355[72] = 16'hffd8;
  assign literal_9355[73] = 16'hffe5;
  assign literal_9355[74] = 16'hfff3;
  assign literal_9355[75] = 16'h0000;
  assign literal_9355[76] = 16'h0000;
  assign literal_9355[77] = 16'h0000;
  assign literal_9355[78] = 16'h0000;
  assign literal_9355[79] = 16'h0000;
  assign literal_9355[80] = 16'h0000;
  assign literal_9355[81] = 16'h0077;
  assign literal_9355[82] = 16'h07f3;
  assign literal_9355[83] = 16'h1fea;
  assign literal_9355[84] = 16'hff94;
  assign literal_9355[85] = 16'hffa2;
  assign literal_9355[86] = 16'hffc0;
  assign literal_9355[87] = 16'hffcc;
  assign literal_9355[88] = 16'hffd9;
  assign literal_9355[89] = 16'hffe6;
  assign literal_9355[90] = 16'hfff4;
  assign literal_9355[91] = 16'h0000;
  assign literal_9355[92] = 16'h0000;
  assign literal_9355[93] = 16'h0000;
  assign literal_9355[94] = 16'h0000;
  assign literal_9355[95] = 16'h0000;
  assign literal_9355[96] = 16'h0000;
  assign literal_9355[97] = 16'h0079;
  assign literal_9355[98] = 16'h07f4;
  assign literal_9355[99] = 16'h1fed;
  assign literal_9355[100] = 16'hffa0;
  assign literal_9355[101] = 16'hffb5;
  assign literal_9355[102] = 16'hffc1;
  assign literal_9355[103] = 16'hffcd;
  assign literal_9355[104] = 16'hffda;
  assign literal_9355[105] = 16'hffe7;
  assign literal_9355[106] = 16'hfff5;
  assign literal_9355[107] = 16'h0000;
  assign literal_9355[108] = 16'h0000;
  assign literal_9355[109] = 16'h0000;
  assign literal_9355[110] = 16'h0000;
  assign literal_9355[111] = 16'h0000;
  assign literal_9355[112] = 16'h0000;
  assign literal_9355[113] = 16'h00f7;
  assign literal_9355[114] = 16'h07f5;
  assign literal_9355[115] = 16'h3fe1;
  assign literal_9355[116] = 16'hffa1;
  assign literal_9355[117] = 16'hffb6;
  assign literal_9355[118] = 16'hffc2;
  assign literal_9355[119] = 16'hffce;
  assign literal_9355[120] = 16'hffdb;
  assign literal_9355[121] = 16'hffe8;
  assign literal_9355[122] = 16'hfff6;
  assign literal_9355[123] = 16'h0000;
  assign literal_9355[124] = 16'h0000;
  assign literal_9355[125] = 16'h0000;
  assign literal_9355[126] = 16'h0000;
  assign literal_9355[127] = 16'h0000;
  assign literal_9355[128] = 16'h0000;
  assign literal_9355[129] = 16'h00f8;
  assign literal_9355[130] = 16'h0ff3;
  assign literal_9355[131] = 16'hff92;
  assign literal_9355[132] = 16'hffad;
  assign literal_9355[133] = 16'hffb7;
  assign literal_9355[134] = 16'hffc3;
  assign literal_9355[135] = 16'hffcf;
  assign literal_9355[136] = 16'hffdc;
  assign literal_9355[137] = 16'hffe9;
  assign literal_9355[138] = 16'hfff7;
  assign literal_9355[139] = 16'h0000;
  assign literal_9355[140] = 16'h0000;
  assign literal_9355[141] = 16'h0000;
  assign literal_9355[142] = 16'h0000;
  assign literal_9355[143] = 16'h0000;
  assign literal_9355[144] = 16'h0000;
  assign literal_9355[145] = 16'h00f9;
  assign literal_9355[146] = 16'h1fe9;
  assign literal_9355[147] = 16'hff95;
  assign literal_9355[148] = 16'hffae;
  assign literal_9355[149] = 16'hffb8;
  assign literal_9355[150] = 16'hffc4;
  assign literal_9355[151] = 16'hffd0;
  assign literal_9355[152] = 16'hffdd;
  assign literal_9355[153] = 16'hffea;
  assign literal_9355[154] = 16'hfff8;
  assign literal_9355[155] = 16'h0000;
  assign literal_9355[156] = 16'h0000;
  assign literal_9355[157] = 16'h0000;
  assign literal_9355[158] = 16'h0000;
  assign literal_9355[159] = 16'h0000;
  assign literal_9355[160] = 16'h0000;
  assign literal_9355[161] = 16'h01f6;
  assign literal_9355[162] = 16'h1fec;
  assign literal_9355[163] = 16'hffa5;
  assign literal_9355[164] = 16'hffaf;
  assign literal_9355[165] = 16'hffb9;
  assign literal_9355[166] = 16'hffc5;
  assign literal_9355[167] = 16'hffd1;
  assign literal_9355[168] = 16'hffde;
  assign literal_9355[169] = 16'hffeb;
  assign literal_9355[170] = 16'hfff9;
  assign literal_9355[171] = 16'h0000;
  assign literal_9355[172] = 16'h0000;
  assign literal_9355[173] = 16'h0000;
  assign literal_9355[174] = 16'h0000;
  assign literal_9355[175] = 16'h0000;
  assign literal_9355[176] = 16'h0000;
  assign literal_9355[177] = 16'h01f7;
  assign literal_9355[178] = 16'h1fee;
  assign literal_9355[179] = 16'hffa6;
  assign literal_9355[180] = 16'hffb0;
  assign literal_9355[181] = 16'hffba;
  assign literal_9355[182] = 16'hffc6;
  assign literal_9355[183] = 16'hffd2;
  assign literal_9355[184] = 16'hffdf;
  assign literal_9355[185] = 16'hffec;
  assign literal_9355[186] = 16'hfffa;
  assign literal_9355[187] = 16'h0000;
  assign literal_9355[188] = 16'h0000;
  assign literal_9355[189] = 16'h0000;
  assign literal_9355[190] = 16'h0000;
  assign literal_9355[191] = 16'h0000;
  assign literal_9355[192] = 16'h0000;
  assign literal_9355[193] = 16'h03f4;
  assign literal_9355[194] = 16'h1fef;
  assign literal_9355[195] = 16'hffa7;
  assign literal_9355[196] = 16'hffb1;
  assign literal_9355[197] = 16'hffbb;
  assign literal_9355[198] = 16'hffc7;
  assign literal_9355[199] = 16'hffd3;
  assign literal_9355[200] = 16'hffe0;
  assign literal_9355[201] = 16'hffed;
  assign literal_9355[202] = 16'hfffb;
  assign literal_9355[203] = 16'h0000;
  assign literal_9355[204] = 16'h0000;
  assign literal_9355[205] = 16'h0000;
  assign literal_9355[206] = 16'h0000;
  assign literal_9355[207] = 16'h0000;
  assign literal_9355[208] = 16'h0000;
  assign literal_9355[209] = 16'h03f5;
  assign literal_9355[210] = 16'h3fe2;
  assign literal_9355[211] = 16'hffaa;
  assign literal_9355[212] = 16'hffb2;
  assign literal_9355[213] = 16'hffbc;
  assign literal_9355[214] = 16'hffc8;
  assign literal_9355[215] = 16'hffd4;
  assign literal_9355[216] = 16'hffe1;
  assign literal_9355[217] = 16'hffee;
  assign literal_9355[218] = 16'hfffc;
  assign literal_9355[219] = 16'h0000;
  assign literal_9355[220] = 16'h0000;
  assign literal_9355[221] = 16'h0000;
  assign literal_9355[222] = 16'h0000;
  assign literal_9355[223] = 16'h0000;
  assign literal_9355[224] = 16'h0000;
  assign literal_9355[225] = 16'h03f6;
  assign literal_9355[226] = 16'h7fc7;
  assign literal_9355[227] = 16'hffab;
  assign literal_9355[228] = 16'hffb3;
  assign literal_9355[229] = 16'hffbd;
  assign literal_9355[230] = 16'hffc9;
  assign literal_9355[231] = 16'hffd5;
  assign literal_9355[232] = 16'hffe2;
  assign literal_9355[233] = 16'hffef;
  assign literal_9355[234] = 16'hfffd;
  assign literal_9355[235] = 16'h0000;
  assign literal_9355[236] = 16'h0000;
  assign literal_9355[237] = 16'h0000;
  assign literal_9355[238] = 16'h0000;
  assign literal_9355[239] = 16'h0000;
  assign literal_9355[240] = 16'h01f8;
  assign literal_9355[241] = 16'h07f6;
  assign literal_9355[242] = 16'hffa4;
  assign literal_9355[243] = 16'hffac;
  assign literal_9355[244] = 16'hffb4;
  assign literal_9355[245] = 16'hffbe;
  assign literal_9355[246] = 16'hffca;
  assign literal_9355[247] = 16'hffd6;
  assign literal_9355[248] = 16'hffe3;
  assign literal_9355[249] = 16'hfff0;
  assign literal_9355[250] = 16'hfffe;
  assign literal_9355[251] = 16'h0000;
  wire [15:0] literal_9356[0:251];
  assign literal_9356[0] = 16'h000c;
  assign literal_9356[1] = 16'h0000;
  assign literal_9356[2] = 16'h0001;
  assign literal_9356[3] = 16'h0004;
  assign literal_9356[4] = 16'h000b;
  assign literal_9356[5] = 16'h001a;
  assign literal_9356[6] = 16'h0079;
  assign literal_9356[7] = 16'h01f9;
  assign literal_9356[8] = 16'hff9c;
  assign literal_9356[9] = 16'hff9f;
  assign literal_9356[10] = 16'hffa0;
  assign literal_9356[11] = 16'h0000;
  assign literal_9356[12] = 16'h0000;
  assign literal_9356[13] = 16'h0000;
  assign literal_9356[14] = 16'h0000;
  assign literal_9356[15] = 16'h0000;
  assign literal_9356[16] = 16'h0000;
  assign literal_9356[17] = 16'h000a;
  assign literal_9356[18] = 16'h001c;
  assign literal_9356[19] = 16'h007a;
  assign literal_9356[20] = 16'h01f5;
  assign literal_9356[21] = 16'h03f4;
  assign literal_9356[22] = 16'h07f8;
  assign literal_9356[23] = 16'hff95;
  assign literal_9356[24] = 16'hffa1;
  assign literal_9356[25] = 16'hffa2;
  assign literal_9356[26] = 16'hffad;
  assign literal_9356[27] = 16'h0000;
  assign literal_9356[28] = 16'h0000;
  assign literal_9356[29] = 16'h0000;
  assign literal_9356[30] = 16'h0000;
  assign literal_9356[31] = 16'h0000;
  assign literal_9356[32] = 16'h0000;
  assign literal_9356[33] = 16'h001b;
  assign literal_9356[34] = 16'h00f8;
  assign literal_9356[35] = 16'h03f7;
  assign literal_9356[36] = 16'h0ff4;
  assign literal_9356[37] = 16'h3fdc;
  assign literal_9356[38] = 16'hff9d;
  assign literal_9356[39] = 16'hff90;
  assign literal_9356[40] = 16'hffac;
  assign literal_9356[41] = 16'hffe3;
  assign literal_9356[42] = 16'hfff1;
  assign literal_9356[43] = 16'h0000;
  assign literal_9356[44] = 16'h0000;
  assign literal_9356[45] = 16'h0000;
  assign literal_9356[46] = 16'h0000;
  assign literal_9356[47] = 16'h0000;
  assign literal_9356[48] = 16'h0000;
  assign literal_9356[49] = 16'h003a;
  assign literal_9356[50] = 16'h01f6;
  assign literal_9356[51] = 16'h07f7;
  assign literal_9356[52] = 16'h3fde;
  assign literal_9356[53] = 16'hff8e;
  assign literal_9356[54] = 16'hff94;
  assign literal_9356[55] = 16'hffc9;
  assign literal_9356[56] = 16'hffd6;
  assign literal_9356[57] = 16'hffe4;
  assign literal_9356[58] = 16'hfff2;
  assign literal_9356[59] = 16'h0000;
  assign literal_9356[60] = 16'h0000;
  assign literal_9356[61] = 16'h0000;
  assign literal_9356[62] = 16'h0000;
  assign literal_9356[63] = 16'h0000;
  assign literal_9356[64] = 16'h0000;
  assign literal_9356[65] = 16'h003b;
  assign literal_9356[66] = 16'h03f6;
  assign literal_9356[67] = 16'h3fdd;
  assign literal_9356[68] = 16'hff8f;
  assign literal_9356[69] = 16'hffa5;
  assign literal_9356[70] = 16'hffa6;
  assign literal_9356[71] = 16'hffca;
  assign literal_9356[72] = 16'hffd7;
  assign literal_9356[73] = 16'hffe5;
  assign literal_9356[74] = 16'hfff3;
  assign literal_9356[75] = 16'h0000;
  assign literal_9356[76] = 16'h0000;
  assign literal_9356[77] = 16'h0000;
  assign literal_9356[78] = 16'h0000;
  assign literal_9356[79] = 16'h0000;
  assign literal_9356[80] = 16'h0000;
  assign literal_9356[81] = 16'h0078;
  assign literal_9356[82] = 16'h03f9;
  assign literal_9356[83] = 16'h3fdf;
  assign literal_9356[84] = 16'hff96;
  assign literal_9356[85] = 16'hffab;
  assign literal_9356[86] = 16'hffa9;
  assign literal_9356[87] = 16'hffcb;
  assign literal_9356[88] = 16'hffd8;
  assign literal_9356[89] = 16'hffe6;
  assign literal_9356[90] = 16'hfff4;
  assign literal_9356[91] = 16'h0000;
  assign literal_9356[92] = 16'h0000;
  assign literal_9356[93] = 16'h0000;
  assign literal_9356[94] = 16'h0000;
  assign literal_9356[95] = 16'h0000;
  assign literal_9356[96] = 16'h0000;
  assign literal_9356[97] = 16'h007b;
  assign literal_9356[98] = 16'h0ff2;
  assign literal_9356[99] = 16'h7fc5;
  assign literal_9356[100] = 16'hff97;
  assign literal_9356[101] = 16'hffb5;
  assign literal_9356[102] = 16'hffbf;
  assign literal_9356[103] = 16'hffcc;
  assign literal_9356[104] = 16'hffd9;
  assign literal_9356[105] = 16'hffe7;
  assign literal_9356[106] = 16'hfff5;
  assign literal_9356[107] = 16'h0000;
  assign literal_9356[108] = 16'h0000;
  assign literal_9356[109] = 16'h0000;
  assign literal_9356[110] = 16'h0000;
  assign literal_9356[111] = 16'h0000;
  assign literal_9356[112] = 16'h0000;
  assign literal_9356[113] = 16'h00f9;
  assign literal_9356[114] = 16'h0ff5;
  assign literal_9356[115] = 16'hff8c;
  assign literal_9356[116] = 16'hff98;
  assign literal_9356[117] = 16'hffb6;
  assign literal_9356[118] = 16'hffc0;
  assign literal_9356[119] = 16'hffcd;
  assign literal_9356[120] = 16'hffda;
  assign literal_9356[121] = 16'hffe8;
  assign literal_9356[122] = 16'hfff6;
  assign literal_9356[123] = 16'h0000;
  assign literal_9356[124] = 16'h0000;
  assign literal_9356[125] = 16'h0000;
  assign literal_9356[126] = 16'h0000;
  assign literal_9356[127] = 16'h0000;
  assign literal_9356[128] = 16'h0000;
  assign literal_9356[129] = 16'h01f4;
  assign literal_9356[130] = 16'h1fec;
  assign literal_9356[131] = 16'hff9e;
  assign literal_9356[132] = 16'hffa3;
  assign literal_9356[133] = 16'hffb7;
  assign literal_9356[134] = 16'hffc1;
  assign literal_9356[135] = 16'hffce;
  assign literal_9356[136] = 16'hffdb;
  assign literal_9356[137] = 16'hffe9;
  assign literal_9356[138] = 16'hfff7;
  assign literal_9356[139] = 16'h0000;
  assign literal_9356[140] = 16'h0000;
  assign literal_9356[141] = 16'h0000;
  assign literal_9356[142] = 16'h0000;
  assign literal_9356[143] = 16'h0000;
  assign literal_9356[144] = 16'h0000;
  assign literal_9356[145] = 16'h01f7;
  assign literal_9356[146] = 16'h3fe0;
  assign literal_9356[147] = 16'hff91;
  assign literal_9356[148] = 16'hffa4;
  assign literal_9356[149] = 16'hffb8;
  assign literal_9356[150] = 16'hffc2;
  assign literal_9356[151] = 16'hffcf;
  assign literal_9356[152] = 16'hffdc;
  assign literal_9356[153] = 16'hffea;
  assign literal_9356[154] = 16'hfff8;
  assign literal_9356[155] = 16'h0000;
  assign literal_9356[156] = 16'h0000;
  assign literal_9356[157] = 16'h0000;
  assign literal_9356[158] = 16'h0000;
  assign literal_9356[159] = 16'h0000;
  assign literal_9356[160] = 16'h0000;
  assign literal_9356[161] = 16'h01f8;
  assign literal_9356[162] = 16'h3fe1;
  assign literal_9356[163] = 16'hff92;
  assign literal_9356[164] = 16'hffa7;
  assign literal_9356[165] = 16'hffb9;
  assign literal_9356[166] = 16'hffc3;
  assign literal_9356[167] = 16'hffd0;
  assign literal_9356[168] = 16'hffdd;
  assign literal_9356[169] = 16'hffeb;
  assign literal_9356[170] = 16'hfff9;
  assign literal_9356[171] = 16'h0000;
  assign literal_9356[172] = 16'h0000;
  assign literal_9356[173] = 16'h0000;
  assign literal_9356[174] = 16'h0000;
  assign literal_9356[175] = 16'h0000;
  assign literal_9356[176] = 16'h0000;
  assign literal_9356[177] = 16'h03f5;
  assign literal_9356[178] = 16'h7fc4;
  assign literal_9356[179] = 16'hff93;
  assign literal_9356[180] = 16'hffa8;
  assign literal_9356[181] = 16'hffba;
  assign literal_9356[182] = 16'hffc4;
  assign literal_9356[183] = 16'hffd1;
  assign literal_9356[184] = 16'hffde;
  assign literal_9356[185] = 16'hffec;
  assign literal_9356[186] = 16'hfffa;
  assign literal_9356[187] = 16'h0000;
  assign literal_9356[188] = 16'h0000;
  assign literal_9356[189] = 16'h0000;
  assign literal_9356[190] = 16'h0000;
  assign literal_9356[191] = 16'h0000;
  assign literal_9356[192] = 16'h0000;
  assign literal_9356[193] = 16'h03f8;
  assign literal_9356[194] = 16'hff8d;
  assign literal_9356[195] = 16'hff99;
  assign literal_9356[196] = 16'hffb1;
  assign literal_9356[197] = 16'hffbb;
  assign literal_9356[198] = 16'hffc5;
  assign literal_9356[199] = 16'hffd2;
  assign literal_9356[200] = 16'hffdf;
  assign literal_9356[201] = 16'hffed;
  assign literal_9356[202] = 16'hfffb;
  assign literal_9356[203] = 16'h0000;
  assign literal_9356[204] = 16'h0000;
  assign literal_9356[205] = 16'h0000;
  assign literal_9356[206] = 16'h0000;
  assign literal_9356[207] = 16'h0000;
  assign literal_9356[208] = 16'h0000;
  assign literal_9356[209] = 16'h03fa;
  assign literal_9356[210] = 16'hff9a;
  assign literal_9356[211] = 16'hffaa;
  assign literal_9356[212] = 16'hffb2;
  assign literal_9356[213] = 16'hffbc;
  assign literal_9356[214] = 16'hffc6;
  assign literal_9356[215] = 16'hffd3;
  assign literal_9356[216] = 16'hffe0;
  assign literal_9356[217] = 16'hffee;
  assign literal_9356[218] = 16'hfffc;
  assign literal_9356[219] = 16'h0000;
  assign literal_9356[220] = 16'h0000;
  assign literal_9356[221] = 16'h0000;
  assign literal_9356[222] = 16'h0000;
  assign literal_9356[223] = 16'h0000;
  assign literal_9356[224] = 16'h0000;
  assign literal_9356[225] = 16'h07f6;
  assign literal_9356[226] = 16'hff9b;
  assign literal_9356[227] = 16'hffaf;
  assign literal_9356[228] = 16'hffb3;
  assign literal_9356[229] = 16'hffbd;
  assign literal_9356[230] = 16'hffc7;
  assign literal_9356[231] = 16'hffd4;
  assign literal_9356[232] = 16'hffe1;
  assign literal_9356[233] = 16'hffef;
  assign literal_9356[234] = 16'hfffd;
  assign literal_9356[235] = 16'h0000;
  assign literal_9356[236] = 16'h0000;
  assign literal_9356[237] = 16'h0000;
  assign literal_9356[238] = 16'h0000;
  assign literal_9356[239] = 16'h0000;
  assign literal_9356[240] = 16'h0ff3;
  assign literal_9356[241] = 16'h1fed;
  assign literal_9356[242] = 16'hffae;
  assign literal_9356[243] = 16'hffb0;
  assign literal_9356[244] = 16'hffb4;
  assign literal_9356[245] = 16'hffbe;
  assign literal_9356[246] = 16'hffc8;
  assign literal_9356[247] = 16'hffd5;
  assign literal_9356[248] = 16'hffe2;
  assign literal_9356[249] = 16'hfff0;
  assign literal_9356[250] = 16'hfffe;
  assign literal_9356[251] = 16'h0000;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [2:0] p1_huff_code__1_squeezed_squeezed_comb;
  wire [9:0] p1_row0_comb[0:7];
  wire [9:0] p1_row1_comb[0:7];
  wire [9:0] p1_array_concat_8413_comb[0:15];
  wire [9:0] p1_row2_comb[0:7];
  wire [9:0] p1_array_concat_8416_comb[0:23];
  wire [9:0] p1_row3_comb[0:7];
  wire [2:0] p1_idx_u8__4_squeezed_comb;
  wire [9:0] p1_array_concat_8419_comb[0:31];
  wire [9:0] p1_row4_comb[0:7];
  wire [2:0] p1_idx_u8__5_squeezed_comb;
  wire [9:0] p1_array_concat_8422_comb[0:39];
  wire [9:0] p1_row5_comb[0:7];
  wire [2:0] p1_idx_u8__6_squeezed_comb;
  wire [7:0] p1_idx_u8__1_comb;
  wire [7:0] p1_idx_u8__3_comb;
  wire [7:0] p1_idx_u8__5_comb;
  wire [7:0] p1_idx_u8__7_comb;
  wire [7:0] p1_idx_u8__9_comb;
  wire [7:0] p1_idx_u8__11_comb;
  wire [7:0] p1_idx_u8__13_comb;
  wire [9:0] p1_array_concat_8428_comb[0:47];
  wire [9:0] p1_row6_comb[0:7];
  wire [2:0] p1_idx_u8__7_squeezed_comb;
  wire [6:0] p1_add_8431_comb;
  wire [7:0] p1_actual_index__1_comb;
  wire [6:0] p1_add_8546_comb;
  wire [7:0] p1_actual_index__3_comb;
  wire [5:0] p1_add_8529_comb;
  wire [7:0] p1_actual_index__5_comb;
  wire [6:0] p1_add_8513_comb;
  wire [7:0] p1_actual_index__7_comb;
  wire [7:0] p1_actual_index__9_comb;
  wire [6:0] p1_add_8464_comb;
  wire [7:0] p1_actual_index__11_comb;
  wire [7:0] p1_actual_index__13_comb;
  wire [7:0] p1_idx_u8__15_comb;
  wire [3:0] p1_huff_code__1_squeezed__1_comb;
  wire [7:0] p1_idx_u8__17_comb;
  wire [7:0] p1_idx_u8__19_comb;
  wire [7:0] p1_idx_u8__21_comb;
  wire [7:0] p1_idx_u8__23_comb;
  wire [7:0] p1_idx_u8__25_comb;
  wire [7:0] p1_idx_u8__27_comb;
  wire [7:0] p1_idx_u8__29_comb;
  wire [7:0] p1_idx_u8__31_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__2_comb;
  wire [7:0] p1_idx_u8__33_comb;
  wire [7:0] p1_idx_u8__35_comb;
  wire [7:0] p1_idx_u8__37_comb;
  wire [7:0] p1_idx_u8__39_comb;
  wire [7:0] p1_idx_u8__41_comb;
  wire [7:0] p1_idx_u8__43_comb;
  wire [7:0] p1_idx_u8__45_comb;
  wire [7:0] p1_idx_u8__47_comb;
  wire [7:0] p1_idx_u8__49_comb;
  wire [7:0] p1_idx_u8__51_comb;
  wire [7:0] p1_idx_u8__53_comb;
  wire [7:0] p1_idx_u8__55_comb;
  wire [7:0] p1_idx_u8__57_comb;
  wire [7:0] p1_idx_u8__59_comb;
  wire [7:0] p1_idx_u8__61_comb;
  wire [9:0] p1_array_concat_8435_comb[0:55];
  wire [9:0] p1_row7_comb[0:7];
  wire [5:0] p1_add_8440_comb;
  wire [4:0] p1_add_8483_comb;
  wire [7:0] p1_actual_index__15_comb;
  wire [3:0] p1_add_8649_comb;
  wire [7:0] p1_actual_index__17_comb;
  wire [6:0] p1_add_8651_comb;
  wire [7:0] p1_actual_index__19_comb;
  wire [5:0] p1_add_8653_comb;
  wire [7:0] p1_actual_index__21_comb;
  wire [6:0] p1_add_8655_comb;
  wire [7:0] p1_actual_index__23_comb;
  wire [4:0] p1_add_8657_comb;
  wire [7:0] p1_actual_index__25_comb;
  wire [6:0] p1_add_8659_comb;
  wire [7:0] p1_actual_index__27_comb;
  wire [5:0] p1_add_8661_comb;
  wire [7:0] p1_actual_index__29_comb;
  wire [6:0] p1_add_8663_comb;
  wire [7:0] p1_actual_index__31_comb;
  wire [2:0] p1_add_8665_comb;
  wire [7:0] p1_actual_index__33_comb;
  wire [6:0] p1_add_8667_comb;
  wire [7:0] p1_actual_index__35_comb;
  wire [5:0] p1_add_8669_comb;
  wire [7:0] p1_actual_index__37_comb;
  wire [6:0] p1_add_8671_comb;
  wire [7:0] p1_actual_index__39_comb;
  wire [4:0] p1_add_8673_comb;
  wire [7:0] p1_actual_index__41_comb;
  wire [6:0] p1_add_8675_comb;
  wire [7:0] p1_actual_index__43_comb;
  wire [5:0] p1_add_8677_comb;
  wire [7:0] p1_actual_index__45_comb;
  wire [6:0] p1_add_8679_comb;
  wire [7:0] p1_actual_index__47_comb;
  wire [3:0] p1_add_8681_comb;
  wire [7:0] p1_actual_index__49_comb;
  wire [6:0] p1_add_8683_comb;
  wire [7:0] p1_actual_index__51_comb;
  wire [5:0] p1_add_8685_comb;
  wire [7:0] p1_actual_index__53_comb;
  wire [6:0] p1_add_8687_comb;
  wire [7:0] p1_actual_index__55_comb;
  wire [4:0] p1_add_8689_comb;
  wire [7:0] p1_actual_index__57_comb;
  wire [6:0] p1_add_8691_comb;
  wire [7:0] p1_actual_index__59_comb;
  wire [5:0] p1_add_8693_comb;
  wire [7:0] p1_actual_index__61_comb;
  wire [6:0] p1_add_8695_comb;
  wire [9:0] p1_flat_comb[0:63];
  wire [7:0] p1_actual_index__14_comb;
  wire [7:0] p1_actual_index__2_comb;
  wire [7:0] p1_actual_index__4_comb;
  wire [7:0] p1_actual_index__6_comb;
  wire [7:0] p1_actual_index__10_comb;
  wire [7:0] p1_actual_index__12_comb;
  wire [7:0] p1_actual_index__8_comb;
  wire [7:0] p1_actual_index__16_comb;
  wire [7:0] p1_actual_index__18_comb;
  wire [7:0] p1_actual_index__20_comb;
  wire [7:0] p1_actual_index__22_comb;
  wire [7:0] p1_actual_index__24_comb;
  wire [7:0] p1_actual_index__26_comb;
  wire [7:0] p1_actual_index__28_comb;
  wire [7:0] p1_actual_index__30_comb;
  wire [7:0] p1_actual_index__32_comb;
  wire [7:0] p1_actual_index__34_comb;
  wire [7:0] p1_actual_index__36_comb;
  wire [7:0] p1_actual_index__38_comb;
  wire [7:0] p1_actual_index__40_comb;
  wire [7:0] p1_actual_index__42_comb;
  wire [7:0] p1_actual_index__44_comb;
  wire [7:0] p1_actual_index__46_comb;
  wire [7:0] p1_actual_index__48_comb;
  wire [7:0] p1_actual_index__50_comb;
  wire [7:0] p1_actual_index__52_comb;
  wire [7:0] p1_actual_index__54_comb;
  wire [7:0] p1_actual_index__56_comb;
  wire [7:0] p1_actual_index__58_comb;
  wire [7:0] p1_actual_index__60_comb;
  wire [7:0] p1_actual_index__62_comb;
  wire [9:0] p1_and_8459_comb;
  wire [9:0] p1_and_8590_comb;
  wire [9:0] p1_and_8592_comb;
  wire [9:0] p1_and_8587_comb;
  wire [9:0] p1_and_8580_comb;
  wire [9:0] p1_and_8573_comb;
  wire [9:0] p1_and_8562_comb;
  wire [9:0] p1_and_8553_comb;
  wire [9:0] p1_and_8543_comb;
  wire [9:0] p1_and_8516_comb;
  wire [9:0] p1_and_8507_comb;
  wire [9:0] p1_and_8499_comb;
  wire [9:0] p1_and_8467_comb;
  wire p1_eq_8470_comb;
  wire [9:0] p1_and_8471_comb;
  wire p1_ne_8595_comb;
  wire p1_ne_8596_comb;
  wire p1_ne_8594_comb;
  wire p1_ne_8589_comb;
  wire p1_ne_8582_comb;
  wire p1_ne_8575_comb;
  wire p1_ne_8564_comb;
  wire p1_ne_8555_comb;
  wire [9:0] p1_and_8519_comb;
  wire p1_ne_8526_comb;
  wire p1_ne_8518_comb;
  wire p1_ne_8509_comb;
  wire p1_ne_8479_comb;
  wire [9:0] p1_value_comb;
  wire [1:0] p1_idx_u8__1_squeezed_comb;
  wire p1_eq_8482_comb;
  wire p1_not_8597_comb;
  wire p1_eq_8527_comb;
  wire [7:0] p1_bin_value__1_comb;
  wire [7:0] p1_flipped_comb;
  wire [1:0] p1_sel_8490_comb;
  wire [1:0] p1_sign_ext_8491_comb;
  wire p1_and_9119_comb;
  wire [7:0] p1_code_list_comb;
  assign p1_huff_code__1_squeezed_squeezed_comb = 3'h1;
  assign p1_row0_comb[0] = p0_matrix[3'h0][0];
  assign p1_row0_comb[1] = p0_matrix[3'h0][1];
  assign p1_row0_comb[2] = p0_matrix[3'h0][2];
  assign p1_row0_comb[3] = p0_matrix[3'h0][3];
  assign p1_row0_comb[4] = p0_matrix[3'h0][4];
  assign p1_row0_comb[5] = p0_matrix[3'h0][5];
  assign p1_row0_comb[6] = p0_matrix[3'h0][6];
  assign p1_row0_comb[7] = p0_matrix[3'h0][7];
  assign p1_row1_comb[0] = p0_matrix[p1_huff_code__1_squeezed_squeezed_comb][0];
  assign p1_row1_comb[1] = p0_matrix[p1_huff_code__1_squeezed_squeezed_comb][1];
  assign p1_row1_comb[2] = p0_matrix[p1_huff_code__1_squeezed_squeezed_comb][2];
  assign p1_row1_comb[3] = p0_matrix[p1_huff_code__1_squeezed_squeezed_comb][3];
  assign p1_row1_comb[4] = p0_matrix[p1_huff_code__1_squeezed_squeezed_comb][4];
  assign p1_row1_comb[5] = p0_matrix[p1_huff_code__1_squeezed_squeezed_comb][5];
  assign p1_row1_comb[6] = p0_matrix[p1_huff_code__1_squeezed_squeezed_comb][6];
  assign p1_row1_comb[7] = p0_matrix[p1_huff_code__1_squeezed_squeezed_comb][7];
  assign p1_array_concat_8413_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_8413_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_8413_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_8413_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_8413_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_8413_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_8413_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_8413_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_8413_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_8413_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_8413_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_8413_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_8413_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_8413_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_8413_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_8413_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_8416_comb[0] = p1_array_concat_8413_comb[0];
  assign p1_array_concat_8416_comb[1] = p1_array_concat_8413_comb[1];
  assign p1_array_concat_8416_comb[2] = p1_array_concat_8413_comb[2];
  assign p1_array_concat_8416_comb[3] = p1_array_concat_8413_comb[3];
  assign p1_array_concat_8416_comb[4] = p1_array_concat_8413_comb[4];
  assign p1_array_concat_8416_comb[5] = p1_array_concat_8413_comb[5];
  assign p1_array_concat_8416_comb[6] = p1_array_concat_8413_comb[6];
  assign p1_array_concat_8416_comb[7] = p1_array_concat_8413_comb[7];
  assign p1_array_concat_8416_comb[8] = p1_array_concat_8413_comb[8];
  assign p1_array_concat_8416_comb[9] = p1_array_concat_8413_comb[9];
  assign p1_array_concat_8416_comb[10] = p1_array_concat_8413_comb[10];
  assign p1_array_concat_8416_comb[11] = p1_array_concat_8413_comb[11];
  assign p1_array_concat_8416_comb[12] = p1_array_concat_8413_comb[12];
  assign p1_array_concat_8416_comb[13] = p1_array_concat_8413_comb[13];
  assign p1_array_concat_8416_comb[14] = p1_array_concat_8413_comb[14];
  assign p1_array_concat_8416_comb[15] = p1_array_concat_8413_comb[15];
  assign p1_array_concat_8416_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_8416_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_8416_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_8416_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_8416_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_8416_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_8416_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_8416_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_idx_u8__4_squeezed_comb = 3'h4;
  assign p1_array_concat_8419_comb[0] = p1_array_concat_8416_comb[0];
  assign p1_array_concat_8419_comb[1] = p1_array_concat_8416_comb[1];
  assign p1_array_concat_8419_comb[2] = p1_array_concat_8416_comb[2];
  assign p1_array_concat_8419_comb[3] = p1_array_concat_8416_comb[3];
  assign p1_array_concat_8419_comb[4] = p1_array_concat_8416_comb[4];
  assign p1_array_concat_8419_comb[5] = p1_array_concat_8416_comb[5];
  assign p1_array_concat_8419_comb[6] = p1_array_concat_8416_comb[6];
  assign p1_array_concat_8419_comb[7] = p1_array_concat_8416_comb[7];
  assign p1_array_concat_8419_comb[8] = p1_array_concat_8416_comb[8];
  assign p1_array_concat_8419_comb[9] = p1_array_concat_8416_comb[9];
  assign p1_array_concat_8419_comb[10] = p1_array_concat_8416_comb[10];
  assign p1_array_concat_8419_comb[11] = p1_array_concat_8416_comb[11];
  assign p1_array_concat_8419_comb[12] = p1_array_concat_8416_comb[12];
  assign p1_array_concat_8419_comb[13] = p1_array_concat_8416_comb[13];
  assign p1_array_concat_8419_comb[14] = p1_array_concat_8416_comb[14];
  assign p1_array_concat_8419_comb[15] = p1_array_concat_8416_comb[15];
  assign p1_array_concat_8419_comb[16] = p1_array_concat_8416_comb[16];
  assign p1_array_concat_8419_comb[17] = p1_array_concat_8416_comb[17];
  assign p1_array_concat_8419_comb[18] = p1_array_concat_8416_comb[18];
  assign p1_array_concat_8419_comb[19] = p1_array_concat_8416_comb[19];
  assign p1_array_concat_8419_comb[20] = p1_array_concat_8416_comb[20];
  assign p1_array_concat_8419_comb[21] = p1_array_concat_8416_comb[21];
  assign p1_array_concat_8419_comb[22] = p1_array_concat_8416_comb[22];
  assign p1_array_concat_8419_comb[23] = p1_array_concat_8416_comb[23];
  assign p1_array_concat_8419_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_8419_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_8419_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_8419_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_8419_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_8419_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_8419_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_8419_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[p1_idx_u8__4_squeezed_comb][0];
  assign p1_row4_comb[1] = p0_matrix[p1_idx_u8__4_squeezed_comb][1];
  assign p1_row4_comb[2] = p0_matrix[p1_idx_u8__4_squeezed_comb][2];
  assign p1_row4_comb[3] = p0_matrix[p1_idx_u8__4_squeezed_comb][3];
  assign p1_row4_comb[4] = p0_matrix[p1_idx_u8__4_squeezed_comb][4];
  assign p1_row4_comb[5] = p0_matrix[p1_idx_u8__4_squeezed_comb][5];
  assign p1_row4_comb[6] = p0_matrix[p1_idx_u8__4_squeezed_comb][6];
  assign p1_row4_comb[7] = p0_matrix[p1_idx_u8__4_squeezed_comb][7];
  assign p1_idx_u8__5_squeezed_comb = 3'h5;
  assign p1_array_concat_8422_comb[0] = p1_array_concat_8419_comb[0];
  assign p1_array_concat_8422_comb[1] = p1_array_concat_8419_comb[1];
  assign p1_array_concat_8422_comb[2] = p1_array_concat_8419_comb[2];
  assign p1_array_concat_8422_comb[3] = p1_array_concat_8419_comb[3];
  assign p1_array_concat_8422_comb[4] = p1_array_concat_8419_comb[4];
  assign p1_array_concat_8422_comb[5] = p1_array_concat_8419_comb[5];
  assign p1_array_concat_8422_comb[6] = p1_array_concat_8419_comb[6];
  assign p1_array_concat_8422_comb[7] = p1_array_concat_8419_comb[7];
  assign p1_array_concat_8422_comb[8] = p1_array_concat_8419_comb[8];
  assign p1_array_concat_8422_comb[9] = p1_array_concat_8419_comb[9];
  assign p1_array_concat_8422_comb[10] = p1_array_concat_8419_comb[10];
  assign p1_array_concat_8422_comb[11] = p1_array_concat_8419_comb[11];
  assign p1_array_concat_8422_comb[12] = p1_array_concat_8419_comb[12];
  assign p1_array_concat_8422_comb[13] = p1_array_concat_8419_comb[13];
  assign p1_array_concat_8422_comb[14] = p1_array_concat_8419_comb[14];
  assign p1_array_concat_8422_comb[15] = p1_array_concat_8419_comb[15];
  assign p1_array_concat_8422_comb[16] = p1_array_concat_8419_comb[16];
  assign p1_array_concat_8422_comb[17] = p1_array_concat_8419_comb[17];
  assign p1_array_concat_8422_comb[18] = p1_array_concat_8419_comb[18];
  assign p1_array_concat_8422_comb[19] = p1_array_concat_8419_comb[19];
  assign p1_array_concat_8422_comb[20] = p1_array_concat_8419_comb[20];
  assign p1_array_concat_8422_comb[21] = p1_array_concat_8419_comb[21];
  assign p1_array_concat_8422_comb[22] = p1_array_concat_8419_comb[22];
  assign p1_array_concat_8422_comb[23] = p1_array_concat_8419_comb[23];
  assign p1_array_concat_8422_comb[24] = p1_array_concat_8419_comb[24];
  assign p1_array_concat_8422_comb[25] = p1_array_concat_8419_comb[25];
  assign p1_array_concat_8422_comb[26] = p1_array_concat_8419_comb[26];
  assign p1_array_concat_8422_comb[27] = p1_array_concat_8419_comb[27];
  assign p1_array_concat_8422_comb[28] = p1_array_concat_8419_comb[28];
  assign p1_array_concat_8422_comb[29] = p1_array_concat_8419_comb[29];
  assign p1_array_concat_8422_comb[30] = p1_array_concat_8419_comb[30];
  assign p1_array_concat_8422_comb[31] = p1_array_concat_8419_comb[31];
  assign p1_array_concat_8422_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_8422_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_8422_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_8422_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_8422_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_8422_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_8422_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_8422_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[p1_idx_u8__5_squeezed_comb][0];
  assign p1_row5_comb[1] = p0_matrix[p1_idx_u8__5_squeezed_comb][1];
  assign p1_row5_comb[2] = p0_matrix[p1_idx_u8__5_squeezed_comb][2];
  assign p1_row5_comb[3] = p0_matrix[p1_idx_u8__5_squeezed_comb][3];
  assign p1_row5_comb[4] = p0_matrix[p1_idx_u8__5_squeezed_comb][4];
  assign p1_row5_comb[5] = p0_matrix[p1_idx_u8__5_squeezed_comb][5];
  assign p1_row5_comb[6] = p0_matrix[p1_idx_u8__5_squeezed_comb][6];
  assign p1_row5_comb[7] = p0_matrix[p1_idx_u8__5_squeezed_comb][7];
  assign p1_idx_u8__6_squeezed_comb = 3'h6;
  assign p1_idx_u8__1_comb = 8'h01;
  assign p1_idx_u8__3_comb = 8'h03;
  assign p1_idx_u8__5_comb = 8'h05;
  assign p1_idx_u8__7_comb = 8'h07;
  assign p1_idx_u8__9_comb = 8'h09;
  assign p1_idx_u8__11_comb = 8'h0b;
  assign p1_idx_u8__13_comb = 8'h0d;
  assign p1_array_concat_8428_comb[0] = p1_array_concat_8422_comb[0];
  assign p1_array_concat_8428_comb[1] = p1_array_concat_8422_comb[1];
  assign p1_array_concat_8428_comb[2] = p1_array_concat_8422_comb[2];
  assign p1_array_concat_8428_comb[3] = p1_array_concat_8422_comb[3];
  assign p1_array_concat_8428_comb[4] = p1_array_concat_8422_comb[4];
  assign p1_array_concat_8428_comb[5] = p1_array_concat_8422_comb[5];
  assign p1_array_concat_8428_comb[6] = p1_array_concat_8422_comb[6];
  assign p1_array_concat_8428_comb[7] = p1_array_concat_8422_comb[7];
  assign p1_array_concat_8428_comb[8] = p1_array_concat_8422_comb[8];
  assign p1_array_concat_8428_comb[9] = p1_array_concat_8422_comb[9];
  assign p1_array_concat_8428_comb[10] = p1_array_concat_8422_comb[10];
  assign p1_array_concat_8428_comb[11] = p1_array_concat_8422_comb[11];
  assign p1_array_concat_8428_comb[12] = p1_array_concat_8422_comb[12];
  assign p1_array_concat_8428_comb[13] = p1_array_concat_8422_comb[13];
  assign p1_array_concat_8428_comb[14] = p1_array_concat_8422_comb[14];
  assign p1_array_concat_8428_comb[15] = p1_array_concat_8422_comb[15];
  assign p1_array_concat_8428_comb[16] = p1_array_concat_8422_comb[16];
  assign p1_array_concat_8428_comb[17] = p1_array_concat_8422_comb[17];
  assign p1_array_concat_8428_comb[18] = p1_array_concat_8422_comb[18];
  assign p1_array_concat_8428_comb[19] = p1_array_concat_8422_comb[19];
  assign p1_array_concat_8428_comb[20] = p1_array_concat_8422_comb[20];
  assign p1_array_concat_8428_comb[21] = p1_array_concat_8422_comb[21];
  assign p1_array_concat_8428_comb[22] = p1_array_concat_8422_comb[22];
  assign p1_array_concat_8428_comb[23] = p1_array_concat_8422_comb[23];
  assign p1_array_concat_8428_comb[24] = p1_array_concat_8422_comb[24];
  assign p1_array_concat_8428_comb[25] = p1_array_concat_8422_comb[25];
  assign p1_array_concat_8428_comb[26] = p1_array_concat_8422_comb[26];
  assign p1_array_concat_8428_comb[27] = p1_array_concat_8422_comb[27];
  assign p1_array_concat_8428_comb[28] = p1_array_concat_8422_comb[28];
  assign p1_array_concat_8428_comb[29] = p1_array_concat_8422_comb[29];
  assign p1_array_concat_8428_comb[30] = p1_array_concat_8422_comb[30];
  assign p1_array_concat_8428_comb[31] = p1_array_concat_8422_comb[31];
  assign p1_array_concat_8428_comb[32] = p1_array_concat_8422_comb[32];
  assign p1_array_concat_8428_comb[33] = p1_array_concat_8422_comb[33];
  assign p1_array_concat_8428_comb[34] = p1_array_concat_8422_comb[34];
  assign p1_array_concat_8428_comb[35] = p1_array_concat_8422_comb[35];
  assign p1_array_concat_8428_comb[36] = p1_array_concat_8422_comb[36];
  assign p1_array_concat_8428_comb[37] = p1_array_concat_8422_comb[37];
  assign p1_array_concat_8428_comb[38] = p1_array_concat_8422_comb[38];
  assign p1_array_concat_8428_comb[39] = p1_array_concat_8422_comb[39];
  assign p1_array_concat_8428_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_8428_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_8428_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_8428_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_8428_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_8428_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_8428_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_8428_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[p1_idx_u8__6_squeezed_comb][0];
  assign p1_row6_comb[1] = p0_matrix[p1_idx_u8__6_squeezed_comb][1];
  assign p1_row6_comb[2] = p0_matrix[p1_idx_u8__6_squeezed_comb][2];
  assign p1_row6_comb[3] = p0_matrix[p1_idx_u8__6_squeezed_comb][3];
  assign p1_row6_comb[4] = p0_matrix[p1_idx_u8__6_squeezed_comb][4];
  assign p1_row6_comb[5] = p0_matrix[p1_idx_u8__6_squeezed_comb][5];
  assign p1_row6_comb[6] = p0_matrix[p1_idx_u8__6_squeezed_comb][6];
  assign p1_row6_comb[7] = p0_matrix[p1_idx_u8__6_squeezed_comb][7];
  assign p1_idx_u8__7_squeezed_comb = 3'h7;
  assign p1_add_8431_comb = p0_start_pix[7:1] + 7'h07;
  assign p1_actual_index__1_comb = p0_start_pix + p1_idx_u8__1_comb;
  assign p1_add_8546_comb = p0_start_pix[7:1] + 7'h01;
  assign p1_actual_index__3_comb = p0_start_pix + p1_idx_u8__3_comb;
  assign p1_add_8529_comb = p0_start_pix[7:2] + 6'h01;
  assign p1_actual_index__5_comb = p0_start_pix + p1_idx_u8__5_comb;
  assign p1_add_8513_comb = p0_start_pix[7:1] + 7'h03;
  assign p1_actual_index__7_comb = p0_start_pix + p1_idx_u8__7_comb;
  assign p1_actual_index__9_comb = p0_start_pix + p1_idx_u8__9_comb;
  assign p1_add_8464_comb = p0_start_pix[7:1] + 7'h05;
  assign p1_actual_index__11_comb = p0_start_pix + p1_idx_u8__11_comb;
  assign p1_actual_index__13_comb = p0_start_pix + p1_idx_u8__13_comb;
  assign p1_idx_u8__15_comb = 8'h0f;
  assign p1_huff_code__1_squeezed__1_comb = 4'h1;
  assign p1_idx_u8__17_comb = 8'h11;
  assign p1_idx_u8__19_comb = 8'h13;
  assign p1_idx_u8__21_comb = 8'h15;
  assign p1_idx_u8__23_comb = 8'h17;
  assign p1_idx_u8__25_comb = 8'h19;
  assign p1_idx_u8__27_comb = 8'h1b;
  assign p1_idx_u8__29_comb = 8'h1d;
  assign p1_idx_u8__31_comb = 8'h1f;
  assign p1_huff_code__1_squeezed_squeezed__2_comb = 3'h1;
  assign p1_idx_u8__33_comb = 8'h21;
  assign p1_idx_u8__35_comb = 8'h23;
  assign p1_idx_u8__37_comb = 8'h25;
  assign p1_idx_u8__39_comb = 8'h27;
  assign p1_idx_u8__41_comb = 8'h29;
  assign p1_idx_u8__43_comb = 8'h2b;
  assign p1_idx_u8__45_comb = 8'h2d;
  assign p1_idx_u8__47_comb = 8'h2f;
  assign p1_idx_u8__49_comb = 8'h31;
  assign p1_idx_u8__51_comb = 8'h33;
  assign p1_idx_u8__53_comb = 8'h35;
  assign p1_idx_u8__55_comb = 8'h37;
  assign p1_idx_u8__57_comb = 8'h39;
  assign p1_idx_u8__59_comb = 8'h3b;
  assign p1_idx_u8__61_comb = 8'h3d;
  assign p1_array_concat_8435_comb[0] = p1_array_concat_8428_comb[0];
  assign p1_array_concat_8435_comb[1] = p1_array_concat_8428_comb[1];
  assign p1_array_concat_8435_comb[2] = p1_array_concat_8428_comb[2];
  assign p1_array_concat_8435_comb[3] = p1_array_concat_8428_comb[3];
  assign p1_array_concat_8435_comb[4] = p1_array_concat_8428_comb[4];
  assign p1_array_concat_8435_comb[5] = p1_array_concat_8428_comb[5];
  assign p1_array_concat_8435_comb[6] = p1_array_concat_8428_comb[6];
  assign p1_array_concat_8435_comb[7] = p1_array_concat_8428_comb[7];
  assign p1_array_concat_8435_comb[8] = p1_array_concat_8428_comb[8];
  assign p1_array_concat_8435_comb[9] = p1_array_concat_8428_comb[9];
  assign p1_array_concat_8435_comb[10] = p1_array_concat_8428_comb[10];
  assign p1_array_concat_8435_comb[11] = p1_array_concat_8428_comb[11];
  assign p1_array_concat_8435_comb[12] = p1_array_concat_8428_comb[12];
  assign p1_array_concat_8435_comb[13] = p1_array_concat_8428_comb[13];
  assign p1_array_concat_8435_comb[14] = p1_array_concat_8428_comb[14];
  assign p1_array_concat_8435_comb[15] = p1_array_concat_8428_comb[15];
  assign p1_array_concat_8435_comb[16] = p1_array_concat_8428_comb[16];
  assign p1_array_concat_8435_comb[17] = p1_array_concat_8428_comb[17];
  assign p1_array_concat_8435_comb[18] = p1_array_concat_8428_comb[18];
  assign p1_array_concat_8435_comb[19] = p1_array_concat_8428_comb[19];
  assign p1_array_concat_8435_comb[20] = p1_array_concat_8428_comb[20];
  assign p1_array_concat_8435_comb[21] = p1_array_concat_8428_comb[21];
  assign p1_array_concat_8435_comb[22] = p1_array_concat_8428_comb[22];
  assign p1_array_concat_8435_comb[23] = p1_array_concat_8428_comb[23];
  assign p1_array_concat_8435_comb[24] = p1_array_concat_8428_comb[24];
  assign p1_array_concat_8435_comb[25] = p1_array_concat_8428_comb[25];
  assign p1_array_concat_8435_comb[26] = p1_array_concat_8428_comb[26];
  assign p1_array_concat_8435_comb[27] = p1_array_concat_8428_comb[27];
  assign p1_array_concat_8435_comb[28] = p1_array_concat_8428_comb[28];
  assign p1_array_concat_8435_comb[29] = p1_array_concat_8428_comb[29];
  assign p1_array_concat_8435_comb[30] = p1_array_concat_8428_comb[30];
  assign p1_array_concat_8435_comb[31] = p1_array_concat_8428_comb[31];
  assign p1_array_concat_8435_comb[32] = p1_array_concat_8428_comb[32];
  assign p1_array_concat_8435_comb[33] = p1_array_concat_8428_comb[33];
  assign p1_array_concat_8435_comb[34] = p1_array_concat_8428_comb[34];
  assign p1_array_concat_8435_comb[35] = p1_array_concat_8428_comb[35];
  assign p1_array_concat_8435_comb[36] = p1_array_concat_8428_comb[36];
  assign p1_array_concat_8435_comb[37] = p1_array_concat_8428_comb[37];
  assign p1_array_concat_8435_comb[38] = p1_array_concat_8428_comb[38];
  assign p1_array_concat_8435_comb[39] = p1_array_concat_8428_comb[39];
  assign p1_array_concat_8435_comb[40] = p1_array_concat_8428_comb[40];
  assign p1_array_concat_8435_comb[41] = p1_array_concat_8428_comb[41];
  assign p1_array_concat_8435_comb[42] = p1_array_concat_8428_comb[42];
  assign p1_array_concat_8435_comb[43] = p1_array_concat_8428_comb[43];
  assign p1_array_concat_8435_comb[44] = p1_array_concat_8428_comb[44];
  assign p1_array_concat_8435_comb[45] = p1_array_concat_8428_comb[45];
  assign p1_array_concat_8435_comb[46] = p1_array_concat_8428_comb[46];
  assign p1_array_concat_8435_comb[47] = p1_array_concat_8428_comb[47];
  assign p1_array_concat_8435_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_8435_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_8435_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_8435_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_8435_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_8435_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_8435_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_8435_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[p1_idx_u8__7_squeezed_comb][0];
  assign p1_row7_comb[1] = p0_matrix[p1_idx_u8__7_squeezed_comb][1];
  assign p1_row7_comb[2] = p0_matrix[p1_idx_u8__7_squeezed_comb][2];
  assign p1_row7_comb[3] = p0_matrix[p1_idx_u8__7_squeezed_comb][3];
  assign p1_row7_comb[4] = p0_matrix[p1_idx_u8__7_squeezed_comb][4];
  assign p1_row7_comb[5] = p0_matrix[p1_idx_u8__7_squeezed_comb][5];
  assign p1_row7_comb[6] = p0_matrix[p1_idx_u8__7_squeezed_comb][6];
  assign p1_row7_comb[7] = p0_matrix[p1_idx_u8__7_squeezed_comb][7];
  assign p1_add_8440_comb = p0_start_pix[7:2] + 6'h03;
  assign p1_add_8483_comb = p0_start_pix[7:3] + 5'h01;
  assign p1_actual_index__15_comb = p0_start_pix + p1_idx_u8__15_comb;
  assign p1_add_8649_comb = p0_start_pix[7:4] + p1_huff_code__1_squeezed__1_comb;
  assign p1_actual_index__17_comb = p0_start_pix + p1_idx_u8__17_comb;
  assign p1_add_8651_comb = p0_start_pix[7:1] + 7'h09;
  assign p1_actual_index__19_comb = p0_start_pix + p1_idx_u8__19_comb;
  assign p1_add_8653_comb = p0_start_pix[7:2] + 6'h05;
  assign p1_actual_index__21_comb = p0_start_pix + p1_idx_u8__21_comb;
  assign p1_add_8655_comb = p0_start_pix[7:1] + 7'h0b;
  assign p1_actual_index__23_comb = p0_start_pix + p1_idx_u8__23_comb;
  assign p1_add_8657_comb = p0_start_pix[7:3] + 5'h03;
  assign p1_actual_index__25_comb = p0_start_pix + p1_idx_u8__25_comb;
  assign p1_add_8659_comb = p0_start_pix[7:1] + 7'h0d;
  assign p1_actual_index__27_comb = p0_start_pix + p1_idx_u8__27_comb;
  assign p1_add_8661_comb = p0_start_pix[7:2] + 6'h07;
  assign p1_actual_index__29_comb = p0_start_pix + p1_idx_u8__29_comb;
  assign p1_add_8663_comb = p0_start_pix[7:1] + 7'h0f;
  assign p1_actual_index__31_comb = p0_start_pix + p1_idx_u8__31_comb;
  assign p1_add_8665_comb = p0_start_pix[7:5] + p1_huff_code__1_squeezed_squeezed__2_comb;
  assign p1_actual_index__33_comb = p0_start_pix + p1_idx_u8__33_comb;
  assign p1_add_8667_comb = p0_start_pix[7:1] + 7'h11;
  assign p1_actual_index__35_comb = p0_start_pix + p1_idx_u8__35_comb;
  assign p1_add_8669_comb = p0_start_pix[7:2] + 6'h09;
  assign p1_actual_index__37_comb = p0_start_pix + p1_idx_u8__37_comb;
  assign p1_add_8671_comb = p0_start_pix[7:1] + 7'h13;
  assign p1_actual_index__39_comb = p0_start_pix + p1_idx_u8__39_comb;
  assign p1_add_8673_comb = p0_start_pix[7:3] + 5'h05;
  assign p1_actual_index__41_comb = p0_start_pix + p1_idx_u8__41_comb;
  assign p1_add_8675_comb = p0_start_pix[7:1] + 7'h15;
  assign p1_actual_index__43_comb = p0_start_pix + p1_idx_u8__43_comb;
  assign p1_add_8677_comb = p0_start_pix[7:2] + 6'h0b;
  assign p1_actual_index__45_comb = p0_start_pix + p1_idx_u8__45_comb;
  assign p1_add_8679_comb = p0_start_pix[7:1] + 7'h17;
  assign p1_actual_index__47_comb = p0_start_pix + p1_idx_u8__47_comb;
  assign p1_add_8681_comb = p0_start_pix[7:4] + 4'h3;
  assign p1_actual_index__49_comb = p0_start_pix + p1_idx_u8__49_comb;
  assign p1_add_8683_comb = p0_start_pix[7:1] + 7'h19;
  assign p1_actual_index__51_comb = p0_start_pix + p1_idx_u8__51_comb;
  assign p1_add_8685_comb = p0_start_pix[7:2] + 6'h0d;
  assign p1_actual_index__53_comb = p0_start_pix + p1_idx_u8__53_comb;
  assign p1_add_8687_comb = p0_start_pix[7:1] + 7'h1b;
  assign p1_actual_index__55_comb = p0_start_pix + p1_idx_u8__55_comb;
  assign p1_add_8689_comb = p0_start_pix[7:3] + 5'h07;
  assign p1_actual_index__57_comb = p0_start_pix + p1_idx_u8__57_comb;
  assign p1_add_8691_comb = p0_start_pix[7:1] + 7'h1d;
  assign p1_actual_index__59_comb = p0_start_pix + p1_idx_u8__59_comb;
  assign p1_add_8693_comb = p0_start_pix[7:2] + 6'h0f;
  assign p1_actual_index__61_comb = p0_start_pix + p1_idx_u8__61_comb;
  assign p1_add_8695_comb = p0_start_pix[7:1] + 7'h1f;
  assign p1_flat_comb[0] = p1_array_concat_8435_comb[0];
  assign p1_flat_comb[1] = p1_array_concat_8435_comb[1];
  assign p1_flat_comb[2] = p1_array_concat_8435_comb[2];
  assign p1_flat_comb[3] = p1_array_concat_8435_comb[3];
  assign p1_flat_comb[4] = p1_array_concat_8435_comb[4];
  assign p1_flat_comb[5] = p1_array_concat_8435_comb[5];
  assign p1_flat_comb[6] = p1_array_concat_8435_comb[6];
  assign p1_flat_comb[7] = p1_array_concat_8435_comb[7];
  assign p1_flat_comb[8] = p1_array_concat_8435_comb[8];
  assign p1_flat_comb[9] = p1_array_concat_8435_comb[9];
  assign p1_flat_comb[10] = p1_array_concat_8435_comb[10];
  assign p1_flat_comb[11] = p1_array_concat_8435_comb[11];
  assign p1_flat_comb[12] = p1_array_concat_8435_comb[12];
  assign p1_flat_comb[13] = p1_array_concat_8435_comb[13];
  assign p1_flat_comb[14] = p1_array_concat_8435_comb[14];
  assign p1_flat_comb[15] = p1_array_concat_8435_comb[15];
  assign p1_flat_comb[16] = p1_array_concat_8435_comb[16];
  assign p1_flat_comb[17] = p1_array_concat_8435_comb[17];
  assign p1_flat_comb[18] = p1_array_concat_8435_comb[18];
  assign p1_flat_comb[19] = p1_array_concat_8435_comb[19];
  assign p1_flat_comb[20] = p1_array_concat_8435_comb[20];
  assign p1_flat_comb[21] = p1_array_concat_8435_comb[21];
  assign p1_flat_comb[22] = p1_array_concat_8435_comb[22];
  assign p1_flat_comb[23] = p1_array_concat_8435_comb[23];
  assign p1_flat_comb[24] = p1_array_concat_8435_comb[24];
  assign p1_flat_comb[25] = p1_array_concat_8435_comb[25];
  assign p1_flat_comb[26] = p1_array_concat_8435_comb[26];
  assign p1_flat_comb[27] = p1_array_concat_8435_comb[27];
  assign p1_flat_comb[28] = p1_array_concat_8435_comb[28];
  assign p1_flat_comb[29] = p1_array_concat_8435_comb[29];
  assign p1_flat_comb[30] = p1_array_concat_8435_comb[30];
  assign p1_flat_comb[31] = p1_array_concat_8435_comb[31];
  assign p1_flat_comb[32] = p1_array_concat_8435_comb[32];
  assign p1_flat_comb[33] = p1_array_concat_8435_comb[33];
  assign p1_flat_comb[34] = p1_array_concat_8435_comb[34];
  assign p1_flat_comb[35] = p1_array_concat_8435_comb[35];
  assign p1_flat_comb[36] = p1_array_concat_8435_comb[36];
  assign p1_flat_comb[37] = p1_array_concat_8435_comb[37];
  assign p1_flat_comb[38] = p1_array_concat_8435_comb[38];
  assign p1_flat_comb[39] = p1_array_concat_8435_comb[39];
  assign p1_flat_comb[40] = p1_array_concat_8435_comb[40];
  assign p1_flat_comb[41] = p1_array_concat_8435_comb[41];
  assign p1_flat_comb[42] = p1_array_concat_8435_comb[42];
  assign p1_flat_comb[43] = p1_array_concat_8435_comb[43];
  assign p1_flat_comb[44] = p1_array_concat_8435_comb[44];
  assign p1_flat_comb[45] = p1_array_concat_8435_comb[45];
  assign p1_flat_comb[46] = p1_array_concat_8435_comb[46];
  assign p1_flat_comb[47] = p1_array_concat_8435_comb[47];
  assign p1_flat_comb[48] = p1_array_concat_8435_comb[48];
  assign p1_flat_comb[49] = p1_array_concat_8435_comb[49];
  assign p1_flat_comb[50] = p1_array_concat_8435_comb[50];
  assign p1_flat_comb[51] = p1_array_concat_8435_comb[51];
  assign p1_flat_comb[52] = p1_array_concat_8435_comb[52];
  assign p1_flat_comb[53] = p1_array_concat_8435_comb[53];
  assign p1_flat_comb[54] = p1_array_concat_8435_comb[54];
  assign p1_flat_comb[55] = p1_array_concat_8435_comb[55];
  assign p1_flat_comb[56] = p1_row7_comb[0];
  assign p1_flat_comb[57] = p1_row7_comb[1];
  assign p1_flat_comb[58] = p1_row7_comb[2];
  assign p1_flat_comb[59] = p1_row7_comb[3];
  assign p1_flat_comb[60] = p1_row7_comb[4];
  assign p1_flat_comb[61] = p1_row7_comb[5];
  assign p1_flat_comb[62] = p1_row7_comb[6];
  assign p1_flat_comb[63] = p1_row7_comb[7];
  assign p1_actual_index__14_comb = {p1_add_8431_comb, p0_start_pix[0]};
  assign p1_actual_index__2_comb = {p1_add_8546_comb, p0_start_pix[0]};
  assign p1_actual_index__4_comb = {p1_add_8529_comb, p0_start_pix[1:0]};
  assign p1_actual_index__6_comb = {p1_add_8513_comb, p0_start_pix[0]};
  assign p1_actual_index__10_comb = {p1_add_8464_comb, p0_start_pix[0]};
  assign p1_actual_index__12_comb = {p1_add_8440_comb, p0_start_pix[1:0]};
  assign p1_actual_index__8_comb = {p1_add_8483_comb, p0_start_pix[2:0]};
  assign p1_actual_index__16_comb = {p1_add_8649_comb, p0_start_pix[3:0]};
  assign p1_actual_index__18_comb = {p1_add_8651_comb, p0_start_pix[0]};
  assign p1_actual_index__20_comb = {p1_add_8653_comb, p0_start_pix[1:0]};
  assign p1_actual_index__22_comb = {p1_add_8655_comb, p0_start_pix[0]};
  assign p1_actual_index__24_comb = {p1_add_8657_comb, p0_start_pix[2:0]};
  assign p1_actual_index__26_comb = {p1_add_8659_comb, p0_start_pix[0]};
  assign p1_actual_index__28_comb = {p1_add_8661_comb, p0_start_pix[1:0]};
  assign p1_actual_index__30_comb = {p1_add_8663_comb, p0_start_pix[0]};
  assign p1_actual_index__32_comb = {p1_add_8665_comb, p0_start_pix[4:0]};
  assign p1_actual_index__34_comb = {p1_add_8667_comb, p0_start_pix[0]};
  assign p1_actual_index__36_comb = {p1_add_8669_comb, p0_start_pix[1:0]};
  assign p1_actual_index__38_comb = {p1_add_8671_comb, p0_start_pix[0]};
  assign p1_actual_index__40_comb = {p1_add_8673_comb, p0_start_pix[2:0]};
  assign p1_actual_index__42_comb = {p1_add_8675_comb, p0_start_pix[0]};
  assign p1_actual_index__44_comb = {p1_add_8677_comb, p0_start_pix[1:0]};
  assign p1_actual_index__46_comb = {p1_add_8679_comb, p0_start_pix[0]};
  assign p1_actual_index__48_comb = {p1_add_8681_comb, p0_start_pix[3:0]};
  assign p1_actual_index__50_comb = {p1_add_8683_comb, p0_start_pix[0]};
  assign p1_actual_index__52_comb = {p1_add_8685_comb, p0_start_pix[1:0]};
  assign p1_actual_index__54_comb = {p1_add_8687_comb, p0_start_pix[0]};
  assign p1_actual_index__56_comb = {p1_add_8689_comb, p0_start_pix[2:0]};
  assign p1_actual_index__58_comb = {p1_add_8691_comb, p0_start_pix[0]};
  assign p1_actual_index__60_comb = {p1_add_8693_comb, p0_start_pix[1:0]};
  assign p1_actual_index__62_comb = {p1_add_8695_comb, p0_start_pix[0]};
  assign p1_and_8459_comb = p1_flat_comb[p1_actual_index__14_comb > 8'h3f ? 6'h3f : p1_actual_index__14_comb[5:0]] & {10{~(p1_add_8431_comb[5] | p1_add_8431_comb[6])}};
  assign p1_and_8590_comb = p1_flat_comb[p0_start_pix > 8'h3f ? 6'h3f : p0_start_pix[5:0]] & {10{~(p0_start_pix[6] | p0_start_pix[7])}};
  assign p1_and_8592_comb = p1_flat_comb[p1_actual_index__1_comb > 8'h3f ? 6'h3f : p1_actual_index__1_comb[5:0]] & {10{~(p1_actual_index__1_comb[6] | p1_actual_index__1_comb[7])}};
  assign p1_and_8587_comb = p1_flat_comb[p1_actual_index__2_comb > 8'h3f ? 6'h3f : p1_actual_index__2_comb[5:0]] & {10{~(p1_add_8546_comb[5] | p1_add_8546_comb[6])}};
  assign p1_and_8580_comb = p1_flat_comb[p1_actual_index__3_comb > 8'h3f ? 6'h3f : p1_actual_index__3_comb[5:0]] & {10{~(p1_actual_index__3_comb[6] | p1_actual_index__3_comb[7])}};
  assign p1_and_8573_comb = p1_flat_comb[p1_actual_index__4_comb > 8'h3f ? 6'h3f : p1_actual_index__4_comb[5:0]] & {10{~(p1_add_8529_comb[4] | p1_add_8529_comb[5])}};
  assign p1_and_8562_comb = p1_flat_comb[p1_actual_index__5_comb > 8'h3f ? 6'h3f : p1_actual_index__5_comb[5:0]] & {10{~(p1_actual_index__5_comb[6] | p1_actual_index__5_comb[7])}};
  assign p1_and_8553_comb = p1_flat_comb[p1_actual_index__6_comb > 8'h3f ? 6'h3f : p1_actual_index__6_comb[5:0]] & {10{~(p1_add_8513_comb[5] | p1_add_8513_comb[6])}};
  assign p1_and_8543_comb = p1_flat_comb[p1_actual_index__7_comb > 8'h3f ? 6'h3f : p1_actual_index__7_comb[5:0]] & {10{~(p1_actual_index__7_comb[6] | p1_actual_index__7_comb[7])}};
  assign p1_and_8516_comb = p1_flat_comb[p1_actual_index__9_comb > 8'h3f ? 6'h3f : p1_actual_index__9_comb[5:0]] & {10{~(p1_actual_index__9_comb[6] | p1_actual_index__9_comb[7])}};
  assign p1_and_8507_comb = p1_flat_comb[p1_actual_index__10_comb > 8'h3f ? 6'h3f : p1_actual_index__10_comb[5:0]] & {10{~(p1_add_8464_comb[5] | p1_add_8464_comb[6])}};
  assign p1_and_8499_comb = p1_flat_comb[p1_actual_index__11_comb > 8'h3f ? 6'h3f : p1_actual_index__11_comb[5:0]] & {10{~(p1_actual_index__11_comb[6] | p1_actual_index__11_comb[7])}};
  assign p1_and_8467_comb = p1_flat_comb[p1_actual_index__13_comb > 8'h3f ? 6'h3f : p1_actual_index__13_comb[5:0]] & {10{~(p1_actual_index__13_comb[6] | p1_actual_index__13_comb[7])}};
  assign p1_eq_8470_comb = p1_and_8459_comb == 10'h000;
  assign p1_and_8471_comb = p1_flat_comb[p1_actual_index__12_comb > 8'h3f ? 6'h3f : p1_actual_index__12_comb[5:0]] & {10{~(p1_add_8440_comb[4] | p1_add_8440_comb[5])}};
  assign p1_ne_8595_comb = p1_and_8590_comb != 10'h000;
  assign p1_ne_8596_comb = p1_and_8592_comb != 10'h000;
  assign p1_ne_8594_comb = p1_and_8587_comb != 10'h000;
  assign p1_ne_8589_comb = p1_and_8580_comb != 10'h000;
  assign p1_ne_8582_comb = p1_and_8573_comb != 10'h000;
  assign p1_ne_8575_comb = p1_and_8562_comb != 10'h000;
  assign p1_ne_8564_comb = p1_and_8553_comb != 10'h000;
  assign p1_ne_8555_comb = p1_and_8543_comb != 10'h000;
  assign p1_and_8519_comb = p1_flat_comb[p1_actual_index__8_comb > 8'h3f ? 6'h3f : p1_actual_index__8_comb[5:0]] & {10{~(p1_add_8483_comb[3] | p1_add_8483_comb[4])}};
  assign p1_ne_8526_comb = p1_and_8516_comb != 10'h000;
  assign p1_ne_8518_comb = p1_and_8507_comb != 10'h000;
  assign p1_ne_8509_comb = p1_and_8499_comb != 10'h000;
  assign p1_ne_8479_comb = p1_and_8467_comb != 10'h000;
  assign p1_value_comb = p0_matrix[3'h0][3'h0];
  assign p1_idx_u8__1_squeezed_comb = 2'h1;
  assign p1_eq_8482_comb = p1_and_8471_comb == 10'h000;
  assign p1_not_8597_comb = ~p1_ne_8595_comb;
  assign p1_eq_8527_comb = p1_and_8519_comb == 10'h000;
  assign p1_bin_value__1_comb = p1_value_comb[7:0];
  assign p1_flipped_comb = 8'hff;
  assign p1_sel_8490_comb = p1_ne_8479_comb ? p1_idx_u8__1_squeezed_comb : {1'h1, p1_eq_8470_comb};
  assign p1_sign_ext_8491_comb = {2{p1_eq_8482_comb}};
  assign p1_and_9119_comb = p1_not_8597_comb & ~p1_ne_8596_comb & ~p1_ne_8594_comb & ~p1_ne_8589_comb & ~p1_ne_8582_comb & ~p1_ne_8575_comb & ~p1_ne_8564_comb & ~p1_ne_8555_comb & p1_eq_8527_comb & ~p1_ne_8526_comb & ~p1_ne_8518_comb & ~p1_ne_8509_comb & p1_eq_8482_comb & ~p1_ne_8479_comb & p1_eq_8470_comb & (p1_flat_comb[p1_actual_index__15_comb > 8'h3f ? 6'h3f : p1_actual_index__15_comb[5:0]] & {10{~(p1_actual_index__15_comb[6] | p1_actual_index__15_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__16_comb > 8'h3f ? 6'h3f : p1_actual_index__16_comb[5:0]] & {10{~(p1_add_8649_comb[2] | p1_add_8649_comb[3])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__17_comb > 8'h3f ? 6'h3f : p1_actual_index__17_comb[5:0]] & {10{~(p1_actual_index__17_comb[6] | p1_actual_index__17_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__18_comb > 8'h3f ? 6'h3f : p1_actual_index__18_comb[5:0]] & {10{~(p1_add_8651_comb[5] | p1_add_8651_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__19_comb > 8'h3f ? 6'h3f : p1_actual_index__19_comb[5:0]] & {10{~(p1_actual_index__19_comb[6] | p1_actual_index__19_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__20_comb > 8'h3f ? 6'h3f : p1_actual_index__20_comb[5:0]] & {10{~(p1_add_8653_comb[4] | p1_add_8653_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__21_comb > 8'h3f ? 6'h3f : p1_actual_index__21_comb[5:0]] & {10{~(p1_actual_index__21_comb[6] | p1_actual_index__21_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__22_comb > 8'h3f ? 6'h3f : p1_actual_index__22_comb[5:0]] & {10{~(p1_add_8655_comb[5] | p1_add_8655_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__23_comb > 8'h3f ? 6'h3f : p1_actual_index__23_comb[5:0]] & {10{~(p1_actual_index__23_comb[6] | p1_actual_index__23_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__24_comb > 8'h3f ? 6'h3f : p1_actual_index__24_comb[5:0]] & {10{~(p1_add_8657_comb[3] | p1_add_8657_comb[4])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__25_comb > 8'h3f ? 6'h3f : p1_actual_index__25_comb[5:0]] & {10{~(p1_actual_index__25_comb[6] | p1_actual_index__25_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__26_comb > 8'h3f ? 6'h3f : p1_actual_index__26_comb[5:0]] & {10{~(p1_add_8659_comb[5] | p1_add_8659_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__27_comb > 8'h3f ? 6'h3f : p1_actual_index__27_comb[5:0]] & {10{~(p1_actual_index__27_comb[6] | p1_actual_index__27_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__28_comb > 8'h3f ? 6'h3f : p1_actual_index__28_comb[5:0]] & {10{~(p1_add_8661_comb[4] | p1_add_8661_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__29_comb > 8'h3f ? 6'h3f : p1_actual_index__29_comb[5:0]] & {10{~(p1_actual_index__29_comb[6] | p1_actual_index__29_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__30_comb > 8'h3f ? 6'h3f : p1_actual_index__30_comb[5:0]] & {10{~(p1_add_8663_comb[5] | p1_add_8663_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__31_comb > 8'h3f ? 6'h3f : p1_actual_index__31_comb[5:0]] & {10{~(p1_actual_index__31_comb[6] | p1_actual_index__31_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__32_comb > 8'h3f ? 6'h3f : p1_actual_index__32_comb[5:0]] & {10{~(p1_add_8665_comb[1] | p1_add_8665_comb[2])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__33_comb > 8'h3f ? 6'h3f : p1_actual_index__33_comb[5:0]] & {10{~(p1_actual_index__33_comb[6] | p1_actual_index__33_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__34_comb > 8'h3f ? 6'h3f : p1_actual_index__34_comb[5:0]] & {10{~(p1_add_8667_comb[5] | p1_add_8667_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__35_comb > 8'h3f ? 6'h3f : p1_actual_index__35_comb[5:0]] & {10{~(p1_actual_index__35_comb[6] | p1_actual_index__35_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__36_comb > 8'h3f ? 6'h3f : p1_actual_index__36_comb[5:0]] & {10{~(p1_add_8669_comb[4] | p1_add_8669_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__37_comb > 8'h3f ? 6'h3f : p1_actual_index__37_comb[5:0]] & {10{~(p1_actual_index__37_comb[6] | p1_actual_index__37_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__38_comb > 8'h3f ? 6'h3f : p1_actual_index__38_comb[5:0]] & {10{~(p1_add_8671_comb[5] | p1_add_8671_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__39_comb > 8'h3f ? 6'h3f : p1_actual_index__39_comb[5:0]] & {10{~(p1_actual_index__39_comb[6] | p1_actual_index__39_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__40_comb > 8'h3f ? 6'h3f : p1_actual_index__40_comb[5:0]] & {10{~(p1_add_8673_comb[3] | p1_add_8673_comb[4])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__41_comb > 8'h3f ? 6'h3f : p1_actual_index__41_comb[5:0]] & {10{~(p1_actual_index__41_comb[6] | p1_actual_index__41_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__42_comb > 8'h3f ? 6'h3f : p1_actual_index__42_comb[5:0]] & {10{~(p1_add_8675_comb[5] | p1_add_8675_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__43_comb > 8'h3f ? 6'h3f : p1_actual_index__43_comb[5:0]] & {10{~(p1_actual_index__43_comb[6] | p1_actual_index__43_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__44_comb > 8'h3f ? 6'h3f : p1_actual_index__44_comb[5:0]] & {10{~(p1_add_8677_comb[4] | p1_add_8677_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__45_comb > 8'h3f ? 6'h3f : p1_actual_index__45_comb[5:0]] & {10{~(p1_actual_index__45_comb[6] | p1_actual_index__45_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__46_comb > 8'h3f ? 6'h3f : p1_actual_index__46_comb[5:0]] & {10{~(p1_add_8679_comb[5] | p1_add_8679_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__47_comb > 8'h3f ? 6'h3f : p1_actual_index__47_comb[5:0]] & {10{~(p1_actual_index__47_comb[6] | p1_actual_index__47_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__48_comb > 8'h3f ? 6'h3f : p1_actual_index__48_comb[5:0]] & {10{~(p1_add_8681_comb[2] | p1_add_8681_comb[3])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__49_comb > 8'h3f ? 6'h3f : p1_actual_index__49_comb[5:0]] & {10{~(p1_actual_index__49_comb[6] | p1_actual_index__49_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__50_comb > 8'h3f ? 6'h3f : p1_actual_index__50_comb[5:0]] & {10{~(p1_add_8683_comb[5] | p1_add_8683_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__51_comb > 8'h3f ? 6'h3f : p1_actual_index__51_comb[5:0]] & {10{~(p1_actual_index__51_comb[6] | p1_actual_index__51_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__52_comb > 8'h3f ? 6'h3f : p1_actual_index__52_comb[5:0]] & {10{~(p1_add_8685_comb[4] | p1_add_8685_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__53_comb > 8'h3f ? 6'h3f : p1_actual_index__53_comb[5:0]] & {10{~(p1_actual_index__53_comb[6] | p1_actual_index__53_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__54_comb > 8'h3f ? 6'h3f : p1_actual_index__54_comb[5:0]] & {10{~(p1_add_8687_comb[5] | p1_add_8687_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__55_comb > 8'h3f ? 6'h3f : p1_actual_index__55_comb[5:0]] & {10{~(p1_actual_index__55_comb[6] | p1_actual_index__55_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__56_comb > 8'h3f ? 6'h3f : p1_actual_index__56_comb[5:0]] & {10{~(p1_add_8689_comb[3] | p1_add_8689_comb[4])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__57_comb > 8'h3f ? 6'h3f : p1_actual_index__57_comb[5:0]] & {10{~(p1_actual_index__57_comb[6] | p1_actual_index__57_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__58_comb > 8'h3f ? 6'h3f : p1_actual_index__58_comb[5:0]] & {10{~(p1_add_8691_comb[5] | p1_add_8691_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__59_comb > 8'h3f ? 6'h3f : p1_actual_index__59_comb[5:0]] & {10{~(p1_actual_index__59_comb[6] | p1_actual_index__59_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__60_comb > 8'h3f ? 6'h3f : p1_actual_index__60_comb[5:0]] & {10{~(p1_add_8693_comb[4] | p1_add_8693_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__61_comb > 8'h3f ? 6'h3f : p1_actual_index__61_comb[5:0]] & {10{~(p1_actual_index__61_comb[6] | p1_actual_index__61_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__62_comb > 8'h3f ? 6'h3f : p1_actual_index__62_comb[5:0]] & {10{~(p1_add_8695_comb[5] | p1_add_8695_comb[6])}}) == 10'h000;
  assign p1_code_list_comb = p1_value_comb == 10'h000 ? p1_flipped_comb : p1_bin_value__1_comb;

  // Registers for pipe stage 1:
  reg p1_is_luminance;
  reg [9:0] p1_and_8459;
  reg [9:0] p1_and_8467;
  reg [9:0] p1_and_8471;
  reg [1:0] p1_sel_8490;
  reg [1:0] p1_sign_ext_8491;
  reg [9:0] p1_and_8499;
  reg [9:0] p1_and_8507;
  reg p1_ne_8509;
  reg [9:0] p1_and_8516;
  reg p1_ne_8518;
  reg [9:0] p1_and_8519;
  reg p1_ne_8526;
  reg p1_eq_8527;
  reg [9:0] p1_and_8543;
  reg [9:0] p1_and_8553;
  reg p1_ne_8555;
  reg [9:0] p1_and_8562;
  reg p1_ne_8564;
  reg [9:0] p1_and_8573;
  reg p1_ne_8575;
  reg [9:0] p1_and_8580;
  reg p1_ne_8582;
  reg [9:0] p1_and_8587;
  reg p1_ne_8589;
  reg [9:0] p1_and_8590;
  reg [9:0] p1_and_8592;
  reg p1_ne_8594;
  reg p1_ne_8595;
  reg p1_ne_8596;
  reg p1_not_8597;
  reg p1_and_9119;
  reg [7:0] p1_code_list;
  always @ (posedge clk) begin
    p1_is_luminance <= p0_is_luminance;
    p1_and_8459 <= p1_and_8459_comb;
    p1_and_8467 <= p1_and_8467_comb;
    p1_and_8471 <= p1_and_8471_comb;
    p1_sel_8490 <= p1_sel_8490_comb;
    p1_sign_ext_8491 <= p1_sign_ext_8491_comb;
    p1_and_8499 <= p1_and_8499_comb;
    p1_and_8507 <= p1_and_8507_comb;
    p1_ne_8509 <= p1_ne_8509_comb;
    p1_and_8516 <= p1_and_8516_comb;
    p1_ne_8518 <= p1_ne_8518_comb;
    p1_and_8519 <= p1_and_8519_comb;
    p1_ne_8526 <= p1_ne_8526_comb;
    p1_eq_8527 <= p1_eq_8527_comb;
    p1_and_8543 <= p1_and_8543_comb;
    p1_and_8553 <= p1_and_8553_comb;
    p1_ne_8555 <= p1_ne_8555_comb;
    p1_and_8562 <= p1_and_8562_comb;
    p1_ne_8564 <= p1_ne_8564_comb;
    p1_and_8573 <= p1_and_8573_comb;
    p1_ne_8575 <= p1_ne_8575_comb;
    p1_and_8580 <= p1_and_8580_comb;
    p1_ne_8582 <= p1_ne_8582_comb;
    p1_and_8587 <= p1_and_8587_comb;
    p1_ne_8589 <= p1_ne_8589_comb;
    p1_and_8590 <= p1_and_8590_comb;
    p1_and_8592 <= p1_and_8592_comb;
    p1_ne_8594 <= p1_ne_8594_comb;
    p1_ne_8595 <= p1_ne_8595_comb;
    p1_ne_8596 <= p1_ne_8596_comb;
    p1_not_8597 <= p1_not_8597_comb;
    p1_and_9119 <= p1_and_9119_comb;
    p1_code_list <= p1_code_list_comb;
  end

  // ===== Pipe stage 2:
  wire [2:0] p2_huff_code__1_squeezed_squeezed__1_comb;
  wire [2:0] p2_and_9203_comb;
  wire [3:0] p2_idx_u8__4_squeezed__2_comb;
  wire [3:0] p2_sel_9212_comb;
  wire [3:0] p2_sel_9216_comb;
  assign p2_huff_code__1_squeezed_squeezed__1_comb = 3'h1;
  assign p2_and_9203_comb = (p1_ne_8526 ? p2_huff_code__1_squeezed_squeezed__1_comb : (p1_ne_8518 ? 3'h2 : (p1_ne_8509 ? 3'h3 : {1'h1, p1_sel_8490 & p1_sign_ext_8491}))) & {3{p1_eq_8527}};
  assign p2_idx_u8__4_squeezed__2_comb = 4'h4;
  assign p2_sel_9212_comb = p1_ne_8582 ? p2_idx_u8__4_squeezed__2_comb : (p1_ne_8575 ? 4'h5 : (p1_ne_8564 ? 4'h6 : (p1_ne_8555 ? 4'h7 : {1'h1, p2_and_9203_comb})));
  assign p2_sel_9216_comb = p1_ne_8594 ? 4'h2 : (p1_ne_8589 ? 4'h3 : p2_sel_9212_comb);

  // Registers for pipe stage 2:
  reg p2_is_luminance;
  reg [9:0] p2_and_8459;
  reg [9:0] p2_and_8467;
  reg [9:0] p2_and_8471;
  reg [9:0] p2_and_8499;
  reg [9:0] p2_and_8507;
  reg [9:0] p2_and_8516;
  reg [9:0] p2_and_8519;
  reg [9:0] p2_and_8543;
  reg [9:0] p2_and_8553;
  reg [9:0] p2_and_8562;
  reg [9:0] p2_and_8573;
  reg [9:0] p2_and_8580;
  reg [9:0] p2_and_8587;
  reg [9:0] p2_and_8590;
  reg [9:0] p2_and_8592;
  reg p2_ne_8595;
  reg p2_ne_8596;
  reg [3:0] p2_sel_9216;
  reg p2_not_8597;
  reg p2_and_9119;
  reg [7:0] p2_code_list;
  always @ (posedge clk) begin
    p2_is_luminance <= p1_is_luminance;
    p2_and_8459 <= p1_and_8459;
    p2_and_8467 <= p1_and_8467;
    p2_and_8471 <= p1_and_8471;
    p2_and_8499 <= p1_and_8499;
    p2_and_8507 <= p1_and_8507;
    p2_and_8516 <= p1_and_8516;
    p2_and_8519 <= p1_and_8519;
    p2_and_8543 <= p1_and_8543;
    p2_and_8553 <= p1_and_8553;
    p2_and_8562 <= p1_and_8562;
    p2_and_8573 <= p1_and_8573;
    p2_and_8580 <= p1_and_8580;
    p2_and_8587 <= p1_and_8587;
    p2_and_8590 <= p1_and_8590;
    p2_and_8592 <= p1_and_8592;
    p2_ne_8595 <= p1_ne_8595;
    p2_ne_8596 <= p1_ne_8596;
    p2_sel_9216 <= p2_sel_9216_comb;
    p2_not_8597 <= p1_not_8597;
    p2_and_9119 <= p1_and_9119;
    p2_code_list <= p1_code_list;
  end

  // ===== Pipe stage 3:
  wire [3:0] p3_huff_code__1_squeezed_comb;
  wire [3:0] p3_sel_9262_comb;
  wire [3:0] p3_run_comb;
  wire [9:0] p3_value__1_comb;
  wire [7:0] p3_bin_value__2_comb;
  wire [7:0] p3_bin_value__3_comb;
  wire [7:0] p3_value_abs_comb;
  wire [1:0] p3_idx_u8__1_squeezed__1_comb;
  wire [1:0] p3_idx_u8__2_squeezed_comb;
  wire [1:0] p3_idx_u8__3_squeezed_comb;
  wire p3_eq_9299_comb;
  wire [7:0] p3_flipped__1_comb;
  wire [2:0] p3_idx_u8__4_squeezed__1_comb;
  wire [7:0] p3_Code_list_comb;
  wire [2:0] p3_sel_9288_comb;
  wire [2:0] p3_idx_u8__5_squeezed__1_comb;
  wire p3_or_reduce_9291_comb;
  wire [2:0] p3_sel_9292_comb;
  wire p3_or_reduce_9293_comb;
  wire p3_bit_slice_9294_comb;
  wire p3_ne_9296_comb;
  wire [7:0] p3_sel_9310_comb;
  wire [3:0] p3_sel_9311_comb;
  assign p3_huff_code__1_squeezed_comb = 4'h1;
  assign p3_sel_9262_comb = p2_ne_8596 ? p3_huff_code__1_squeezed_comb : p2_sel_9216;
  assign p3_run_comb = p3_sel_9262_comb & {4{p2_not_8597}};
  assign p3_value__1_comb = p3_run_comb == 4'h0 ? p2_and_8590 : (p3_run_comb == 4'h1 ? p2_and_8592 : (p3_run_comb == 4'h2 ? p2_and_8587 : (p3_run_comb == 4'h3 ? p2_and_8580 : (p3_run_comb == 4'h4 ? p2_and_8573 : (p3_run_comb == 4'h5 ? p2_and_8562 : (p3_run_comb == 4'h6 ? p2_and_8553 : (p3_run_comb == 4'h7 ? p2_and_8543 : (p3_run_comb == 4'h8 ? p2_and_8519 : (p3_run_comb == 4'h9 ? p2_and_8516 : (p3_run_comb == 4'ha ? p2_and_8507 : (p3_run_comb == 4'hb ? p2_and_8499 : (p3_run_comb == 4'hc ? p2_and_8471 : (p3_run_comb == 4'hd ? p2_and_8467 : (p3_run_comb == 4'he ? p2_and_8459 : 10'h000))))))))))))));
  assign p3_bin_value__2_comb = p3_value__1_comb[7:0];
  assign p3_bin_value__3_comb = -p3_bin_value__2_comb;
  assign p3_value_abs_comb = p3_value__1_comb[9] ? p3_bin_value__3_comb : p3_bin_value__2_comb;
  assign p3_idx_u8__1_squeezed__1_comb = 2'h1;
  assign p3_idx_u8__2_squeezed_comb = 2'h2;
  assign p3_idx_u8__3_squeezed_comb = 2'h3;
  assign p3_eq_9299_comb = p3_run_comb == 4'hf;
  assign p3_flipped__1_comb = ~p3_bin_value__3_comb;
  assign p3_idx_u8__4_squeezed__1_comb = 3'h4;
  assign p3_Code_list_comb = $signed(p3_value__1_comb) <= $signed(10'h000) ? p3_flipped__1_comb : p3_bin_value__2_comb;
  assign p3_sel_9288_comb = |p3_value_abs_comb[7:3] ? p3_idx_u8__4_squeezed__1_comb : {1'h0, |p3_value_abs_comb[7:2] ? p3_idx_u8__3_squeezed_comb : (|p3_value_abs_comb[7:1] ? p3_idx_u8__2_squeezed_comb : p3_idx_u8__1_squeezed__1_comb)};
  assign p3_idx_u8__5_squeezed__1_comb = 3'h5;
  assign p3_or_reduce_9291_comb = |p3_value_abs_comb[7:5];
  assign p3_sel_9292_comb = |p3_value_abs_comb[7:4] ? p3_idx_u8__5_squeezed__1_comb : p3_sel_9288_comb;
  assign p3_or_reduce_9293_comb = |p3_value_abs_comb[7:6];
  assign p3_bit_slice_9294_comb = p3_value_abs_comb[7];
  assign p3_ne_9296_comb = p3_value_abs_comb != 8'h00;
  assign p3_sel_9310_comb = p2_and_9119 ? p2_code_list : p3_Code_list_comb & {8{~p3_eq_9299_comb}};
  assign p3_sel_9311_comb = p2_and_9119 ? 4'hf : p3_sel_9262_comb & {4{~(p3_eq_9299_comb | p2_ne_8595)}};

  // Registers for pipe stage 3:
  reg p3_is_luminance;
  reg [3:0] p3_run;
  reg p3_or_reduce_9291;
  reg [2:0] p3_sel_9292;
  reg p3_or_reduce_9293;
  reg p3_bit_slice_9294;
  reg p3_ne_9296;
  reg p3_eq_9299;
  reg p3_and_9119;
  reg [7:0] p3_sel_9310;
  reg [3:0] p3_sel_9311;
  always @ (posedge clk) begin
    p3_is_luminance <= p2_is_luminance;
    p3_run <= p3_run_comb;
    p3_or_reduce_9291 <= p3_or_reduce_9291_comb;
    p3_sel_9292 <= p3_sel_9292_comb;
    p3_or_reduce_9293 <= p3_or_reduce_9293_comb;
    p3_bit_slice_9294 <= p3_bit_slice_9294_comb;
    p3_ne_9296 <= p3_ne_9296_comb;
    p3_eq_9299 <= p3_eq_9299_comb;
    p3_and_9119 <= p2_and_9119;
    p3_sel_9310 <= p3_sel_9310_comb;
    p3_sel_9311 <= p3_sel_9311_comb;
  end

  // ===== Pipe stage 4:
  wire [2:0] p4_idx_u8__6_squeezed__1_comb;
  wire [2:0] p4_idx_u8__7_squeezed__1_comb;
  wire [3:0] p4_idx_u8__8_squeezed_comb;
  wire [7:0] p4_Code_size_comb;
  wire [2:0] p4_huff_code__1_squeezed_squeezed__3_comb;
  wire [2:0] p4_idx_u8__4_squeezed__3_comb;
  wire [7:0] p4_run_size_str_u8_comb;
  wire [1:0] p4_idx_u8__1_squeezed__2_comb;
  wire [1:0] p4_idx_u8__2_squeezed__1_comb;
  wire [2:0] p4_sel_9357_comb;
  wire [3:0] p4_Code_size_squeezed_comb;
  wire [3:0] p4_idx_u8__4_squeezed__4_comb;
  wire p4_or_9369_comb;
  wire [4:0] p4_Huffman_length_squeezed_comb;
  wire [15:0] p4_Huffman_code_full_comb;
  wire [43:0] p4_tuple_9384_comb;
  assign p4_idx_u8__6_squeezed__1_comb = 3'h6;
  assign p4_idx_u8__7_squeezed__1_comb = 3'h7;
  assign p4_idx_u8__8_squeezed_comb = 4'h8;
  assign p4_Code_size_comb = {4'h0, p3_bit_slice_9294 ? p4_idx_u8__8_squeezed_comb : {1'h0, p3_or_reduce_9293 ? p4_idx_u8__7_squeezed__1_comb : (p3_or_reduce_9291 ? p4_idx_u8__6_squeezed__1_comb : p3_sel_9292)}} & {8{p3_ne_9296}};
  assign p4_huff_code__1_squeezed_squeezed__3_comb = 3'h1;
  assign p4_idx_u8__4_squeezed__3_comb = 3'h4;
  assign p4_run_size_str_u8_comb = {p3_run, 4'h0} | p4_Code_size_comb;
  assign p4_idx_u8__1_squeezed__2_comb = 2'h1;
  assign p4_idx_u8__2_squeezed__1_comb = 2'h2;
  assign p4_sel_9357_comb = p3_is_luminance ? p4_idx_u8__4_squeezed__3_comb : p4_huff_code__1_squeezed_squeezed__3_comb;
  assign p4_Code_size_squeezed_comb = p4_Code_size_comb[3:0];
  assign p4_idx_u8__4_squeezed__4_comb = 4'h4;
  assign p4_or_9369_comb = p3_and_9119 | p3_eq_9299;
  assign p4_Huffman_length_squeezed_comb = p3_is_luminance ? literal_9352[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_9350[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_Huffman_code_full_comb = p3_is_luminance ? literal_9356[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_9355[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_tuple_9384_comb = {p4_or_9369_comb ? {12'h000, {{1{p4_sel_9357_comb[2]}}, p4_sel_9357_comb}} : p4_Huffman_code_full_comb, {3'h0, p4_or_9369_comb ? {2'h0, p3_is_luminance ? p4_idx_u8__2_squeezed__1_comb : p4_idx_u8__1_squeezed__2_comb, 1'h0} : p4_Huffman_length_squeezed_comb}, p3_sel_9310, {4'h0, p3_eq_9299 ? p4_idx_u8__4_squeezed__4_comb : p4_Code_size_squeezed_comb} & {8{~p3_and_9119}}, p3_sel_9311};

  // Registers for pipe stage 4:
  reg [43:0] p4_tuple_9384;
  always @ (posedge clk) begin
    p4_tuple_9384 <= p4_tuple_9384_comb;
  end
  assign out = p4_tuple_9384;
endmodule
