module dct_1d_u8(
  input wire clk,
  input wire [63:0] x,
  output wire [63:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [15:0] smul16b_8b_x_9b (input reg [7:0] lhs, input reg [8:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [15:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul16b_8b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_8b (input reg [7:0] lhs, input reg [7:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_6b (input reg [7:0] lhs, input reg [5:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [23:0] umul24b_24b_x_7b (input reg [23:0] lhs, input reg [6:0] rhs);
    begin
      umul24b_24b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [7:0] x_unflattened[0:7];
  assign x_unflattened[0] = x[7:0];
  assign x_unflattened[1] = x[15:8];
  assign x_unflattened[2] = x[23:16];
  assign x_unflattened[3] = x[31:24];
  assign x_unflattened[4] = x[39:32];
  assign x_unflattened[5] = x[47:40];
  assign x_unflattened[6] = x[55:48];
  assign x_unflattened[7] = x[63:56];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_x[0:7];
  always @ (posedge clk) begin
    p0_x[0] <= x_unflattened[0];
    p0_x[1] <= x_unflattened[1];
    p0_x[2] <= x_unflattened[2];
    p0_x[3] <= x_unflattened[3];
    p0_x[4] <= x_unflattened[4];
    p0_x[5] <= x_unflattened[5];
    p0_x[6] <= x_unflattened[6];
    p0_x[7] <= x_unflattened[7];
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_array_index_5918_comb;
  wire [7:0] p1_array_index_5919_comb;
  wire [7:0] p1_array_index_5920_comb;
  wire [7:0] p1_array_index_5921_comb;
  wire [7:0] p1_array_index_5922_comb;
  wire [7:0] p1_array_index_5923_comb;
  wire [7:0] p1_array_index_5924_comb;
  wire [7:0] p1_array_index_5925_comb;
  wire [7:0] p1_concat_5950_comb;
  wire [7:0] p1_concat_5952_comb;
  wire [7:0] p1_concat_5954_comb;
  wire [7:0] p1_concat_5956_comb;
  wire [7:0] p1_concat_5959_comb;
  wire [7:0] p1_concat_5961_comb;
  wire [7:0] p1_concat_5965_comb;
  wire [7:0] p1_concat_5967_comb;
  wire [15:0] p1_smul_3303_NarrowedMult__comb;
  wire [15:0] p1_smul_3302_NarrowedMult__comb;
  wire [15:0] p1_smul_3297_NarrowedMult__comb;
  wire [15:0] p1_smul_3296_NarrowedMult__comb;
  wire [15:0] p1_smul_3287_NarrowedMult__comb;
  wire [15:0] p1_smul_3285_NarrowedMult__comb;
  wire [15:0] p1_smul_3282_NarrowedMult__comb;
  wire [15:0] p1_smul_3280_NarrowedMult__comb;
  wire [15:0] p1_smul_3270_NarrowedMult__comb;
  wire [15:0] p1_smul_3268_NarrowedMult__comb;
  wire [15:0] p1_smul_3267_NarrowedMult__comb;
  wire [15:0] p1_smul_3265_NarrowedMult__comb;
  wire [15:0] p1_smul_3253_NarrowedMult__comb;
  wire [15:0] p1_smul_3252_NarrowedMult__comb;
  wire [15:0] p1_smul_3251_NarrowedMult__comb;
  wire [15:0] p1_smul_3250_NarrowedMult__comb;
  wire [14:0] p1_smul_3301_NarrowedMult__comb;
  wire [13:0] p1_smul_3317_NarrowedMult__comb;
  wire [13:0] p1_smul_3319_NarrowedMult__comb;
  wire [14:0] p1_smul_3298_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6018_comb;
  wire [13:0] p1_smul_3378_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6020_comb;
  wire [14:0] p1_smul_3284_NarrowedMult__comb;
  wire [14:0] p1_smul_3283_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6023_comb;
  wire [13:0] p1_smul_3398_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6025_comb;
  wire [14:0] p1_smul_3271_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6035_comb;
  wire [13:0] p1_smul_3445_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6037_comb;
  wire [14:0] p1_bit_slice_6038_comb;
  wire [13:0] p1_smul_3455_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6040_comb;
  wire [14:0] p1_smul_3264_NarrowedMult__comb;
  wire [13:0] p1_smul_3506_NarrowedMult__comb;
  wire [14:0] p1_smul_3254_NarrowedMult__comb;
  wire [14:0] p1_smul_3249_NarrowedMult__comb;
  wire [13:0] p1_smul_3534_NarrowedMult__comb;
  wire [16:0] p1_add_6054_comb;
  wire [16:0] p1_add_6059_comb;
  wire [14:0] p1_smul_3294_NarrowedMult__comb;
  wire [14:0] p1_smul_3293_NarrowedMult__comb;
  wire [14:0] p1_smul_3290_NarrowedMult__comb;
  wire [14:0] p1_smul_3289_NarrowedMult__comb;
  wire [15:0] p1_smul_3279_NarrowedMult__comb;
  wire [15:0] p1_smul_3278_NarrowedMult__comb;
  wire [15:0] p1_smul_3277_NarrowedMult__comb;
  wire [15:0] p1_smul_3276_NarrowedMult__comb;
  wire [15:0] p1_smul_3275_NarrowedMult__comb;
  wire [15:0] p1_smul_3274_NarrowedMult__comb;
  wire [15:0] p1_smul_3273_NarrowedMult__comb;
  wire [15:0] p1_smul_3272_NarrowedMult__comb;
  wire [14:0] p1_smul_3263_NarrowedMult__comb;
  wire [14:0] p1_smul_3261_NarrowedMult__comb;
  wire [14:0] p1_smul_3258_NarrowedMult__comb;
  wire [14:0] p1_smul_3256_NarrowedMult__comb;
  wire [16:0] p1_add_6102_comb;
  wire [16:0] p1_add_6103_comb;
  wire [15:0] p1_bit_slice_6106_comb;
  wire [15:0] p1_add_6107_comb;
  wire [15:0] p1_add_6108_comb;
  wire [15:0] p1_bit_slice_6109_comb;
  wire [13:0] p1_smul_3295_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6111_comb;
  wire [13:0] p1_bit_slice_6112_comb;
  wire [13:0] p1_smul_3292_NarrowedMult__comb;
  wire [13:0] p1_smul_3291_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6115_comb;
  wire [13:0] p1_bit_slice_6116_comb;
  wire [13:0] p1_smul_3288_NarrowedMult__comb;
  wire [15:0] p1_add_6118_comb;
  wire [15:0] p1_add_6120_comb;
  wire [15:0] p1_add_6122_comb;
  wire [15:0] p1_add_6124_comb;
  wire [15:0] p1_add_6134_comb;
  wire [15:0] p1_add_6136_comb;
  wire [15:0] p1_add_6138_comb;
  wire [15:0] p1_add_6140_comb;
  wire [13:0] p1_bit_slice_6142_comb;
  wire [13:0] p1_smul_3262_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6144_comb;
  wire [13:0] p1_smul_3260_NarrowedMult__comb;
  wire [13:0] p1_smul_3259_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6147_comb;
  wire [13:0] p1_smul_3257_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6149_comb;
  wire [15:0] p1_add_6150_comb;
  wire [15:0] p1_bit_slice_6151_comb;
  wire [15:0] p1_bit_slice_6152_comb;
  wire [15:0] p1_add_6153_comb;
  wire [16:0] p1_concat_6174_comb;
  wire [16:0] p1_concat_6175_comb;
  wire [16:0] p1_concat_6176_comb;
  wire [16:0] p1_concat_6177_comb;
  wire [16:0] p1_add_6178_comb;
  wire [16:0] p1_add_6179_comb;
  wire [16:0] p1_add_6180_comb;
  wire [16:0] p1_add_6181_comb;
  wire [16:0] p1_concat_6182_comb;
  wire [16:0] p1_concat_6183_comb;
  wire [16:0] p1_concat_6184_comb;
  wire [16:0] p1_concat_6185_comb;
  wire [8:0] p1_add_6198_comb;
  wire [8:0] p1_add_6199_comb;
  wire [8:0] p1_add_6200_comb;
  wire [8:0] p1_add_6201_comb;
  wire [23:0] p1_add_6202_comb;
  wire [23:0] p1_add_6204_comb;
  wire [14:0] p1_add_6206_comb;
  wire [14:0] p1_add_6208_comb;
  wire [14:0] p1_add_6210_comb;
  wire [14:0] p1_add_6212_comb;
  wire [24:0] p1_sum__101_comb;
  wire [24:0] p1_sum__102_comb;
  wire [24:0] p1_sum__103_comb;
  wire [24:0] p1_sum__104_comb;
  wire [24:0] p1_sum__97_comb;
  wire [24:0] p1_sum__98_comb;
  wire [24:0] p1_sum__99_comb;
  wire [24:0] p1_sum__100_comb;
  wire [24:0] p1_sum__93_comb;
  wire [24:0] p1_sum__94_comb;
  wire [24:0] p1_sum__95_comb;
  wire [24:0] p1_sum__96_comb;
  wire [14:0] p1_add_6226_comb;
  wire [14:0] p1_add_6228_comb;
  wire [14:0] p1_add_6230_comb;
  wire [14:0] p1_add_6232_comb;
  wire [23:0] p1_add_6234_comb;
  wire [23:0] p1_add_6236_comb;
  wire [24:0] p1_sum__83_comb;
  wire [24:0] p1_sum__84_comb;
  wire [15:0] p1_concat_6244_comb;
  wire [15:0] p1_concat_6245_comb;
  wire [15:0] p1_concat_6246_comb;
  wire [15:0] p1_concat_6247_comb;
  wire [24:0] p1_sum__79_comb;
  wire [24:0] p1_sum__80_comb;
  wire [24:0] p1_sum__77_comb;
  wire [24:0] p1_sum__78_comb;
  wire [24:0] p1_sum__75_comb;
  wire [24:0] p1_sum__76_comb;
  wire [15:0] p1_concat_6254_comb;
  wire [15:0] p1_concat_6255_comb;
  wire [15:0] p1_concat_6256_comb;
  wire [15:0] p1_concat_6257_comb;
  wire [24:0] p1_sum__71_comb;
  wire [24:0] p1_sum__72_comb;
  wire [23:0] p1_add_6260_comb;
  wire [23:0] p1_add_6261_comb;
  wire [24:0] p1_sum__70_comb;
  wire [24:0] p1_sum__68_comb;
  wire [24:0] p1_sum__67_comb;
  wire [24:0] p1_sum__66_comb;
  wire [24:0] p1_sum__64_comb;
  wire [23:0] p1_add_6280_comb;
  wire [24:0] p1_add_6282_comb;
  wire [23:0] p1_add_6283_comb;
  wire [23:0] p1_add_6284_comb;
  wire [24:0] p1_add_6285_comb;
  wire [24:0] p1_add_6286_comb;
  wire [24:0] p1_add_6287_comb;
  wire [23:0] p1_add_6288_comb;
  wire [23:0] p1_add_6289_comb;
  wire [24:0] p1_add_6290_comb;
  wire [23:0] p1_umul_2792_NarrowedMult__comb;
  wire [23:0] p1_add_6295_comb;
  wire [23:0] p1_add_6303_comb;
  wire [8:0] p1_clipped__16_comb;
  wire [8:0] p1_clipped__17_comb;
  wire [8:0] p1_clipped__18_comb;
  wire [8:0] p1_clipped__19_comb;
  wire [8:0] p1_clipped__20_comb;
  wire [8:0] p1_clipped__21_comb;
  wire [8:0] p1_clipped__22_comb;
  wire [8:0] p1_clipped__23_comb;
  wire [9:0] p1_add_6387_comb;
  wire [9:0] p1_add_6388_comb;
  wire [9:0] p1_add_6389_comb;
  wire [9:0] p1_add_6390_comb;
  wire [9:0] p1_add_6391_comb;
  wire [9:0] p1_add_6392_comb;
  wire [9:0] p1_add_6393_comb;
  wire [9:0] p1_add_6394_comb;
  wire [1:0] p1_bit_slice_6395_comb;
  wire [1:0] p1_bit_slice_6396_comb;
  wire [1:0] p1_bit_slice_6397_comb;
  wire [1:0] p1_bit_slice_6398_comb;
  wire [1:0] p1_bit_slice_6399_comb;
  wire [1:0] p1_bit_slice_6400_comb;
  wire [1:0] p1_bit_slice_6401_comb;
  wire [1:0] p1_bit_slice_6402_comb;
  wire [2:0] p1_add_6419_comb;
  wire [2:0] p1_add_6420_comb;
  wire [2:0] p1_add_6421_comb;
  wire [2:0] p1_add_6422_comb;
  wire [2:0] p1_add_6423_comb;
  wire [2:0] p1_add_6424_comb;
  wire [2:0] p1_add_6425_comb;
  wire [2:0] p1_add_6426_comb;
  wire [7:0] p1_clipped__8_comb;
  wire [7:0] p1_clipped__9_comb;
  wire [7:0] p1_clipped__10_comb;
  wire [7:0] p1_clipped__11_comb;
  wire [7:0] p1_clipped__12_comb;
  wire [7:0] p1_clipped__13_comb;
  wire [7:0] p1_clipped__14_comb;
  wire [7:0] p1_clipped__15_comb;
  wire [7:0] p1_result_comb[0:7];
  assign p1_array_index_5918_comb = p0_x[3'h0];
  assign p1_array_index_5919_comb = p0_x[3'h1];
  assign p1_array_index_5920_comb = p0_x[3'h6];
  assign p1_array_index_5921_comb = p0_x[3'h7];
  assign p1_array_index_5922_comb = p0_x[3'h2];
  assign p1_array_index_5923_comb = p0_x[3'h5];
  assign p1_array_index_5924_comb = p0_x[3'h3];
  assign p1_array_index_5925_comb = p0_x[3'h4];
  assign p1_concat_5950_comb = {~p1_array_index_5918_comb[7], p1_array_index_5918_comb[6:0]};
  assign p1_concat_5952_comb = {~p1_array_index_5919_comb[7], p1_array_index_5919_comb[6:0]};
  assign p1_concat_5954_comb = {~p1_array_index_5920_comb[7], p1_array_index_5920_comb[6:0]};
  assign p1_concat_5956_comb = {~p1_array_index_5921_comb[7], p1_array_index_5921_comb[6:0]};
  assign p1_concat_5959_comb = {~p1_array_index_5922_comb[7], p1_array_index_5922_comb[6:0]};
  assign p1_concat_5961_comb = {~p1_array_index_5923_comb[7], p1_array_index_5923_comb[6:0]};
  assign p1_concat_5965_comb = {~p1_array_index_5924_comb[7], p1_array_index_5924_comb[6:0]};
  assign p1_concat_5967_comb = {~p1_array_index_5925_comb[7], p1_array_index_5925_comb[6:0]};
  assign p1_smul_3303_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5950_comb, 9'h0fb);
  assign p1_smul_3302_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5952_comb, 9'h0d5);
  assign p1_smul_3297_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5954_comb, 9'h12b);
  assign p1_smul_3296_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5956_comb, 9'h105);
  assign p1_smul_3287_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5950_comb, 9'h0d5);
  assign p1_smul_3285_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5959_comb, 9'h105);
  assign p1_smul_3282_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5961_comb, 9'h0fb);
  assign p1_smul_3280_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5956_comb, 9'h12b);
  assign p1_smul_3270_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5952_comb, 9'h105);
  assign p1_smul_3268_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5965_comb, 9'h0d5);
  assign p1_smul_3267_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5967_comb, 9'h0d5);
  assign p1_smul_3265_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5954_comb, 9'h105);
  assign p1_smul_3253_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5959_comb, 9'h0d5);
  assign p1_smul_3252_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5965_comb, 9'h105);
  assign p1_smul_3251_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5967_comb, 9'h105);
  assign p1_smul_3250_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5961_comb, 9'h0d5);
  assign p1_smul_3301_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5959_comb, 8'h47);
  assign p1_smul_3317_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5965_comb, 6'h19);
  assign p1_smul_3319_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5967_comb, 6'h27);
  assign p1_smul_3298_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5961_comb, 8'hb9);
  assign p1_bit_slice_6018_comb = p1_smul_3287_NarrowedMult__comb[15:1];
  assign p1_smul_3378_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5952_comb, 6'h27);
  assign p1_bit_slice_6020_comb = p1_smul_3285_NarrowedMult__comb[15:1];
  assign p1_smul_3284_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5965_comb, 8'hb9);
  assign p1_smul_3283_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5967_comb, 8'h47);
  assign p1_bit_slice_6023_comb = p1_smul_3282_NarrowedMult__comb[15:1];
  assign p1_smul_3398_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5954_comb, 6'h19);
  assign p1_bit_slice_6025_comb = p1_smul_3280_NarrowedMult__comb[15:1];
  assign p1_smul_3271_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5950_comb, 8'h47);
  assign p1_bit_slice_6035_comb = p1_smul_3270_NarrowedMult__comb[15:1];
  assign p1_smul_3445_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5959_comb, 6'h27);
  assign p1_bit_slice_6037_comb = p1_smul_3268_NarrowedMult__comb[15:1];
  assign p1_bit_slice_6038_comb = p1_smul_3267_NarrowedMult__comb[15:1];
  assign p1_smul_3455_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5961_comb, 6'h27);
  assign p1_bit_slice_6040_comb = p1_smul_3265_NarrowedMult__comb[15:1];
  assign p1_smul_3264_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5956_comb, 8'h47);
  assign p1_smul_3506_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5950_comb, 6'h19);
  assign p1_smul_3254_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5952_comb, 8'hb9);
  assign p1_smul_3249_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5954_comb, 8'hb9);
  assign p1_smul_3534_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5956_comb, 6'h19);
  assign p1_add_6054_comb = {{1{p1_smul_3303_NarrowedMult__comb[15]}}, p1_smul_3303_NarrowedMult__comb} + {{1{p1_smul_3302_NarrowedMult__comb[15]}}, p1_smul_3302_NarrowedMult__comb};
  assign p1_add_6059_comb = {{1{p1_smul_3297_NarrowedMult__comb[15]}}, p1_smul_3297_NarrowedMult__comb} + {{1{p1_smul_3296_NarrowedMult__comb[15]}}, p1_smul_3296_NarrowedMult__comb};
  assign p1_smul_3294_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5952_comb, 7'h31);
  assign p1_smul_3293_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5959_comb, 7'h4f);
  assign p1_smul_3290_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5961_comb, 7'h4f);
  assign p1_smul_3289_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5954_comb, 7'h31);
  assign p1_smul_3279_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5950_comb, 9'h0b5);
  assign p1_smul_3278_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5952_comb, 9'h14b);
  assign p1_smul_3277_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5959_comb, 9'h14b);
  assign p1_smul_3276_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5965_comb, 9'h0b5);
  assign p1_smul_3275_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5967_comb, 9'h0b5);
  assign p1_smul_3274_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5961_comb, 9'h14b);
  assign p1_smul_3273_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5954_comb, 9'h14b);
  assign p1_smul_3272_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5956_comb, 9'h0b5);
  assign p1_smul_3263_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5950_comb, 7'h31);
  assign p1_smul_3261_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5959_comb, 7'h31);
  assign p1_smul_3258_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5961_comb, 7'h31);
  assign p1_smul_3256_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5956_comb, 7'h31);
  assign p1_add_6102_comb = {{1{p1_smul_3253_NarrowedMult__comb[15]}}, p1_smul_3253_NarrowedMult__comb} + {{1{p1_smul_3252_NarrowedMult__comb[15]}}, p1_smul_3252_NarrowedMult__comb};
  assign p1_add_6103_comb = {{1{p1_smul_3251_NarrowedMult__comb[15]}}, p1_smul_3251_NarrowedMult__comb} + {{1{p1_smul_3250_NarrowedMult__comb[15]}}, p1_smul_3250_NarrowedMult__comb};
  assign p1_bit_slice_6106_comb = p1_add_6054_comb[16:1];
  assign p1_add_6107_comb = {{1{p1_smul_3301_NarrowedMult__comb[14]}}, p1_smul_3301_NarrowedMult__comb} + {{2{p1_smul_3317_NarrowedMult__comb[13]}}, p1_smul_3317_NarrowedMult__comb};
  assign p1_add_6108_comb = {{2{p1_smul_3319_NarrowedMult__comb[13]}}, p1_smul_3319_NarrowedMult__comb} + {{1{p1_smul_3298_NarrowedMult__comb[14]}}, p1_smul_3298_NarrowedMult__comb};
  assign p1_bit_slice_6109_comb = p1_add_6059_comb[16:1];
  assign p1_smul_3295_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5950_comb, 7'h3b);
  assign p1_bit_slice_6111_comb = p1_smul_3294_NarrowedMult__comb[14:1];
  assign p1_bit_slice_6112_comb = p1_smul_3293_NarrowedMult__comb[14:1];
  assign p1_smul_3292_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5965_comb, 7'h45);
  assign p1_smul_3291_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5967_comb, 7'h45);
  assign p1_bit_slice_6115_comb = p1_smul_3290_NarrowedMult__comb[14:1];
  assign p1_bit_slice_6116_comb = p1_smul_3289_NarrowedMult__comb[14:1];
  assign p1_smul_3288_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5956_comb, 7'h3b);
  assign p1_add_6118_comb = {{1{p1_bit_slice_6018_comb[14]}}, p1_bit_slice_6018_comb} + {{2{p1_smul_3378_NarrowedMult__comb[13]}}, p1_smul_3378_NarrowedMult__comb};
  assign p1_add_6120_comb = {{1{p1_bit_slice_6020_comb[14]}}, p1_bit_slice_6020_comb} + {{1{p1_smul_3284_NarrowedMult__comb[14]}}, p1_smul_3284_NarrowedMult__comb};
  assign p1_add_6122_comb = {{1{p1_smul_3283_NarrowedMult__comb[14]}}, p1_smul_3283_NarrowedMult__comb} + {{1{p1_bit_slice_6023_comb[14]}}, p1_bit_slice_6023_comb};
  assign p1_add_6124_comb = {{2{p1_smul_3398_NarrowedMult__comb[13]}}, p1_smul_3398_NarrowedMult__comb} + {{1{p1_bit_slice_6025_comb[14]}}, p1_bit_slice_6025_comb};
  assign p1_add_6134_comb = {{1{p1_smul_3271_NarrowedMult__comb[14]}}, p1_smul_3271_NarrowedMult__comb} + {{1{p1_bit_slice_6035_comb[14]}}, p1_bit_slice_6035_comb};
  assign p1_add_6136_comb = {{2{p1_smul_3445_NarrowedMult__comb[13]}}, p1_smul_3445_NarrowedMult__comb} + {{1{p1_bit_slice_6037_comb[14]}}, p1_bit_slice_6037_comb};
  assign p1_add_6138_comb = {{1{p1_bit_slice_6038_comb[14]}}, p1_bit_slice_6038_comb} + {{2{p1_smul_3455_NarrowedMult__comb[13]}}, p1_smul_3455_NarrowedMult__comb};
  assign p1_add_6140_comb = {{1{p1_bit_slice_6040_comb[14]}}, p1_bit_slice_6040_comb} + {{1{p1_smul_3264_NarrowedMult__comb[14]}}, p1_smul_3264_NarrowedMult__comb};
  assign p1_bit_slice_6142_comb = p1_smul_3263_NarrowedMult__comb[14:1];
  assign p1_smul_3262_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5952_comb, 7'h45);
  assign p1_bit_slice_6144_comb = p1_smul_3261_NarrowedMult__comb[14:1];
  assign p1_smul_3260_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5965_comb, 7'h3b);
  assign p1_smul_3259_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5967_comb, 7'h3b);
  assign p1_bit_slice_6147_comb = p1_smul_3258_NarrowedMult__comb[14:1];
  assign p1_smul_3257_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5954_comb, 7'h45);
  assign p1_bit_slice_6149_comb = p1_smul_3256_NarrowedMult__comb[14:1];
  assign p1_add_6150_comb = {{2{p1_smul_3506_NarrowedMult__comb[13]}}, p1_smul_3506_NarrowedMult__comb} + {{1{p1_smul_3254_NarrowedMult__comb[14]}}, p1_smul_3254_NarrowedMult__comb};
  assign p1_bit_slice_6151_comb = p1_add_6102_comb[16:1];
  assign p1_bit_slice_6152_comb = p1_add_6103_comb[16:1];
  assign p1_add_6153_comb = {{1{p1_smul_3249_NarrowedMult__comb[14]}}, p1_smul_3249_NarrowedMult__comb} + {{2{p1_smul_3534_NarrowedMult__comb[13]}}, p1_smul_3534_NarrowedMult__comb};
  assign p1_concat_6174_comb = {p1_add_6118_comb, p1_smul_3287_NarrowedMult__comb[0]};
  assign p1_concat_6175_comb = {p1_add_6120_comb, p1_smul_3285_NarrowedMult__comb[0]};
  assign p1_concat_6176_comb = {p1_add_6122_comb, p1_smul_3282_NarrowedMult__comb[0]};
  assign p1_concat_6177_comb = {p1_add_6124_comb, p1_smul_3280_NarrowedMult__comb[0]};
  assign p1_add_6178_comb = {{1{p1_smul_3279_NarrowedMult__comb[15]}}, p1_smul_3279_NarrowedMult__comb} + {{1{p1_smul_3278_NarrowedMult__comb[15]}}, p1_smul_3278_NarrowedMult__comb};
  assign p1_add_6179_comb = {{1{p1_smul_3277_NarrowedMult__comb[15]}}, p1_smul_3277_NarrowedMult__comb} + {{1{p1_smul_3276_NarrowedMult__comb[15]}}, p1_smul_3276_NarrowedMult__comb};
  assign p1_add_6180_comb = {{1{p1_smul_3275_NarrowedMult__comb[15]}}, p1_smul_3275_NarrowedMult__comb} + {{1{p1_smul_3274_NarrowedMult__comb[15]}}, p1_smul_3274_NarrowedMult__comb};
  assign p1_add_6181_comb = {{1{p1_smul_3273_NarrowedMult__comb[15]}}, p1_smul_3273_NarrowedMult__comb} + {{1{p1_smul_3272_NarrowedMult__comb[15]}}, p1_smul_3272_NarrowedMult__comb};
  assign p1_concat_6182_comb = {p1_add_6134_comb, p1_smul_3270_NarrowedMult__comb[0]};
  assign p1_concat_6183_comb = {p1_add_6136_comb, p1_smul_3268_NarrowedMult__comb[0]};
  assign p1_concat_6184_comb = {p1_add_6138_comb, p1_smul_3267_NarrowedMult__comb[0]};
  assign p1_concat_6185_comb = {p1_add_6140_comb, p1_smul_3265_NarrowedMult__comb[0]};
  assign p1_add_6198_comb = {{1{p1_concat_5950_comb[7]}}, p1_concat_5950_comb} + {{1{p1_concat_5952_comb[7]}}, p1_concat_5952_comb};
  assign p1_add_6199_comb = {{1{p1_concat_5959_comb[7]}}, p1_concat_5959_comb} + {{1{p1_concat_5965_comb[7]}}, p1_concat_5965_comb};
  assign p1_add_6200_comb = {{1{p1_concat_5967_comb[7]}}, p1_concat_5967_comb} + {{1{p1_concat_5961_comb[7]}}, p1_concat_5961_comb};
  assign p1_add_6201_comb = {{1{p1_concat_5954_comb[7]}}, p1_concat_5954_comb} + {{1{p1_concat_5956_comb[7]}}, p1_concat_5956_comb};
  assign p1_add_6202_comb = {{8{p1_bit_slice_6106_comb[15]}}, p1_bit_slice_6106_comb} + {{8{p1_add_6107_comb[15]}}, p1_add_6107_comb};
  assign p1_add_6204_comb = {{8{p1_add_6108_comb[15]}}, p1_add_6108_comb} + {{8{p1_bit_slice_6109_comb[15]}}, p1_bit_slice_6109_comb};
  assign p1_add_6206_comb = {{1{p1_smul_3295_NarrowedMult__comb[13]}}, p1_smul_3295_NarrowedMult__comb} + {{1{p1_bit_slice_6111_comb[13]}}, p1_bit_slice_6111_comb};
  assign p1_add_6208_comb = {{1{p1_bit_slice_6112_comb[13]}}, p1_bit_slice_6112_comb} + {{1{p1_smul_3292_NarrowedMult__comb[13]}}, p1_smul_3292_NarrowedMult__comb};
  assign p1_add_6210_comb = {{1{p1_smul_3291_NarrowedMult__comb[13]}}, p1_smul_3291_NarrowedMult__comb} + {{1{p1_bit_slice_6115_comb[13]}}, p1_bit_slice_6115_comb};
  assign p1_add_6212_comb = {{1{p1_bit_slice_6116_comb[13]}}, p1_bit_slice_6116_comb} + {{1{p1_smul_3288_NarrowedMult__comb[13]}}, p1_smul_3288_NarrowedMult__comb};
  assign p1_sum__101_comb = {{8{p1_concat_6174_comb[16]}}, p1_concat_6174_comb};
  assign p1_sum__102_comb = {{8{p1_concat_6175_comb[16]}}, p1_concat_6175_comb};
  assign p1_sum__103_comb = {{8{p1_concat_6176_comb[16]}}, p1_concat_6176_comb};
  assign p1_sum__104_comb = {{8{p1_concat_6177_comb[16]}}, p1_concat_6177_comb};
  assign p1_sum__97_comb = {{8{p1_add_6178_comb[16]}}, p1_add_6178_comb};
  assign p1_sum__98_comb = {{8{p1_add_6179_comb[16]}}, p1_add_6179_comb};
  assign p1_sum__99_comb = {{8{p1_add_6180_comb[16]}}, p1_add_6180_comb};
  assign p1_sum__100_comb = {{8{p1_add_6181_comb[16]}}, p1_add_6181_comb};
  assign p1_sum__93_comb = {{8{p1_concat_6182_comb[16]}}, p1_concat_6182_comb};
  assign p1_sum__94_comb = {{8{p1_concat_6183_comb[16]}}, p1_concat_6183_comb};
  assign p1_sum__95_comb = {{8{p1_concat_6184_comb[16]}}, p1_concat_6184_comb};
  assign p1_sum__96_comb = {{8{p1_concat_6185_comb[16]}}, p1_concat_6185_comb};
  assign p1_add_6226_comb = {{1{p1_bit_slice_6142_comb[13]}}, p1_bit_slice_6142_comb} + {{1{p1_smul_3262_NarrowedMult__comb[13]}}, p1_smul_3262_NarrowedMult__comb};
  assign p1_add_6228_comb = {{1{p1_bit_slice_6144_comb[13]}}, p1_bit_slice_6144_comb} + {{1{p1_smul_3260_NarrowedMult__comb[13]}}, p1_smul_3260_NarrowedMult__comb};
  assign p1_add_6230_comb = {{1{p1_smul_3259_NarrowedMult__comb[13]}}, p1_smul_3259_NarrowedMult__comb} + {{1{p1_bit_slice_6147_comb[13]}}, p1_bit_slice_6147_comb};
  assign p1_add_6232_comb = {{1{p1_smul_3257_NarrowedMult__comb[13]}}, p1_smul_3257_NarrowedMult__comb} + {{1{p1_bit_slice_6149_comb[13]}}, p1_bit_slice_6149_comb};
  assign p1_add_6234_comb = {{8{p1_add_6150_comb[15]}}, p1_add_6150_comb} + {{8{p1_bit_slice_6151_comb[15]}}, p1_bit_slice_6151_comb};
  assign p1_add_6236_comb = {{8{p1_bit_slice_6152_comb[15]}}, p1_bit_slice_6152_comb} + {{8{p1_add_6153_comb[15]}}, p1_add_6153_comb};
  assign p1_sum__83_comb = {p1_add_6202_comb, p1_add_6054_comb[0]};
  assign p1_sum__84_comb = {p1_add_6204_comb, p1_add_6059_comb[0]};
  assign p1_concat_6244_comb = {p1_add_6206_comb, p1_smul_3294_NarrowedMult__comb[0]};
  assign p1_concat_6245_comb = {p1_add_6208_comb, p1_smul_3293_NarrowedMult__comb[0]};
  assign p1_concat_6246_comb = {p1_add_6210_comb, p1_smul_3290_NarrowedMult__comb[0]};
  assign p1_concat_6247_comb = {p1_add_6212_comb, p1_smul_3289_NarrowedMult__comb[0]};
  assign p1_sum__79_comb = p1_sum__101_comb + p1_sum__102_comb;
  assign p1_sum__80_comb = p1_sum__103_comb + p1_sum__104_comb;
  assign p1_sum__77_comb = p1_sum__97_comb + p1_sum__98_comb;
  assign p1_sum__78_comb = p1_sum__99_comb + p1_sum__100_comb;
  assign p1_sum__75_comb = p1_sum__93_comb + p1_sum__94_comb;
  assign p1_sum__76_comb = p1_sum__95_comb + p1_sum__96_comb;
  assign p1_concat_6254_comb = {p1_add_6226_comb, p1_smul_3263_NarrowedMult__comb[0]};
  assign p1_concat_6255_comb = {p1_add_6228_comb, p1_smul_3261_NarrowedMult__comb[0]};
  assign p1_concat_6256_comb = {p1_add_6230_comb, p1_smul_3258_NarrowedMult__comb[0]};
  assign p1_concat_6257_comb = {p1_add_6232_comb, p1_smul_3256_NarrowedMult__comb[0]};
  assign p1_sum__71_comb = {p1_add_6234_comb, p1_add_6102_comb[0]};
  assign p1_sum__72_comb = {p1_add_6236_comb, p1_add_6103_comb[0]};
  assign p1_add_6260_comb = {{15{p1_add_6198_comb[8]}}, p1_add_6198_comb} + {{15{p1_add_6199_comb[8]}}, p1_add_6199_comb};
  assign p1_add_6261_comb = {{15{p1_add_6200_comb[8]}}, p1_add_6200_comb} + {{15{p1_add_6201_comb[8]}}, p1_add_6201_comb};
  assign p1_sum__70_comb = p1_sum__83_comb + p1_sum__84_comb;
  assign p1_sum__68_comb = p1_sum__79_comb + p1_sum__80_comb;
  assign p1_sum__67_comb = p1_sum__77_comb + p1_sum__78_comb;
  assign p1_sum__66_comb = p1_sum__75_comb + p1_sum__76_comb;
  assign p1_sum__64_comb = p1_sum__71_comb + p1_sum__72_comb;
  assign p1_add_6280_comb = p1_add_6260_comb + p1_add_6261_comb;
  assign p1_add_6282_comb = p1_sum__70_comb + 25'h000_0001;
  assign p1_add_6283_comb = {{8{p1_concat_6244_comb[15]}}, p1_concat_6244_comb} + {{8{p1_concat_6245_comb[15]}}, p1_concat_6245_comb};
  assign p1_add_6284_comb = {{8{p1_concat_6246_comb[15]}}, p1_concat_6246_comb} + {{8{p1_concat_6247_comb[15]}}, p1_concat_6247_comb};
  assign p1_add_6285_comb = p1_sum__68_comb + 25'h000_0001;
  assign p1_add_6286_comb = p1_sum__67_comb + 25'h000_0001;
  assign p1_add_6287_comb = p1_sum__66_comb + 25'h000_0001;
  assign p1_add_6288_comb = {{8{p1_concat_6254_comb[15]}}, p1_concat_6254_comb} + {{8{p1_concat_6255_comb[15]}}, p1_concat_6255_comb};
  assign p1_add_6289_comb = {{8{p1_concat_6256_comb[15]}}, p1_concat_6256_comb} + {{8{p1_concat_6257_comb[15]}}, p1_concat_6257_comb};
  assign p1_add_6290_comb = p1_sum__64_comb + 25'h000_0001;
  assign p1_umul_2792_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_6280_comb, 7'h5b);
  assign p1_add_6295_comb = p1_add_6283_comb + p1_add_6284_comb;
  assign p1_add_6303_comb = p1_add_6288_comb + p1_add_6289_comb;
  assign p1_clipped__16_comb = $signed(p1_umul_2792_NarrowedMult__comb) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_umul_2792_NarrowedMult__comb) > $signed(24'h00_7fff) ? 9'h0ff : p1_umul_2792_NarrowedMult__comb[15:7]);
  assign p1_clipped__17_comb = $signed(p1_add_6282_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_6282_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_6282_comb[16:8]);
  assign p1_clipped__18_comb = $signed(p1_add_6295_comb) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_6295_comb) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_6295_comb[15:7]);
  assign p1_clipped__19_comb = $signed(p1_add_6285_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_6285_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_6285_comb[16:8]);
  assign p1_clipped__20_comb = $signed(p1_add_6286_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_6286_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_6286_comb[16:8]);
  assign p1_clipped__21_comb = $signed(p1_add_6287_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_6287_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_6287_comb[16:8]);
  assign p1_clipped__22_comb = $signed(p1_add_6303_comb) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_6303_comb) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_6303_comb[15:7]);
  assign p1_clipped__23_comb = $signed(p1_add_6290_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_6290_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_6290_comb[16:8]);
  assign p1_add_6387_comb = {{1{p1_clipped__16_comb[8]}}, p1_clipped__16_comb} + 10'h001;
  assign p1_add_6388_comb = {{1{p1_clipped__17_comb[8]}}, p1_clipped__17_comb} + 10'h001;
  assign p1_add_6389_comb = {{1{p1_clipped__18_comb[8]}}, p1_clipped__18_comb} + 10'h001;
  assign p1_add_6390_comb = {{1{p1_clipped__19_comb[8]}}, p1_clipped__19_comb} + 10'h001;
  assign p1_add_6391_comb = {{1{p1_clipped__20_comb[8]}}, p1_clipped__20_comb} + 10'h001;
  assign p1_add_6392_comb = {{1{p1_clipped__21_comb[8]}}, p1_clipped__21_comb} + 10'h001;
  assign p1_add_6393_comb = {{1{p1_clipped__22_comb[8]}}, p1_clipped__22_comb} + 10'h001;
  assign p1_add_6394_comb = {{1{p1_clipped__23_comb[8]}}, p1_clipped__23_comb} + 10'h001;
  assign p1_bit_slice_6395_comb = p1_add_6387_comb[9:8];
  assign p1_bit_slice_6396_comb = p1_add_6388_comb[9:8];
  assign p1_bit_slice_6397_comb = p1_add_6389_comb[9:8];
  assign p1_bit_slice_6398_comb = p1_add_6390_comb[9:8];
  assign p1_bit_slice_6399_comb = p1_add_6391_comb[9:8];
  assign p1_bit_slice_6400_comb = p1_add_6392_comb[9:8];
  assign p1_bit_slice_6401_comb = p1_add_6393_comb[9:8];
  assign p1_bit_slice_6402_comb = p1_add_6394_comb[9:8];
  assign p1_add_6419_comb = {{1{p1_bit_slice_6395_comb[1]}}, p1_bit_slice_6395_comb} + 3'h1;
  assign p1_add_6420_comb = {{1{p1_bit_slice_6396_comb[1]}}, p1_bit_slice_6396_comb} + 3'h1;
  assign p1_add_6421_comb = {{1{p1_bit_slice_6397_comb[1]}}, p1_bit_slice_6397_comb} + 3'h1;
  assign p1_add_6422_comb = {{1{p1_bit_slice_6398_comb[1]}}, p1_bit_slice_6398_comb} + 3'h1;
  assign p1_add_6423_comb = {{1{p1_bit_slice_6399_comb[1]}}, p1_bit_slice_6399_comb} + 3'h1;
  assign p1_add_6424_comb = {{1{p1_bit_slice_6400_comb[1]}}, p1_bit_slice_6400_comb} + 3'h1;
  assign p1_add_6425_comb = {{1{p1_bit_slice_6401_comb[1]}}, p1_bit_slice_6401_comb} + 3'h1;
  assign p1_add_6426_comb = {{1{p1_bit_slice_6402_comb[1]}}, p1_bit_slice_6402_comb} + 3'h1;
  assign p1_clipped__8_comb = p1_add_6419_comb[1] ? 8'hff : {p1_add_6419_comb[0], p1_add_6387_comb[7:1]};
  assign p1_clipped__9_comb = p1_add_6420_comb[1] ? 8'hff : {p1_add_6420_comb[0], p1_add_6388_comb[7:1]};
  assign p1_clipped__10_comb = p1_add_6421_comb[1] ? 8'hff : {p1_add_6421_comb[0], p1_add_6389_comb[7:1]};
  assign p1_clipped__11_comb = p1_add_6422_comb[1] ? 8'hff : {p1_add_6422_comb[0], p1_add_6390_comb[7:1]};
  assign p1_clipped__12_comb = p1_add_6423_comb[1] ? 8'hff : {p1_add_6423_comb[0], p1_add_6391_comb[7:1]};
  assign p1_clipped__13_comb = p1_add_6424_comb[1] ? 8'hff : {p1_add_6424_comb[0], p1_add_6392_comb[7:1]};
  assign p1_clipped__14_comb = p1_add_6425_comb[1] ? 8'hff : {p1_add_6425_comb[0], p1_add_6393_comb[7:1]};
  assign p1_clipped__15_comb = p1_add_6426_comb[1] ? 8'hff : {p1_add_6426_comb[0], p1_add_6394_comb[7:1]};
  assign p1_result_comb[0] = p1_clipped__8_comb;
  assign p1_result_comb[1] = p1_clipped__9_comb;
  assign p1_result_comb[2] = p1_clipped__10_comb;
  assign p1_result_comb[3] = p1_clipped__11_comb;
  assign p1_result_comb[4] = p1_clipped__12_comb;
  assign p1_result_comb[5] = p1_clipped__13_comb;
  assign p1_result_comb[6] = p1_clipped__14_comb;
  assign p1_result_comb[7] = p1_clipped__15_comb;

  // Registers for pipe stage 1:
  reg [7:0] p1_result[0:7];
  always @ (posedge clk) begin
    p1_result[0] <= p1_result_comb[0];
    p1_result[1] <= p1_result_comb[1];
    p1_result[2] <= p1_result_comb[2];
    p1_result[3] <= p1_result_comb[3];
    p1_result[4] <= p1_result_comb[4];
    p1_result[5] <= p1_result_comb[5];
    p1_result[6] <= p1_result_comb[6];
    p1_result[7] <= p1_result_comb[7];
  end
  assign out = {p1_result[7], p1_result[6], p1_result[5], p1_result[4], p1_result[3], p1_result[2], p1_result[1], p1_result[0]};
endmodule
