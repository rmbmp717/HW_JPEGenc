module Huffman_ACenc(
  input wire clk,
  input wire [511:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [35:0] out
);
  wire [7:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[7:0];
  assign matrix_unflattened[0][1] = matrix[15:8];
  assign matrix_unflattened[0][2] = matrix[23:16];
  assign matrix_unflattened[0][3] = matrix[31:24];
  assign matrix_unflattened[0][4] = matrix[39:32];
  assign matrix_unflattened[0][5] = matrix[47:40];
  assign matrix_unflattened[0][6] = matrix[55:48];
  assign matrix_unflattened[0][7] = matrix[63:56];
  assign matrix_unflattened[1][0] = matrix[71:64];
  assign matrix_unflattened[1][1] = matrix[79:72];
  assign matrix_unflattened[1][2] = matrix[87:80];
  assign matrix_unflattened[1][3] = matrix[95:88];
  assign matrix_unflattened[1][4] = matrix[103:96];
  assign matrix_unflattened[1][5] = matrix[111:104];
  assign matrix_unflattened[1][6] = matrix[119:112];
  assign matrix_unflattened[1][7] = matrix[127:120];
  assign matrix_unflattened[2][0] = matrix[135:128];
  assign matrix_unflattened[2][1] = matrix[143:136];
  assign matrix_unflattened[2][2] = matrix[151:144];
  assign matrix_unflattened[2][3] = matrix[159:152];
  assign matrix_unflattened[2][4] = matrix[167:160];
  assign matrix_unflattened[2][5] = matrix[175:168];
  assign matrix_unflattened[2][6] = matrix[183:176];
  assign matrix_unflattened[2][7] = matrix[191:184];
  assign matrix_unflattened[3][0] = matrix[199:192];
  assign matrix_unflattened[3][1] = matrix[207:200];
  assign matrix_unflattened[3][2] = matrix[215:208];
  assign matrix_unflattened[3][3] = matrix[223:216];
  assign matrix_unflattened[3][4] = matrix[231:224];
  assign matrix_unflattened[3][5] = matrix[239:232];
  assign matrix_unflattened[3][6] = matrix[247:240];
  assign matrix_unflattened[3][7] = matrix[255:248];
  assign matrix_unflattened[4][0] = matrix[263:256];
  assign matrix_unflattened[4][1] = matrix[271:264];
  assign matrix_unflattened[4][2] = matrix[279:272];
  assign matrix_unflattened[4][3] = matrix[287:280];
  assign matrix_unflattened[4][4] = matrix[295:288];
  assign matrix_unflattened[4][5] = matrix[303:296];
  assign matrix_unflattened[4][6] = matrix[311:304];
  assign matrix_unflattened[4][7] = matrix[319:312];
  assign matrix_unflattened[5][0] = matrix[327:320];
  assign matrix_unflattened[5][1] = matrix[335:328];
  assign matrix_unflattened[5][2] = matrix[343:336];
  assign matrix_unflattened[5][3] = matrix[351:344];
  assign matrix_unflattened[5][4] = matrix[359:352];
  assign matrix_unflattened[5][5] = matrix[367:360];
  assign matrix_unflattened[5][6] = matrix[375:368];
  assign matrix_unflattened[5][7] = matrix[383:376];
  assign matrix_unflattened[6][0] = matrix[391:384];
  assign matrix_unflattened[6][1] = matrix[399:392];
  assign matrix_unflattened[6][2] = matrix[407:400];
  assign matrix_unflattened[6][3] = matrix[415:408];
  assign matrix_unflattened[6][4] = matrix[423:416];
  assign matrix_unflattened[6][5] = matrix[431:424];
  assign matrix_unflattened[6][6] = matrix[439:432];
  assign matrix_unflattened[6][7] = matrix[447:440];
  assign matrix_unflattened[7][0] = matrix[455:448];
  assign matrix_unflattened[7][1] = matrix[463:456];
  assign matrix_unflattened[7][2] = matrix[471:464];
  assign matrix_unflattened[7][3] = matrix[479:472];
  assign matrix_unflattened[7][4] = matrix[487:480];
  assign matrix_unflattened[7][5] = matrix[495:488];
  assign matrix_unflattened[7][6] = matrix[503:496];
  assign matrix_unflattened[7][7] = matrix[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_array_index_4670_comb;
  wire [7:0] p1_array_index_4674_comb;
  wire p1_eq_4677_comb;
  wire [7:0] p1_array_index_4678_comb;
  wire p1_ne_4680_comb;
  wire p1_eq_4683_comb;
  wire [7:0] p1_array_index_4690_comb;
  wire [7:0] p1_array_index_4696_comb;
  wire p1_ne_4698_comb;
  wire [7:0] p1_array_index_4703_comb;
  wire p1_ne_4705_comb;
  wire [2:0] p1_sel_4706_comb;
  wire [7:0] p1_array_index_4708_comb;
  wire p1_ne_4710_comb;
  wire p1_eq_4713_comb;
  wire [7:0] p1_array_index_4720_comb;
  wire [7:0] p1_array_index_4726_comb;
  wire p1_ne_4728_comb;
  wire [7:0] p1_array_index_4733_comb;
  wire p1_ne_4735_comb;
  wire [3:0] p1_sel_4736_comb;
  wire [7:0] p1_array_index_4740_comb;
  wire p1_ne_4742_comb;
  wire [7:0] p1_array_index_4747_comb;
  wire p1_ne_4749_comb;
  wire [7:0] p1_array_index_4756_comb;
  wire p1_ne_4758_comb;
  wire [7:0] p1_array_index_4761_comb;
  wire [7:0] p1_array_index_4763_comb;
  wire p1_ne_4765_comb;
  wire p1_ne_4768_comb;
  wire p1_ne_4769_comb;
  wire [3:0] p1_sel_4770_comb;
  wire [3:0] p1_sel_4773_comb;
  wire [3:0] p1_run_comb;
  wire [7:0] p1_array_index_4872_comb;
  wire [7:0] p1_value_comb;
  wire p1_and_5030_comb;
  wire p1_eq_5031_comb;
  wire [7:0] p1_code_list_comb;
  wire [35:0] p1_tuple_5049_comb;
  assign p1_array_index_4670_comb = p0_matrix[3'h1][3'h7];
  assign p1_array_index_4674_comb = p0_matrix[3'h1][3'h6];
  assign p1_eq_4677_comb = p1_array_index_4670_comb == 8'h00;
  assign p1_array_index_4678_comb = p0_matrix[3'h1][3'h5];
  assign p1_ne_4680_comb = p1_array_index_4674_comb != 8'h00;
  assign p1_eq_4683_comb = p1_array_index_4678_comb == 8'h00;
  assign p1_array_index_4690_comb = p0_matrix[3'h1][3'h4];
  assign p1_array_index_4696_comb = p0_matrix[3'h1][3'h3];
  assign p1_ne_4698_comb = p1_array_index_4690_comb != 8'h00;
  assign p1_array_index_4703_comb = p0_matrix[3'h1][3'h2];
  assign p1_ne_4705_comb = p1_array_index_4696_comb != 8'h00;
  assign p1_sel_4706_comb = p1_ne_4698_comb ? 3'h3 : {1'h1, (p1_ne_4680_comb ? 2'h1 : {1'h1, p1_eq_4677_comb}) & {2{p1_eq_4683_comb}}};
  assign p1_array_index_4708_comb = p0_matrix[3'h1][3'h1];
  assign p1_ne_4710_comb = p1_array_index_4703_comb != 8'h00;
  assign p1_eq_4713_comb = p1_array_index_4708_comb == 8'h00;
  assign p1_array_index_4720_comb = p0_matrix[3'h1][3'h0];
  assign p1_array_index_4726_comb = p0_matrix[3'h0][3'h7];
  assign p1_ne_4728_comb = p1_array_index_4720_comb != 8'h00;
  assign p1_array_index_4733_comb = p0_matrix[3'h0][3'h6];
  assign p1_ne_4735_comb = p1_array_index_4726_comb != 8'h00;
  assign p1_sel_4736_comb = p1_ne_4728_comb ? 4'h7 : {1'h1, (p1_ne_4710_comb ? 3'h1 : (p1_ne_4705_comb ? 3'h2 : p1_sel_4706_comb)) & {3{p1_eq_4713_comb}}};
  assign p1_array_index_4740_comb = p0_matrix[3'h0][3'h5];
  assign p1_ne_4742_comb = p1_array_index_4733_comb != 8'h00;
  assign p1_array_index_4747_comb = p0_matrix[3'h0][3'h4];
  assign p1_ne_4749_comb = p1_array_index_4740_comb != 8'h00;
  assign p1_array_index_4756_comb = p0_matrix[3'h0][3'h3];
  assign p1_ne_4758_comb = p1_array_index_4747_comb != 8'h00;
  assign p1_array_index_4761_comb = p0_matrix[3'h0][3'h1];
  assign p1_array_index_4763_comb = p0_matrix[3'h0][3'h2];
  assign p1_ne_4765_comb = p1_array_index_4756_comb != 8'h00;
  assign p1_ne_4768_comb = p1_array_index_4761_comb != 8'h00;
  assign p1_ne_4769_comb = p1_array_index_4763_comb != 8'h00;
  assign p1_sel_4770_comb = p1_ne_4765_comb ? 4'h2 : (p1_ne_4758_comb ? 4'h3 : (p1_ne_4749_comb ? 4'h4 : (p1_ne_4742_comb ? 4'h5 : (p1_ne_4735_comb ? 4'h6 : p1_sel_4736_comb))));
  assign p1_sel_4773_comb = p1_ne_4769_comb ? 4'h1 : p1_sel_4770_comb;
  assign p1_run_comb = p1_sel_4773_comb & {4{~p1_ne_4768_comb}};
  assign p1_array_index_4872_comb = p0_matrix[3'h2][3'h0];
  assign p1_value_comb = p1_run_comb == 4'h0 ? p1_array_index_4761_comb : (p1_run_comb == 4'h1 ? p1_array_index_4763_comb : (p1_run_comb == 4'h2 ? p1_array_index_4756_comb : (p1_run_comb == 4'h3 ? p1_array_index_4747_comb : (p1_run_comb == 4'h4 ? p1_array_index_4740_comb : (p1_run_comb == 4'h5 ? p1_array_index_4733_comb : (p1_run_comb == 4'h6 ? p1_array_index_4726_comb : (p1_run_comb == 4'h7 ? p1_array_index_4720_comb : (p1_run_comb == 4'h8 ? p1_array_index_4708_comb : (p1_run_comb == 4'h9 ? p1_array_index_4703_comb : (p1_run_comb == 4'ha ? p1_array_index_4696_comb : (p1_run_comb == 4'hb ? p1_array_index_4690_comb : (p1_run_comb == 4'hc ? p1_array_index_4678_comb : (p1_run_comb == 4'hd ? p1_array_index_4674_comb : (p1_run_comb == 4'he ? p1_array_index_4670_comb : p1_array_index_4872_comb))))))))))))));
  assign p1_and_5030_comb = ~p1_ne_4768_comb & ~p1_ne_4769_comb & ~p1_ne_4765_comb & ~p1_ne_4758_comb & ~p1_ne_4749_comb & ~p1_ne_4742_comb & ~p1_ne_4735_comb & ~p1_ne_4728_comb & p1_eq_4713_comb & ~p1_ne_4710_comb & ~p1_ne_4705_comb & ~p1_ne_4698_comb & p1_eq_4683_comb & ~p1_ne_4680_comb & p1_eq_4677_comb & p1_array_index_4872_comb == 8'h00 & p0_matrix[3'h2][3'h1] == 8'h00 & p0_matrix[3'h2][3'h2] == 8'h00 & p0_matrix[3'h2][3'h3] == 8'h00 & p0_matrix[3'h2][3'h4] == 8'h00 & p0_matrix[3'h2][3'h5] == 8'h00 & p0_matrix[3'h2][3'h6] == 8'h00 & p0_matrix[3'h2][3'h7] == 8'h00 & p0_matrix[3'h3][3'h0] == 8'h00 & p0_matrix[3'h3][3'h1] == 8'h00 & p0_matrix[3'h3][3'h2] == 8'h00 & p0_matrix[3'h3][3'h3] == 8'h00 & p0_matrix[3'h3][3'h4] == 8'h00 & p0_matrix[3'h3][3'h5] == 8'h00 & p0_matrix[3'h3][3'h6] == 8'h00 & p0_matrix[3'h3][3'h7] == 8'h00 & p0_matrix[3'h4][3'h0] == 8'h00 & p0_matrix[3'h4][3'h1] == 8'h00 & p0_matrix[3'h4][3'h2] == 8'h00 & p0_matrix[3'h4][3'h3] == 8'h00 & p0_matrix[3'h4][3'h4] == 8'h00 & p0_matrix[3'h4][3'h5] == 8'h00 & p0_matrix[3'h4][3'h6] == 8'h00 & p0_matrix[3'h4][3'h7] == 8'h00 & p0_matrix[3'h5][3'h0] == 8'h00 & p0_matrix[3'h5][3'h1] == 8'h00 & p0_matrix[3'h5][3'h2] == 8'h00 & p0_matrix[3'h5][3'h3] == 8'h00 & p0_matrix[3'h5][3'h4] == 8'h00 & p0_matrix[3'h5][3'h5] == 8'h00 & p0_matrix[3'h5][3'h6] == 8'h00 & p0_matrix[3'h5][3'h7] == 8'h00 & p0_matrix[3'h6][3'h0] == 8'h00 & p0_matrix[3'h6][3'h1] == 8'h00 & p0_matrix[3'h6][3'h2] == 8'h00 & p0_matrix[3'h6][3'h3] == 8'h00 & p0_matrix[3'h6][3'h4] == 8'h00 & p0_matrix[3'h6][3'h5] == 8'h00 & p0_matrix[3'h6][3'h6] == 8'h00 & p0_matrix[3'h6][3'h7] == 8'h00 & p0_matrix[3'h7][3'h0] == 8'h00 & p0_matrix[3'h7][3'h1] == 8'h00 & p0_matrix[3'h7][3'h2] == 8'h00 & p0_matrix[3'h7][3'h3] == 8'h00 & p0_matrix[3'h7][3'h4] == 8'h00 & p0_matrix[3'h7][3'h5] == 8'h00 & p0_matrix[3'h7][3'h6] == 8'h00 & p0_matrix[3'h7][3'h7] == 8'h00;
  assign p1_eq_5031_comb = p1_run_comb == 4'hf;
  assign p1_code_list_comb = ~((|p1_value_comb[7:1]) | p1_value_comb[0]) ? 8'hff : p1_value_comb;
  assign p1_tuple_5049_comb = {{15'h0000, ~(p1_and_5030_comb | p1_eq_5031_comb)}, p1_and_5030_comb ? p0_start_pix : 8'h02, p1_code_list_comb & {8{~(p1_and_5030_comb | p1_eq_5031_comb)}}, p1_sel_4773_comb & {4{~(p1_and_5030_comb | p1_eq_5031_comb | p1_ne_4768_comb)}}};

  // Registers for pipe stage 1:
  reg [35:0] p1_tuple_5049;
  always @ (posedge clk) begin
    p1_tuple_5049 <= p1_tuple_5049_comb;
  end
  assign out = p1_tuple_5049;
endmodule
