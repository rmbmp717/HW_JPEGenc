module Huffman_ACenc(
  input wire clk,
  input wire [511:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [35:0] out
);
  wire [4:0] literal_6170[0:161];
  assign literal_6170[0] = 5'h02;
  assign literal_6170[1] = 5'h02;
  assign literal_6170[2] = 5'h03;
  assign literal_6170[3] = 5'h03;
  assign literal_6170[4] = 5'h04;
  assign literal_6170[5] = 5'h05;
  assign literal_6170[6] = 5'h05;
  assign literal_6170[7] = 5'h06;
  assign literal_6170[8] = 5'h06;
  assign literal_6170[9] = 5'h06;
  assign literal_6170[10] = 5'h07;
  assign literal_6170[11] = 5'h07;
  assign literal_6170[12] = 5'h07;
  assign literal_6170[13] = 5'h07;
  assign literal_6170[14] = 5'h07;
  assign literal_6170[15] = 5'h08;
  assign literal_6170[16] = 5'h08;
  assign literal_6170[17] = 5'h08;
  assign literal_6170[18] = 5'h08;
  assign literal_6170[19] = 5'h08;
  assign literal_6170[20] = 5'h09;
  assign literal_6170[21] = 5'h09;
  assign literal_6170[22] = 5'h09;
  assign literal_6170[23] = 5'h09;
  assign literal_6170[24] = 5'h0a;
  assign literal_6170[25] = 5'h0a;
  assign literal_6170[26] = 5'h0a;
  assign literal_6170[27] = 5'h0a;
  assign literal_6170[28] = 5'h0a;
  assign literal_6170[29] = 5'h0b;
  assign literal_6170[30] = 5'h0b;
  assign literal_6170[31] = 5'h0b;
  assign literal_6170[32] = 5'h0b;
  assign literal_6170[33] = 5'h0b;
  assign literal_6170[34] = 5'h0b;
  assign literal_6170[35] = 5'h0c;
  assign literal_6170[36] = 5'h0c;
  assign literal_6170[37] = 5'h0c;
  assign literal_6170[38] = 5'h0c;
  assign literal_6170[39] = 5'h0d;
  assign literal_6170[40] = 5'h0d;
  assign literal_6170[41] = 5'h0d;
  assign literal_6170[42] = 5'h0d;
  assign literal_6170[43] = 5'h0d;
  assign literal_6170[44] = 5'h0d;
  assign literal_6170[45] = 5'h0d;
  assign literal_6170[46] = 5'h0d;
  assign literal_6170[47] = 5'h0e;
  assign literal_6170[48] = 5'h0e;
  assign literal_6170[49] = 5'h0e;
  assign literal_6170[50] = 5'h0f;
  assign literal_6170[51] = 5'h0f;
  assign literal_6170[52] = 5'h0f;
  assign literal_6170[53] = 5'h10;
  assign literal_6170[54] = 5'h10;
  assign literal_6170[55] = 5'h10;
  assign literal_6170[56] = 5'h10;
  assign literal_6170[57] = 5'h10;
  assign literal_6170[58] = 5'h10;
  assign literal_6170[59] = 5'h10;
  assign literal_6170[60] = 5'h10;
  assign literal_6170[61] = 5'h10;
  assign literal_6170[62] = 5'h10;
  assign literal_6170[63] = 5'h10;
  assign literal_6170[64] = 5'h10;
  assign literal_6170[65] = 5'h10;
  assign literal_6170[66] = 5'h10;
  assign literal_6170[67] = 5'h10;
  assign literal_6170[68] = 5'h10;
  assign literal_6170[69] = 5'h10;
  assign literal_6170[70] = 5'h10;
  assign literal_6170[71] = 5'h10;
  assign literal_6170[72] = 5'h10;
  assign literal_6170[73] = 5'h10;
  assign literal_6170[74] = 5'h10;
  assign literal_6170[75] = 5'h10;
  assign literal_6170[76] = 5'h10;
  assign literal_6170[77] = 5'h10;
  assign literal_6170[78] = 5'h10;
  assign literal_6170[79] = 5'h10;
  assign literal_6170[80] = 5'h10;
  assign literal_6170[81] = 5'h10;
  assign literal_6170[82] = 5'h10;
  assign literal_6170[83] = 5'h10;
  assign literal_6170[84] = 5'h10;
  assign literal_6170[85] = 5'h10;
  assign literal_6170[86] = 5'h10;
  assign literal_6170[87] = 5'h10;
  assign literal_6170[88] = 5'h10;
  assign literal_6170[89] = 5'h10;
  assign literal_6170[90] = 5'h10;
  assign literal_6170[91] = 5'h10;
  assign literal_6170[92] = 5'h10;
  assign literal_6170[93] = 5'h10;
  assign literal_6170[94] = 5'h10;
  assign literal_6170[95] = 5'h10;
  assign literal_6170[96] = 5'h10;
  assign literal_6170[97] = 5'h10;
  assign literal_6170[98] = 5'h10;
  assign literal_6170[99] = 5'h10;
  assign literal_6170[100] = 5'h10;
  assign literal_6170[101] = 5'h10;
  assign literal_6170[102] = 5'h10;
  assign literal_6170[103] = 5'h10;
  assign literal_6170[104] = 5'h10;
  assign literal_6170[105] = 5'h10;
  assign literal_6170[106] = 5'h10;
  assign literal_6170[107] = 5'h10;
  assign literal_6170[108] = 5'h10;
  assign literal_6170[109] = 5'h10;
  assign literal_6170[110] = 5'h10;
  assign literal_6170[111] = 5'h10;
  assign literal_6170[112] = 5'h10;
  assign literal_6170[113] = 5'h10;
  assign literal_6170[114] = 5'h10;
  assign literal_6170[115] = 5'h10;
  assign literal_6170[116] = 5'h10;
  assign literal_6170[117] = 5'h10;
  assign literal_6170[118] = 5'h10;
  assign literal_6170[119] = 5'h10;
  assign literal_6170[120] = 5'h10;
  assign literal_6170[121] = 5'h10;
  assign literal_6170[122] = 5'h10;
  assign literal_6170[123] = 5'h10;
  assign literal_6170[124] = 5'h10;
  assign literal_6170[125] = 5'h10;
  assign literal_6170[126] = 5'h10;
  assign literal_6170[127] = 5'h10;
  assign literal_6170[128] = 5'h10;
  assign literal_6170[129] = 5'h10;
  assign literal_6170[130] = 5'h10;
  assign literal_6170[131] = 5'h10;
  assign literal_6170[132] = 5'h10;
  assign literal_6170[133] = 5'h10;
  assign literal_6170[134] = 5'h10;
  assign literal_6170[135] = 5'h10;
  assign literal_6170[136] = 5'h10;
  assign literal_6170[137] = 5'h10;
  assign literal_6170[138] = 5'h10;
  assign literal_6170[139] = 5'h10;
  assign literal_6170[140] = 5'h10;
  assign literal_6170[141] = 5'h10;
  assign literal_6170[142] = 5'h10;
  assign literal_6170[143] = 5'h10;
  assign literal_6170[144] = 5'h10;
  assign literal_6170[145] = 5'h10;
  assign literal_6170[146] = 5'h10;
  assign literal_6170[147] = 5'h10;
  assign literal_6170[148] = 5'h10;
  assign literal_6170[149] = 5'h10;
  assign literal_6170[150] = 5'h10;
  assign literal_6170[151] = 5'h10;
  assign literal_6170[152] = 5'h10;
  assign literal_6170[153] = 5'h10;
  assign literal_6170[154] = 5'h10;
  assign literal_6170[155] = 5'h10;
  assign literal_6170[156] = 5'h10;
  assign literal_6170[157] = 5'h10;
  assign literal_6170[158] = 5'h10;
  assign literal_6170[159] = 5'h10;
  assign literal_6170[160] = 5'h10;
  assign literal_6170[161] = 5'h10;
  wire [15:0] AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[0:161];
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[0] = 16'h0000;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[1] = 16'h0001;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[2] = 16'h0004;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[3] = 16'h0005;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[4] = 16'h000c;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[5] = 16'h001a;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[6] = 16'h001b;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[7] = 16'h0038;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[8] = 16'h0039;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[9] = 16'h003a;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[10] = 16'h0076;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[11] = 16'h0077;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[12] = 16'h0078;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[13] = 16'h0079;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[14] = 16'h007a;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[15] = 16'h00f6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[16] = 16'h00f7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[17] = 16'h00f8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[18] = 16'h00f9;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[19] = 16'h00fa;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[20] = 16'h01f6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[21] = 16'h01f7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[22] = 16'h01f8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[23] = 16'h01f9;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[24] = 16'h03f4;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[25] = 16'h03f5;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[26] = 16'h03f6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[27] = 16'h03f7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[28] = 16'h03f8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[29] = 16'h07f2;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[30] = 16'h07f3;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[31] = 16'h07f4;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[32] = 16'h07f5;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[33] = 16'h07f6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[34] = 16'h07f7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[35] = 16'h0ff0;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[36] = 16'h0ff1;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[37] = 16'h0ff2;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[38] = 16'h0ff3;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[39] = 16'h1fe8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[40] = 16'h1fe9;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[41] = 16'h1fea;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[42] = 16'h1feb;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[43] = 16'h1fec;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[44] = 16'h1fed;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[45] = 16'h1fee;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[46] = 16'h1fef;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[47] = 16'h3fe0;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[48] = 16'h3fe1;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[49] = 16'h3fe2;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[50] = 16'h7fc6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[51] = 16'h7fc7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[52] = 16'h7fc8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[53] = 16'hff92;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[54] = 16'hff93;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[55] = 16'hff94;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[56] = 16'hff95;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[57] = 16'hff96;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[58] = 16'hff97;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[59] = 16'hff98;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[60] = 16'hff99;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[61] = 16'hff9a;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[62] = 16'hff9b;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[63] = 16'hff9c;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[64] = 16'hff9d;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[65] = 16'hff9e;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[66] = 16'hff9f;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[67] = 16'hffa0;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[68] = 16'hffa1;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[69] = 16'hffa2;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[70] = 16'hffa3;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[71] = 16'hffa4;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[72] = 16'hffa5;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[73] = 16'hffa6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[74] = 16'hffa7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[75] = 16'hffa8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[76] = 16'hffa9;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[77] = 16'hffaa;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[78] = 16'hffab;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[79] = 16'hffac;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[80] = 16'hffad;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[81] = 16'hffae;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[82] = 16'hffaf;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[83] = 16'hffb0;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[84] = 16'hffb1;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[85] = 16'hffb2;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[86] = 16'hffb3;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[87] = 16'hffb4;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[88] = 16'hffb5;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[89] = 16'hffb6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[90] = 16'hffb7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[91] = 16'hffb8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[92] = 16'hffb9;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[93] = 16'hffba;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[94] = 16'hffbb;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[95] = 16'hffbc;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[96] = 16'hffbd;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[97] = 16'hffbe;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[98] = 16'hffbf;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[99] = 16'hffc0;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[100] = 16'hffc1;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[101] = 16'hffc2;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[102] = 16'hffc3;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[103] = 16'hffc4;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[104] = 16'hffc5;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[105] = 16'hffc6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[106] = 16'hffc7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[107] = 16'hffc8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[108] = 16'hffc9;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[109] = 16'hffca;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[110] = 16'hffcb;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[111] = 16'hffcc;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[112] = 16'hffcd;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[113] = 16'hffce;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[114] = 16'hffcf;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[115] = 16'hffd0;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[116] = 16'hffd1;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[117] = 16'hffd2;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[118] = 16'hffd3;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[119] = 16'hffd4;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[120] = 16'hffd5;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[121] = 16'hffd6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[122] = 16'hffd7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[123] = 16'hffd8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[124] = 16'hffd9;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[125] = 16'hffda;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[126] = 16'hffdb;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[127] = 16'hffdc;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[128] = 16'hffdd;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[129] = 16'hffde;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[130] = 16'hffdf;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[131] = 16'hffe0;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[132] = 16'hffe1;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[133] = 16'hffe2;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[134] = 16'hffe3;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[135] = 16'hffe4;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[136] = 16'hffe5;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[137] = 16'hffe6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[138] = 16'hffe7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[139] = 16'hffe8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[140] = 16'hffe9;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[141] = 16'hffea;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[142] = 16'hffeb;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[143] = 16'hffec;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[144] = 16'hffed;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[145] = 16'hffee;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[146] = 16'hffef;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[147] = 16'hfff0;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[148] = 16'hfff1;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[149] = 16'hfff2;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[150] = 16'hfff3;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[151] = 16'hfff4;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[152] = 16'hfff5;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[153] = 16'hfff6;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[154] = 16'hfff7;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[155] = 16'hfff8;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[156] = 16'hfff9;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[157] = 16'hfffa;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[158] = 16'hfffb;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[159] = 16'hfffc;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[160] = 16'hfffd;
  assign AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[161] = 16'hfffe;
  wire [15:0] AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[0:161];
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[0] = 16'h0000;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[1] = 16'h0001;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[2] = 16'h0004;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[3] = 16'h000a;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[4] = 16'h000b;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[5] = 16'h000c;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[6] = 16'h001a;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[7] = 16'h001b;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[8] = 16'h001c;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[9] = 16'h003a;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[10] = 16'h003b;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[11] = 16'h0078;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[12] = 16'h0079;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[13] = 16'h007a;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[14] = 16'h007b;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[15] = 16'h00f8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[16] = 16'h00f9;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[17] = 16'h01f4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[18] = 16'h01f5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[19] = 16'h01f6;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[20] = 16'h01f7;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[21] = 16'h01f8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[22] = 16'h01f9;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[23] = 16'h03f4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[24] = 16'h03f5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[25] = 16'h03f6;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[26] = 16'h03f7;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[27] = 16'h03f8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[28] = 16'h03f9;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[29] = 16'h03fa;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[30] = 16'h07f6;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[31] = 16'h07f7;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[32] = 16'h07f8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[33] = 16'h0ff2;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[34] = 16'h0ff3;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[35] = 16'h0ff4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[36] = 16'h0ff5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[37] = 16'h3fd4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[38] = 16'h3fd5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[39] = 16'hff5c;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[40] = 16'hff5d;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[41] = 16'hff5e;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[42] = 16'hff5f;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[43] = 16'h7fc0;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[44] = 16'h7fc1;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[45] = 16'hff84;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[46] = 16'hff85;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[47] = 16'hff8c;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[48] = 16'hff8d;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[49] = 16'hff8e;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[50] = 16'hff8f;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[51] = 16'hff90;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[52] = 16'hff91;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[53] = 16'hff92;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[54] = 16'hff93;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[55] = 16'hff94;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[56] = 16'hff95;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[57] = 16'hff96;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[58] = 16'hff97;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[59] = 16'hff98;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[60] = 16'hff99;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[61] = 16'hff9a;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[62] = 16'hff9b;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[63] = 16'hff9c;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[64] = 16'hff9d;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[65] = 16'hff9e;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[66] = 16'hff9f;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[67] = 16'hffa0;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[68] = 16'hffa1;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[69] = 16'hffa2;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[70] = 16'hffa3;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[71] = 16'hffa4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[72] = 16'hffa5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[73] = 16'hffa6;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[74] = 16'hffa7;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[75] = 16'hffa8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[76] = 16'hffa9;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[77] = 16'hffaa;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[78] = 16'hffab;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[79] = 16'hffac;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[80] = 16'hffad;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[81] = 16'hffae;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[82] = 16'hffaf;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[83] = 16'hffb0;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[84] = 16'hffb1;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[85] = 16'hffb2;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[86] = 16'hffb3;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[87] = 16'hffb4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[88] = 16'hffb5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[89] = 16'hffb6;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[90] = 16'hffb7;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[91] = 16'hffb8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[92] = 16'hffb9;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[93] = 16'hffba;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[94] = 16'hffbb;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[95] = 16'hffbc;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[96] = 16'hffbd;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[97] = 16'hffbe;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[98] = 16'hffbf;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[99] = 16'hffc0;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[100] = 16'hffc1;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[101] = 16'hffc2;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[102] = 16'hffc3;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[103] = 16'hffc4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[104] = 16'hffc5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[105] = 16'hffc6;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[106] = 16'hffc7;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[107] = 16'hffc8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[108] = 16'hffc9;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[109] = 16'hffca;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[110] = 16'hffcb;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[111] = 16'hffcc;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[112] = 16'hffcd;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[113] = 16'hffce;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[114] = 16'hffcf;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[115] = 16'hffd0;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[116] = 16'hffd1;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[117] = 16'hffd2;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[118] = 16'hffd3;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[119] = 16'hffd4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[120] = 16'hffd5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[121] = 16'hffd6;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[122] = 16'hffd7;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[123] = 16'hffd8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[124] = 16'hffd9;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[125] = 16'hffda;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[126] = 16'hffdb;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[127] = 16'hffdc;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[128] = 16'hffdd;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[129] = 16'hffde;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[130] = 16'hffdf;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[131] = 16'hffe0;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[132] = 16'hffe1;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[133] = 16'hffe2;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[134] = 16'hffe3;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[135] = 16'hffe4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[136] = 16'hffe5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[137] = 16'hffe6;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[138] = 16'hffe7;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[139] = 16'hffe8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[140] = 16'hffe9;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[141] = 16'hffea;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[142] = 16'hffeb;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[143] = 16'hffec;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[144] = 16'hffed;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[145] = 16'hffee;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[146] = 16'hffef;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[147] = 16'hfff0;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[148] = 16'hfff1;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[149] = 16'hfff2;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[150] = 16'hfff3;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[151] = 16'hfff4;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[152] = 16'hfff5;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[153] = 16'hfff6;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[154] = 16'hfff7;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[155] = 16'hfff8;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[156] = 16'hfff9;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[157] = 16'hfffa;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[158] = 16'hfffb;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[159] = 16'hfffc;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[160] = 16'hfffd;
  assign AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[161] = 16'hfffe;
  wire [7:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[7:0];
  assign matrix_unflattened[0][1] = matrix[15:8];
  assign matrix_unflattened[0][2] = matrix[23:16];
  assign matrix_unflattened[0][3] = matrix[31:24];
  assign matrix_unflattened[0][4] = matrix[39:32];
  assign matrix_unflattened[0][5] = matrix[47:40];
  assign matrix_unflattened[0][6] = matrix[55:48];
  assign matrix_unflattened[0][7] = matrix[63:56];
  assign matrix_unflattened[1][0] = matrix[71:64];
  assign matrix_unflattened[1][1] = matrix[79:72];
  assign matrix_unflattened[1][2] = matrix[87:80];
  assign matrix_unflattened[1][3] = matrix[95:88];
  assign matrix_unflattened[1][4] = matrix[103:96];
  assign matrix_unflattened[1][5] = matrix[111:104];
  assign matrix_unflattened[1][6] = matrix[119:112];
  assign matrix_unflattened[1][7] = matrix[127:120];
  assign matrix_unflattened[2][0] = matrix[135:128];
  assign matrix_unflattened[2][1] = matrix[143:136];
  assign matrix_unflattened[2][2] = matrix[151:144];
  assign matrix_unflattened[2][3] = matrix[159:152];
  assign matrix_unflattened[2][4] = matrix[167:160];
  assign matrix_unflattened[2][5] = matrix[175:168];
  assign matrix_unflattened[2][6] = matrix[183:176];
  assign matrix_unflattened[2][7] = matrix[191:184];
  assign matrix_unflattened[3][0] = matrix[199:192];
  assign matrix_unflattened[3][1] = matrix[207:200];
  assign matrix_unflattened[3][2] = matrix[215:208];
  assign matrix_unflattened[3][3] = matrix[223:216];
  assign matrix_unflattened[3][4] = matrix[231:224];
  assign matrix_unflattened[3][5] = matrix[239:232];
  assign matrix_unflattened[3][6] = matrix[247:240];
  assign matrix_unflattened[3][7] = matrix[255:248];
  assign matrix_unflattened[4][0] = matrix[263:256];
  assign matrix_unflattened[4][1] = matrix[271:264];
  assign matrix_unflattened[4][2] = matrix[279:272];
  assign matrix_unflattened[4][3] = matrix[287:280];
  assign matrix_unflattened[4][4] = matrix[295:288];
  assign matrix_unflattened[4][5] = matrix[303:296];
  assign matrix_unflattened[4][6] = matrix[311:304];
  assign matrix_unflattened[4][7] = matrix[319:312];
  assign matrix_unflattened[5][0] = matrix[327:320];
  assign matrix_unflattened[5][1] = matrix[335:328];
  assign matrix_unflattened[5][2] = matrix[343:336];
  assign matrix_unflattened[5][3] = matrix[351:344];
  assign matrix_unflattened[5][4] = matrix[359:352];
  assign matrix_unflattened[5][5] = matrix[367:360];
  assign matrix_unflattened[5][6] = matrix[375:368];
  assign matrix_unflattened[5][7] = matrix[383:376];
  assign matrix_unflattened[6][0] = matrix[391:384];
  assign matrix_unflattened[6][1] = matrix[399:392];
  assign matrix_unflattened[6][2] = matrix[407:400];
  assign matrix_unflattened[6][3] = matrix[415:408];
  assign matrix_unflattened[6][4] = matrix[423:416];
  assign matrix_unflattened[6][5] = matrix[431:424];
  assign matrix_unflattened[6][6] = matrix[439:432];
  assign matrix_unflattened[6][7] = matrix[447:440];
  assign matrix_unflattened[7][0] = matrix[455:448];
  assign matrix_unflattened[7][1] = matrix[463:456];
  assign matrix_unflattened[7][2] = matrix[471:464];
  assign matrix_unflattened[7][3] = matrix[479:472];
  assign matrix_unflattened[7][4] = matrix[487:480];
  assign matrix_unflattened[7][5] = matrix[495:488];
  assign matrix_unflattened[7][6] = matrix[503:496];
  assign matrix_unflattened[7][7] = matrix[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_row0_comb[0:7];
  wire [7:0] p1_row1_comb[0:7];
  wire [7:0] p1_array_concat_5303_comb[0:15];
  wire [7:0] p1_row2_comb[0:7];
  wire [7:0] p1_array_concat_5306_comb[0:23];
  wire [7:0] p1_row3_comb[0:7];
  wire [2:0] p1_idx_u8__4_squeezed_comb;
  wire [7:0] p1_idx_u8__1_comb;
  wire [7:0] p1_array_concat_5310_comb[0:31];
  wire [7:0] p1_row4_comb[0:7];
  wire [2:0] p1_idx_u8__5_squeezed_comb;
  wire [7:0] p1_si_u8__1_comb;
  wire [7:0] p1_array_concat_5314_comb[0:39];
  wire [7:0] p1_row5_comb[0:7];
  wire [2:0] p1_idx_u8__6_squeezed_comb;
  wire [7:0] p1_idx_u8__13_comb;
  wire [7:0] p1_array_concat_5320_comb[0:47];
  wire [7:0] p1_row6_comb[0:7];
  wire [2:0] p1_idx_u8__7_squeezed_comb;
  wire [6:0] p1_add_5323_comb;
  wire [7:0] p1_actual_index__13_comb;
  wire [7:0] p1_array_concat_5327_comb[0:55];
  wire [7:0] p1_row7_comb[0:7];
  wire [5:0] p1_add_5332_comb;
  wire [7:0] p1_flat_comb[0:63];
  wire [7:0] p1_actual_index__14_comb;
  wire [7:0] p1_idx_u8__11_comb;
  wire [7:0] p1_actual_index__12_comb;
  wire [7:0] p1_idx_u8__2_comb;
  wire [7:0] p1_idx_u8__3_comb;
  wire [7:0] p1_idx_u8__5_comb;
  wire [7:0] p1_idx_u8__7_comb;
  wire [7:0] p1_idx_u8__9_comb;
  wire [7:0] p1_actual_index__11_comb;
  wire [7:0] p1_and_5351_comb;
  wire [7:0] p1_actual_index__1_comb;
  wire [6:0] p1_add_5445_comb;
  wire [7:0] p1_actual_index__3_comb;
  wire [5:0] p1_add_5428_comb;
  wire [7:0] p1_actual_index__5_comb;
  wire [6:0] p1_add_5409_comb;
  wire [7:0] p1_actual_index__7_comb;
  wire [7:0] p1_actual_index__9_comb;
  wire [6:0] p1_add_5356_comb;
  wire [7:0] p1_idx_u8__15_comb;
  wire [7:0] p1_idx_u8__17_comb;
  wire [7:0] p1_idx_u8__19_comb;
  wire [7:0] p1_idx_u8__21_comb;
  wire [7:0] p1_idx_u8__23_comb;
  wire [7:0] p1_idx_u8__25_comb;
  wire [7:0] p1_idx_u8__27_comb;
  wire [7:0] p1_idx_u8__29_comb;
  wire [7:0] p1_idx_u8__31_comb;
  wire [7:0] p1_idx_u8__33_comb;
  wire [7:0] p1_idx_u8__35_comb;
  wire [7:0] p1_idx_u8__37_comb;
  wire [7:0] p1_idx_u8__39_comb;
  wire [7:0] p1_idx_u8__41_comb;
  wire [7:0] p1_idx_u8__43_comb;
  wire [7:0] p1_idx_u8__45_comb;
  wire [7:0] p1_idx_u8__47_comb;
  wire [7:0] p1_idx_u8__49_comb;
  wire [7:0] p1_idx_u8__51_comb;
  wire [7:0] p1_idx_u8__53_comb;
  wire [7:0] p1_idx_u8__55_comb;
  wire [7:0] p1_idx_u8__57_comb;
  wire [7:0] p1_idx_u8__59_comb;
  wire [7:0] p1_idx_u8__61_comb;
  wire [7:0] p1_and_5359_comb;
  wire p1_eq_5362_comb;
  wire [7:0] p1_and_5363_comb;
  wire [4:0] p1_add_5375_comb;
  wire [7:0] p1_actual_index__15_comb;
  wire [3:0] p1_add_5548_comb;
  wire [7:0] p1_actual_index__17_comb;
  wire [6:0] p1_add_5550_comb;
  wire [7:0] p1_actual_index__19_comb;
  wire [5:0] p1_add_5552_comb;
  wire [7:0] p1_actual_index__21_comb;
  wire [6:0] p1_add_5554_comb;
  wire [7:0] p1_actual_index__23_comb;
  wire [4:0] p1_add_5556_comb;
  wire [7:0] p1_actual_index__25_comb;
  wire [6:0] p1_add_5558_comb;
  wire [7:0] p1_actual_index__27_comb;
  wire [5:0] p1_add_5560_comb;
  wire [7:0] p1_actual_index__29_comb;
  wire [6:0] p1_add_5562_comb;
  wire [7:0] p1_actual_index__31_comb;
  wire [2:0] p1_add_5564_comb;
  wire [7:0] p1_actual_index__33_comb;
  wire [6:0] p1_add_5566_comb;
  wire [7:0] p1_actual_index__35_comb;
  wire [5:0] p1_add_5568_comb;
  wire [7:0] p1_actual_index__37_comb;
  wire [6:0] p1_add_5570_comb;
  wire [7:0] p1_actual_index__39_comb;
  wire [4:0] p1_add_5572_comb;
  wire [7:0] p1_actual_index__41_comb;
  wire [6:0] p1_add_5574_comb;
  wire [7:0] p1_actual_index__43_comb;
  wire [5:0] p1_add_5576_comb;
  wire [7:0] p1_actual_index__45_comb;
  wire [6:0] p1_add_5578_comb;
  wire [7:0] p1_actual_index__47_comb;
  wire [3:0] p1_add_5580_comb;
  wire [7:0] p1_actual_index__49_comb;
  wire [6:0] p1_add_5582_comb;
  wire [7:0] p1_actual_index__51_comb;
  wire [5:0] p1_add_5584_comb;
  wire [7:0] p1_actual_index__53_comb;
  wire [6:0] p1_add_5586_comb;
  wire [7:0] p1_actual_index__55_comb;
  wire [4:0] p1_add_5588_comb;
  wire [7:0] p1_actual_index__57_comb;
  wire [6:0] p1_add_5590_comb;
  wire [7:0] p1_actual_index__59_comb;
  wire [5:0] p1_add_5592_comb;
  wire [7:0] p1_actual_index__61_comb;
  wire [6:0] p1_add_5594_comb;
  wire p1_ne_5371_comb;
  wire [1:0] p1_idx_u8__1_squeezed_comb;
  wire p1_eq_5374_comb;
  wire [7:0] p1_actual_index__2_comb;
  wire [7:0] p1_actual_index__4_comb;
  wire [7:0] p1_actual_index__6_comb;
  wire [7:0] p1_actual_index__10_comb;
  wire [7:0] p1_actual_index__8_comb;
  wire [7:0] p1_actual_index__16_comb;
  wire [7:0] p1_actual_index__18_comb;
  wire [7:0] p1_actual_index__20_comb;
  wire [7:0] p1_actual_index__22_comb;
  wire [7:0] p1_actual_index__24_comb;
  wire [7:0] p1_actual_index__26_comb;
  wire [7:0] p1_actual_index__28_comb;
  wire [7:0] p1_actual_index__30_comb;
  wire [7:0] p1_actual_index__32_comb;
  wire [7:0] p1_actual_index__34_comb;
  wire [7:0] p1_actual_index__36_comb;
  wire [7:0] p1_actual_index__38_comb;
  wire [7:0] p1_actual_index__40_comb;
  wire [7:0] p1_actual_index__42_comb;
  wire [7:0] p1_actual_index__44_comb;
  wire [7:0] p1_actual_index__46_comb;
  wire [7:0] p1_actual_index__48_comb;
  wire [7:0] p1_actual_index__50_comb;
  wire [7:0] p1_actual_index__52_comb;
  wire [7:0] p1_actual_index__54_comb;
  wire [7:0] p1_actual_index__56_comb;
  wire [7:0] p1_actual_index__58_comb;
  wire [7:0] p1_actual_index__60_comb;
  wire [7:0] p1_actual_index__62_comb;
  wire [7:0] p1_and_5391_comb;
  wire [7:0] p1_and_5489_comb;
  wire [7:0] p1_and_5491_comb;
  wire [7:0] p1_and_5486_comb;
  wire [7:0] p1_and_5479_comb;
  wire [7:0] p1_and_5472_comb;
  wire [7:0] p1_and_5461_comb;
  wire [7:0] p1_and_5452_comb;
  wire [7:0] p1_and_5442_comb;
  wire [7:0] p1_and_5412_comb;
  wire [7:0] p1_and_5401_comb;
  wire p1_ne_5403_comb;
  wire p1_ne_5494_comb;
  wire p1_ne_5495_comb;
  wire p1_ne_5493_comb;
  wire p1_ne_5488_comb;
  wire p1_ne_5481_comb;
  wire p1_ne_5474_comb;
  wire p1_ne_5463_comb;
  wire p1_ne_5454_comb;
  wire [7:0] p1_and_5417_comb;
  wire p1_ne_5424_comb;
  wire p1_ne_5414_comb;
  wire [2:0] p1_sel_5415_comb;
  wire p1_not_5496_comb;
  wire p1_eq_5426_comb;
  wire [2:0] p1_sel_5425_comb;
  wire p1_and_6016_comb;
  assign p1_row0_comb[0] = p0_matrix[3'h0][0];
  assign p1_row0_comb[1] = p0_matrix[3'h0][1];
  assign p1_row0_comb[2] = p0_matrix[3'h0][2];
  assign p1_row0_comb[3] = p0_matrix[3'h0][3];
  assign p1_row0_comb[4] = p0_matrix[3'h0][4];
  assign p1_row0_comb[5] = p0_matrix[3'h0][5];
  assign p1_row0_comb[6] = p0_matrix[3'h0][6];
  assign p1_row0_comb[7] = p0_matrix[3'h0][7];
  assign p1_row1_comb[0] = p0_matrix[3'h1][0];
  assign p1_row1_comb[1] = p0_matrix[3'h1][1];
  assign p1_row1_comb[2] = p0_matrix[3'h1][2];
  assign p1_row1_comb[3] = p0_matrix[3'h1][3];
  assign p1_row1_comb[4] = p0_matrix[3'h1][4];
  assign p1_row1_comb[5] = p0_matrix[3'h1][5];
  assign p1_row1_comb[6] = p0_matrix[3'h1][6];
  assign p1_row1_comb[7] = p0_matrix[3'h1][7];
  assign p1_array_concat_5303_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_5303_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_5303_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_5303_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_5303_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_5303_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_5303_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_5303_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_5303_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_5303_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_5303_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_5303_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_5303_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_5303_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_5303_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_5303_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_5306_comb[0] = p1_array_concat_5303_comb[0];
  assign p1_array_concat_5306_comb[1] = p1_array_concat_5303_comb[1];
  assign p1_array_concat_5306_comb[2] = p1_array_concat_5303_comb[2];
  assign p1_array_concat_5306_comb[3] = p1_array_concat_5303_comb[3];
  assign p1_array_concat_5306_comb[4] = p1_array_concat_5303_comb[4];
  assign p1_array_concat_5306_comb[5] = p1_array_concat_5303_comb[5];
  assign p1_array_concat_5306_comb[6] = p1_array_concat_5303_comb[6];
  assign p1_array_concat_5306_comb[7] = p1_array_concat_5303_comb[7];
  assign p1_array_concat_5306_comb[8] = p1_array_concat_5303_comb[8];
  assign p1_array_concat_5306_comb[9] = p1_array_concat_5303_comb[9];
  assign p1_array_concat_5306_comb[10] = p1_array_concat_5303_comb[10];
  assign p1_array_concat_5306_comb[11] = p1_array_concat_5303_comb[11];
  assign p1_array_concat_5306_comb[12] = p1_array_concat_5303_comb[12];
  assign p1_array_concat_5306_comb[13] = p1_array_concat_5303_comb[13];
  assign p1_array_concat_5306_comb[14] = p1_array_concat_5303_comb[14];
  assign p1_array_concat_5306_comb[15] = p1_array_concat_5303_comb[15];
  assign p1_array_concat_5306_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_5306_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_5306_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_5306_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_5306_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_5306_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_5306_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_5306_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_idx_u8__4_squeezed_comb = 3'h4;
  assign p1_idx_u8__1_comb = 8'h01;
  assign p1_array_concat_5310_comb[0] = p1_array_concat_5306_comb[0];
  assign p1_array_concat_5310_comb[1] = p1_array_concat_5306_comb[1];
  assign p1_array_concat_5310_comb[2] = p1_array_concat_5306_comb[2];
  assign p1_array_concat_5310_comb[3] = p1_array_concat_5306_comb[3];
  assign p1_array_concat_5310_comb[4] = p1_array_concat_5306_comb[4];
  assign p1_array_concat_5310_comb[5] = p1_array_concat_5306_comb[5];
  assign p1_array_concat_5310_comb[6] = p1_array_concat_5306_comb[6];
  assign p1_array_concat_5310_comb[7] = p1_array_concat_5306_comb[7];
  assign p1_array_concat_5310_comb[8] = p1_array_concat_5306_comb[8];
  assign p1_array_concat_5310_comb[9] = p1_array_concat_5306_comb[9];
  assign p1_array_concat_5310_comb[10] = p1_array_concat_5306_comb[10];
  assign p1_array_concat_5310_comb[11] = p1_array_concat_5306_comb[11];
  assign p1_array_concat_5310_comb[12] = p1_array_concat_5306_comb[12];
  assign p1_array_concat_5310_comb[13] = p1_array_concat_5306_comb[13];
  assign p1_array_concat_5310_comb[14] = p1_array_concat_5306_comb[14];
  assign p1_array_concat_5310_comb[15] = p1_array_concat_5306_comb[15];
  assign p1_array_concat_5310_comb[16] = p1_array_concat_5306_comb[16];
  assign p1_array_concat_5310_comb[17] = p1_array_concat_5306_comb[17];
  assign p1_array_concat_5310_comb[18] = p1_array_concat_5306_comb[18];
  assign p1_array_concat_5310_comb[19] = p1_array_concat_5306_comb[19];
  assign p1_array_concat_5310_comb[20] = p1_array_concat_5306_comb[20];
  assign p1_array_concat_5310_comb[21] = p1_array_concat_5306_comb[21];
  assign p1_array_concat_5310_comb[22] = p1_array_concat_5306_comb[22];
  assign p1_array_concat_5310_comb[23] = p1_array_concat_5306_comb[23];
  assign p1_array_concat_5310_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_5310_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_5310_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_5310_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_5310_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_5310_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_5310_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_5310_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[p1_idx_u8__4_squeezed_comb][0];
  assign p1_row4_comb[1] = p0_matrix[p1_idx_u8__4_squeezed_comb][1];
  assign p1_row4_comb[2] = p0_matrix[p1_idx_u8__4_squeezed_comb][2];
  assign p1_row4_comb[3] = p0_matrix[p1_idx_u8__4_squeezed_comb][3];
  assign p1_row4_comb[4] = p0_matrix[p1_idx_u8__4_squeezed_comb][4];
  assign p1_row4_comb[5] = p0_matrix[p1_idx_u8__4_squeezed_comb][5];
  assign p1_row4_comb[6] = p0_matrix[p1_idx_u8__4_squeezed_comb][6];
  assign p1_row4_comb[7] = p0_matrix[p1_idx_u8__4_squeezed_comb][7];
  assign p1_idx_u8__5_squeezed_comb = 3'h5;
  assign p1_si_u8__1_comb = p0_start_pix + p1_idx_u8__1_comb;
  assign p1_array_concat_5314_comb[0] = p1_array_concat_5310_comb[0];
  assign p1_array_concat_5314_comb[1] = p1_array_concat_5310_comb[1];
  assign p1_array_concat_5314_comb[2] = p1_array_concat_5310_comb[2];
  assign p1_array_concat_5314_comb[3] = p1_array_concat_5310_comb[3];
  assign p1_array_concat_5314_comb[4] = p1_array_concat_5310_comb[4];
  assign p1_array_concat_5314_comb[5] = p1_array_concat_5310_comb[5];
  assign p1_array_concat_5314_comb[6] = p1_array_concat_5310_comb[6];
  assign p1_array_concat_5314_comb[7] = p1_array_concat_5310_comb[7];
  assign p1_array_concat_5314_comb[8] = p1_array_concat_5310_comb[8];
  assign p1_array_concat_5314_comb[9] = p1_array_concat_5310_comb[9];
  assign p1_array_concat_5314_comb[10] = p1_array_concat_5310_comb[10];
  assign p1_array_concat_5314_comb[11] = p1_array_concat_5310_comb[11];
  assign p1_array_concat_5314_comb[12] = p1_array_concat_5310_comb[12];
  assign p1_array_concat_5314_comb[13] = p1_array_concat_5310_comb[13];
  assign p1_array_concat_5314_comb[14] = p1_array_concat_5310_comb[14];
  assign p1_array_concat_5314_comb[15] = p1_array_concat_5310_comb[15];
  assign p1_array_concat_5314_comb[16] = p1_array_concat_5310_comb[16];
  assign p1_array_concat_5314_comb[17] = p1_array_concat_5310_comb[17];
  assign p1_array_concat_5314_comb[18] = p1_array_concat_5310_comb[18];
  assign p1_array_concat_5314_comb[19] = p1_array_concat_5310_comb[19];
  assign p1_array_concat_5314_comb[20] = p1_array_concat_5310_comb[20];
  assign p1_array_concat_5314_comb[21] = p1_array_concat_5310_comb[21];
  assign p1_array_concat_5314_comb[22] = p1_array_concat_5310_comb[22];
  assign p1_array_concat_5314_comb[23] = p1_array_concat_5310_comb[23];
  assign p1_array_concat_5314_comb[24] = p1_array_concat_5310_comb[24];
  assign p1_array_concat_5314_comb[25] = p1_array_concat_5310_comb[25];
  assign p1_array_concat_5314_comb[26] = p1_array_concat_5310_comb[26];
  assign p1_array_concat_5314_comb[27] = p1_array_concat_5310_comb[27];
  assign p1_array_concat_5314_comb[28] = p1_array_concat_5310_comb[28];
  assign p1_array_concat_5314_comb[29] = p1_array_concat_5310_comb[29];
  assign p1_array_concat_5314_comb[30] = p1_array_concat_5310_comb[30];
  assign p1_array_concat_5314_comb[31] = p1_array_concat_5310_comb[31];
  assign p1_array_concat_5314_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_5314_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_5314_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_5314_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_5314_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_5314_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_5314_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_5314_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[p1_idx_u8__5_squeezed_comb][0];
  assign p1_row5_comb[1] = p0_matrix[p1_idx_u8__5_squeezed_comb][1];
  assign p1_row5_comb[2] = p0_matrix[p1_idx_u8__5_squeezed_comb][2];
  assign p1_row5_comb[3] = p0_matrix[p1_idx_u8__5_squeezed_comb][3];
  assign p1_row5_comb[4] = p0_matrix[p1_idx_u8__5_squeezed_comb][4];
  assign p1_row5_comb[5] = p0_matrix[p1_idx_u8__5_squeezed_comb][5];
  assign p1_row5_comb[6] = p0_matrix[p1_idx_u8__5_squeezed_comb][6];
  assign p1_row5_comb[7] = p0_matrix[p1_idx_u8__5_squeezed_comb][7];
  assign p1_idx_u8__6_squeezed_comb = 3'h6;
  assign p1_idx_u8__13_comb = 8'h0d;
  assign p1_array_concat_5320_comb[0] = p1_array_concat_5314_comb[0];
  assign p1_array_concat_5320_comb[1] = p1_array_concat_5314_comb[1];
  assign p1_array_concat_5320_comb[2] = p1_array_concat_5314_comb[2];
  assign p1_array_concat_5320_comb[3] = p1_array_concat_5314_comb[3];
  assign p1_array_concat_5320_comb[4] = p1_array_concat_5314_comb[4];
  assign p1_array_concat_5320_comb[5] = p1_array_concat_5314_comb[5];
  assign p1_array_concat_5320_comb[6] = p1_array_concat_5314_comb[6];
  assign p1_array_concat_5320_comb[7] = p1_array_concat_5314_comb[7];
  assign p1_array_concat_5320_comb[8] = p1_array_concat_5314_comb[8];
  assign p1_array_concat_5320_comb[9] = p1_array_concat_5314_comb[9];
  assign p1_array_concat_5320_comb[10] = p1_array_concat_5314_comb[10];
  assign p1_array_concat_5320_comb[11] = p1_array_concat_5314_comb[11];
  assign p1_array_concat_5320_comb[12] = p1_array_concat_5314_comb[12];
  assign p1_array_concat_5320_comb[13] = p1_array_concat_5314_comb[13];
  assign p1_array_concat_5320_comb[14] = p1_array_concat_5314_comb[14];
  assign p1_array_concat_5320_comb[15] = p1_array_concat_5314_comb[15];
  assign p1_array_concat_5320_comb[16] = p1_array_concat_5314_comb[16];
  assign p1_array_concat_5320_comb[17] = p1_array_concat_5314_comb[17];
  assign p1_array_concat_5320_comb[18] = p1_array_concat_5314_comb[18];
  assign p1_array_concat_5320_comb[19] = p1_array_concat_5314_comb[19];
  assign p1_array_concat_5320_comb[20] = p1_array_concat_5314_comb[20];
  assign p1_array_concat_5320_comb[21] = p1_array_concat_5314_comb[21];
  assign p1_array_concat_5320_comb[22] = p1_array_concat_5314_comb[22];
  assign p1_array_concat_5320_comb[23] = p1_array_concat_5314_comb[23];
  assign p1_array_concat_5320_comb[24] = p1_array_concat_5314_comb[24];
  assign p1_array_concat_5320_comb[25] = p1_array_concat_5314_comb[25];
  assign p1_array_concat_5320_comb[26] = p1_array_concat_5314_comb[26];
  assign p1_array_concat_5320_comb[27] = p1_array_concat_5314_comb[27];
  assign p1_array_concat_5320_comb[28] = p1_array_concat_5314_comb[28];
  assign p1_array_concat_5320_comb[29] = p1_array_concat_5314_comb[29];
  assign p1_array_concat_5320_comb[30] = p1_array_concat_5314_comb[30];
  assign p1_array_concat_5320_comb[31] = p1_array_concat_5314_comb[31];
  assign p1_array_concat_5320_comb[32] = p1_array_concat_5314_comb[32];
  assign p1_array_concat_5320_comb[33] = p1_array_concat_5314_comb[33];
  assign p1_array_concat_5320_comb[34] = p1_array_concat_5314_comb[34];
  assign p1_array_concat_5320_comb[35] = p1_array_concat_5314_comb[35];
  assign p1_array_concat_5320_comb[36] = p1_array_concat_5314_comb[36];
  assign p1_array_concat_5320_comb[37] = p1_array_concat_5314_comb[37];
  assign p1_array_concat_5320_comb[38] = p1_array_concat_5314_comb[38];
  assign p1_array_concat_5320_comb[39] = p1_array_concat_5314_comb[39];
  assign p1_array_concat_5320_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_5320_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_5320_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_5320_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_5320_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_5320_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_5320_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_5320_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[p1_idx_u8__6_squeezed_comb][0];
  assign p1_row6_comb[1] = p0_matrix[p1_idx_u8__6_squeezed_comb][1];
  assign p1_row6_comb[2] = p0_matrix[p1_idx_u8__6_squeezed_comb][2];
  assign p1_row6_comb[3] = p0_matrix[p1_idx_u8__6_squeezed_comb][3];
  assign p1_row6_comb[4] = p0_matrix[p1_idx_u8__6_squeezed_comb][4];
  assign p1_row6_comb[5] = p0_matrix[p1_idx_u8__6_squeezed_comb][5];
  assign p1_row6_comb[6] = p0_matrix[p1_idx_u8__6_squeezed_comb][6];
  assign p1_row6_comb[7] = p0_matrix[p1_idx_u8__6_squeezed_comb][7];
  assign p1_idx_u8__7_squeezed_comb = 3'h7;
  assign p1_add_5323_comb = p1_si_u8__1_comb[7:1] + 7'h07;
  assign p1_actual_index__13_comb = p1_si_u8__1_comb + p1_idx_u8__13_comb;
  assign p1_array_concat_5327_comb[0] = p1_array_concat_5320_comb[0];
  assign p1_array_concat_5327_comb[1] = p1_array_concat_5320_comb[1];
  assign p1_array_concat_5327_comb[2] = p1_array_concat_5320_comb[2];
  assign p1_array_concat_5327_comb[3] = p1_array_concat_5320_comb[3];
  assign p1_array_concat_5327_comb[4] = p1_array_concat_5320_comb[4];
  assign p1_array_concat_5327_comb[5] = p1_array_concat_5320_comb[5];
  assign p1_array_concat_5327_comb[6] = p1_array_concat_5320_comb[6];
  assign p1_array_concat_5327_comb[7] = p1_array_concat_5320_comb[7];
  assign p1_array_concat_5327_comb[8] = p1_array_concat_5320_comb[8];
  assign p1_array_concat_5327_comb[9] = p1_array_concat_5320_comb[9];
  assign p1_array_concat_5327_comb[10] = p1_array_concat_5320_comb[10];
  assign p1_array_concat_5327_comb[11] = p1_array_concat_5320_comb[11];
  assign p1_array_concat_5327_comb[12] = p1_array_concat_5320_comb[12];
  assign p1_array_concat_5327_comb[13] = p1_array_concat_5320_comb[13];
  assign p1_array_concat_5327_comb[14] = p1_array_concat_5320_comb[14];
  assign p1_array_concat_5327_comb[15] = p1_array_concat_5320_comb[15];
  assign p1_array_concat_5327_comb[16] = p1_array_concat_5320_comb[16];
  assign p1_array_concat_5327_comb[17] = p1_array_concat_5320_comb[17];
  assign p1_array_concat_5327_comb[18] = p1_array_concat_5320_comb[18];
  assign p1_array_concat_5327_comb[19] = p1_array_concat_5320_comb[19];
  assign p1_array_concat_5327_comb[20] = p1_array_concat_5320_comb[20];
  assign p1_array_concat_5327_comb[21] = p1_array_concat_5320_comb[21];
  assign p1_array_concat_5327_comb[22] = p1_array_concat_5320_comb[22];
  assign p1_array_concat_5327_comb[23] = p1_array_concat_5320_comb[23];
  assign p1_array_concat_5327_comb[24] = p1_array_concat_5320_comb[24];
  assign p1_array_concat_5327_comb[25] = p1_array_concat_5320_comb[25];
  assign p1_array_concat_5327_comb[26] = p1_array_concat_5320_comb[26];
  assign p1_array_concat_5327_comb[27] = p1_array_concat_5320_comb[27];
  assign p1_array_concat_5327_comb[28] = p1_array_concat_5320_comb[28];
  assign p1_array_concat_5327_comb[29] = p1_array_concat_5320_comb[29];
  assign p1_array_concat_5327_comb[30] = p1_array_concat_5320_comb[30];
  assign p1_array_concat_5327_comb[31] = p1_array_concat_5320_comb[31];
  assign p1_array_concat_5327_comb[32] = p1_array_concat_5320_comb[32];
  assign p1_array_concat_5327_comb[33] = p1_array_concat_5320_comb[33];
  assign p1_array_concat_5327_comb[34] = p1_array_concat_5320_comb[34];
  assign p1_array_concat_5327_comb[35] = p1_array_concat_5320_comb[35];
  assign p1_array_concat_5327_comb[36] = p1_array_concat_5320_comb[36];
  assign p1_array_concat_5327_comb[37] = p1_array_concat_5320_comb[37];
  assign p1_array_concat_5327_comb[38] = p1_array_concat_5320_comb[38];
  assign p1_array_concat_5327_comb[39] = p1_array_concat_5320_comb[39];
  assign p1_array_concat_5327_comb[40] = p1_array_concat_5320_comb[40];
  assign p1_array_concat_5327_comb[41] = p1_array_concat_5320_comb[41];
  assign p1_array_concat_5327_comb[42] = p1_array_concat_5320_comb[42];
  assign p1_array_concat_5327_comb[43] = p1_array_concat_5320_comb[43];
  assign p1_array_concat_5327_comb[44] = p1_array_concat_5320_comb[44];
  assign p1_array_concat_5327_comb[45] = p1_array_concat_5320_comb[45];
  assign p1_array_concat_5327_comb[46] = p1_array_concat_5320_comb[46];
  assign p1_array_concat_5327_comb[47] = p1_array_concat_5320_comb[47];
  assign p1_array_concat_5327_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_5327_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_5327_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_5327_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_5327_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_5327_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_5327_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_5327_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[p1_idx_u8__7_squeezed_comb][0];
  assign p1_row7_comb[1] = p0_matrix[p1_idx_u8__7_squeezed_comb][1];
  assign p1_row7_comb[2] = p0_matrix[p1_idx_u8__7_squeezed_comb][2];
  assign p1_row7_comb[3] = p0_matrix[p1_idx_u8__7_squeezed_comb][3];
  assign p1_row7_comb[4] = p0_matrix[p1_idx_u8__7_squeezed_comb][4];
  assign p1_row7_comb[5] = p0_matrix[p1_idx_u8__7_squeezed_comb][5];
  assign p1_row7_comb[6] = p0_matrix[p1_idx_u8__7_squeezed_comb][6];
  assign p1_row7_comb[7] = p0_matrix[p1_idx_u8__7_squeezed_comb][7];
  assign p1_add_5332_comb = p1_si_u8__1_comb[7:2] + 6'h03;
  assign p1_flat_comb[0] = p1_array_concat_5327_comb[0];
  assign p1_flat_comb[1] = p1_array_concat_5327_comb[1];
  assign p1_flat_comb[2] = p1_array_concat_5327_comb[2];
  assign p1_flat_comb[3] = p1_array_concat_5327_comb[3];
  assign p1_flat_comb[4] = p1_array_concat_5327_comb[4];
  assign p1_flat_comb[5] = p1_array_concat_5327_comb[5];
  assign p1_flat_comb[6] = p1_array_concat_5327_comb[6];
  assign p1_flat_comb[7] = p1_array_concat_5327_comb[7];
  assign p1_flat_comb[8] = p1_array_concat_5327_comb[8];
  assign p1_flat_comb[9] = p1_array_concat_5327_comb[9];
  assign p1_flat_comb[10] = p1_array_concat_5327_comb[10];
  assign p1_flat_comb[11] = p1_array_concat_5327_comb[11];
  assign p1_flat_comb[12] = p1_array_concat_5327_comb[12];
  assign p1_flat_comb[13] = p1_array_concat_5327_comb[13];
  assign p1_flat_comb[14] = p1_array_concat_5327_comb[14];
  assign p1_flat_comb[15] = p1_array_concat_5327_comb[15];
  assign p1_flat_comb[16] = p1_array_concat_5327_comb[16];
  assign p1_flat_comb[17] = p1_array_concat_5327_comb[17];
  assign p1_flat_comb[18] = p1_array_concat_5327_comb[18];
  assign p1_flat_comb[19] = p1_array_concat_5327_comb[19];
  assign p1_flat_comb[20] = p1_array_concat_5327_comb[20];
  assign p1_flat_comb[21] = p1_array_concat_5327_comb[21];
  assign p1_flat_comb[22] = p1_array_concat_5327_comb[22];
  assign p1_flat_comb[23] = p1_array_concat_5327_comb[23];
  assign p1_flat_comb[24] = p1_array_concat_5327_comb[24];
  assign p1_flat_comb[25] = p1_array_concat_5327_comb[25];
  assign p1_flat_comb[26] = p1_array_concat_5327_comb[26];
  assign p1_flat_comb[27] = p1_array_concat_5327_comb[27];
  assign p1_flat_comb[28] = p1_array_concat_5327_comb[28];
  assign p1_flat_comb[29] = p1_array_concat_5327_comb[29];
  assign p1_flat_comb[30] = p1_array_concat_5327_comb[30];
  assign p1_flat_comb[31] = p1_array_concat_5327_comb[31];
  assign p1_flat_comb[32] = p1_array_concat_5327_comb[32];
  assign p1_flat_comb[33] = p1_array_concat_5327_comb[33];
  assign p1_flat_comb[34] = p1_array_concat_5327_comb[34];
  assign p1_flat_comb[35] = p1_array_concat_5327_comb[35];
  assign p1_flat_comb[36] = p1_array_concat_5327_comb[36];
  assign p1_flat_comb[37] = p1_array_concat_5327_comb[37];
  assign p1_flat_comb[38] = p1_array_concat_5327_comb[38];
  assign p1_flat_comb[39] = p1_array_concat_5327_comb[39];
  assign p1_flat_comb[40] = p1_array_concat_5327_comb[40];
  assign p1_flat_comb[41] = p1_array_concat_5327_comb[41];
  assign p1_flat_comb[42] = p1_array_concat_5327_comb[42];
  assign p1_flat_comb[43] = p1_array_concat_5327_comb[43];
  assign p1_flat_comb[44] = p1_array_concat_5327_comb[44];
  assign p1_flat_comb[45] = p1_array_concat_5327_comb[45];
  assign p1_flat_comb[46] = p1_array_concat_5327_comb[46];
  assign p1_flat_comb[47] = p1_array_concat_5327_comb[47];
  assign p1_flat_comb[48] = p1_array_concat_5327_comb[48];
  assign p1_flat_comb[49] = p1_array_concat_5327_comb[49];
  assign p1_flat_comb[50] = p1_array_concat_5327_comb[50];
  assign p1_flat_comb[51] = p1_array_concat_5327_comb[51];
  assign p1_flat_comb[52] = p1_array_concat_5327_comb[52];
  assign p1_flat_comb[53] = p1_array_concat_5327_comb[53];
  assign p1_flat_comb[54] = p1_array_concat_5327_comb[54];
  assign p1_flat_comb[55] = p1_array_concat_5327_comb[55];
  assign p1_flat_comb[56] = p1_row7_comb[0];
  assign p1_flat_comb[57] = p1_row7_comb[1];
  assign p1_flat_comb[58] = p1_row7_comb[2];
  assign p1_flat_comb[59] = p1_row7_comb[3];
  assign p1_flat_comb[60] = p1_row7_comb[4];
  assign p1_flat_comb[61] = p1_row7_comb[5];
  assign p1_flat_comb[62] = p1_row7_comb[6];
  assign p1_flat_comb[63] = p1_row7_comb[7];
  assign p1_actual_index__14_comb = {p1_add_5323_comb, p1_si_u8__1_comb[0]};
  assign p1_idx_u8__11_comb = 8'h0b;
  assign p1_actual_index__12_comb = {p1_add_5332_comb, p1_si_u8__1_comb[1:0]};
  assign p1_idx_u8__2_comb = 8'h01;
  assign p1_idx_u8__3_comb = 8'h03;
  assign p1_idx_u8__5_comb = 8'h05;
  assign p1_idx_u8__7_comb = 8'h07;
  assign p1_idx_u8__9_comb = 8'h09;
  assign p1_actual_index__11_comb = p1_si_u8__1_comb + p1_idx_u8__11_comb;
  assign p1_and_5351_comb = p1_flat_comb[p1_actual_index__14_comb > 8'h3f ? 6'h3f : p1_actual_index__14_comb[5:0]] & {8{~(p1_add_5323_comb[5] | p1_add_5323_comb[6])}};
  assign p1_actual_index__1_comb = p1_si_u8__1_comb + p1_idx_u8__2_comb;
  assign p1_add_5445_comb = p1_si_u8__1_comb[7:1] + 7'h01;
  assign p1_actual_index__3_comb = p1_si_u8__1_comb + p1_idx_u8__3_comb;
  assign p1_add_5428_comb = p1_si_u8__1_comb[7:2] + 6'h01;
  assign p1_actual_index__5_comb = p1_si_u8__1_comb + p1_idx_u8__5_comb;
  assign p1_add_5409_comb = p1_si_u8__1_comb[7:1] + 7'h03;
  assign p1_actual_index__7_comb = p1_si_u8__1_comb + p1_idx_u8__7_comb;
  assign p1_actual_index__9_comb = p1_si_u8__1_comb + p1_idx_u8__9_comb;
  assign p1_add_5356_comb = p1_si_u8__1_comb[7:1] + 7'h05;
  assign p1_idx_u8__15_comb = 8'h0f;
  assign p1_idx_u8__17_comb = 8'h11;
  assign p1_idx_u8__19_comb = 8'h13;
  assign p1_idx_u8__21_comb = 8'h15;
  assign p1_idx_u8__23_comb = 8'h17;
  assign p1_idx_u8__25_comb = 8'h19;
  assign p1_idx_u8__27_comb = 8'h1b;
  assign p1_idx_u8__29_comb = 8'h1d;
  assign p1_idx_u8__31_comb = 8'h1f;
  assign p1_idx_u8__33_comb = 8'h21;
  assign p1_idx_u8__35_comb = 8'h23;
  assign p1_idx_u8__37_comb = 8'h25;
  assign p1_idx_u8__39_comb = 8'h27;
  assign p1_idx_u8__41_comb = 8'h29;
  assign p1_idx_u8__43_comb = 8'h2b;
  assign p1_idx_u8__45_comb = 8'h2d;
  assign p1_idx_u8__47_comb = 8'h2f;
  assign p1_idx_u8__49_comb = 8'h31;
  assign p1_idx_u8__51_comb = 8'h33;
  assign p1_idx_u8__53_comb = 8'h35;
  assign p1_idx_u8__55_comb = 8'h37;
  assign p1_idx_u8__57_comb = 8'h39;
  assign p1_idx_u8__59_comb = 8'h3b;
  assign p1_idx_u8__61_comb = 8'h3d;
  assign p1_and_5359_comb = p1_flat_comb[p1_actual_index__13_comb > 8'h3f ? 6'h3f : p1_actual_index__13_comb[5:0]] & {8{~(p1_actual_index__13_comb[6] | p1_actual_index__13_comb[7])}};
  assign p1_eq_5362_comb = p1_and_5351_comb == 8'h00;
  assign p1_and_5363_comb = p1_flat_comb[p1_actual_index__12_comb > 8'h3f ? 6'h3f : p1_actual_index__12_comb[5:0]] & {8{~(p1_add_5332_comb[4] | p1_add_5332_comb[5])}};
  assign p1_add_5375_comb = p1_si_u8__1_comb[7:3] + 5'h01;
  assign p1_actual_index__15_comb = p1_si_u8__1_comb + p1_idx_u8__15_comb;
  assign p1_add_5548_comb = p1_si_u8__1_comb[7:4] + 4'h1;
  assign p1_actual_index__17_comb = p1_si_u8__1_comb + p1_idx_u8__17_comb;
  assign p1_add_5550_comb = p1_si_u8__1_comb[7:1] + 7'h09;
  assign p1_actual_index__19_comb = p1_si_u8__1_comb + p1_idx_u8__19_comb;
  assign p1_add_5552_comb = p1_si_u8__1_comb[7:2] + 6'h05;
  assign p1_actual_index__21_comb = p1_si_u8__1_comb + p1_idx_u8__21_comb;
  assign p1_add_5554_comb = p1_si_u8__1_comb[7:1] + 7'h0b;
  assign p1_actual_index__23_comb = p1_si_u8__1_comb + p1_idx_u8__23_comb;
  assign p1_add_5556_comb = p1_si_u8__1_comb[7:3] + 5'h03;
  assign p1_actual_index__25_comb = p1_si_u8__1_comb + p1_idx_u8__25_comb;
  assign p1_add_5558_comb = p1_si_u8__1_comb[7:1] + 7'h0d;
  assign p1_actual_index__27_comb = p1_si_u8__1_comb + p1_idx_u8__27_comb;
  assign p1_add_5560_comb = p1_si_u8__1_comb[7:2] + 6'h07;
  assign p1_actual_index__29_comb = p1_si_u8__1_comb + p1_idx_u8__29_comb;
  assign p1_add_5562_comb = p1_si_u8__1_comb[7:1] + 7'h0f;
  assign p1_actual_index__31_comb = p1_si_u8__1_comb + p1_idx_u8__31_comb;
  assign p1_add_5564_comb = p1_si_u8__1_comb[7:5] + 3'h1;
  assign p1_actual_index__33_comb = p1_si_u8__1_comb + p1_idx_u8__33_comb;
  assign p1_add_5566_comb = p1_si_u8__1_comb[7:1] + 7'h11;
  assign p1_actual_index__35_comb = p1_si_u8__1_comb + p1_idx_u8__35_comb;
  assign p1_add_5568_comb = p1_si_u8__1_comb[7:2] + 6'h09;
  assign p1_actual_index__37_comb = p1_si_u8__1_comb + p1_idx_u8__37_comb;
  assign p1_add_5570_comb = p1_si_u8__1_comb[7:1] + 7'h13;
  assign p1_actual_index__39_comb = p1_si_u8__1_comb + p1_idx_u8__39_comb;
  assign p1_add_5572_comb = p1_si_u8__1_comb[7:3] + 5'h05;
  assign p1_actual_index__41_comb = p1_si_u8__1_comb + p1_idx_u8__41_comb;
  assign p1_add_5574_comb = p1_si_u8__1_comb[7:1] + 7'h15;
  assign p1_actual_index__43_comb = p1_si_u8__1_comb + p1_idx_u8__43_comb;
  assign p1_add_5576_comb = p1_si_u8__1_comb[7:2] + 6'h0b;
  assign p1_actual_index__45_comb = p1_si_u8__1_comb + p1_idx_u8__45_comb;
  assign p1_add_5578_comb = p1_si_u8__1_comb[7:1] + 7'h17;
  assign p1_actual_index__47_comb = p1_si_u8__1_comb + p1_idx_u8__47_comb;
  assign p1_add_5580_comb = p1_si_u8__1_comb[7:4] + 4'h3;
  assign p1_actual_index__49_comb = p1_si_u8__1_comb + p1_idx_u8__49_comb;
  assign p1_add_5582_comb = p1_si_u8__1_comb[7:1] + 7'h19;
  assign p1_actual_index__51_comb = p1_si_u8__1_comb + p1_idx_u8__51_comb;
  assign p1_add_5584_comb = p1_si_u8__1_comb[7:2] + 6'h0d;
  assign p1_actual_index__53_comb = p1_si_u8__1_comb + p1_idx_u8__53_comb;
  assign p1_add_5586_comb = p1_si_u8__1_comb[7:1] + 7'h1b;
  assign p1_actual_index__55_comb = p1_si_u8__1_comb + p1_idx_u8__55_comb;
  assign p1_add_5588_comb = p1_si_u8__1_comb[7:3] + 5'h07;
  assign p1_actual_index__57_comb = p1_si_u8__1_comb + p1_idx_u8__57_comb;
  assign p1_add_5590_comb = p1_si_u8__1_comb[7:1] + 7'h1d;
  assign p1_actual_index__59_comb = p1_si_u8__1_comb + p1_idx_u8__59_comb;
  assign p1_add_5592_comb = p1_si_u8__1_comb[7:2] + 6'h0f;
  assign p1_actual_index__61_comb = p1_si_u8__1_comb + p1_idx_u8__61_comb;
  assign p1_add_5594_comb = p1_si_u8__1_comb[7:1] + 7'h1f;
  assign p1_ne_5371_comb = p1_and_5359_comb != 8'h00;
  assign p1_idx_u8__1_squeezed_comb = 2'h1;
  assign p1_eq_5374_comb = p1_and_5363_comb == 8'h00;
  assign p1_actual_index__2_comb = {p1_add_5445_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__4_comb = {p1_add_5428_comb, p1_si_u8__1_comb[1:0]};
  assign p1_actual_index__6_comb = {p1_add_5409_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__10_comb = {p1_add_5356_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__8_comb = {p1_add_5375_comb, p1_si_u8__1_comb[2:0]};
  assign p1_actual_index__16_comb = {p1_add_5548_comb, p1_si_u8__1_comb[3:0]};
  assign p1_actual_index__18_comb = {p1_add_5550_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__20_comb = {p1_add_5552_comb, p1_si_u8__1_comb[1:0]};
  assign p1_actual_index__22_comb = {p1_add_5554_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__24_comb = {p1_add_5556_comb, p1_si_u8__1_comb[2:0]};
  assign p1_actual_index__26_comb = {p1_add_5558_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__28_comb = {p1_add_5560_comb, p1_si_u8__1_comb[1:0]};
  assign p1_actual_index__30_comb = {p1_add_5562_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__32_comb = {p1_add_5564_comb, p1_si_u8__1_comb[4:0]};
  assign p1_actual_index__34_comb = {p1_add_5566_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__36_comb = {p1_add_5568_comb, p1_si_u8__1_comb[1:0]};
  assign p1_actual_index__38_comb = {p1_add_5570_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__40_comb = {p1_add_5572_comb, p1_si_u8__1_comb[2:0]};
  assign p1_actual_index__42_comb = {p1_add_5574_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__44_comb = {p1_add_5576_comb, p1_si_u8__1_comb[1:0]};
  assign p1_actual_index__46_comb = {p1_add_5578_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__48_comb = {p1_add_5580_comb, p1_si_u8__1_comb[3:0]};
  assign p1_actual_index__50_comb = {p1_add_5582_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__52_comb = {p1_add_5584_comb, p1_si_u8__1_comb[1:0]};
  assign p1_actual_index__54_comb = {p1_add_5586_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__56_comb = {p1_add_5588_comb, p1_si_u8__1_comb[2:0]};
  assign p1_actual_index__58_comb = {p1_add_5590_comb, p1_si_u8__1_comb[0]};
  assign p1_actual_index__60_comb = {p1_add_5592_comb, p1_si_u8__1_comb[1:0]};
  assign p1_actual_index__62_comb = {p1_add_5594_comb, p1_si_u8__1_comb[0]};
  assign p1_and_5391_comb = p1_flat_comb[p1_actual_index__11_comb > 8'h3f ? 6'h3f : p1_actual_index__11_comb[5:0]] & {8{~(p1_actual_index__11_comb[6] | p1_actual_index__11_comb[7])}};
  assign p1_and_5489_comb = p1_flat_comb[p1_si_u8__1_comb > 8'h3f ? 6'h3f : p1_si_u8__1_comb[5:0]] & {8{~(p1_si_u8__1_comb[6] | p1_si_u8__1_comb[7])}};
  assign p1_and_5491_comb = p1_flat_comb[p1_actual_index__1_comb > 8'h3f ? 6'h3f : p1_actual_index__1_comb[5:0]] & {8{~(p1_actual_index__1_comb[6] | p1_actual_index__1_comb[7])}};
  assign p1_and_5486_comb = p1_flat_comb[p1_actual_index__2_comb > 8'h3f ? 6'h3f : p1_actual_index__2_comb[5:0]] & {8{~(p1_add_5445_comb[5] | p1_add_5445_comb[6])}};
  assign p1_and_5479_comb = p1_flat_comb[p1_actual_index__3_comb > 8'h3f ? 6'h3f : p1_actual_index__3_comb[5:0]] & {8{~(p1_actual_index__3_comb[6] | p1_actual_index__3_comb[7])}};
  assign p1_and_5472_comb = p1_flat_comb[p1_actual_index__4_comb > 8'h3f ? 6'h3f : p1_actual_index__4_comb[5:0]] & {8{~(p1_add_5428_comb[4] | p1_add_5428_comb[5])}};
  assign p1_and_5461_comb = p1_flat_comb[p1_actual_index__5_comb > 8'h3f ? 6'h3f : p1_actual_index__5_comb[5:0]] & {8{~(p1_actual_index__5_comb[6] | p1_actual_index__5_comb[7])}};
  assign p1_and_5452_comb = p1_flat_comb[p1_actual_index__6_comb > 8'h3f ? 6'h3f : p1_actual_index__6_comb[5:0]] & {8{~(p1_add_5409_comb[5] | p1_add_5409_comb[6])}};
  assign p1_and_5442_comb = p1_flat_comb[p1_actual_index__7_comb > 8'h3f ? 6'h3f : p1_actual_index__7_comb[5:0]] & {8{~(p1_actual_index__7_comb[6] | p1_actual_index__7_comb[7])}};
  assign p1_and_5412_comb = p1_flat_comb[p1_actual_index__9_comb > 8'h3f ? 6'h3f : p1_actual_index__9_comb[5:0]] & {8{~(p1_actual_index__9_comb[6] | p1_actual_index__9_comb[7])}};
  assign p1_and_5401_comb = p1_flat_comb[p1_actual_index__10_comb > 8'h3f ? 6'h3f : p1_actual_index__10_comb[5:0]] & {8{~(p1_add_5356_comb[5] | p1_add_5356_comb[6])}};
  assign p1_ne_5403_comb = p1_and_5391_comb != 8'h00;
  assign p1_ne_5494_comb = p1_and_5489_comb != 8'h00;
  assign p1_ne_5495_comb = p1_and_5491_comb != 8'h00;
  assign p1_ne_5493_comb = p1_and_5486_comb != 8'h00;
  assign p1_ne_5488_comb = p1_and_5479_comb != 8'h00;
  assign p1_ne_5481_comb = p1_and_5472_comb != 8'h00;
  assign p1_ne_5474_comb = p1_and_5461_comb != 8'h00;
  assign p1_ne_5463_comb = p1_and_5452_comb != 8'h00;
  assign p1_ne_5454_comb = p1_and_5442_comb != 8'h00;
  assign p1_and_5417_comb = p1_flat_comb[p1_actual_index__8_comb > 8'h3f ? 6'h3f : p1_actual_index__8_comb[5:0]] & {8{~(p1_add_5375_comb[3] | p1_add_5375_comb[4])}};
  assign p1_ne_5424_comb = p1_and_5412_comb != 8'h00;
  assign p1_ne_5414_comb = p1_and_5401_comb != 8'h00;
  assign p1_sel_5415_comb = p1_ne_5403_comb ? 3'h3 : {1'h1, (p1_ne_5371_comb ? p1_idx_u8__1_squeezed_comb : {1'h1, p1_eq_5362_comb}) & {2{p1_eq_5374_comb}}};
  assign p1_not_5496_comb = ~p1_ne_5494_comb;
  assign p1_eq_5426_comb = p1_and_5417_comb == 8'h00;
  assign p1_sel_5425_comb = p1_ne_5414_comb ? 3'h2 : p1_sel_5415_comb;
  assign p1_and_6016_comb = p1_not_5496_comb & ~p1_ne_5495_comb & ~p1_ne_5493_comb & ~p1_ne_5488_comb & ~p1_ne_5481_comb & ~p1_ne_5474_comb & ~p1_ne_5463_comb & ~p1_ne_5454_comb & p1_eq_5426_comb & ~p1_ne_5424_comb & ~p1_ne_5414_comb & ~p1_ne_5403_comb & p1_eq_5374_comb & ~p1_ne_5371_comb & p1_eq_5362_comb & (p1_flat_comb[p1_actual_index__15_comb > 8'h3f ? 6'h3f : p1_actual_index__15_comb[5:0]] & {8{~(p1_actual_index__15_comb[6] | p1_actual_index__15_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__16_comb > 8'h3f ? 6'h3f : p1_actual_index__16_comb[5:0]] & {8{~(p1_add_5548_comb[2] | p1_add_5548_comb[3])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__17_comb > 8'h3f ? 6'h3f : p1_actual_index__17_comb[5:0]] & {8{~(p1_actual_index__17_comb[6] | p1_actual_index__17_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__18_comb > 8'h3f ? 6'h3f : p1_actual_index__18_comb[5:0]] & {8{~(p1_add_5550_comb[5] | p1_add_5550_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__19_comb > 8'h3f ? 6'h3f : p1_actual_index__19_comb[5:0]] & {8{~(p1_actual_index__19_comb[6] | p1_actual_index__19_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__20_comb > 8'h3f ? 6'h3f : p1_actual_index__20_comb[5:0]] & {8{~(p1_add_5552_comb[4] | p1_add_5552_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__21_comb > 8'h3f ? 6'h3f : p1_actual_index__21_comb[5:0]] & {8{~(p1_actual_index__21_comb[6] | p1_actual_index__21_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__22_comb > 8'h3f ? 6'h3f : p1_actual_index__22_comb[5:0]] & {8{~(p1_add_5554_comb[5] | p1_add_5554_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__23_comb > 8'h3f ? 6'h3f : p1_actual_index__23_comb[5:0]] & {8{~(p1_actual_index__23_comb[6] | p1_actual_index__23_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__24_comb > 8'h3f ? 6'h3f : p1_actual_index__24_comb[5:0]] & {8{~(p1_add_5556_comb[3] | p1_add_5556_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__25_comb > 8'h3f ? 6'h3f : p1_actual_index__25_comb[5:0]] & {8{~(p1_actual_index__25_comb[6] | p1_actual_index__25_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__26_comb > 8'h3f ? 6'h3f : p1_actual_index__26_comb[5:0]] & {8{~(p1_add_5558_comb[5] | p1_add_5558_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__27_comb > 8'h3f ? 6'h3f : p1_actual_index__27_comb[5:0]] & {8{~(p1_actual_index__27_comb[6] | p1_actual_index__27_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__28_comb > 8'h3f ? 6'h3f : p1_actual_index__28_comb[5:0]] & {8{~(p1_add_5560_comb[4] | p1_add_5560_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__29_comb > 8'h3f ? 6'h3f : p1_actual_index__29_comb[5:0]] & {8{~(p1_actual_index__29_comb[6] | p1_actual_index__29_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__30_comb > 8'h3f ? 6'h3f : p1_actual_index__30_comb[5:0]] & {8{~(p1_add_5562_comb[5] | p1_add_5562_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__31_comb > 8'h3f ? 6'h3f : p1_actual_index__31_comb[5:0]] & {8{~(p1_actual_index__31_comb[6] | p1_actual_index__31_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__32_comb > 8'h3f ? 6'h3f : p1_actual_index__32_comb[5:0]] & {8{~(p1_add_5564_comb[1] | p1_add_5564_comb[2])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__33_comb > 8'h3f ? 6'h3f : p1_actual_index__33_comb[5:0]] & {8{~(p1_actual_index__33_comb[6] | p1_actual_index__33_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__34_comb > 8'h3f ? 6'h3f : p1_actual_index__34_comb[5:0]] & {8{~(p1_add_5566_comb[5] | p1_add_5566_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__35_comb > 8'h3f ? 6'h3f : p1_actual_index__35_comb[5:0]] & {8{~(p1_actual_index__35_comb[6] | p1_actual_index__35_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__36_comb > 8'h3f ? 6'h3f : p1_actual_index__36_comb[5:0]] & {8{~(p1_add_5568_comb[4] | p1_add_5568_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__37_comb > 8'h3f ? 6'h3f : p1_actual_index__37_comb[5:0]] & {8{~(p1_actual_index__37_comb[6] | p1_actual_index__37_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__38_comb > 8'h3f ? 6'h3f : p1_actual_index__38_comb[5:0]] & {8{~(p1_add_5570_comb[5] | p1_add_5570_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__39_comb > 8'h3f ? 6'h3f : p1_actual_index__39_comb[5:0]] & {8{~(p1_actual_index__39_comb[6] | p1_actual_index__39_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__40_comb > 8'h3f ? 6'h3f : p1_actual_index__40_comb[5:0]] & {8{~(p1_add_5572_comb[3] | p1_add_5572_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__41_comb > 8'h3f ? 6'h3f : p1_actual_index__41_comb[5:0]] & {8{~(p1_actual_index__41_comb[6] | p1_actual_index__41_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__42_comb > 8'h3f ? 6'h3f : p1_actual_index__42_comb[5:0]] & {8{~(p1_add_5574_comb[5] | p1_add_5574_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__43_comb > 8'h3f ? 6'h3f : p1_actual_index__43_comb[5:0]] & {8{~(p1_actual_index__43_comb[6] | p1_actual_index__43_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__44_comb > 8'h3f ? 6'h3f : p1_actual_index__44_comb[5:0]] & {8{~(p1_add_5576_comb[4] | p1_add_5576_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__45_comb > 8'h3f ? 6'h3f : p1_actual_index__45_comb[5:0]] & {8{~(p1_actual_index__45_comb[6] | p1_actual_index__45_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__46_comb > 8'h3f ? 6'h3f : p1_actual_index__46_comb[5:0]] & {8{~(p1_add_5578_comb[5] | p1_add_5578_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__47_comb > 8'h3f ? 6'h3f : p1_actual_index__47_comb[5:0]] & {8{~(p1_actual_index__47_comb[6] | p1_actual_index__47_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__48_comb > 8'h3f ? 6'h3f : p1_actual_index__48_comb[5:0]] & {8{~(p1_add_5580_comb[2] | p1_add_5580_comb[3])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__49_comb > 8'h3f ? 6'h3f : p1_actual_index__49_comb[5:0]] & {8{~(p1_actual_index__49_comb[6] | p1_actual_index__49_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__50_comb > 8'h3f ? 6'h3f : p1_actual_index__50_comb[5:0]] & {8{~(p1_add_5582_comb[5] | p1_add_5582_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__51_comb > 8'h3f ? 6'h3f : p1_actual_index__51_comb[5:0]] & {8{~(p1_actual_index__51_comb[6] | p1_actual_index__51_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__52_comb > 8'h3f ? 6'h3f : p1_actual_index__52_comb[5:0]] & {8{~(p1_add_5584_comb[4] | p1_add_5584_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__53_comb > 8'h3f ? 6'h3f : p1_actual_index__53_comb[5:0]] & {8{~(p1_actual_index__53_comb[6] | p1_actual_index__53_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__54_comb > 8'h3f ? 6'h3f : p1_actual_index__54_comb[5:0]] & {8{~(p1_add_5586_comb[5] | p1_add_5586_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__55_comb > 8'h3f ? 6'h3f : p1_actual_index__55_comb[5:0]] & {8{~(p1_actual_index__55_comb[6] | p1_actual_index__55_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__56_comb > 8'h3f ? 6'h3f : p1_actual_index__56_comb[5:0]] & {8{~(p1_add_5588_comb[3] | p1_add_5588_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__57_comb > 8'h3f ? 6'h3f : p1_actual_index__57_comb[5:0]] & {8{~(p1_actual_index__57_comb[6] | p1_actual_index__57_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__58_comb > 8'h3f ? 6'h3f : p1_actual_index__58_comb[5:0]] & {8{~(p1_add_5590_comb[5] | p1_add_5590_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__59_comb > 8'h3f ? 6'h3f : p1_actual_index__59_comb[5:0]] & {8{~(p1_actual_index__59_comb[6] | p1_actual_index__59_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__60_comb > 8'h3f ? 6'h3f : p1_actual_index__60_comb[5:0]] & {8{~(p1_add_5592_comb[4] | p1_add_5592_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__61_comb > 8'h3f ? 6'h3f : p1_actual_index__61_comb[5:0]] & {8{~(p1_actual_index__61_comb[6] | p1_actual_index__61_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__62_comb > 8'h3f ? 6'h3f : p1_actual_index__62_comb[5:0]] & {8{~(p1_add_5594_comb[5] | p1_add_5594_comb[6])}}) == 8'h00;

  // Registers for pipe stage 1:
  reg [7:0] p1_start_pix;
  reg p1_is_luminance;
  reg [7:0] p1_and_5351;
  reg [7:0] p1_and_5359;
  reg [7:0] p1_and_5363;
  reg [7:0] p1_and_5391;
  reg [7:0] p1_and_5401;
  reg [7:0] p1_and_5412;
  reg [7:0] p1_and_5417;
  reg p1_ne_5424;
  reg [2:0] p1_sel_5425;
  reg p1_eq_5426;
  reg [7:0] p1_and_5442;
  reg [7:0] p1_and_5452;
  reg p1_ne_5454;
  reg [7:0] p1_and_5461;
  reg p1_ne_5463;
  reg [7:0] p1_and_5472;
  reg p1_ne_5474;
  reg [7:0] p1_and_5479;
  reg p1_ne_5481;
  reg [7:0] p1_and_5486;
  reg p1_ne_5488;
  reg [7:0] p1_and_5489;
  reg [7:0] p1_and_5491;
  reg p1_ne_5493;
  reg p1_ne_5494;
  reg p1_ne_5495;
  reg p1_not_5496;
  reg p1_and_6016;
  always @ (posedge clk) begin
    p1_start_pix <= p0_start_pix;
    p1_is_luminance <= p0_is_luminance;
    p1_and_5351 <= p1_and_5351_comb;
    p1_and_5359 <= p1_and_5359_comb;
    p1_and_5363 <= p1_and_5363_comb;
    p1_and_5391 <= p1_and_5391_comb;
    p1_and_5401 <= p1_and_5401_comb;
    p1_and_5412 <= p1_and_5412_comb;
    p1_and_5417 <= p1_and_5417_comb;
    p1_ne_5424 <= p1_ne_5424_comb;
    p1_sel_5425 <= p1_sel_5425_comb;
    p1_eq_5426 <= p1_eq_5426_comb;
    p1_and_5442 <= p1_and_5442_comb;
    p1_and_5452 <= p1_and_5452_comb;
    p1_ne_5454 <= p1_ne_5454_comb;
    p1_and_5461 <= p1_and_5461_comb;
    p1_ne_5463 <= p1_ne_5463_comb;
    p1_and_5472 <= p1_and_5472_comb;
    p1_ne_5474 <= p1_ne_5474_comb;
    p1_and_5479 <= p1_and_5479_comb;
    p1_ne_5481 <= p1_ne_5481_comb;
    p1_and_5486 <= p1_and_5486_comb;
    p1_ne_5488 <= p1_ne_5488_comb;
    p1_and_5489 <= p1_and_5489_comb;
    p1_and_5491 <= p1_and_5491_comb;
    p1_ne_5493 <= p1_ne_5493_comb;
    p1_ne_5494 <= p1_ne_5494_comb;
    p1_ne_5495 <= p1_ne_5495_comb;
    p1_not_5496 <= p1_not_5496_comb;
    p1_and_6016 <= p1_and_6016_comb;
  end

  // ===== Pipe stage 2:
  wire [3:0] p2_sel_6086_comb;
  wire [3:0] p2_sel_6092_comb;
  wire [3:0] p2_sel_6096_comb;
  wire [3:0] p2_run_comb;
  wire [7:0] p2_value_comb;
  wire p2_eq_6116_comb;
  wire [1:0] p2_idx_u8__1_squeezed__1_comb;
  wire [1:0] p2_idx_u8__2_squeezed_comb;
  wire [1:0] p2_idx_u8__3_squeezed_comb;
  wire [3:0] p2_add_6113_comb;
  wire [1:0] p2_sel_6109_comb;
  wire [3:0] p2_run_u8__1_comb;
  wire [3:0] p2_and_6120_comb;
  assign p2_sel_6086_comb = p1_ne_5463 ? 4'h6 : (p1_ne_5454 ? 4'h7 : {1'h1, (p1_ne_5424 ? 3'h1 : p1_sel_5425) & {3{p1_eq_5426}}});
  assign p2_sel_6092_comb = p1_ne_5488 ? 4'h3 : (p1_ne_5481 ? 4'h4 : (p1_ne_5474 ? 4'h5 : p2_sel_6086_comb));
  assign p2_sel_6096_comb = p1_ne_5495 ? 4'h1 : (p1_ne_5493 ? 4'h2 : p2_sel_6092_comb);
  assign p2_run_comb = p2_sel_6096_comb & {4{p1_not_5496}};
  assign p2_value_comb = p2_run_comb == 4'h0 ? p1_and_5489 : (p2_run_comb == 4'h1 ? p1_and_5491 : (p2_run_comb == 4'h2 ? p1_and_5486 : (p2_run_comb == 4'h3 ? p1_and_5479 : (p2_run_comb == 4'h4 ? p1_and_5472 : (p2_run_comb == 4'h5 ? p1_and_5461 : (p2_run_comb == 4'h6 ? p1_and_5452 : (p2_run_comb == 4'h7 ? p1_and_5442 : (p2_run_comb == 4'h8 ? p1_and_5417 : (p2_run_comb == 4'h9 ? p1_and_5412 : (p2_run_comb == 4'ha ? p1_and_5401 : (p2_run_comb == 4'hb ? p1_and_5391 : (p2_run_comb == 4'hc ? p1_and_5363 : (p2_run_comb == 4'hd ? p1_and_5359 : (p2_run_comb == 4'he ? p1_and_5351 : 8'h00))))))))))))));
  assign p2_eq_6116_comb = p2_run_comb == 4'hf;
  assign p2_idx_u8__1_squeezed__1_comb = 2'h1;
  assign p2_idx_u8__2_squeezed_comb = 2'h2;
  assign p2_idx_u8__3_squeezed_comb = 2'h3;
  assign p2_add_6113_comb = p2_sel_6092_comb + 4'h7;
  assign p2_sel_6109_comb = |p2_value_comb[7:2] ? p2_idx_u8__3_squeezed_comb : (|p2_value_comb[7:1] ? p2_idx_u8__2_squeezed_comb : p2_idx_u8__1_squeezed__1_comb);
  assign p2_run_u8__1_comb = p2_run_comb < 4'ha ? p2_run_comb : p2_add_6113_comb;
  assign p2_and_6120_comb = p2_sel_6096_comb & {4{~(p1_and_6016 | p2_eq_6116_comb | p1_ne_5494)}};

  // Registers for pipe stage 2:
  reg [7:0] p2_start_pix;
  reg p2_is_luminance;
  reg [7:0] p2_value;
  reg [1:0] p2_sel_6109;
  reg [3:0] p2_run_u8__1;
  reg p2_and_6016;
  reg p2_eq_6116;
  reg [3:0] p2_and_6120;
  always @ (posedge clk) begin
    p2_start_pix <= p1_start_pix;
    p2_is_luminance <= p1_is_luminance;
    p2_value <= p2_value_comb;
    p2_sel_6109 <= p2_sel_6109_comb;
    p2_run_u8__1 <= p2_run_u8__1_comb;
    p2_and_6016 <= p1_and_6016;
    p2_eq_6116 <= p2_eq_6116_comb;
    p2_and_6120 <= p2_and_6120_comb;
  end

  // ===== Pipe stage 3:
  wire [2:0] p3_idx_u8__4_squeezed__1_comb;
  wire [2:0] p3_idx_u8__5_squeezed__1_comb;
  wire [2:0] p3_idx_u8__6_squeezed__1_comb;
  wire [2:0] p3_idx_u8__7_squeezed__1_comb;
  wire [2:0] p3_sel_6155_comb;
  wire [3:0] p3_idx_u8__8_squeezed_comb;
  wire p3_eq_6160_comb;
  wire [7:0] p3_size__1_comb;
  wire [7:0] p3_idx_u8__48_comb;
  wire [7:0] p3_run_size_str_u8_comb;
  wire [4:0] p3_idx_u8__16_squeezed_comb;
  wire [4:0] p3_huffman_length_squeezed_comb;
  wire [4:0] p3_idx_u8__2_squeezed__1_comb;
  wire [7:0] p3_flipped_comb;
  wire [15:0] p3_huffman_code_full_comb;
  wire [7:0] p3_code_list_comb;
  wire [35:0] p3_tuple_6193_comb;
  assign p3_idx_u8__4_squeezed__1_comb = 3'h4;
  assign p3_idx_u8__5_squeezed__1_comb = 3'h5;
  assign p3_idx_u8__6_squeezed__1_comb = 3'h6;
  assign p3_idx_u8__7_squeezed__1_comb = 3'h7;
  assign p3_sel_6155_comb = |p2_value[7:6] ? p3_idx_u8__7_squeezed__1_comb : (|p2_value[7:5] ? p3_idx_u8__6_squeezed__1_comb : (|p2_value[7:4] ? p3_idx_u8__5_squeezed__1_comb : (|p2_value[7:3] ? p3_idx_u8__4_squeezed__1_comb : {1'h0, p2_sel_6109})));
  assign p3_idx_u8__8_squeezed_comb = 4'h8;
  assign p3_eq_6160_comb = p2_value == 8'h00;
  assign p3_size__1_comb = {4'h0, p2_value[7] ? p3_idx_u8__8_squeezed_comb : {1'h0, p3_sel_6155_comb}} & {8{~p3_eq_6160_comb}};
  assign p3_idx_u8__48_comb = 8'h30;
  assign p3_run_size_str_u8_comb = {p2_run_u8__1, 4'h0} | p3_size__1_comb | p3_idx_u8__48_comb;
  assign p3_idx_u8__16_squeezed_comb = 5'h10;
  assign p3_huffman_length_squeezed_comb = p2_is_luminance ? p3_idx_u8__16_squeezed_comb : literal_6170[p3_run_size_str_u8_comb > 8'ha1 ? 8'ha1 : p3_run_size_str_u8_comb];
  assign p3_idx_u8__2_squeezed__1_comb = 5'h02;
  assign p3_flipped_comb = 8'hff;
  assign p3_huffman_code_full_comb = p2_is_luminance ? AC_LUMINANCE_SIZE_TO_CODE_tuple_idx_0[p3_run_size_str_u8_comb > 8'ha1 ? 8'ha1 : p3_run_size_str_u8_comb] : AC_CHROMINANCE_SIZE_TO_CODE_tuple_idx_0[p3_run_size_str_u8_comb > 8'ha1 ? 8'ha1 : p3_run_size_str_u8_comb];
  assign p3_code_list_comb = p3_eq_6160_comb ? p3_flipped_comb : p2_value;
  assign p3_tuple_6193_comb = {p3_huffman_code_full_comb & {16{~(p2_and_6016 | p2_eq_6116)}}, p2_and_6016 ? p2_start_pix : {3'h0, p2_eq_6116 ? p3_idx_u8__2_squeezed__1_comb : p3_huffman_length_squeezed_comb}, p3_code_list_comb & {8{~(p2_and_6016 | p2_eq_6116)}}, p2_and_6120};

  // Registers for pipe stage 3:
  reg [35:0] p3_tuple_6193;
  always @ (posedge clk) begin
    p3_tuple_6193 <= p3_tuple_6193_comb;
  end
  assign out = p3_tuple_6193;
endmodule
