module dct_1d_s10(
  input wire clk,
  input wire [79:0] x,
  output wire [79:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [15:0] smul16b_8b_x_9b (input reg [7:0] lhs, input reg [8:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [15:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul16b_8b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_8b (input reg [7:0] lhs, input reg [7:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_6b (input reg [7:0] lhs, input reg [5:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [23:0] umul24b_24b_x_7b (input reg [23:0] lhs, input reg [6:0] rhs);
    begin
      umul24b_24b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [9:0] x_unflattened[0:7];
  assign x_unflattened[0] = x[9:0];
  assign x_unflattened[1] = x[19:10];
  assign x_unflattened[2] = x[29:20];
  assign x_unflattened[3] = x[39:30];
  assign x_unflattened[4] = x[49:40];
  assign x_unflattened[5] = x[59:50];
  assign x_unflattened[6] = x[69:60];
  assign x_unflattened[7] = x[79:70];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_x[0:7];
  always @ (posedge clk) begin
    p0_x[0] <= x_unflattened[0];
    p0_x[1] <= x_unflattened[1];
    p0_x[2] <= x_unflattened[2];
    p0_x[3] <= x_unflattened[3];
    p0_x[4] <= x_unflattened[4];
    p0_x[5] <= x_unflattened[5];
    p0_x[6] <= x_unflattened[6];
    p0_x[7] <= x_unflattened[7];
  end

  // ===== Pipe stage 1:
  wire [9:0] p1_array_index_5947_comb;
  wire [9:0] p1_array_index_5948_comb;
  wire [9:0] p1_array_index_5949_comb;
  wire [9:0] p1_array_index_5950_comb;
  wire [9:0] p1_array_index_5951_comb;
  wire [9:0] p1_array_index_5952_comb;
  wire [9:0] p1_array_index_5953_comb;
  wire [9:0] p1_array_index_5954_comb;
  wire [7:0] p1_concat_5979_comb;
  wire [7:0] p1_concat_5981_comb;
  wire [7:0] p1_concat_5983_comb;
  wire [7:0] p1_concat_5985_comb;
  wire [7:0] p1_concat_5988_comb;
  wire [7:0] p1_concat_5990_comb;
  wire [7:0] p1_concat_5994_comb;
  wire [7:0] p1_concat_5996_comb;
  wire [15:0] p1_smul_3316_NarrowedMult__comb;
  wire [15:0] p1_smul_3315_NarrowedMult__comb;
  wire [15:0] p1_smul_3310_NarrowedMult__comb;
  wire [15:0] p1_smul_3309_NarrowedMult__comb;
  wire [15:0] p1_smul_3300_NarrowedMult__comb;
  wire [15:0] p1_smul_3298_NarrowedMult__comb;
  wire [15:0] p1_smul_3295_NarrowedMult__comb;
  wire [15:0] p1_smul_3293_NarrowedMult__comb;
  wire [15:0] p1_smul_3283_NarrowedMult__comb;
  wire [15:0] p1_smul_3281_NarrowedMult__comb;
  wire [15:0] p1_smul_3280_NarrowedMult__comb;
  wire [15:0] p1_smul_3278_NarrowedMult__comb;
  wire [15:0] p1_smul_3266_NarrowedMult__comb;
  wire [15:0] p1_smul_3265_NarrowedMult__comb;
  wire [15:0] p1_smul_3264_NarrowedMult__comb;
  wire [15:0] p1_smul_3263_NarrowedMult__comb;
  wire [14:0] p1_smul_3307_NarrowedMult__comb;
  wire [14:0] p1_smul_3306_NarrowedMult__comb;
  wire [14:0] p1_smul_3303_NarrowedMult__comb;
  wire [14:0] p1_smul_3302_NarrowedMult__comb;
  wire [15:0] p1_smul_3292_NarrowedMult__comb;
  wire [15:0] p1_smul_3291_NarrowedMult__comb;
  wire [15:0] p1_smul_3290_NarrowedMult__comb;
  wire [15:0] p1_smul_3289_NarrowedMult__comb;
  wire [15:0] p1_smul_3288_NarrowedMult__comb;
  wire [15:0] p1_smul_3287_NarrowedMult__comb;
  wire [15:0] p1_smul_3286_NarrowedMult__comb;
  wire [15:0] p1_smul_3285_NarrowedMult__comb;
  wire [14:0] p1_smul_3276_NarrowedMult__comb;
  wire [14:0] p1_smul_3274_NarrowedMult__comb;
  wire [14:0] p1_smul_3271_NarrowedMult__comb;
  wire [14:0] p1_smul_3269_NarrowedMult__comb;
  wire [14:0] p1_smul_3314_NarrowedMult__comb;
  wire [13:0] p1_smul_3330_NarrowedMult__comb;
  wire [13:0] p1_smul_3332_NarrowedMult__comb;
  wire [14:0] p1_smul_3311_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6047_comb;
  wire [13:0] p1_smul_3391_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6049_comb;
  wire [14:0] p1_smul_3297_NarrowedMult__comb;
  wire [14:0] p1_smul_3296_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6052_comb;
  wire [13:0] p1_smul_3411_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6054_comb;
  wire [14:0] p1_smul_3284_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6064_comb;
  wire [13:0] p1_smul_3458_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6066_comb;
  wire [14:0] p1_bit_slice_6067_comb;
  wire [13:0] p1_smul_3468_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6069_comb;
  wire [14:0] p1_smul_3277_NarrowedMult__comb;
  wire [13:0] p1_smul_3519_NarrowedMult__comb;
  wire [14:0] p1_smul_3267_NarrowedMult__comb;
  wire [14:0] p1_smul_3262_NarrowedMult__comb;
  wire [13:0] p1_smul_3547_NarrowedMult__comb;
  wire [13:0] p1_smul_3308_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6140_comb;
  wire [13:0] p1_bit_slice_6141_comb;
  wire [13:0] p1_smul_3305_NarrowedMult__comb;
  wire [13:0] p1_smul_3304_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6144_comb;
  wire [13:0] p1_bit_slice_6145_comb;
  wire [13:0] p1_smul_3301_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6171_comb;
  wire [13:0] p1_smul_3275_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6173_comb;
  wire [13:0] p1_smul_3273_NarrowedMult__comb;
  wire [13:0] p1_smul_3272_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6176_comb;
  wire [13:0] p1_smul_3270_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6178_comb;
  wire [8:0] p1_add_6227_comb;
  wire [8:0] p1_add_6228_comb;
  wire [8:0] p1_add_6229_comb;
  wire [8:0] p1_add_6230_comb;
  wire [16:0] p1_add_6083_comb;
  wire [16:0] p1_add_6088_comb;
  wire [16:0] p1_add_6131_comb;
  wire [16:0] p1_add_6132_comb;
  wire [16:0] p1_add_6207_comb;
  wire [16:0] p1_add_6208_comb;
  wire [16:0] p1_add_6209_comb;
  wire [16:0] p1_add_6210_comb;
  wire [15:0] p1_bit_slice_6135_comb;
  wire [15:0] p1_add_6136_comb;
  wire [15:0] p1_add_6137_comb;
  wire [15:0] p1_bit_slice_6138_comb;
  wire [15:0] p1_add_6147_comb;
  wire [15:0] p1_add_6149_comb;
  wire [15:0] p1_add_6151_comb;
  wire [15:0] p1_add_6153_comb;
  wire [15:0] p1_add_6163_comb;
  wire [15:0] p1_add_6165_comb;
  wire [15:0] p1_add_6167_comb;
  wire [15:0] p1_add_6169_comb;
  wire [15:0] p1_add_6179_comb;
  wire [15:0] p1_bit_slice_6180_comb;
  wire [15:0] p1_bit_slice_6181_comb;
  wire [15:0] p1_add_6182_comb;
  wire [14:0] p1_add_6233_comb;
  wire [14:0] p1_add_6235_comb;
  wire [14:0] p1_add_6237_comb;
  wire [14:0] p1_add_6239_comb;
  wire [24:0] p1_sum__97_comb;
  wire [24:0] p1_sum__98_comb;
  wire [24:0] p1_sum__99_comb;
  wire [24:0] p1_sum__100_comb;
  wire [14:0] p1_add_6245_comb;
  wire [14:0] p1_add_6247_comb;
  wire [14:0] p1_add_6249_comb;
  wire [14:0] p1_add_6251_comb;
  wire [23:0] p1_add_6269_comb;
  wire [23:0] p1_add_6270_comb;
  wire [23:0] p1_sign_ext_6191_comb;
  wire [23:0] p1_sign_ext_6192_comb;
  wire [23:0] p1_sign_ext_6193_comb;
  wire [23:0] p1_sign_ext_6194_comb;
  wire [16:0] p1_concat_6203_comb;
  wire [16:0] p1_concat_6204_comb;
  wire [16:0] p1_concat_6205_comb;
  wire [16:0] p1_concat_6206_comb;
  wire [16:0] p1_concat_6211_comb;
  wire [16:0] p1_concat_6212_comb;
  wire [16:0] p1_concat_6213_comb;
  wire [16:0] p1_concat_6214_comb;
  wire [23:0] p1_sign_ext_6223_comb;
  wire [23:0] p1_sign_ext_6224_comb;
  wire [23:0] p1_sign_ext_6225_comb;
  wire [23:0] p1_sign_ext_6226_comb;
  wire p1_bit_slice_6231_comb;
  wire p1_bit_slice_6232_comb;
  wire p1_bit_slice_6253_comb;
  wire p1_bit_slice_6254_comb;
  wire [15:0] p1_concat_6259_comb;
  wire [15:0] p1_concat_6260_comb;
  wire [15:0] p1_concat_6261_comb;
  wire [15:0] p1_concat_6262_comb;
  wire [24:0] p1_sum__77_comb;
  wire [24:0] p1_sum__78_comb;
  wire [15:0] p1_concat_6265_comb;
  wire [15:0] p1_concat_6266_comb;
  wire [15:0] p1_concat_6267_comb;
  wire [15:0] p1_concat_6268_comb;
  wire [23:0] p1_add_6271_comb;
  assign p1_array_index_5947_comb = p0_x[3'h0];
  assign p1_array_index_5948_comb = p0_x[3'h1];
  assign p1_array_index_5949_comb = p0_x[3'h6];
  assign p1_array_index_5950_comb = p0_x[3'h7];
  assign p1_array_index_5951_comb = p0_x[3'h2];
  assign p1_array_index_5952_comb = p0_x[3'h5];
  assign p1_array_index_5953_comb = p0_x[3'h3];
  assign p1_array_index_5954_comb = p0_x[3'h4];
  assign p1_concat_5979_comb = {~p1_array_index_5947_comb[7], p1_array_index_5947_comb[6:0]};
  assign p1_concat_5981_comb = {~p1_array_index_5948_comb[7], p1_array_index_5948_comb[6:0]};
  assign p1_concat_5983_comb = {~p1_array_index_5949_comb[7], p1_array_index_5949_comb[6:0]};
  assign p1_concat_5985_comb = {~p1_array_index_5950_comb[7], p1_array_index_5950_comb[6:0]};
  assign p1_concat_5988_comb = {~p1_array_index_5951_comb[7], p1_array_index_5951_comb[6:0]};
  assign p1_concat_5990_comb = {~p1_array_index_5952_comb[7], p1_array_index_5952_comb[6:0]};
  assign p1_concat_5994_comb = {~p1_array_index_5953_comb[7], p1_array_index_5953_comb[6:0]};
  assign p1_concat_5996_comb = {~p1_array_index_5954_comb[7], p1_array_index_5954_comb[6:0]};
  assign p1_smul_3316_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5979_comb, 9'h0fb);
  assign p1_smul_3315_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5981_comb, 9'h0d5);
  assign p1_smul_3310_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5983_comb, 9'h12b);
  assign p1_smul_3309_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5985_comb, 9'h105);
  assign p1_smul_3300_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5979_comb, 9'h0d5);
  assign p1_smul_3298_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5988_comb, 9'h105);
  assign p1_smul_3295_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5990_comb, 9'h0fb);
  assign p1_smul_3293_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5985_comb, 9'h12b);
  assign p1_smul_3283_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5981_comb, 9'h105);
  assign p1_smul_3281_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5994_comb, 9'h0d5);
  assign p1_smul_3280_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5996_comb, 9'h0d5);
  assign p1_smul_3278_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5983_comb, 9'h105);
  assign p1_smul_3266_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5988_comb, 9'h0d5);
  assign p1_smul_3265_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5994_comb, 9'h105);
  assign p1_smul_3264_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5996_comb, 9'h105);
  assign p1_smul_3263_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5990_comb, 9'h0d5);
  assign p1_smul_3307_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5981_comb, 7'h31);
  assign p1_smul_3306_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5988_comb, 7'h4f);
  assign p1_smul_3303_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5990_comb, 7'h4f);
  assign p1_smul_3302_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5983_comb, 7'h31);
  assign p1_smul_3292_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5979_comb, 9'h0b5);
  assign p1_smul_3291_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5981_comb, 9'h14b);
  assign p1_smul_3290_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5988_comb, 9'h14b);
  assign p1_smul_3289_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5994_comb, 9'h0b5);
  assign p1_smul_3288_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5996_comb, 9'h0b5);
  assign p1_smul_3287_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5990_comb, 9'h14b);
  assign p1_smul_3286_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5983_comb, 9'h14b);
  assign p1_smul_3285_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5985_comb, 9'h0b5);
  assign p1_smul_3276_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5979_comb, 7'h31);
  assign p1_smul_3274_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5988_comb, 7'h31);
  assign p1_smul_3271_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5990_comb, 7'h31);
  assign p1_smul_3269_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5985_comb, 7'h31);
  assign p1_smul_3314_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5988_comb, 8'h47);
  assign p1_smul_3330_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5994_comb, 6'h19);
  assign p1_smul_3332_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5996_comb, 6'h27);
  assign p1_smul_3311_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5990_comb, 8'hb9);
  assign p1_bit_slice_6047_comb = p1_smul_3300_NarrowedMult__comb[15:1];
  assign p1_smul_3391_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5981_comb, 6'h27);
  assign p1_bit_slice_6049_comb = p1_smul_3298_NarrowedMult__comb[15:1];
  assign p1_smul_3297_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5994_comb, 8'hb9);
  assign p1_smul_3296_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5996_comb, 8'h47);
  assign p1_bit_slice_6052_comb = p1_smul_3295_NarrowedMult__comb[15:1];
  assign p1_smul_3411_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5983_comb, 6'h19);
  assign p1_bit_slice_6054_comb = p1_smul_3293_NarrowedMult__comb[15:1];
  assign p1_smul_3284_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5979_comb, 8'h47);
  assign p1_bit_slice_6064_comb = p1_smul_3283_NarrowedMult__comb[15:1];
  assign p1_smul_3458_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5988_comb, 6'h27);
  assign p1_bit_slice_6066_comb = p1_smul_3281_NarrowedMult__comb[15:1];
  assign p1_bit_slice_6067_comb = p1_smul_3280_NarrowedMult__comb[15:1];
  assign p1_smul_3468_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5990_comb, 6'h27);
  assign p1_bit_slice_6069_comb = p1_smul_3278_NarrowedMult__comb[15:1];
  assign p1_smul_3277_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5985_comb, 8'h47);
  assign p1_smul_3519_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5979_comb, 6'h19);
  assign p1_smul_3267_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5981_comb, 8'hb9);
  assign p1_smul_3262_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5983_comb, 8'hb9);
  assign p1_smul_3547_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5985_comb, 6'h19);
  assign p1_smul_3308_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5979_comb, 7'h3b);
  assign p1_bit_slice_6140_comb = p1_smul_3307_NarrowedMult__comb[14:1];
  assign p1_bit_slice_6141_comb = p1_smul_3306_NarrowedMult__comb[14:1];
  assign p1_smul_3305_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5994_comb, 7'h45);
  assign p1_smul_3304_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5996_comb, 7'h45);
  assign p1_bit_slice_6144_comb = p1_smul_3303_NarrowedMult__comb[14:1];
  assign p1_bit_slice_6145_comb = p1_smul_3302_NarrowedMult__comb[14:1];
  assign p1_smul_3301_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5985_comb, 7'h3b);
  assign p1_bit_slice_6171_comb = p1_smul_3276_NarrowedMult__comb[14:1];
  assign p1_smul_3275_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5981_comb, 7'h45);
  assign p1_bit_slice_6173_comb = p1_smul_3274_NarrowedMult__comb[14:1];
  assign p1_smul_3273_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5994_comb, 7'h3b);
  assign p1_smul_3272_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5996_comb, 7'h3b);
  assign p1_bit_slice_6176_comb = p1_smul_3271_NarrowedMult__comb[14:1];
  assign p1_smul_3270_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5983_comb, 7'h45);
  assign p1_bit_slice_6178_comb = p1_smul_3269_NarrowedMult__comb[14:1];
  assign p1_add_6227_comb = {{1{p1_concat_5979_comb[7]}}, p1_concat_5979_comb} + {{1{p1_concat_5981_comb[7]}}, p1_concat_5981_comb};
  assign p1_add_6228_comb = {{1{p1_concat_5988_comb[7]}}, p1_concat_5988_comb} + {{1{p1_concat_5994_comb[7]}}, p1_concat_5994_comb};
  assign p1_add_6229_comb = {{1{p1_concat_5996_comb[7]}}, p1_concat_5996_comb} + {{1{p1_concat_5990_comb[7]}}, p1_concat_5990_comb};
  assign p1_add_6230_comb = {{1{p1_concat_5983_comb[7]}}, p1_concat_5983_comb} + {{1{p1_concat_5985_comb[7]}}, p1_concat_5985_comb};
  assign p1_add_6083_comb = {{1{p1_smul_3316_NarrowedMult__comb[15]}}, p1_smul_3316_NarrowedMult__comb} + {{1{p1_smul_3315_NarrowedMult__comb[15]}}, p1_smul_3315_NarrowedMult__comb};
  assign p1_add_6088_comb = {{1{p1_smul_3310_NarrowedMult__comb[15]}}, p1_smul_3310_NarrowedMult__comb} + {{1{p1_smul_3309_NarrowedMult__comb[15]}}, p1_smul_3309_NarrowedMult__comb};
  assign p1_add_6131_comb = {{1{p1_smul_3266_NarrowedMult__comb[15]}}, p1_smul_3266_NarrowedMult__comb} + {{1{p1_smul_3265_NarrowedMult__comb[15]}}, p1_smul_3265_NarrowedMult__comb};
  assign p1_add_6132_comb = {{1{p1_smul_3264_NarrowedMult__comb[15]}}, p1_smul_3264_NarrowedMult__comb} + {{1{p1_smul_3263_NarrowedMult__comb[15]}}, p1_smul_3263_NarrowedMult__comb};
  assign p1_add_6207_comb = {{1{p1_smul_3292_NarrowedMult__comb[15]}}, p1_smul_3292_NarrowedMult__comb} + {{1{p1_smul_3291_NarrowedMult__comb[15]}}, p1_smul_3291_NarrowedMult__comb};
  assign p1_add_6208_comb = {{1{p1_smul_3290_NarrowedMult__comb[15]}}, p1_smul_3290_NarrowedMult__comb} + {{1{p1_smul_3289_NarrowedMult__comb[15]}}, p1_smul_3289_NarrowedMult__comb};
  assign p1_add_6209_comb = {{1{p1_smul_3288_NarrowedMult__comb[15]}}, p1_smul_3288_NarrowedMult__comb} + {{1{p1_smul_3287_NarrowedMult__comb[15]}}, p1_smul_3287_NarrowedMult__comb};
  assign p1_add_6210_comb = {{1{p1_smul_3286_NarrowedMult__comb[15]}}, p1_smul_3286_NarrowedMult__comb} + {{1{p1_smul_3285_NarrowedMult__comb[15]}}, p1_smul_3285_NarrowedMult__comb};
  assign p1_bit_slice_6135_comb = p1_add_6083_comb[16:1];
  assign p1_add_6136_comb = {{1{p1_smul_3314_NarrowedMult__comb[14]}}, p1_smul_3314_NarrowedMult__comb} + {{2{p1_smul_3330_NarrowedMult__comb[13]}}, p1_smul_3330_NarrowedMult__comb};
  assign p1_add_6137_comb = {{2{p1_smul_3332_NarrowedMult__comb[13]}}, p1_smul_3332_NarrowedMult__comb} + {{1{p1_smul_3311_NarrowedMult__comb[14]}}, p1_smul_3311_NarrowedMult__comb};
  assign p1_bit_slice_6138_comb = p1_add_6088_comb[16:1];
  assign p1_add_6147_comb = {{1{p1_bit_slice_6047_comb[14]}}, p1_bit_slice_6047_comb} + {{2{p1_smul_3391_NarrowedMult__comb[13]}}, p1_smul_3391_NarrowedMult__comb};
  assign p1_add_6149_comb = {{1{p1_bit_slice_6049_comb[14]}}, p1_bit_slice_6049_comb} + {{1{p1_smul_3297_NarrowedMult__comb[14]}}, p1_smul_3297_NarrowedMult__comb};
  assign p1_add_6151_comb = {{1{p1_smul_3296_NarrowedMult__comb[14]}}, p1_smul_3296_NarrowedMult__comb} + {{1{p1_bit_slice_6052_comb[14]}}, p1_bit_slice_6052_comb};
  assign p1_add_6153_comb = {{2{p1_smul_3411_NarrowedMult__comb[13]}}, p1_smul_3411_NarrowedMult__comb} + {{1{p1_bit_slice_6054_comb[14]}}, p1_bit_slice_6054_comb};
  assign p1_add_6163_comb = {{1{p1_smul_3284_NarrowedMult__comb[14]}}, p1_smul_3284_NarrowedMult__comb} + {{1{p1_bit_slice_6064_comb[14]}}, p1_bit_slice_6064_comb};
  assign p1_add_6165_comb = {{2{p1_smul_3458_NarrowedMult__comb[13]}}, p1_smul_3458_NarrowedMult__comb} + {{1{p1_bit_slice_6066_comb[14]}}, p1_bit_slice_6066_comb};
  assign p1_add_6167_comb = {{1{p1_bit_slice_6067_comb[14]}}, p1_bit_slice_6067_comb} + {{2{p1_smul_3468_NarrowedMult__comb[13]}}, p1_smul_3468_NarrowedMult__comb};
  assign p1_add_6169_comb = {{1{p1_bit_slice_6069_comb[14]}}, p1_bit_slice_6069_comb} + {{1{p1_smul_3277_NarrowedMult__comb[14]}}, p1_smul_3277_NarrowedMult__comb};
  assign p1_add_6179_comb = {{2{p1_smul_3519_NarrowedMult__comb[13]}}, p1_smul_3519_NarrowedMult__comb} + {{1{p1_smul_3267_NarrowedMult__comb[14]}}, p1_smul_3267_NarrowedMult__comb};
  assign p1_bit_slice_6180_comb = p1_add_6131_comb[16:1];
  assign p1_bit_slice_6181_comb = p1_add_6132_comb[16:1];
  assign p1_add_6182_comb = {{1{p1_smul_3262_NarrowedMult__comb[14]}}, p1_smul_3262_NarrowedMult__comb} + {{2{p1_smul_3547_NarrowedMult__comb[13]}}, p1_smul_3547_NarrowedMult__comb};
  assign p1_add_6233_comb = {{1{p1_smul_3308_NarrowedMult__comb[13]}}, p1_smul_3308_NarrowedMult__comb} + {{1{p1_bit_slice_6140_comb[13]}}, p1_bit_slice_6140_comb};
  assign p1_add_6235_comb = {{1{p1_bit_slice_6141_comb[13]}}, p1_bit_slice_6141_comb} + {{1{p1_smul_3305_NarrowedMult__comb[13]}}, p1_smul_3305_NarrowedMult__comb};
  assign p1_add_6237_comb = {{1{p1_smul_3304_NarrowedMult__comb[13]}}, p1_smul_3304_NarrowedMult__comb} + {{1{p1_bit_slice_6144_comb[13]}}, p1_bit_slice_6144_comb};
  assign p1_add_6239_comb = {{1{p1_bit_slice_6145_comb[13]}}, p1_bit_slice_6145_comb} + {{1{p1_smul_3301_NarrowedMult__comb[13]}}, p1_smul_3301_NarrowedMult__comb};
  assign p1_sum__97_comb = {{8{p1_add_6207_comb[16]}}, p1_add_6207_comb};
  assign p1_sum__98_comb = {{8{p1_add_6208_comb[16]}}, p1_add_6208_comb};
  assign p1_sum__99_comb = {{8{p1_add_6209_comb[16]}}, p1_add_6209_comb};
  assign p1_sum__100_comb = {{8{p1_add_6210_comb[16]}}, p1_add_6210_comb};
  assign p1_add_6245_comb = {{1{p1_bit_slice_6171_comb[13]}}, p1_bit_slice_6171_comb} + {{1{p1_smul_3275_NarrowedMult__comb[13]}}, p1_smul_3275_NarrowedMult__comb};
  assign p1_add_6247_comb = {{1{p1_bit_slice_6173_comb[13]}}, p1_bit_slice_6173_comb} + {{1{p1_smul_3273_NarrowedMult__comb[13]}}, p1_smul_3273_NarrowedMult__comb};
  assign p1_add_6249_comb = {{1{p1_smul_3272_NarrowedMult__comb[13]}}, p1_smul_3272_NarrowedMult__comb} + {{1{p1_bit_slice_6176_comb[13]}}, p1_bit_slice_6176_comb};
  assign p1_add_6251_comb = {{1{p1_smul_3270_NarrowedMult__comb[13]}}, p1_smul_3270_NarrowedMult__comb} + {{1{p1_bit_slice_6178_comb[13]}}, p1_bit_slice_6178_comb};
  assign p1_add_6269_comb = {{15{p1_add_6227_comb[8]}}, p1_add_6227_comb} + {{15{p1_add_6228_comb[8]}}, p1_add_6228_comb};
  assign p1_add_6270_comb = {{15{p1_add_6229_comb[8]}}, p1_add_6229_comb} + {{15{p1_add_6230_comb[8]}}, p1_add_6230_comb};
  assign p1_sign_ext_6191_comb = {{8{p1_bit_slice_6135_comb[15]}}, p1_bit_slice_6135_comb};
  assign p1_sign_ext_6192_comb = {{8{p1_add_6136_comb[15]}}, p1_add_6136_comb};
  assign p1_sign_ext_6193_comb = {{8{p1_add_6137_comb[15]}}, p1_add_6137_comb};
  assign p1_sign_ext_6194_comb = {{8{p1_bit_slice_6138_comb[15]}}, p1_bit_slice_6138_comb};
  assign p1_concat_6203_comb = {p1_add_6147_comb, p1_smul_3300_NarrowedMult__comb[0]};
  assign p1_concat_6204_comb = {p1_add_6149_comb, p1_smul_3298_NarrowedMult__comb[0]};
  assign p1_concat_6205_comb = {p1_add_6151_comb, p1_smul_3295_NarrowedMult__comb[0]};
  assign p1_concat_6206_comb = {p1_add_6153_comb, p1_smul_3293_NarrowedMult__comb[0]};
  assign p1_concat_6211_comb = {p1_add_6163_comb, p1_smul_3283_NarrowedMult__comb[0]};
  assign p1_concat_6212_comb = {p1_add_6165_comb, p1_smul_3281_NarrowedMult__comb[0]};
  assign p1_concat_6213_comb = {p1_add_6167_comb, p1_smul_3280_NarrowedMult__comb[0]};
  assign p1_concat_6214_comb = {p1_add_6169_comb, p1_smul_3278_NarrowedMult__comb[0]};
  assign p1_sign_ext_6223_comb = {{8{p1_add_6179_comb[15]}}, p1_add_6179_comb};
  assign p1_sign_ext_6224_comb = {{8{p1_bit_slice_6180_comb[15]}}, p1_bit_slice_6180_comb};
  assign p1_sign_ext_6225_comb = {{8{p1_bit_slice_6181_comb[15]}}, p1_bit_slice_6181_comb};
  assign p1_sign_ext_6226_comb = {{8{p1_add_6182_comb[15]}}, p1_add_6182_comb};
  assign p1_bit_slice_6231_comb = p1_add_6083_comb[0];
  assign p1_bit_slice_6232_comb = p1_add_6088_comb[0];
  assign p1_bit_slice_6253_comb = p1_add_6131_comb[0];
  assign p1_bit_slice_6254_comb = p1_add_6132_comb[0];
  assign p1_concat_6259_comb = {p1_add_6233_comb, p1_smul_3307_NarrowedMult__comb[0]};
  assign p1_concat_6260_comb = {p1_add_6235_comb, p1_smul_3306_NarrowedMult__comb[0]};
  assign p1_concat_6261_comb = {p1_add_6237_comb, p1_smul_3303_NarrowedMult__comb[0]};
  assign p1_concat_6262_comb = {p1_add_6239_comb, p1_smul_3302_NarrowedMult__comb[0]};
  assign p1_sum__77_comb = p1_sum__97_comb + p1_sum__98_comb;
  assign p1_sum__78_comb = p1_sum__99_comb + p1_sum__100_comb;
  assign p1_concat_6265_comb = {p1_add_6245_comb, p1_smul_3276_NarrowedMult__comb[0]};
  assign p1_concat_6266_comb = {p1_add_6247_comb, p1_smul_3274_NarrowedMult__comb[0]};
  assign p1_concat_6267_comb = {p1_add_6249_comb, p1_smul_3271_NarrowedMult__comb[0]};
  assign p1_concat_6268_comb = {p1_add_6251_comb, p1_smul_3269_NarrowedMult__comb[0]};
  assign p1_add_6271_comb = p1_add_6269_comb + p1_add_6270_comb;

  // Registers for pipe stage 1:
  reg [23:0] p1_sign_ext_6191;
  reg [23:0] p1_sign_ext_6192;
  reg [23:0] p1_sign_ext_6193;
  reg [23:0] p1_sign_ext_6194;
  reg [16:0] p1_concat_6203;
  reg [16:0] p1_concat_6204;
  reg [16:0] p1_concat_6205;
  reg [16:0] p1_concat_6206;
  reg [16:0] p1_concat_6211;
  reg [16:0] p1_concat_6212;
  reg [16:0] p1_concat_6213;
  reg [16:0] p1_concat_6214;
  reg [23:0] p1_sign_ext_6223;
  reg [23:0] p1_sign_ext_6224;
  reg [23:0] p1_sign_ext_6225;
  reg [23:0] p1_sign_ext_6226;
  reg p1_bit_slice_6231;
  reg p1_bit_slice_6232;
  reg p1_bit_slice_6253;
  reg p1_bit_slice_6254;
  reg [15:0] p1_concat_6259;
  reg [15:0] p1_concat_6260;
  reg [15:0] p1_concat_6261;
  reg [15:0] p1_concat_6262;
  reg [24:0] p1_sum__77;
  reg [24:0] p1_sum__78;
  reg [15:0] p1_concat_6265;
  reg [15:0] p1_concat_6266;
  reg [15:0] p1_concat_6267;
  reg [15:0] p1_concat_6268;
  reg [23:0] p1_add_6271;
  always @ (posedge clk) begin
    p1_sign_ext_6191 <= p1_sign_ext_6191_comb;
    p1_sign_ext_6192 <= p1_sign_ext_6192_comb;
    p1_sign_ext_6193 <= p1_sign_ext_6193_comb;
    p1_sign_ext_6194 <= p1_sign_ext_6194_comb;
    p1_concat_6203 <= p1_concat_6203_comb;
    p1_concat_6204 <= p1_concat_6204_comb;
    p1_concat_6205 <= p1_concat_6205_comb;
    p1_concat_6206 <= p1_concat_6206_comb;
    p1_concat_6211 <= p1_concat_6211_comb;
    p1_concat_6212 <= p1_concat_6212_comb;
    p1_concat_6213 <= p1_concat_6213_comb;
    p1_concat_6214 <= p1_concat_6214_comb;
    p1_sign_ext_6223 <= p1_sign_ext_6223_comb;
    p1_sign_ext_6224 <= p1_sign_ext_6224_comb;
    p1_sign_ext_6225 <= p1_sign_ext_6225_comb;
    p1_sign_ext_6226 <= p1_sign_ext_6226_comb;
    p1_bit_slice_6231 <= p1_bit_slice_6231_comb;
    p1_bit_slice_6232 <= p1_bit_slice_6232_comb;
    p1_bit_slice_6253 <= p1_bit_slice_6253_comb;
    p1_bit_slice_6254 <= p1_bit_slice_6254_comb;
    p1_concat_6259 <= p1_concat_6259_comb;
    p1_concat_6260 <= p1_concat_6260_comb;
    p1_concat_6261 <= p1_concat_6261_comb;
    p1_concat_6262 <= p1_concat_6262_comb;
    p1_sum__77 <= p1_sum__77_comb;
    p1_sum__78 <= p1_sum__78_comb;
    p1_concat_6265 <= p1_concat_6265_comb;
    p1_concat_6266 <= p1_concat_6266_comb;
    p1_concat_6267 <= p1_concat_6267_comb;
    p1_concat_6268 <= p1_concat_6268_comb;
    p1_add_6271 <= p1_add_6271_comb;
  end

  // ===== Pipe stage 2:
  wire [23:0] p2_add_6334_comb;
  wire [23:0] p2_add_6335_comb;
  wire [24:0] p2_sum__101_comb;
  wire [24:0] p2_sum__102_comb;
  wire [24:0] p2_sum__103_comb;
  wire [24:0] p2_sum__104_comb;
  wire [24:0] p2_sum__93_comb;
  wire [24:0] p2_sum__94_comb;
  wire [24:0] p2_sum__95_comb;
  wire [24:0] p2_sum__96_comb;
  wire [23:0] p2_add_6344_comb;
  wire [23:0] p2_add_6345_comb;
  wire [24:0] p2_sum__67_comb;
  wire [24:0] p2_sum__83_comb;
  wire [24:0] p2_sum__84_comb;
  wire [24:0] p2_sum__79_comb;
  wire [24:0] p2_sum__80_comb;
  wire [24:0] p2_sum__75_comb;
  wire [24:0] p2_sum__76_comb;
  wire [24:0] p2_sum__71_comb;
  wire [24:0] p2_sum__72_comb;
  wire [23:0] p2_add_6374_comb;
  wire [23:0] p2_add_6375_comb;
  wire [24:0] p2_add_6377_comb;
  wire [23:0] p2_add_6379_comb;
  wire [23:0] p2_add_6380_comb;
  wire [24:0] p2_sum__70_comb;
  wire [24:0] p2_sum__68_comb;
  wire [24:0] p2_sum__66_comb;
  wire [24:0] p2_sum__64_comb;
  wire [23:0] p2_umul_2805_NarrowedMult__comb;
  wire [23:0] p2_add_6386_comb;
  wire [23:0] p2_add_6394_comb;
  wire [24:0] p2_add_6373_comb;
  wire [24:0] p2_add_6376_comb;
  wire [24:0] p2_add_6378_comb;
  wire [24:0] p2_add_6381_comb;
  wire [8:0] p2_clipped__16_comb;
  wire [8:0] p2_clipped__18_comb;
  wire [8:0] p2_clipped__20_comb;
  wire [8:0] p2_clipped__22_comb;
  wire [8:0] p2_clipped__17_comb;
  wire [8:0] p2_clipped__19_comb;
  wire [8:0] p2_clipped__21_comb;
  wire [8:0] p2_clipped__23_comb;
  wire [9:0] p2_add_6474_comb;
  wire [9:0] p2_add_6475_comb;
  wire [9:0] p2_add_6476_comb;
  wire [9:0] p2_add_6477_comb;
  wire [9:0] p2_sign_ext_6464_comb;
  wire [9:0] p2_sign_ext_6467_comb;
  wire [9:0] p2_sign_ext_6470_comb;
  wire [9:0] p2_sign_ext_6473_comb;
  wire [1:0] p2_bit_slice_6478_comb;
  wire [1:0] p2_bit_slice_6479_comb;
  wire [1:0] p2_bit_slice_6480_comb;
  wire [1:0] p2_bit_slice_6481_comb;
  wire [6:0] p2_bit_slice_6482_comb;
  wire [6:0] p2_bit_slice_6483_comb;
  wire [6:0] p2_bit_slice_6484_comb;
  wire [6:0] p2_bit_slice_6485_comb;
  assign p2_add_6334_comb = p1_sign_ext_6191 + p1_sign_ext_6192;
  assign p2_add_6335_comb = p1_sign_ext_6193 + p1_sign_ext_6194;
  assign p2_sum__101_comb = {{8{p1_concat_6203[16]}}, p1_concat_6203};
  assign p2_sum__102_comb = {{8{p1_concat_6204[16]}}, p1_concat_6204};
  assign p2_sum__103_comb = {{8{p1_concat_6205[16]}}, p1_concat_6205};
  assign p2_sum__104_comb = {{8{p1_concat_6206[16]}}, p1_concat_6206};
  assign p2_sum__93_comb = {{8{p1_concat_6211[16]}}, p1_concat_6211};
  assign p2_sum__94_comb = {{8{p1_concat_6212[16]}}, p1_concat_6212};
  assign p2_sum__95_comb = {{8{p1_concat_6213[16]}}, p1_concat_6213};
  assign p2_sum__96_comb = {{8{p1_concat_6214[16]}}, p1_concat_6214};
  assign p2_add_6344_comb = p1_sign_ext_6223 + p1_sign_ext_6224;
  assign p2_add_6345_comb = p1_sign_ext_6225 + p1_sign_ext_6226;
  assign p2_sum__67_comb = p1_sum__77 + p1_sum__78;
  assign p2_sum__83_comb = {p2_add_6334_comb, p1_bit_slice_6231};
  assign p2_sum__84_comb = {p2_add_6335_comb, p1_bit_slice_6232};
  assign p2_sum__79_comb = p2_sum__101_comb + p2_sum__102_comb;
  assign p2_sum__80_comb = p2_sum__103_comb + p2_sum__104_comb;
  assign p2_sum__75_comb = p2_sum__93_comb + p2_sum__94_comb;
  assign p2_sum__76_comb = p2_sum__95_comb + p2_sum__96_comb;
  assign p2_sum__71_comb = {p2_add_6344_comb, p1_bit_slice_6253};
  assign p2_sum__72_comb = {p2_add_6345_comb, p1_bit_slice_6254};
  assign p2_add_6374_comb = {{8{p1_concat_6259[15]}}, p1_concat_6259} + {{8{p1_concat_6260[15]}}, p1_concat_6260};
  assign p2_add_6375_comb = {{8{p1_concat_6261[15]}}, p1_concat_6261} + {{8{p1_concat_6262[15]}}, p1_concat_6262};
  assign p2_add_6377_comb = p2_sum__67_comb + 25'h000_0001;
  assign p2_add_6379_comb = {{8{p1_concat_6265[15]}}, p1_concat_6265} + {{8{p1_concat_6266[15]}}, p1_concat_6266};
  assign p2_add_6380_comb = {{8{p1_concat_6267[15]}}, p1_concat_6267} + {{8{p1_concat_6268[15]}}, p1_concat_6268};
  assign p2_sum__70_comb = p2_sum__83_comb + p2_sum__84_comb;
  assign p2_sum__68_comb = p2_sum__79_comb + p2_sum__80_comb;
  assign p2_sum__66_comb = p2_sum__75_comb + p2_sum__76_comb;
  assign p2_sum__64_comb = p2_sum__71_comb + p2_sum__72_comb;
  assign p2_umul_2805_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_6271, 7'h5b);
  assign p2_add_6386_comb = p2_add_6374_comb + p2_add_6375_comb;
  assign p2_add_6394_comb = p2_add_6379_comb + p2_add_6380_comb;
  assign p2_add_6373_comb = p2_sum__70_comb + 25'h000_0001;
  assign p2_add_6376_comb = p2_sum__68_comb + 25'h000_0001;
  assign p2_add_6378_comb = p2_sum__66_comb + 25'h000_0001;
  assign p2_add_6381_comb = p2_sum__64_comb + 25'h000_0001;
  assign p2_clipped__16_comb = $signed(p2_umul_2805_NarrowedMult__comb) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_umul_2805_NarrowedMult__comb) > $signed(24'h00_7fff) ? 9'h0ff : p2_umul_2805_NarrowedMult__comb[15:7]);
  assign p2_clipped__18_comb = $signed(p2_add_6386_comb) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6386_comb) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6386_comb[15:7]);
  assign p2_clipped__20_comb = $signed(p2_add_6377_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6377_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6377_comb[16:8]);
  assign p2_clipped__22_comb = $signed(p2_add_6394_comb) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6394_comb) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6394_comb[15:7]);
  assign p2_clipped__17_comb = $signed(p2_add_6373_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6373_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6373_comb[16:8]);
  assign p2_clipped__19_comb = $signed(p2_add_6376_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6376_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6376_comb[16:8]);
  assign p2_clipped__21_comb = $signed(p2_add_6378_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6378_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6378_comb[16:8]);
  assign p2_clipped__23_comb = $signed(p2_add_6381_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6381_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6381_comb[16:8]);
  assign p2_add_6474_comb = {{1{p2_clipped__16_comb[8]}}, p2_clipped__16_comb} + 10'h001;
  assign p2_add_6475_comb = {{1{p2_clipped__18_comb[8]}}, p2_clipped__18_comb} + 10'h001;
  assign p2_add_6476_comb = {{1{p2_clipped__20_comb[8]}}, p2_clipped__20_comb} + 10'h001;
  assign p2_add_6477_comb = {{1{p2_clipped__22_comb[8]}}, p2_clipped__22_comb} + 10'h001;
  assign p2_sign_ext_6464_comb = {{1{p2_clipped__17_comb[8]}}, p2_clipped__17_comb};
  assign p2_sign_ext_6467_comb = {{1{p2_clipped__19_comb[8]}}, p2_clipped__19_comb};
  assign p2_sign_ext_6470_comb = {{1{p2_clipped__21_comb[8]}}, p2_clipped__21_comb};
  assign p2_sign_ext_6473_comb = {{1{p2_clipped__23_comb[8]}}, p2_clipped__23_comb};
  assign p2_bit_slice_6478_comb = p2_add_6474_comb[9:8];
  assign p2_bit_slice_6479_comb = p2_add_6475_comb[9:8];
  assign p2_bit_slice_6480_comb = p2_add_6476_comb[9:8];
  assign p2_bit_slice_6481_comb = p2_add_6477_comb[9:8];
  assign p2_bit_slice_6482_comb = p2_add_6474_comb[7:1];
  assign p2_bit_slice_6483_comb = p2_add_6475_comb[7:1];
  assign p2_bit_slice_6484_comb = p2_add_6476_comb[7:1];
  assign p2_bit_slice_6485_comb = p2_add_6477_comb[7:1];

  // Registers for pipe stage 2:
  reg [9:0] p2_sign_ext_6464;
  reg [9:0] p2_sign_ext_6467;
  reg [9:0] p2_sign_ext_6470;
  reg [9:0] p2_sign_ext_6473;
  reg [1:0] p2_bit_slice_6478;
  reg [1:0] p2_bit_slice_6479;
  reg [1:0] p2_bit_slice_6480;
  reg [1:0] p2_bit_slice_6481;
  reg [6:0] p2_bit_slice_6482;
  reg [6:0] p2_bit_slice_6483;
  reg [6:0] p2_bit_slice_6484;
  reg [6:0] p2_bit_slice_6485;
  always @ (posedge clk) begin
    p2_sign_ext_6464 <= p2_sign_ext_6464_comb;
    p2_sign_ext_6467 <= p2_sign_ext_6467_comb;
    p2_sign_ext_6470 <= p2_sign_ext_6470_comb;
    p2_sign_ext_6473 <= p2_sign_ext_6473_comb;
    p2_bit_slice_6478 <= p2_bit_slice_6478_comb;
    p2_bit_slice_6479 <= p2_bit_slice_6479_comb;
    p2_bit_slice_6480 <= p2_bit_slice_6480_comb;
    p2_bit_slice_6481 <= p2_bit_slice_6481_comb;
    p2_bit_slice_6482 <= p2_bit_slice_6482_comb;
    p2_bit_slice_6483 <= p2_bit_slice_6483_comb;
    p2_bit_slice_6484 <= p2_bit_slice_6484_comb;
    p2_bit_slice_6485 <= p2_bit_slice_6485_comb;
  end

  // ===== Pipe stage 3:
  wire [9:0] p3_add_6514_comb;
  wire [9:0] p3_add_6515_comb;
  wire [9:0] p3_add_6516_comb;
  wire [9:0] p3_add_6517_comb;
  wire [1:0] p3_bit_slice_6518_comb;
  wire [1:0] p3_bit_slice_6519_comb;
  wire [1:0] p3_bit_slice_6520_comb;
  wire [1:0] p3_bit_slice_6521_comb;
  wire [2:0] p3_add_6538_comb;
  wire [2:0] p3_add_6539_comb;
  wire [2:0] p3_add_6540_comb;
  wire [2:0] p3_add_6541_comb;
  wire [2:0] p3_add_6542_comb;
  wire [2:0] p3_add_6543_comb;
  wire [2:0] p3_add_6544_comb;
  wire [2:0] p3_add_6545_comb;
  wire p3_clipped__8_squeezed_const_msb_bits_comb;
  wire [8:0] p3_clipped__8_squeezed_comb;
  wire p3_clipped__8_squeezed_const_msb_bits__1_comb;
  wire [8:0] p3_clipped__9_squeezed_comb;
  wire p3_clipped__8_squeezed_const_msb_bits__2_comb;
  wire [8:0] p3_clipped__10_squeezed_comb;
  wire p3_clipped__8_squeezed_const_msb_bits__3_comb;
  wire [8:0] p3_clipped__11_squeezed_comb;
  wire p3_clipped__8_squeezed_const_msb_bits__4_comb;
  wire [8:0] p3_clipped__12_squeezed_comb;
  wire p3_clipped__8_squeezed_const_msb_bits__5_comb;
  wire [8:0] p3_clipped__13_squeezed_comb;
  wire p3_clipped__8_squeezed_const_msb_bits__6_comb;
  wire [8:0] p3_clipped__14_squeezed_comb;
  wire p3_clipped__8_squeezed_const_msb_bits__7_comb;
  wire [8:0] p3_clipped__15_squeezed_comb;
  wire [9:0] p3_clipped__8_comb;
  wire [9:0] p3_clipped__9_comb;
  wire [9:0] p3_clipped__10_comb;
  wire [9:0] p3_clipped__11_comb;
  wire [9:0] p3_clipped__12_comb;
  wire [9:0] p3_clipped__13_comb;
  wire [9:0] p3_clipped__14_comb;
  wire [9:0] p3_clipped__15_comb;
  wire [9:0] p3_result_comb[0:7];
  assign p3_add_6514_comb = p2_sign_ext_6464 + 10'h001;
  assign p3_add_6515_comb = p2_sign_ext_6467 + 10'h001;
  assign p3_add_6516_comb = p2_sign_ext_6470 + 10'h001;
  assign p3_add_6517_comb = p2_sign_ext_6473 + 10'h001;
  assign p3_bit_slice_6518_comb = p3_add_6514_comb[9:8];
  assign p3_bit_slice_6519_comb = p3_add_6515_comb[9:8];
  assign p3_bit_slice_6520_comb = p3_add_6516_comb[9:8];
  assign p3_bit_slice_6521_comb = p3_add_6517_comb[9:8];
  assign p3_add_6538_comb = {{1{p2_bit_slice_6478[1]}}, p2_bit_slice_6478} + 3'h1;
  assign p3_add_6539_comb = {{1{p3_bit_slice_6518_comb[1]}}, p3_bit_slice_6518_comb} + 3'h1;
  assign p3_add_6540_comb = {{1{p2_bit_slice_6479[1]}}, p2_bit_slice_6479} + 3'h1;
  assign p3_add_6541_comb = {{1{p3_bit_slice_6519_comb[1]}}, p3_bit_slice_6519_comb} + 3'h1;
  assign p3_add_6542_comb = {{1{p2_bit_slice_6480[1]}}, p2_bit_slice_6480} + 3'h1;
  assign p3_add_6543_comb = {{1{p3_bit_slice_6520_comb[1]}}, p3_bit_slice_6520_comb} + 3'h1;
  assign p3_add_6544_comb = {{1{p2_bit_slice_6481[1]}}, p2_bit_slice_6481} + 3'h1;
  assign p3_add_6545_comb = {{1{p3_bit_slice_6521_comb[1]}}, p3_bit_slice_6521_comb} + 3'h1;
  assign p3_clipped__8_squeezed_const_msb_bits_comb = 1'h0;
  assign p3_clipped__8_squeezed_comb = p3_add_6538_comb[1] ? 9'h0ff : {p3_add_6538_comb[1:0], p2_bit_slice_6482};
  assign p3_clipped__8_squeezed_const_msb_bits__1_comb = 1'h0;
  assign p3_clipped__9_squeezed_comb = p3_add_6539_comb[1] ? 9'h0ff : {p3_add_6539_comb[1:0], p3_add_6514_comb[7:1]};
  assign p3_clipped__8_squeezed_const_msb_bits__2_comb = 1'h0;
  assign p3_clipped__10_squeezed_comb = p3_add_6540_comb[1] ? 9'h0ff : {p3_add_6540_comb[1:0], p2_bit_slice_6483};
  assign p3_clipped__8_squeezed_const_msb_bits__3_comb = 1'h0;
  assign p3_clipped__11_squeezed_comb = p3_add_6541_comb[1] ? 9'h0ff : {p3_add_6541_comb[1:0], p3_add_6515_comb[7:1]};
  assign p3_clipped__8_squeezed_const_msb_bits__4_comb = 1'h0;
  assign p3_clipped__12_squeezed_comb = p3_add_6542_comb[1] ? 9'h0ff : {p3_add_6542_comb[1:0], p2_bit_slice_6484};
  assign p3_clipped__8_squeezed_const_msb_bits__5_comb = 1'h0;
  assign p3_clipped__13_squeezed_comb = p3_add_6543_comb[1] ? 9'h0ff : {p3_add_6543_comb[1:0], p3_add_6516_comb[7:1]};
  assign p3_clipped__8_squeezed_const_msb_bits__6_comb = 1'h0;
  assign p3_clipped__14_squeezed_comb = p3_add_6544_comb[1] ? 9'h0ff : {p3_add_6544_comb[1:0], p2_bit_slice_6485};
  assign p3_clipped__8_squeezed_const_msb_bits__7_comb = 1'h0;
  assign p3_clipped__15_squeezed_comb = p3_add_6545_comb[1] ? 9'h0ff : {p3_add_6545_comb[1:0], p3_add_6517_comb[7:1]};
  assign p3_clipped__8_comb = {p3_clipped__8_squeezed_const_msb_bits_comb, p3_clipped__8_squeezed_comb};
  assign p3_clipped__9_comb = {p3_clipped__8_squeezed_const_msb_bits__1_comb, p3_clipped__9_squeezed_comb};
  assign p3_clipped__10_comb = {p3_clipped__8_squeezed_const_msb_bits__2_comb, p3_clipped__10_squeezed_comb};
  assign p3_clipped__11_comb = {p3_clipped__8_squeezed_const_msb_bits__3_comb, p3_clipped__11_squeezed_comb};
  assign p3_clipped__12_comb = {p3_clipped__8_squeezed_const_msb_bits__4_comb, p3_clipped__12_squeezed_comb};
  assign p3_clipped__13_comb = {p3_clipped__8_squeezed_const_msb_bits__5_comb, p3_clipped__13_squeezed_comb};
  assign p3_clipped__14_comb = {p3_clipped__8_squeezed_const_msb_bits__6_comb, p3_clipped__14_squeezed_comb};
  assign p3_clipped__15_comb = {p3_clipped__8_squeezed_const_msb_bits__7_comb, p3_clipped__15_squeezed_comb};
  assign p3_result_comb[0] = p3_clipped__8_comb;
  assign p3_result_comb[1] = p3_clipped__9_comb;
  assign p3_result_comb[2] = p3_clipped__10_comb;
  assign p3_result_comb[3] = p3_clipped__11_comb;
  assign p3_result_comb[4] = p3_clipped__12_comb;
  assign p3_result_comb[5] = p3_clipped__13_comb;
  assign p3_result_comb[6] = p3_clipped__14_comb;
  assign p3_result_comb[7] = p3_clipped__15_comb;

  // Registers for pipe stage 3:
  reg [9:0] p3_result[0:7];
  always @ (posedge clk) begin
    p3_result[0] <= p3_result_comb[0];
    p3_result[1] <= p3_result_comb[1];
    p3_result[2] <= p3_result_comb[2];
    p3_result[3] <= p3_result_comb[3];
    p3_result[4] <= p3_result_comb[4];
    p3_result[5] <= p3_result_comb[5];
    p3_result[6] <= p3_result_comb[6];
    p3_result[7] <= p3_result_comb[7];
  end
  assign out = {p3_result[7], p3_result[6], p3_result[5], p3_result[4], p3_result[3], p3_result[2], p3_result[1], p3_result[0]};
endmodule
