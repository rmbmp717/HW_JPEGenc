module zigzag_reorder(
  input wire clk,
  input wire [511:0] matrix,
  output wire [511:0] out
);
  wire [7:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[7:0];
  assign matrix_unflattened[0][1] = matrix[15:8];
  assign matrix_unflattened[0][2] = matrix[23:16];
  assign matrix_unflattened[0][3] = matrix[31:24];
  assign matrix_unflattened[0][4] = matrix[39:32];
  assign matrix_unflattened[0][5] = matrix[47:40];
  assign matrix_unflattened[0][6] = matrix[55:48];
  assign matrix_unflattened[0][7] = matrix[63:56];
  assign matrix_unflattened[1][0] = matrix[71:64];
  assign matrix_unflattened[1][1] = matrix[79:72];
  assign matrix_unflattened[1][2] = matrix[87:80];
  assign matrix_unflattened[1][3] = matrix[95:88];
  assign matrix_unflattened[1][4] = matrix[103:96];
  assign matrix_unflattened[1][5] = matrix[111:104];
  assign matrix_unflattened[1][6] = matrix[119:112];
  assign matrix_unflattened[1][7] = matrix[127:120];
  assign matrix_unflattened[2][0] = matrix[135:128];
  assign matrix_unflattened[2][1] = matrix[143:136];
  assign matrix_unflattened[2][2] = matrix[151:144];
  assign matrix_unflattened[2][3] = matrix[159:152];
  assign matrix_unflattened[2][4] = matrix[167:160];
  assign matrix_unflattened[2][5] = matrix[175:168];
  assign matrix_unflattened[2][6] = matrix[183:176];
  assign matrix_unflattened[2][7] = matrix[191:184];
  assign matrix_unflattened[3][0] = matrix[199:192];
  assign matrix_unflattened[3][1] = matrix[207:200];
  assign matrix_unflattened[3][2] = matrix[215:208];
  assign matrix_unflattened[3][3] = matrix[223:216];
  assign matrix_unflattened[3][4] = matrix[231:224];
  assign matrix_unflattened[3][5] = matrix[239:232];
  assign matrix_unflattened[3][6] = matrix[247:240];
  assign matrix_unflattened[3][7] = matrix[255:248];
  assign matrix_unflattened[4][0] = matrix[263:256];
  assign matrix_unflattened[4][1] = matrix[271:264];
  assign matrix_unflattened[4][2] = matrix[279:272];
  assign matrix_unflattened[4][3] = matrix[287:280];
  assign matrix_unflattened[4][4] = matrix[295:288];
  assign matrix_unflattened[4][5] = matrix[303:296];
  assign matrix_unflattened[4][6] = matrix[311:304];
  assign matrix_unflattened[4][7] = matrix[319:312];
  assign matrix_unflattened[5][0] = matrix[327:320];
  assign matrix_unflattened[5][1] = matrix[335:328];
  assign matrix_unflattened[5][2] = matrix[343:336];
  assign matrix_unflattened[5][3] = matrix[351:344];
  assign matrix_unflattened[5][4] = matrix[359:352];
  assign matrix_unflattened[5][5] = matrix[367:360];
  assign matrix_unflattened[5][6] = matrix[375:368];
  assign matrix_unflattened[5][7] = matrix[383:376];
  assign matrix_unflattened[6][0] = matrix[391:384];
  assign matrix_unflattened[6][1] = matrix[399:392];
  assign matrix_unflattened[6][2] = matrix[407:400];
  assign matrix_unflattened[6][3] = matrix[415:408];
  assign matrix_unflattened[6][4] = matrix[423:416];
  assign matrix_unflattened[6][5] = matrix[431:424];
  assign matrix_unflattened[6][6] = matrix[439:432];
  assign matrix_unflattened[6][7] = matrix[447:440];
  assign matrix_unflattened[7][0] = matrix[455:448];
  assign matrix_unflattened[7][1] = matrix[463:456];
  assign matrix_unflattened[7][2] = matrix[471:464];
  assign matrix_unflattened[7][3] = matrix[479:472];
  assign matrix_unflattened[7][4] = matrix[487:480];
  assign matrix_unflattened[7][5] = matrix[495:488];
  assign matrix_unflattened[7][6] = matrix[503:496];
  assign matrix_unflattened[7][7] = matrix[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_matrix[0:7][0:7];
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_array_1498_comb[0:63];
  assign p1_array_1498_comb[0] = p0_matrix[3'h0][3'h0];
  assign p1_array_1498_comb[1] = p0_matrix[3'h0][3'h1];
  assign p1_array_1498_comb[2] = p0_matrix[3'h1][3'h0];
  assign p1_array_1498_comb[3] = p0_matrix[3'h2][3'h0];
  assign p1_array_1498_comb[4] = p0_matrix[3'h1][3'h1];
  assign p1_array_1498_comb[5] = p0_matrix[3'h0][3'h2];
  assign p1_array_1498_comb[6] = p0_matrix[3'h0][3'h3];
  assign p1_array_1498_comb[7] = p0_matrix[3'h1][3'h2];
  assign p1_array_1498_comb[8] = p0_matrix[3'h2][3'h1];
  assign p1_array_1498_comb[9] = p0_matrix[3'h3][3'h0];
  assign p1_array_1498_comb[10] = p0_matrix[3'h4][3'h0];
  assign p1_array_1498_comb[11] = p0_matrix[3'h3][3'h1];
  assign p1_array_1498_comb[12] = p0_matrix[3'h2][3'h2];
  assign p1_array_1498_comb[13] = p0_matrix[3'h1][3'h3];
  assign p1_array_1498_comb[14] = p0_matrix[3'h0][3'h4];
  assign p1_array_1498_comb[15] = p0_matrix[3'h0][3'h5];
  assign p1_array_1498_comb[16] = p0_matrix[3'h1][3'h4];
  assign p1_array_1498_comb[17] = p0_matrix[3'h2][3'h3];
  assign p1_array_1498_comb[18] = p0_matrix[3'h3][3'h2];
  assign p1_array_1498_comb[19] = p0_matrix[3'h4][3'h1];
  assign p1_array_1498_comb[20] = p0_matrix[3'h5][3'h0];
  assign p1_array_1498_comb[21] = p0_matrix[3'h6][3'h0];
  assign p1_array_1498_comb[22] = p0_matrix[3'h5][3'h1];
  assign p1_array_1498_comb[23] = p0_matrix[3'h4][3'h2];
  assign p1_array_1498_comb[24] = p0_matrix[3'h3][3'h3];
  assign p1_array_1498_comb[25] = p0_matrix[3'h2][3'h4];
  assign p1_array_1498_comb[26] = p0_matrix[3'h1][3'h5];
  assign p1_array_1498_comb[27] = p0_matrix[3'h0][3'h6];
  assign p1_array_1498_comb[28] = p0_matrix[3'h0][3'h7];
  assign p1_array_1498_comb[29] = p0_matrix[3'h1][3'h6];
  assign p1_array_1498_comb[30] = p0_matrix[3'h2][3'h5];
  assign p1_array_1498_comb[31] = p0_matrix[3'h3][3'h4];
  assign p1_array_1498_comb[32] = p0_matrix[3'h4][3'h3];
  assign p1_array_1498_comb[33] = p0_matrix[3'h5][3'h2];
  assign p1_array_1498_comb[34] = p0_matrix[3'h6][3'h1];
  assign p1_array_1498_comb[35] = p0_matrix[3'h7][3'h0];
  assign p1_array_1498_comb[36] = p0_matrix[3'h7][3'h1];
  assign p1_array_1498_comb[37] = p0_matrix[3'h6][3'h2];
  assign p1_array_1498_comb[38] = p0_matrix[3'h5][3'h3];
  assign p1_array_1498_comb[39] = p0_matrix[3'h4][3'h4];
  assign p1_array_1498_comb[40] = p0_matrix[3'h3][3'h5];
  assign p1_array_1498_comb[41] = p0_matrix[3'h2][3'h6];
  assign p1_array_1498_comb[42] = p0_matrix[3'h1][3'h7];
  assign p1_array_1498_comb[43] = p0_matrix[3'h2][3'h7];
  assign p1_array_1498_comb[44] = p0_matrix[3'h3][3'h6];
  assign p1_array_1498_comb[45] = p0_matrix[3'h4][3'h5];
  assign p1_array_1498_comb[46] = p0_matrix[3'h5][3'h4];
  assign p1_array_1498_comb[47] = p0_matrix[3'h6][3'h3];
  assign p1_array_1498_comb[48] = p0_matrix[3'h7][3'h2];
  assign p1_array_1498_comb[49] = p0_matrix[3'h7][3'h3];
  assign p1_array_1498_comb[50] = p0_matrix[3'h6][3'h4];
  assign p1_array_1498_comb[51] = p0_matrix[3'h5][3'h5];
  assign p1_array_1498_comb[52] = p0_matrix[3'h4][3'h6];
  assign p1_array_1498_comb[53] = p0_matrix[3'h3][3'h7];
  assign p1_array_1498_comb[54] = p0_matrix[3'h4][3'h7];
  assign p1_array_1498_comb[55] = p0_matrix[3'h5][3'h6];
  assign p1_array_1498_comb[56] = p0_matrix[3'h6][3'h5];
  assign p1_array_1498_comb[57] = p0_matrix[3'h7][3'h4];
  assign p1_array_1498_comb[58] = p0_matrix[3'h7][3'h5];
  assign p1_array_1498_comb[59] = p0_matrix[3'h6][3'h6];
  assign p1_array_1498_comb[60] = p0_matrix[3'h5][3'h7];
  assign p1_array_1498_comb[61] = p0_matrix[3'h6][3'h7];
  assign p1_array_1498_comb[62] = p0_matrix[3'h7][3'h6];
  assign p1_array_1498_comb[63] = p0_matrix[3'h7][3'h7];

  // Registers for pipe stage 1:
  reg [7:0] p1_array_1498[0:63];
  always @ (posedge clk) begin
    p1_array_1498[0] <= p1_array_1498_comb[0];
    p1_array_1498[1] <= p1_array_1498_comb[1];
    p1_array_1498[2] <= p1_array_1498_comb[2];
    p1_array_1498[3] <= p1_array_1498_comb[3];
    p1_array_1498[4] <= p1_array_1498_comb[4];
    p1_array_1498[5] <= p1_array_1498_comb[5];
    p1_array_1498[6] <= p1_array_1498_comb[6];
    p1_array_1498[7] <= p1_array_1498_comb[7];
    p1_array_1498[8] <= p1_array_1498_comb[8];
    p1_array_1498[9] <= p1_array_1498_comb[9];
    p1_array_1498[10] <= p1_array_1498_comb[10];
    p1_array_1498[11] <= p1_array_1498_comb[11];
    p1_array_1498[12] <= p1_array_1498_comb[12];
    p1_array_1498[13] <= p1_array_1498_comb[13];
    p1_array_1498[14] <= p1_array_1498_comb[14];
    p1_array_1498[15] <= p1_array_1498_comb[15];
    p1_array_1498[16] <= p1_array_1498_comb[16];
    p1_array_1498[17] <= p1_array_1498_comb[17];
    p1_array_1498[18] <= p1_array_1498_comb[18];
    p1_array_1498[19] <= p1_array_1498_comb[19];
    p1_array_1498[20] <= p1_array_1498_comb[20];
    p1_array_1498[21] <= p1_array_1498_comb[21];
    p1_array_1498[22] <= p1_array_1498_comb[22];
    p1_array_1498[23] <= p1_array_1498_comb[23];
    p1_array_1498[24] <= p1_array_1498_comb[24];
    p1_array_1498[25] <= p1_array_1498_comb[25];
    p1_array_1498[26] <= p1_array_1498_comb[26];
    p1_array_1498[27] <= p1_array_1498_comb[27];
    p1_array_1498[28] <= p1_array_1498_comb[28];
    p1_array_1498[29] <= p1_array_1498_comb[29];
    p1_array_1498[30] <= p1_array_1498_comb[30];
    p1_array_1498[31] <= p1_array_1498_comb[31];
    p1_array_1498[32] <= p1_array_1498_comb[32];
    p1_array_1498[33] <= p1_array_1498_comb[33];
    p1_array_1498[34] <= p1_array_1498_comb[34];
    p1_array_1498[35] <= p1_array_1498_comb[35];
    p1_array_1498[36] <= p1_array_1498_comb[36];
    p1_array_1498[37] <= p1_array_1498_comb[37];
    p1_array_1498[38] <= p1_array_1498_comb[38];
    p1_array_1498[39] <= p1_array_1498_comb[39];
    p1_array_1498[40] <= p1_array_1498_comb[40];
    p1_array_1498[41] <= p1_array_1498_comb[41];
    p1_array_1498[42] <= p1_array_1498_comb[42];
    p1_array_1498[43] <= p1_array_1498_comb[43];
    p1_array_1498[44] <= p1_array_1498_comb[44];
    p1_array_1498[45] <= p1_array_1498_comb[45];
    p1_array_1498[46] <= p1_array_1498_comb[46];
    p1_array_1498[47] <= p1_array_1498_comb[47];
    p1_array_1498[48] <= p1_array_1498_comb[48];
    p1_array_1498[49] <= p1_array_1498_comb[49];
    p1_array_1498[50] <= p1_array_1498_comb[50];
    p1_array_1498[51] <= p1_array_1498_comb[51];
    p1_array_1498[52] <= p1_array_1498_comb[52];
    p1_array_1498[53] <= p1_array_1498_comb[53];
    p1_array_1498[54] <= p1_array_1498_comb[54];
    p1_array_1498[55] <= p1_array_1498_comb[55];
    p1_array_1498[56] <= p1_array_1498_comb[56];
    p1_array_1498[57] <= p1_array_1498_comb[57];
    p1_array_1498[58] <= p1_array_1498_comb[58];
    p1_array_1498[59] <= p1_array_1498_comb[59];
    p1_array_1498[60] <= p1_array_1498_comb[60];
    p1_array_1498[61] <= p1_array_1498_comb[61];
    p1_array_1498[62] <= p1_array_1498_comb[62];
    p1_array_1498[63] <= p1_array_1498_comb[63];
  end
  assign out = {p1_array_1498[63], p1_array_1498[62], p1_array_1498[61], p1_array_1498[60], p1_array_1498[59], p1_array_1498[58], p1_array_1498[57], p1_array_1498[56], p1_array_1498[55], p1_array_1498[54], p1_array_1498[53], p1_array_1498[52], p1_array_1498[51], p1_array_1498[50], p1_array_1498[49], p1_array_1498[48], p1_array_1498[47], p1_array_1498[46], p1_array_1498[45], p1_array_1498[44], p1_array_1498[43], p1_array_1498[42], p1_array_1498[41], p1_array_1498[40], p1_array_1498[39], p1_array_1498[38], p1_array_1498[37], p1_array_1498[36], p1_array_1498[35], p1_array_1498[34], p1_array_1498[33], p1_array_1498[32], p1_array_1498[31], p1_array_1498[30], p1_array_1498[29], p1_array_1498[28], p1_array_1498[27], p1_array_1498[26], p1_array_1498[25], p1_array_1498[24], p1_array_1498[23], p1_array_1498[22], p1_array_1498[21], p1_array_1498[20], p1_array_1498[19], p1_array_1498[18], p1_array_1498[17], p1_array_1498[16], p1_array_1498[15], p1_array_1498[14], p1_array_1498[13], p1_array_1498[12], p1_array_1498[11], p1_array_1498[10], p1_array_1498[9], p1_array_1498[8], p1_array_1498[7], p1_array_1498[6], p1_array_1498[5], p1_array_1498[4], p1_array_1498[3], p1_array_1498[2], p1_array_1498[1], p1_array_1498[0]};
endmodule
