module dct_2d_u8(
  input wire clk,
  input wire [511:0] x,
  output wire [511:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [15:0] smul16b_8b_x_8b (input reg [7:0] lhs, input reg [7:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [15:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul16b_8b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_6b (input reg [7:0] lhs, input reg [5:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [16:0] smul17b_8b_x_9b (input reg [7:0] lhs, input reg [8:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [16:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul17b_8b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_7b (input reg [31:0] lhs, input reg [6:0] rhs);
    begin
      umul32b_32b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [7:0] x_unflattened[0:7][0:7];
  assign x_unflattened[0][0] = x[7:0];
  assign x_unflattened[0][1] = x[15:8];
  assign x_unflattened[0][2] = x[23:16];
  assign x_unflattened[0][3] = x[31:24];
  assign x_unflattened[0][4] = x[39:32];
  assign x_unflattened[0][5] = x[47:40];
  assign x_unflattened[0][6] = x[55:48];
  assign x_unflattened[0][7] = x[63:56];
  assign x_unflattened[1][0] = x[71:64];
  assign x_unflattened[1][1] = x[79:72];
  assign x_unflattened[1][2] = x[87:80];
  assign x_unflattened[1][3] = x[95:88];
  assign x_unflattened[1][4] = x[103:96];
  assign x_unflattened[1][5] = x[111:104];
  assign x_unflattened[1][6] = x[119:112];
  assign x_unflattened[1][7] = x[127:120];
  assign x_unflattened[2][0] = x[135:128];
  assign x_unflattened[2][1] = x[143:136];
  assign x_unflattened[2][2] = x[151:144];
  assign x_unflattened[2][3] = x[159:152];
  assign x_unflattened[2][4] = x[167:160];
  assign x_unflattened[2][5] = x[175:168];
  assign x_unflattened[2][6] = x[183:176];
  assign x_unflattened[2][7] = x[191:184];
  assign x_unflattened[3][0] = x[199:192];
  assign x_unflattened[3][1] = x[207:200];
  assign x_unflattened[3][2] = x[215:208];
  assign x_unflattened[3][3] = x[223:216];
  assign x_unflattened[3][4] = x[231:224];
  assign x_unflattened[3][5] = x[239:232];
  assign x_unflattened[3][6] = x[247:240];
  assign x_unflattened[3][7] = x[255:248];
  assign x_unflattened[4][0] = x[263:256];
  assign x_unflattened[4][1] = x[271:264];
  assign x_unflattened[4][2] = x[279:272];
  assign x_unflattened[4][3] = x[287:280];
  assign x_unflattened[4][4] = x[295:288];
  assign x_unflattened[4][5] = x[303:296];
  assign x_unflattened[4][6] = x[311:304];
  assign x_unflattened[4][7] = x[319:312];
  assign x_unflattened[5][0] = x[327:320];
  assign x_unflattened[5][1] = x[335:328];
  assign x_unflattened[5][2] = x[343:336];
  assign x_unflattened[5][3] = x[351:344];
  assign x_unflattened[5][4] = x[359:352];
  assign x_unflattened[5][5] = x[367:360];
  assign x_unflattened[5][6] = x[375:368];
  assign x_unflattened[5][7] = x[383:376];
  assign x_unflattened[6][0] = x[391:384];
  assign x_unflattened[6][1] = x[399:392];
  assign x_unflattened[6][2] = x[407:400];
  assign x_unflattened[6][3] = x[415:408];
  assign x_unflattened[6][4] = x[423:416];
  assign x_unflattened[6][5] = x[431:424];
  assign x_unflattened[6][6] = x[439:432];
  assign x_unflattened[6][7] = x[447:440];
  assign x_unflattened[7][0] = x[455:448];
  assign x_unflattened[7][1] = x[463:456];
  assign x_unflattened[7][2] = x[471:464];
  assign x_unflattened[7][3] = x[479:472];
  assign x_unflattened[7][4] = x[487:480];
  assign x_unflattened[7][5] = x[495:488];
  assign x_unflattened[7][6] = x[503:496];
  assign x_unflattened[7][7] = x[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_x[0:7][0:7];
  always @ (posedge clk) begin
    p0_x[0][0] <= x_unflattened[0][0];
    p0_x[0][1] <= x_unflattened[0][1];
    p0_x[0][2] <= x_unflattened[0][2];
    p0_x[0][3] <= x_unflattened[0][3];
    p0_x[0][4] <= x_unflattened[0][4];
    p0_x[0][5] <= x_unflattened[0][5];
    p0_x[0][6] <= x_unflattened[0][6];
    p0_x[0][7] <= x_unflattened[0][7];
    p0_x[1][0] <= x_unflattened[1][0];
    p0_x[1][1] <= x_unflattened[1][1];
    p0_x[1][2] <= x_unflattened[1][2];
    p0_x[1][3] <= x_unflattened[1][3];
    p0_x[1][4] <= x_unflattened[1][4];
    p0_x[1][5] <= x_unflattened[1][5];
    p0_x[1][6] <= x_unflattened[1][6];
    p0_x[1][7] <= x_unflattened[1][7];
    p0_x[2][0] <= x_unflattened[2][0];
    p0_x[2][1] <= x_unflattened[2][1];
    p0_x[2][2] <= x_unflattened[2][2];
    p0_x[2][3] <= x_unflattened[2][3];
    p0_x[2][4] <= x_unflattened[2][4];
    p0_x[2][5] <= x_unflattened[2][5];
    p0_x[2][6] <= x_unflattened[2][6];
    p0_x[2][7] <= x_unflattened[2][7];
    p0_x[3][0] <= x_unflattened[3][0];
    p0_x[3][1] <= x_unflattened[3][1];
    p0_x[3][2] <= x_unflattened[3][2];
    p0_x[3][3] <= x_unflattened[3][3];
    p0_x[3][4] <= x_unflattened[3][4];
    p0_x[3][5] <= x_unflattened[3][5];
    p0_x[3][6] <= x_unflattened[3][6];
    p0_x[3][7] <= x_unflattened[3][7];
    p0_x[4][0] <= x_unflattened[4][0];
    p0_x[4][1] <= x_unflattened[4][1];
    p0_x[4][2] <= x_unflattened[4][2];
    p0_x[4][3] <= x_unflattened[4][3];
    p0_x[4][4] <= x_unflattened[4][4];
    p0_x[4][5] <= x_unflattened[4][5];
    p0_x[4][6] <= x_unflattened[4][6];
    p0_x[4][7] <= x_unflattened[4][7];
    p0_x[5][0] <= x_unflattened[5][0];
    p0_x[5][1] <= x_unflattened[5][1];
    p0_x[5][2] <= x_unflattened[5][2];
    p0_x[5][3] <= x_unflattened[5][3];
    p0_x[5][4] <= x_unflattened[5][4];
    p0_x[5][5] <= x_unflattened[5][5];
    p0_x[5][6] <= x_unflattened[5][6];
    p0_x[5][7] <= x_unflattened[5][7];
    p0_x[6][0] <= x_unflattened[6][0];
    p0_x[6][1] <= x_unflattened[6][1];
    p0_x[6][2] <= x_unflattened[6][2];
    p0_x[6][3] <= x_unflattened[6][3];
    p0_x[6][4] <= x_unflattened[6][4];
    p0_x[6][5] <= x_unflattened[6][5];
    p0_x[6][6] <= x_unflattened[6][6];
    p0_x[6][7] <= x_unflattened[6][7];
    p0_x[7][0] <= x_unflattened[7][0];
    p0_x[7][1] <= x_unflattened[7][1];
    p0_x[7][2] <= x_unflattened[7][2];
    p0_x[7][3] <= x_unflattened[7][3];
    p0_x[7][4] <= x_unflattened[7][4];
    p0_x[7][5] <= x_unflattened[7][5];
    p0_x[7][6] <= x_unflattened[7][6];
    p0_x[7][7] <= x_unflattened[7][7];
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_array_index_133923_comb;
  wire [7:0] p1_array_index_133924_comb;
  wire [7:0] p1_array_index_133925_comb;
  wire [7:0] p1_array_index_133926_comb;
  wire [7:0] p1_array_index_133927_comb;
  wire [7:0] p1_array_index_133928_comb;
  wire [7:0] p1_array_index_133929_comb;
  wire [7:0] p1_array_index_133930_comb;
  wire [7:0] p1_array_index_133931_comb;
  wire [7:0] p1_array_index_133932_comb;
  wire [7:0] p1_array_index_133933_comb;
  wire [7:0] p1_array_index_133934_comb;
  wire [7:0] p1_array_index_133935_comb;
  wire [7:0] p1_array_index_133936_comb;
  wire [7:0] p1_array_index_133937_comb;
  wire [7:0] p1_array_index_133938_comb;
  wire [7:0] p1_array_index_133939_comb;
  wire [7:0] p1_array_index_133940_comb;
  wire [7:0] p1_array_index_133941_comb;
  wire [7:0] p1_array_index_133942_comb;
  wire [7:0] p1_array_index_133943_comb;
  wire [7:0] p1_array_index_133944_comb;
  wire [7:0] p1_array_index_133945_comb;
  wire [7:0] p1_array_index_133946_comb;
  wire [7:0] p1_array_index_133947_comb;
  wire [7:0] p1_array_index_133948_comb;
  wire [7:0] p1_array_index_133949_comb;
  wire [7:0] p1_array_index_133950_comb;
  wire [7:0] p1_array_index_133951_comb;
  wire [7:0] p1_array_index_133952_comb;
  wire [7:0] p1_array_index_133953_comb;
  wire [7:0] p1_array_index_133954_comb;
  wire [7:0] p1_array_index_133955_comb;
  wire [7:0] p1_array_index_133956_comb;
  wire [7:0] p1_array_index_133957_comb;
  wire [7:0] p1_array_index_133958_comb;
  wire [7:0] p1_array_index_133959_comb;
  wire [7:0] p1_array_index_133960_comb;
  wire [7:0] p1_array_index_133961_comb;
  wire [7:0] p1_array_index_133962_comb;
  wire [7:0] p1_array_index_133963_comb;
  wire [7:0] p1_array_index_133964_comb;
  wire [7:0] p1_array_index_133965_comb;
  wire [7:0] p1_array_index_133966_comb;
  wire [7:0] p1_array_index_133967_comb;
  wire [7:0] p1_array_index_133968_comb;
  wire [7:0] p1_array_index_133969_comb;
  wire [7:0] p1_array_index_133970_comb;
  wire [7:0] p1_array_index_133971_comb;
  wire [7:0] p1_array_index_133972_comb;
  wire [7:0] p1_array_index_133973_comb;
  wire [7:0] p1_array_index_133974_comb;
  wire [7:0] p1_array_index_133975_comb;
  wire [7:0] p1_array_index_133976_comb;
  wire [7:0] p1_array_index_133977_comb;
  wire [7:0] p1_array_index_133978_comb;
  wire [7:0] p1_array_index_133979_comb;
  wire [7:0] p1_array_index_133980_comb;
  wire [7:0] p1_array_index_133981_comb;
  wire [7:0] p1_array_index_133982_comb;
  wire [7:0] p1_array_index_133983_comb;
  wire [7:0] p1_array_index_133984_comb;
  wire [7:0] p1_array_index_133985_comb;
  wire [7:0] p1_array_index_133986_comb;
  wire [7:0] p1_shifted__18_squeezed_comb;
  wire [7:0] p1_shifted__21_squeezed_comb;
  wire [7:0] p1_shifted__42_squeezed_comb;
  wire [7:0] p1_shifted__45_squeezed_comb;
  wire [7:0] p1_shifted__16_squeezed_comb;
  wire [7:0] p1_shifted__17_squeezed_comb;
  wire [7:0] p1_shifted__19_squeezed_comb;
  wire [7:0] p1_shifted__20_squeezed_comb;
  wire [7:0] p1_shifted__22_squeezed_comb;
  wire [7:0] p1_shifted__23_squeezed_comb;
  wire [7:0] p1_shifted__40_squeezed_comb;
  wire [7:0] p1_shifted__41_squeezed_comb;
  wire [7:0] p1_shifted__43_squeezed_comb;
  wire [7:0] p1_shifted__44_squeezed_comb;
  wire [7:0] p1_shifted__46_squeezed_comb;
  wire [7:0] p1_shifted__47_squeezed_comb;
  wire [7:0] p1_shifted__2_squeezed_comb;
  wire [7:0] p1_shifted__5_squeezed_comb;
  wire [7:0] p1_shifted__10_squeezed_comb;
  wire [7:0] p1_shifted__13_squeezed_comb;
  wire [7:0] p1_shifted__26_squeezed_comb;
  wire [7:0] p1_shifted__29_squeezed_comb;
  wire [7:0] p1_shifted__34_squeezed_comb;
  wire [7:0] p1_shifted__37_squeezed_comb;
  wire [7:0] p1_shifted__50_squeezed_comb;
  wire [7:0] p1_shifted__53_squeezed_comb;
  wire [7:0] p1_shifted__58_squeezed_comb;
  wire [7:0] p1_shifted__61_squeezed_comb;
  wire [7:0] p1_shifted_squeezed_comb;
  wire [7:0] p1_shifted__1_squeezed_comb;
  wire [7:0] p1_shifted__3_squeezed_comb;
  wire [7:0] p1_shifted__4_squeezed_comb;
  wire [7:0] p1_shifted__6_squeezed_comb;
  wire [7:0] p1_shifted__7_squeezed_comb;
  wire [7:0] p1_shifted__8_squeezed_comb;
  wire [7:0] p1_shifted__9_squeezed_comb;
  wire [7:0] p1_shifted__11_squeezed_comb;
  wire [7:0] p1_shifted__12_squeezed_comb;
  wire [7:0] p1_shifted__14_squeezed_comb;
  wire [7:0] p1_shifted__15_squeezed_comb;
  wire [7:0] p1_shifted__24_squeezed_comb;
  wire [7:0] p1_shifted__25_squeezed_comb;
  wire [7:0] p1_shifted__27_squeezed_comb;
  wire [7:0] p1_shifted__28_squeezed_comb;
  wire [7:0] p1_shifted__30_squeezed_comb;
  wire [7:0] p1_shifted__31_squeezed_comb;
  wire [7:0] p1_shifted__32_squeezed_comb;
  wire [7:0] p1_shifted__33_squeezed_comb;
  wire [7:0] p1_shifted__35_squeezed_comb;
  wire [7:0] p1_shifted__36_squeezed_comb;
  wire [7:0] p1_shifted__38_squeezed_comb;
  wire [7:0] p1_shifted__39_squeezed_comb;
  wire [7:0] p1_shifted__48_squeezed_comb;
  wire [7:0] p1_shifted__49_squeezed_comb;
  wire [7:0] p1_shifted__51_squeezed_comb;
  wire [7:0] p1_shifted__52_squeezed_comb;
  wire [7:0] p1_shifted__54_squeezed_comb;
  wire [7:0] p1_shifted__55_squeezed_comb;
  wire [7:0] p1_shifted__56_squeezed_comb;
  wire [7:0] p1_shifted__57_squeezed_comb;
  wire [7:0] p1_shifted__59_squeezed_comb;
  wire [7:0] p1_shifted__60_squeezed_comb;
  wire [7:0] p1_shifted__62_squeezed_comb;
  wire [7:0] p1_shifted__63_squeezed_comb;
  wire [15:0] p1_smul_57362_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___8_comb;
  wire [15:0] p1_smul_57368_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___11_comb;
  wire [15:0] p1_smul_57410_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___20_comb;
  wire [15:0] p1_smul_57416_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___23_comb;
  wire [14:0] p1_smul_57486_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___8_comb;
  wire [14:0] p1_smul_57488_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___40_comb;
  wire [14:0] p1_smul_57490_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___41_comb;
  wire [14:0] p1_smul_57492_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___9_comb;
  wire [14:0] p1_smul_57494_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___10_comb;
  wire [14:0] p1_smul_57496_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___42_comb;
  wire [14:0] p1_smul_57498_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___43_comb;
  wire [14:0] p1_smul_57500_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___11_comb;
  wire [14:0] p1_smul_57534_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___20_comb;
  wire [14:0] p1_smul_57536_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___52_comb;
  wire [14:0] p1_smul_57538_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___53_comb;
  wire [14:0] p1_smul_57540_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___21_comb;
  wire [14:0] p1_smul_57542_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___22_comb;
  wire [14:0] p1_smul_57544_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___54_comb;
  wire [14:0] p1_smul_57546_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___55_comb;
  wire [14:0] p1_smul_57548_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___23_comb;
  wire [15:0] p1_smul_57620_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___73_comb;
  wire [15:0] p1_smul_57622_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___74_comb;
  wire [15:0] p1_smul_57668_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___85_comb;
  wire [15:0] p1_smul_57670_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___86_comb;
  wire [15:0] p1_smul_57870_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___104_comb;
  wire [15:0] p1_smul_57884_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___107_comb;
  wire [15:0] p1_smul_57918_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___116_comb;
  wire [15:0] p1_smul_57932_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___119_comb;
  wire [14:0] p1_smul_57998_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___136_comb;
  wire [14:0] p1_smul_58000_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___40_comb;
  wire [14:0] p1_smul_58002_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___137_comb;
  wire [14:0] p1_smul_58004_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___41_comb;
  wire [14:0] p1_smul_58006_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___42_comb;
  wire [14:0] p1_smul_58008_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___138_comb;
  wire [14:0] p1_smul_58010_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___43_comb;
  wire [14:0] p1_smul_58012_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___139_comb;
  wire [14:0] p1_smul_58046_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___148_comb;
  wire [14:0] p1_smul_58048_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___52_comb;
  wire [14:0] p1_smul_58050_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___149_comb;
  wire [14:0] p1_smul_58052_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___53_comb;
  wire [14:0] p1_smul_58054_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___54_comb;
  wire [14:0] p1_smul_58056_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___150_comb;
  wire [14:0] p1_smul_58058_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___55_comb;
  wire [14:0] p1_smul_58060_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___151_comb;
  wire [15:0] p1_smul_58128_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___169_comb;
  wire [15:0] p1_smul_58138_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___170_comb;
  wire [15:0] p1_smul_58176_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___181_comb;
  wire [15:0] p1_smul_58186_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___182_comb;
  wire [15:0] p1_smul_57330_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits__comb;
  wire [15:0] p1_smul_57336_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___3_comb;
  wire [15:0] p1_smul_57346_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___4_comb;
  wire [15:0] p1_smul_57352_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___7_comb;
  wire [15:0] p1_smul_57378_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___12_comb;
  wire [15:0] p1_smul_57384_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___15_comb;
  wire [15:0] p1_smul_57394_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___16_comb;
  wire [15:0] p1_smul_57400_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___19_comb;
  wire [15:0] p1_smul_57426_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___24_comb;
  wire [15:0] p1_smul_57432_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___27_comb;
  wire [15:0] p1_smul_57442_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___28_comb;
  wire [15:0] p1_smul_57448_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___31_comb;
  wire [14:0] p1_smul_57454_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits__comb;
  wire [14:0] p1_smul_57456_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___32_comb;
  wire [14:0] p1_smul_57458_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___33_comb;
  wire [14:0] p1_smul_57460_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___1_comb;
  wire [14:0] p1_smul_57462_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___2_comb;
  wire [14:0] p1_smul_57464_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___34_comb;
  wire [14:0] p1_smul_57466_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___35_comb;
  wire [14:0] p1_smul_57468_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___3_comb;
  wire [14:0] p1_smul_57470_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___4_comb;
  wire [14:0] p1_smul_57472_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___36_comb;
  wire [14:0] p1_smul_57474_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___37_comb;
  wire [14:0] p1_smul_57476_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___5_comb;
  wire [14:0] p1_smul_57478_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___6_comb;
  wire [14:0] p1_smul_57480_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___38_comb;
  wire [14:0] p1_smul_57482_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___39_comb;
  wire [14:0] p1_smul_57484_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___7_comb;
  wire [14:0] p1_smul_57502_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___12_comb;
  wire [14:0] p1_smul_57504_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___44_comb;
  wire [14:0] p1_smul_57506_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___45_comb;
  wire [14:0] p1_smul_57508_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___13_comb;
  wire [14:0] p1_smul_57510_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___14_comb;
  wire [14:0] p1_smul_57512_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___46_comb;
  wire [14:0] p1_smul_57514_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___47_comb;
  wire [14:0] p1_smul_57516_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___15_comb;
  wire [14:0] p1_smul_57518_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___16_comb;
  wire [14:0] p1_smul_57520_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___48_comb;
  wire [14:0] p1_smul_57522_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___49_comb;
  wire [14:0] p1_smul_57524_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___17_comb;
  wire [14:0] p1_smul_57526_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___18_comb;
  wire [14:0] p1_smul_57528_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___50_comb;
  wire [14:0] p1_smul_57530_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___51_comb;
  wire [14:0] p1_smul_57532_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___19_comb;
  wire [14:0] p1_smul_57550_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___24_comb;
  wire [14:0] p1_smul_57552_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___56_comb;
  wire [14:0] p1_smul_57554_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___57_comb;
  wire [14:0] p1_smul_57556_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___25_comb;
  wire [14:0] p1_smul_57558_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___26_comb;
  wire [14:0] p1_smul_57560_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___58_comb;
  wire [14:0] p1_smul_57562_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___59_comb;
  wire [14:0] p1_smul_57564_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___27_comb;
  wire [14:0] p1_smul_57566_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___28_comb;
  wire [14:0] p1_smul_57568_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___60_comb;
  wire [14:0] p1_smul_57570_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___61_comb;
  wire [14:0] p1_smul_57572_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___29_comb;
  wire [14:0] p1_smul_57574_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___30_comb;
  wire [14:0] p1_smul_57576_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___62_comb;
  wire [14:0] p1_smul_57578_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___63_comb;
  wire [14:0] p1_smul_57580_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___31_comb;
  wire [15:0] p1_smul_57588_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___65_comb;
  wire [15:0] p1_smul_57590_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___66_comb;
  wire [15:0] p1_smul_57604_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___69_comb;
  wire [15:0] p1_smul_57606_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___70_comb;
  wire [15:0] p1_smul_57636_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___77_comb;
  wire [15:0] p1_smul_57638_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___78_comb;
  wire [15:0] p1_smul_57652_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___81_comb;
  wire [15:0] p1_smul_57654_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___82_comb;
  wire [15:0] p1_smul_57684_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___89_comb;
  wire [15:0] p1_smul_57686_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___90_comb;
  wire [15:0] p1_smul_57700_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___93_comb;
  wire [15:0] p1_smul_57702_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___94_comb;
  wire [15:0] p1_smul_57838_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___96_comb;
  wire [15:0] p1_smul_57852_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___99_comb;
  wire [15:0] p1_smul_57854_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___100_comb;
  wire [15:0] p1_smul_57868_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___103_comb;
  wire [15:0] p1_smul_57886_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___108_comb;
  wire [15:0] p1_smul_57900_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___111_comb;
  wire [15:0] p1_smul_57902_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___112_comb;
  wire [15:0] p1_smul_57916_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___115_comb;
  wire [15:0] p1_smul_57934_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___120_comb;
  wire [15:0] p1_smul_57948_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___123_comb;
  wire [15:0] p1_smul_57950_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___124_comb;
  wire [15:0] p1_smul_57964_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___127_comb;
  wire [14:0] p1_smul_57966_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___128_comb;
  wire [14:0] p1_smul_57968_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___32_comb;
  wire [14:0] p1_smul_57970_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___129_comb;
  wire [14:0] p1_smul_57972_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___33_comb;
  wire [14:0] p1_smul_57974_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___34_comb;
  wire [14:0] p1_smul_57976_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___130_comb;
  wire [14:0] p1_smul_57978_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___35_comb;
  wire [14:0] p1_smul_57980_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___131_comb;
  wire [14:0] p1_smul_57982_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___132_comb;
  wire [14:0] p1_smul_57984_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___36_comb;
  wire [14:0] p1_smul_57986_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___133_comb;
  wire [14:0] p1_smul_57988_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___37_comb;
  wire [14:0] p1_smul_57990_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___38_comb;
  wire [14:0] p1_smul_57992_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___134_comb;
  wire [14:0] p1_smul_57994_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___39_comb;
  wire [14:0] p1_smul_57996_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___135_comb;
  wire [14:0] p1_smul_58014_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___140_comb;
  wire [14:0] p1_smul_58016_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___44_comb;
  wire [14:0] p1_smul_58018_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___141_comb;
  wire [14:0] p1_smul_58020_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___45_comb;
  wire [14:0] p1_smul_58022_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___46_comb;
  wire [14:0] p1_smul_58024_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___142_comb;
  wire [14:0] p1_smul_58026_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___47_comb;
  wire [14:0] p1_smul_58028_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___143_comb;
  wire [14:0] p1_smul_58030_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___144_comb;
  wire [14:0] p1_smul_58032_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___48_comb;
  wire [14:0] p1_smul_58034_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___145_comb;
  wire [14:0] p1_smul_58036_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___49_comb;
  wire [14:0] p1_smul_58038_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___50_comb;
  wire [14:0] p1_smul_58040_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___146_comb;
  wire [14:0] p1_smul_58042_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___51_comb;
  wire [14:0] p1_smul_58044_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___147_comb;
  wire [14:0] p1_smul_58062_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___152_comb;
  wire [14:0] p1_smul_58064_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___56_comb;
  wire [14:0] p1_smul_58066_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___153_comb;
  wire [14:0] p1_smul_58068_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___57_comb;
  wire [14:0] p1_smul_58070_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___58_comb;
  wire [14:0] p1_smul_58072_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___154_comb;
  wire [14:0] p1_smul_58074_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___59_comb;
  wire [14:0] p1_smul_58076_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___155_comb;
  wire [14:0] p1_smul_58078_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___156_comb;
  wire [14:0] p1_smul_58080_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___60_comb;
  wire [14:0] p1_smul_58082_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___157_comb;
  wire [14:0] p1_smul_58084_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___61_comb;
  wire [14:0] p1_smul_58086_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___62_comb;
  wire [14:0] p1_smul_58088_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___158_comb;
  wire [14:0] p1_smul_58090_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___63_comb;
  wire [14:0] p1_smul_58092_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___159_comb;
  wire [15:0] p1_smul_58096_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___161_comb;
  wire [15:0] p1_smul_58106_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___162_comb;
  wire [15:0] p1_smul_58112_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___165_comb;
  wire [15:0] p1_smul_58122_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___166_comb;
  wire [15:0] p1_smul_58144_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___173_comb;
  wire [15:0] p1_smul_58154_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___174_comb;
  wire [15:0] p1_smul_58160_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___177_comb;
  wire [15:0] p1_smul_58170_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___178_comb;
  wire [15:0] p1_smul_58192_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___185_comb;
  wire [15:0] p1_smul_58202_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___186_comb;
  wire [15:0] p1_smul_58208_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___189_comb;
  wire [15:0] p1_smul_58218_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___190_comb;
  wire [24:0] p1_concat_134899_comb;
  wire [13:0] p1_smul_57364_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___9_comb;
  wire [13:0] p1_smul_57366_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___10_comb;
  wire [24:0] p1_concat_134904_comb;
  wire [24:0] p1_concat_134905_comb;
  wire [13:0] p1_smul_57412_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___21_comb;
  wire [13:0] p1_smul_57414_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___22_comb;
  wire [24:0] p1_concat_134910_comb;
  wire [24:0] p1_concat_134911_comb;
  wire [23:0] p1_concat_134912_comb;
  wire [23:0] p1_concat_134913_comb;
  wire [24:0] p1_concat_134914_comb;
  wire [24:0] p1_concat_134915_comb;
  wire [23:0] p1_concat_134916_comb;
  wire [23:0] p1_concat_134917_comb;
  wire [24:0] p1_concat_134918_comb;
  wire [24:0] p1_concat_134919_comb;
  wire [23:0] p1_concat_134920_comb;
  wire [23:0] p1_concat_134921_comb;
  wire [24:0] p1_concat_134922_comb;
  wire [24:0] p1_concat_134923_comb;
  wire [23:0] p1_concat_134924_comb;
  wire [23:0] p1_concat_134925_comb;
  wire [24:0] p1_concat_134926_comb;
  wire [13:0] p1_smul_57616_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___72_comb;
  wire [24:0] p1_concat_134929_comb;
  wire [24:0] p1_concat_134930_comb;
  wire [13:0] p1_smul_57626_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___75_comb;
  wire [13:0] p1_smul_57664_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___84_comb;
  wire [24:0] p1_concat_134935_comb;
  wire [24:0] p1_concat_134936_comb;
  wire [13:0] p1_smul_57674_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___87_comb;
  wire [24:0] p1_concat_134939_comb;
  wire [13:0] p1_smul_57874_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___105_comb;
  wire [13:0] p1_smul_57880_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___106_comb;
  wire [24:0] p1_concat_134944_comb;
  wire [24:0] p1_concat_134945_comb;
  wire [13:0] p1_smul_57922_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___117_comb;
  wire [13:0] p1_smul_57928_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___118_comb;
  wire [24:0] p1_concat_134950_comb;
  wire [23:0] p1_concat_134951_comb;
  wire [24:0] p1_concat_134952_comb;
  wire [23:0] p1_concat_134953_comb;
  wire [24:0] p1_concat_134954_comb;
  wire [24:0] p1_concat_134955_comb;
  wire [23:0] p1_concat_134956_comb;
  wire [24:0] p1_concat_134957_comb;
  wire [23:0] p1_concat_134958_comb;
  wire [23:0] p1_concat_134959_comb;
  wire [24:0] p1_concat_134960_comb;
  wire [23:0] p1_concat_134961_comb;
  wire [24:0] p1_concat_134962_comb;
  wire [24:0] p1_concat_134963_comb;
  wire [23:0] p1_concat_134964_comb;
  wire [24:0] p1_concat_134965_comb;
  wire [23:0] p1_concat_134966_comb;
  wire [13:0] p1_smul_58126_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___168_comb;
  wire [24:0] p1_concat_134969_comb;
  wire [24:0] p1_concat_134970_comb;
  wire [13:0] p1_smul_58140_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___171_comb;
  wire [13:0] p1_smul_58174_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___180_comb;
  wire [24:0] p1_concat_134975_comb;
  wire [24:0] p1_concat_134976_comb;
  wire [13:0] p1_smul_58188_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___183_comb;
  wire [24:0] p1_concat_135027_comb;
  wire [13:0] p1_smul_57332_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___1_comb;
  wire [13:0] p1_smul_57334_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___2_comb;
  wire [24:0] p1_concat_135032_comb;
  wire [24:0] p1_concat_135033_comb;
  wire [13:0] p1_smul_57348_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___5_comb;
  wire [13:0] p1_smul_57350_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___6_comb;
  wire [24:0] p1_concat_135038_comb;
  wire [24:0] p1_concat_135039_comb;
  wire [13:0] p1_smul_57380_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___13_comb;
  wire [13:0] p1_smul_57382_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___14_comb;
  wire [24:0] p1_concat_135044_comb;
  wire [24:0] p1_concat_135045_comb;
  wire [13:0] p1_smul_57396_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___17_comb;
  wire [13:0] p1_smul_57398_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___18_comb;
  wire [24:0] p1_concat_135050_comb;
  wire [24:0] p1_concat_135051_comb;
  wire [13:0] p1_smul_57428_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___25_comb;
  wire [13:0] p1_smul_57430_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___26_comb;
  wire [24:0] p1_concat_135056_comb;
  wire [24:0] p1_concat_135057_comb;
  wire [13:0] p1_smul_57444_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___29_comb;
  wire [13:0] p1_smul_57446_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___30_comb;
  wire [24:0] p1_concat_135062_comb;
  wire [24:0] p1_concat_135063_comb;
  wire [23:0] p1_concat_135064_comb;
  wire [23:0] p1_concat_135065_comb;
  wire [24:0] p1_concat_135066_comb;
  wire [24:0] p1_concat_135067_comb;
  wire [23:0] p1_concat_135068_comb;
  wire [23:0] p1_concat_135069_comb;
  wire [24:0] p1_concat_135070_comb;
  wire [24:0] p1_concat_135071_comb;
  wire [23:0] p1_concat_135072_comb;
  wire [23:0] p1_concat_135073_comb;
  wire [24:0] p1_concat_135074_comb;
  wire [24:0] p1_concat_135075_comb;
  wire [23:0] p1_concat_135076_comb;
  wire [23:0] p1_concat_135077_comb;
  wire [24:0] p1_concat_135078_comb;
  wire [24:0] p1_concat_135079_comb;
  wire [23:0] p1_concat_135080_comb;
  wire [23:0] p1_concat_135081_comb;
  wire [24:0] p1_concat_135082_comb;
  wire [24:0] p1_concat_135083_comb;
  wire [23:0] p1_concat_135084_comb;
  wire [23:0] p1_concat_135085_comb;
  wire [24:0] p1_concat_135086_comb;
  wire [24:0] p1_concat_135087_comb;
  wire [23:0] p1_concat_135088_comb;
  wire [23:0] p1_concat_135089_comb;
  wire [24:0] p1_concat_135090_comb;
  wire [24:0] p1_concat_135091_comb;
  wire [23:0] p1_concat_135092_comb;
  wire [23:0] p1_concat_135093_comb;
  wire [24:0] p1_concat_135094_comb;
  wire [24:0] p1_concat_135095_comb;
  wire [23:0] p1_concat_135096_comb;
  wire [23:0] p1_concat_135097_comb;
  wire [24:0] p1_concat_135098_comb;
  wire [24:0] p1_concat_135099_comb;
  wire [23:0] p1_concat_135100_comb;
  wire [23:0] p1_concat_135101_comb;
  wire [24:0] p1_concat_135102_comb;
  wire [24:0] p1_concat_135103_comb;
  wire [23:0] p1_concat_135104_comb;
  wire [23:0] p1_concat_135105_comb;
  wire [24:0] p1_concat_135106_comb;
  wire [24:0] p1_concat_135107_comb;
  wire [23:0] p1_concat_135108_comb;
  wire [23:0] p1_concat_135109_comb;
  wire [24:0] p1_concat_135110_comb;
  wire [13:0] p1_smul_57584_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___64_comb;
  wire [24:0] p1_concat_135113_comb;
  wire [24:0] p1_concat_135114_comb;
  wire [13:0] p1_smul_57594_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___67_comb;
  wire [13:0] p1_smul_57600_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___68_comb;
  wire [24:0] p1_concat_135119_comb;
  wire [24:0] p1_concat_135120_comb;
  wire [13:0] p1_smul_57610_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___71_comb;
  wire [13:0] p1_smul_57632_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___76_comb;
  wire [24:0] p1_concat_135125_comb;
  wire [24:0] p1_concat_135126_comb;
  wire [13:0] p1_smul_57642_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___79_comb;
  wire [13:0] p1_smul_57648_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___80_comb;
  wire [24:0] p1_concat_135131_comb;
  wire [24:0] p1_concat_135132_comb;
  wire [13:0] p1_smul_57658_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___83_comb;
  wire [13:0] p1_smul_57680_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___88_comb;
  wire [24:0] p1_concat_135137_comb;
  wire [24:0] p1_concat_135138_comb;
  wire [13:0] p1_smul_57690_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___91_comb;
  wire [13:0] p1_smul_57696_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___92_comb;
  wire [24:0] p1_concat_135143_comb;
  wire [24:0] p1_concat_135144_comb;
  wire [13:0] p1_smul_57706_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___95_comb;
  wire [24:0] p1_concat_135147_comb;
  wire [13:0] p1_smul_57842_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___97_comb;
  wire [13:0] p1_smul_57848_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___98_comb;
  wire [24:0] p1_concat_135152_comb;
  wire [24:0] p1_concat_135153_comb;
  wire [13:0] p1_smul_57858_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___101_comb;
  wire [13:0] p1_smul_57864_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___102_comb;
  wire [24:0] p1_concat_135158_comb;
  wire [24:0] p1_concat_135159_comb;
  wire [13:0] p1_smul_57890_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___109_comb;
  wire [13:0] p1_smul_57896_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___110_comb;
  wire [24:0] p1_concat_135164_comb;
  wire [24:0] p1_concat_135165_comb;
  wire [13:0] p1_smul_57906_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___113_comb;
  wire [13:0] p1_smul_57912_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___114_comb;
  wire [24:0] p1_concat_135170_comb;
  wire [24:0] p1_concat_135171_comb;
  wire [13:0] p1_smul_57938_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___121_comb;
  wire [13:0] p1_smul_57944_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___122_comb;
  wire [24:0] p1_concat_135176_comb;
  wire [24:0] p1_concat_135177_comb;
  wire [13:0] p1_smul_57954_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___125_comb;
  wire [13:0] p1_smul_57960_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___126_comb;
  wire [24:0] p1_concat_135182_comb;
  wire [23:0] p1_concat_135183_comb;
  wire [24:0] p1_concat_135184_comb;
  wire [23:0] p1_concat_135185_comb;
  wire [24:0] p1_concat_135186_comb;
  wire [24:0] p1_concat_135187_comb;
  wire [23:0] p1_concat_135188_comb;
  wire [24:0] p1_concat_135189_comb;
  wire [23:0] p1_concat_135190_comb;
  wire [23:0] p1_concat_135191_comb;
  wire [24:0] p1_concat_135192_comb;
  wire [23:0] p1_concat_135193_comb;
  wire [24:0] p1_concat_135194_comb;
  wire [24:0] p1_concat_135195_comb;
  wire [23:0] p1_concat_135196_comb;
  wire [24:0] p1_concat_135197_comb;
  wire [23:0] p1_concat_135198_comb;
  wire [23:0] p1_concat_135199_comb;
  wire [24:0] p1_concat_135200_comb;
  wire [23:0] p1_concat_135201_comb;
  wire [24:0] p1_concat_135202_comb;
  wire [24:0] p1_concat_135203_comb;
  wire [23:0] p1_concat_135204_comb;
  wire [24:0] p1_concat_135205_comb;
  wire [23:0] p1_concat_135206_comb;
  wire [23:0] p1_concat_135207_comb;
  wire [24:0] p1_concat_135208_comb;
  wire [23:0] p1_concat_135209_comb;
  wire [24:0] p1_concat_135210_comb;
  wire [24:0] p1_concat_135211_comb;
  wire [23:0] p1_concat_135212_comb;
  wire [24:0] p1_concat_135213_comb;
  wire [23:0] p1_concat_135214_comb;
  wire [23:0] p1_concat_135215_comb;
  wire [24:0] p1_concat_135216_comb;
  wire [23:0] p1_concat_135217_comb;
  wire [24:0] p1_concat_135218_comb;
  wire [24:0] p1_concat_135219_comb;
  wire [23:0] p1_concat_135220_comb;
  wire [24:0] p1_concat_135221_comb;
  wire [23:0] p1_concat_135222_comb;
  wire [23:0] p1_concat_135223_comb;
  wire [24:0] p1_concat_135224_comb;
  wire [23:0] p1_concat_135225_comb;
  wire [24:0] p1_concat_135226_comb;
  wire [24:0] p1_concat_135227_comb;
  wire [23:0] p1_concat_135228_comb;
  wire [24:0] p1_concat_135229_comb;
  wire [23:0] p1_concat_135230_comb;
  wire [13:0] p1_smul_58094_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___160_comb;
  wire [24:0] p1_concat_135233_comb;
  wire [24:0] p1_concat_135234_comb;
  wire [13:0] p1_smul_58108_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___163_comb;
  wire [13:0] p1_smul_58110_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___164_comb;
  wire [24:0] p1_concat_135239_comb;
  wire [24:0] p1_concat_135240_comb;
  wire [13:0] p1_smul_58124_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___167_comb;
  wire [13:0] p1_smul_58142_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___172_comb;
  wire [24:0] p1_concat_135245_comb;
  wire [24:0] p1_concat_135246_comb;
  wire [13:0] p1_smul_58156_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___175_comb;
  wire [13:0] p1_smul_58158_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___176_comb;
  wire [24:0] p1_concat_135251_comb;
  wire [24:0] p1_concat_135252_comb;
  wire [13:0] p1_smul_58172_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___179_comb;
  wire [13:0] p1_smul_58190_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___184_comb;
  wire [24:0] p1_concat_135257_comb;
  wire [24:0] p1_concat_135258_comb;
  wire [13:0] p1_smul_58204_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___187_comb;
  wire [13:0] p1_smul_58206_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___188_comb;
  wire [24:0] p1_concat_135263_comb;
  wire [24:0] p1_concat_135264_comb;
  wire [13:0] p1_smul_58220_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___191_comb;
  wire [7:0] p1_smul_57326_TrailingBits___144_comb;
  wire [7:0] p1_smul_57326_TrailingBits___145_comb;
  wire [7:0] p1_smul_57326_TrailingBits___146_comb;
  wire [7:0] p1_smul_57326_TrailingBits___147_comb;
  wire [7:0] p1_smul_57326_TrailingBits___148_comb;
  wire [7:0] p1_smul_57326_TrailingBits___149_comb;
  wire [7:0] p1_smul_57326_TrailingBits___150_comb;
  wire [7:0] p1_smul_57326_TrailingBits___151_comb;
  wire [7:0] p1_smul_57326_TrailingBits___168_comb;
  wire [7:0] p1_smul_57326_TrailingBits___169_comb;
  wire [7:0] p1_smul_57326_TrailingBits___170_comb;
  wire [7:0] p1_smul_57326_TrailingBits___171_comb;
  wire [7:0] p1_smul_57326_TrailingBits___172_comb;
  wire [7:0] p1_smul_57326_TrailingBits___173_comb;
  wire [7:0] p1_smul_57326_TrailingBits___174_comb;
  wire [7:0] p1_smul_57326_TrailingBits___175_comb;
  wire [31:0] p1_prod__135_comb;
  wire [22:0] p1_concat_135317_comb;
  wire [22:0] p1_concat_135318_comb;
  wire [31:0] p1_prod__150_comb;
  wire [31:0] p1_prod__327_comb;
  wire [22:0] p1_concat_135323_comb;
  wire [22:0] p1_concat_135324_comb;
  wire [31:0] p1_prod__342_comb;
  wire [31:0] p1_prod__133_comb;
  wire [31:0] p1_prod__136_comb;
  wire [31:0] p1_prod__140_comb;
  wire [31:0] p1_prod__145_comb;
  wire [31:0] p1_prod__151_comb;
  wire [31:0] p1_prod__158_comb;
  wire [31:0] p1_prod__165_comb;
  wire [31:0] p1_prod__171_comb;
  wire [31:0] p1_prod__325_comb;
  wire [31:0] p1_prod__328_comb;
  wire [31:0] p1_prod__332_comb;
  wire [31:0] p1_prod__337_comb;
  wire [31:0] p1_prod__343_comb;
  wire [31:0] p1_prod__350_comb;
  wire [31:0] p1_prod__357_comb;
  wire [31:0] p1_prod__363_comb;
  wire [22:0] p1_concat_135351_comb;
  wire [31:0] p1_prod__152_comb;
  wire [31:0] p1_prod__159_comb;
  wire [22:0] p1_concat_135356_comb;
  wire [22:0] p1_concat_135357_comb;
  wire [31:0] p1_prod__344_comb;
  wire [31:0] p1_prod__351_comb;
  wire [22:0] p1_concat_135362_comb;
  wire [31:0] p1_prod__148_comb;
  wire [22:0] p1_concat_135365_comb;
  wire [22:0] p1_concat_135366_comb;
  wire [31:0] p1_prod__186_comb;
  wire [31:0] p1_prod__340_comb;
  wire [22:0] p1_concat_135371_comb;
  wire [22:0] p1_concat_135372_comb;
  wire [31:0] p1_prod__378_comb;
  wire [31:0] p1_prod__155_comb;
  wire [31:0] p1_prod__162_comb;
  wire [31:0] p1_prod__169_comb;
  wire [31:0] p1_prod__175_comb;
  wire [31:0] p1_prod__180_comb;
  wire [31:0] p1_prod__184_comb;
  wire [31:0] p1_prod__187_comb;
  wire [31:0] p1_prod__189_comb;
  wire [31:0] p1_prod__347_comb;
  wire [31:0] p1_prod__354_comb;
  wire [31:0] p1_prod__361_comb;
  wire [31:0] p1_prod__367_comb;
  wire [31:0] p1_prod__372_comb;
  wire [31:0] p1_prod__376_comb;
  wire [31:0] p1_prod__379_comb;
  wire [31:0] p1_prod__381_comb;
  wire [22:0] p1_concat_135399_comb;
  wire [31:0] p1_prod__170_comb;
  wire [31:0] p1_prod__190_comb;
  wire [22:0] p1_concat_135404_comb;
  wire [22:0] p1_concat_135405_comb;
  wire [31:0] p1_prod__362_comb;
  wire [31:0] p1_prod__382_comb;
  wire [22:0] p1_concat_135410_comb;
  wire [7:0] p1_smul_57326_TrailingBits___128_comb;
  wire [7:0] p1_smul_57326_TrailingBits___129_comb;
  wire [7:0] p1_smul_57326_TrailingBits___130_comb;
  wire [7:0] p1_smul_57326_TrailingBits___131_comb;
  wire [7:0] p1_smul_57326_TrailingBits___132_comb;
  wire [7:0] p1_smul_57326_TrailingBits___133_comb;
  wire [7:0] p1_smul_57326_TrailingBits___134_comb;
  wire [7:0] p1_smul_57326_TrailingBits___135_comb;
  wire [7:0] p1_smul_57326_TrailingBits___136_comb;
  wire [7:0] p1_smul_57326_TrailingBits___137_comb;
  wire [7:0] p1_smul_57326_TrailingBits___138_comb;
  wire [7:0] p1_smul_57326_TrailingBits___139_comb;
  wire [7:0] p1_smul_57326_TrailingBits___140_comb;
  wire [7:0] p1_smul_57326_TrailingBits___141_comb;
  wire [7:0] p1_smul_57326_TrailingBits___142_comb;
  wire [7:0] p1_smul_57326_TrailingBits___143_comb;
  wire [7:0] p1_smul_57326_TrailingBits___152_comb;
  wire [7:0] p1_smul_57326_TrailingBits___153_comb;
  wire [7:0] p1_smul_57326_TrailingBits___154_comb;
  wire [7:0] p1_smul_57326_TrailingBits___155_comb;
  wire [7:0] p1_smul_57326_TrailingBits___156_comb;
  wire [7:0] p1_smul_57326_TrailingBits___157_comb;
  wire [7:0] p1_smul_57326_TrailingBits___158_comb;
  wire [7:0] p1_smul_57326_TrailingBits___159_comb;
  wire [7:0] p1_smul_57326_TrailingBits___160_comb;
  wire [7:0] p1_smul_57326_TrailingBits___161_comb;
  wire [7:0] p1_smul_57326_TrailingBits___162_comb;
  wire [7:0] p1_smul_57326_TrailingBits___163_comb;
  wire [7:0] p1_smul_57326_TrailingBits___164_comb;
  wire [7:0] p1_smul_57326_TrailingBits___165_comb;
  wire [7:0] p1_smul_57326_TrailingBits___166_comb;
  wire [7:0] p1_smul_57326_TrailingBits___167_comb;
  wire [7:0] p1_smul_57326_TrailingBits___176_comb;
  wire [7:0] p1_smul_57326_TrailingBits___177_comb;
  wire [7:0] p1_smul_57326_TrailingBits___178_comb;
  wire [7:0] p1_smul_57326_TrailingBits___179_comb;
  wire [7:0] p1_smul_57326_TrailingBits___180_comb;
  wire [7:0] p1_smul_57326_TrailingBits___181_comb;
  wire [7:0] p1_smul_57326_TrailingBits___182_comb;
  wire [7:0] p1_smul_57326_TrailingBits___183_comb;
  wire [7:0] p1_smul_57326_TrailingBits___184_comb;
  wire [7:0] p1_smul_57326_TrailingBits___185_comb;
  wire [7:0] p1_smul_57326_TrailingBits___186_comb;
  wire [7:0] p1_smul_57326_TrailingBits___187_comb;
  wire [7:0] p1_smul_57326_TrailingBits___188_comb;
  wire [7:0] p1_smul_57326_TrailingBits___189_comb;
  wire [7:0] p1_smul_57326_TrailingBits___190_comb;
  wire [7:0] p1_smul_57326_TrailingBits___191_comb;
  wire [31:0] p1_prod__10_comb;
  wire [22:0] p1_concat_135557_comb;
  wire [22:0] p1_concat_135558_comb;
  wire [31:0] p1_prod__13_comb;
  wire [31:0] p1_prod__71_comb;
  wire [22:0] p1_concat_135563_comb;
  wire [22:0] p1_concat_135564_comb;
  wire [31:0] p1_prod__86_comb;
  wire [31:0] p1_prod__199_comb;
  wire [22:0] p1_concat_135569_comb;
  wire [22:0] p1_concat_135570_comb;
  wire [31:0] p1_prod__214_comb;
  wire [31:0] p1_prod__263_comb;
  wire [22:0] p1_concat_135575_comb;
  wire [22:0] p1_concat_135576_comb;
  wire [31:0] p1_prod__278_comb;
  wire [31:0] p1_prod__391_comb;
  wire [22:0] p1_concat_135581_comb;
  wire [22:0] p1_concat_135582_comb;
  wire [31:0] p1_prod__406_comb;
  wire [31:0] p1_prod__455_comb;
  wire [22:0] p1_concat_135587_comb;
  wire [22:0] p1_concat_135588_comb;
  wire [31:0] p1_prod__470_comb;
  wire [31:0] p1_prod__16_comb;
  wire [31:0] p1_prod__17_comb;
  wire [31:0] p1_prod__18_comb;
  wire [31:0] p1_prod__19_comb;
  wire [31:0] p1_prod__20_comb;
  wire [31:0] p1_prod__21_comb;
  wire [31:0] p1_prod__22_comb;
  wire [31:0] p1_prod__23_comb;
  wire [31:0] p1_prod__69_comb;
  wire [31:0] p1_prod__72_comb;
  wire [31:0] p1_prod__76_comb;
  wire [31:0] p1_prod__81_comb;
  wire [31:0] p1_prod__87_comb;
  wire [31:0] p1_prod__94_comb;
  wire [31:0] p1_prod__101_comb;
  wire [31:0] p1_prod__107_comb;
  wire [31:0] p1_prod__197_comb;
  wire [31:0] p1_prod__200_comb;
  wire [31:0] p1_prod__204_comb;
  wire [31:0] p1_prod__209_comb;
  wire [31:0] p1_prod__215_comb;
  wire [31:0] p1_prod__222_comb;
  wire [31:0] p1_prod__229_comb;
  wire [31:0] p1_prod__235_comb;
  wire [31:0] p1_prod__261_comb;
  wire [31:0] p1_prod__264_comb;
  wire [31:0] p1_prod__268_comb;
  wire [31:0] p1_prod__273_comb;
  wire [31:0] p1_prod__279_comb;
  wire [31:0] p1_prod__286_comb;
  wire [31:0] p1_prod__293_comb;
  wire [31:0] p1_prod__299_comb;
  wire [31:0] p1_prod__389_comb;
  wire [31:0] p1_prod__392_comb;
  wire [31:0] p1_prod__396_comb;
  wire [31:0] p1_prod__401_comb;
  wire [31:0] p1_prod__407_comb;
  wire [31:0] p1_prod__414_comb;
  wire [31:0] p1_prod__421_comb;
  wire [31:0] p1_prod__427_comb;
  wire [31:0] p1_prod__453_comb;
  wire [31:0] p1_prod__456_comb;
  wire [31:0] p1_prod__460_comb;
  wire [31:0] p1_prod__465_comb;
  wire [31:0] p1_prod__471_comb;
  wire [31:0] p1_prod__478_comb;
  wire [31:0] p1_prod__485_comb;
  wire [31:0] p1_prod__491_comb;
  wire [22:0] p1_concat_135663_comb;
  wire [31:0] p1_prod__27_comb;
  wire [31:0] p1_prod__28_comb;
  wire [22:0] p1_concat_135668_comb;
  wire [22:0] p1_concat_135669_comb;
  wire [31:0] p1_prod__88_comb;
  wire [31:0] p1_prod__95_comb;
  wire [22:0] p1_concat_135674_comb;
  wire [22:0] p1_concat_135675_comb;
  wire [31:0] p1_prod__216_comb;
  wire [31:0] p1_prod__223_comb;
  wire [22:0] p1_concat_135680_comb;
  wire [22:0] p1_concat_135681_comb;
  wire [31:0] p1_prod__280_comb;
  wire [31:0] p1_prod__287_comb;
  wire [22:0] p1_concat_135686_comb;
  wire [22:0] p1_concat_135687_comb;
  wire [31:0] p1_prod__408_comb;
  wire [31:0] p1_prod__415_comb;
  wire [22:0] p1_concat_135692_comb;
  wire [22:0] p1_concat_135693_comb;
  wire [31:0] p1_prod__472_comb;
  wire [31:0] p1_prod__479_comb;
  wire [22:0] p1_concat_135698_comb;
  wire [31:0] p1_prod__40_comb;
  wire [22:0] p1_concat_135701_comb;
  wire [22:0] p1_concat_135702_comb;
  wire [31:0] p1_prod__47_comb;
  wire [31:0] p1_prod__84_comb;
  wire [22:0] p1_concat_135707_comb;
  wire [22:0] p1_concat_135708_comb;
  wire [31:0] p1_prod__122_comb;
  wire [31:0] p1_prod__212_comb;
  wire [22:0] p1_concat_135713_comb;
  wire [22:0] p1_concat_135714_comb;
  wire [31:0] p1_prod__250_comb;
  wire [31:0] p1_prod__276_comb;
  wire [22:0] p1_concat_135719_comb;
  wire [22:0] p1_concat_135720_comb;
  wire [31:0] p1_prod__314_comb;
  wire [31:0] p1_prod__404_comb;
  wire [22:0] p1_concat_135725_comb;
  wire [22:0] p1_concat_135726_comb;
  wire [31:0] p1_prod__442_comb;
  wire [31:0] p1_prod__468_comb;
  wire [22:0] p1_concat_135731_comb;
  wire [22:0] p1_concat_135732_comb;
  wire [31:0] p1_prod__506_comb;
  wire [31:0] p1_prod__48_comb;
  wire [31:0] p1_prod__49_comb;
  wire [31:0] p1_prod__50_comb;
  wire [31:0] p1_prod__51_comb;
  wire [31:0] p1_prod__52_comb;
  wire [31:0] p1_prod__53_comb;
  wire [31:0] p1_prod__54_comb;
  wire [31:0] p1_prod__55_comb;
  wire [31:0] p1_prod__91_comb;
  wire [31:0] p1_prod__98_comb;
  wire [31:0] p1_prod__105_comb;
  wire [31:0] p1_prod__111_comb;
  wire [31:0] p1_prod__116_comb;
  wire [31:0] p1_prod__120_comb;
  wire [31:0] p1_prod__123_comb;
  wire [31:0] p1_prod__125_comb;
  wire [31:0] p1_prod__219_comb;
  wire [31:0] p1_prod__226_comb;
  wire [31:0] p1_prod__233_comb;
  wire [31:0] p1_prod__239_comb;
  wire [31:0] p1_prod__244_comb;
  wire [31:0] p1_prod__248_comb;
  wire [31:0] p1_prod__251_comb;
  wire [31:0] p1_prod__253_comb;
  wire [31:0] p1_prod__283_comb;
  wire [31:0] p1_prod__290_comb;
  wire [31:0] p1_prod__297_comb;
  wire [31:0] p1_prod__303_comb;
  wire [31:0] p1_prod__308_comb;
  wire [31:0] p1_prod__312_comb;
  wire [31:0] p1_prod__315_comb;
  wire [31:0] p1_prod__317_comb;
  wire [31:0] p1_prod__411_comb;
  wire [31:0] p1_prod__418_comb;
  wire [31:0] p1_prod__425_comb;
  wire [31:0] p1_prod__431_comb;
  wire [31:0] p1_prod__436_comb;
  wire [31:0] p1_prod__440_comb;
  wire [31:0] p1_prod__443_comb;
  wire [31:0] p1_prod__445_comb;
  wire [31:0] p1_prod__475_comb;
  wire [31:0] p1_prod__482_comb;
  wire [31:0] p1_prod__489_comb;
  wire [31:0] p1_prod__495_comb;
  wire [31:0] p1_prod__500_comb;
  wire [31:0] p1_prod__504_comb;
  wire [31:0] p1_prod__507_comb;
  wire [31:0] p1_prod__509_comb;
  wire [22:0] p1_concat_135807_comb;
  wire [31:0] p1_prod__57_comb;
  wire [31:0] p1_prod__62_comb;
  wire [22:0] p1_concat_135812_comb;
  wire [22:0] p1_concat_135813_comb;
  wire [31:0] p1_prod__106_comb;
  wire [31:0] p1_prod__126_comb;
  wire [22:0] p1_concat_135818_comb;
  wire [22:0] p1_concat_135819_comb;
  wire [31:0] p1_prod__234_comb;
  wire [31:0] p1_prod__254_comb;
  wire [22:0] p1_concat_135824_comb;
  wire [22:0] p1_concat_135825_comb;
  wire [31:0] p1_prod__298_comb;
  wire [31:0] p1_prod__318_comb;
  wire [22:0] p1_concat_135830_comb;
  wire [22:0] p1_concat_135831_comb;
  wire [31:0] p1_prod__426_comb;
  wire [31:0] p1_prod__446_comb;
  wire [22:0] p1_concat_135836_comb;
  wire [22:0] p1_concat_135837_comb;
  wire [31:0] p1_prod__490_comb;
  wire [31:0] p1_prod__510_comb;
  wire [22:0] p1_concat_135842_comb;
  wire [15:0] p1_shifted__16_comb;
  wire [7:0] p1_smul_57326_TrailingBits___16_comb;
  wire [15:0] p1_shifted__17_comb;
  wire [7:0] p1_smul_57326_TrailingBits___17_comb;
  wire [15:0] p1_shifted__18_comb;
  wire [7:0] p1_smul_57326_TrailingBits___18_comb;
  wire [15:0] p1_shifted__19_comb;
  wire [7:0] p1_smul_57326_TrailingBits___19_comb;
  wire [15:0] p1_shifted__20_comb;
  wire [7:0] p1_smul_57326_TrailingBits___20_comb;
  wire [15:0] p1_shifted__21_comb;
  wire [7:0] p1_smul_57326_TrailingBits___21_comb;
  wire [15:0] p1_shifted__22_comb;
  wire [7:0] p1_smul_57326_TrailingBits___22_comb;
  wire [15:0] p1_shifted__23_comb;
  wire [7:0] p1_smul_57326_TrailingBits___23_comb;
  wire [15:0] p1_shifted__40_comb;
  wire [7:0] p1_smul_57326_TrailingBits___40_comb;
  wire [15:0] p1_shifted__41_comb;
  wire [7:0] p1_smul_57326_TrailingBits___41_comb;
  wire [15:0] p1_shifted__42_comb;
  wire [7:0] p1_smul_57326_TrailingBits___42_comb;
  wire [15:0] p1_shifted__43_comb;
  wire [7:0] p1_smul_57326_TrailingBits___43_comb;
  wire [15:0] p1_shifted__44_comb;
  wire [7:0] p1_smul_57326_TrailingBits___44_comb;
  wire [15:0] p1_shifted__45_comb;
  wire [7:0] p1_smul_57326_TrailingBits___45_comb;
  wire [15:0] p1_shifted__46_comb;
  wire [7:0] p1_smul_57326_TrailingBits___46_comb;
  wire [15:0] p1_shifted__47_comb;
  wire [7:0] p1_smul_57326_TrailingBits___47_comb;
  wire [31:0] p1_or_135911_comb;
  wire [31:0] p1_prod__139_comb;
  wire [31:0] p1_prod__144_comb;
  wire [31:0] p1_or_135918_comb;
  wire [31:0] p1_or_135925_comb;
  wire [31:0] p1_prod__331_comb;
  wire [31:0] p1_prod__336_comb;
  wire [31:0] p1_or_135932_comb;
  wire [31:0] p1_or_135937_comb;
  wire [31:0] p1_or_135944_comb;
  wire [31:0] p1_or_135947_comb;
  wire [31:0] p1_or_135954_comb;
  wire [31:0] p1_or_135957_comb;
  wire [31:0] p1_or_135964_comb;
  wire [31:0] p1_or_135967_comb;
  wire [31:0] p1_or_135974_comb;
  wire [31:0] p1_prod__141_comb;
  wire [31:0] p1_or_135981_comb;
  wire [31:0] p1_or_135984_comb;
  wire [31:0] p1_prod__172_comb;
  wire [31:0] p1_prod__333_comb;
  wire [31:0] p1_or_135995_comb;
  wire [31:0] p1_or_135998_comb;
  wire [31:0] p1_prod__364_comb;
  wire [31:0] p1_or_136021_comb;
  wire [31:0] p1_prod__161_comb;
  wire [31:0] p1_prod__179_comb;
  wire [31:0] p1_or_136032_comb;
  wire [31:0] p1_or_136035_comb;
  wire [31:0] p1_prod__353_comb;
  wire [31:0] p1_prod__371_comb;
  wire [31:0] p1_or_136046_comb;
  wire [31:0] p1_or_136051_comb;
  wire [31:0] p1_or_136056_comb;
  wire [31:0] p1_or_136059_comb;
  wire [31:0] p1_or_136064_comb;
  wire [31:0] p1_or_136071_comb;
  wire [31:0] p1_or_136076_comb;
  wire [31:0] p1_or_136079_comb;
  wire [31:0] p1_or_136084_comb;
  wire [31:0] p1_prod__163_comb;
  wire [31:0] p1_or_136091_comb;
  wire [31:0] p1_or_136098_comb;
  wire [31:0] p1_prod__191_comb;
  wire [31:0] p1_prod__355_comb;
  wire [31:0] p1_or_136105_comb;
  wire [31:0] p1_or_136112_comb;
  wire [31:0] p1_prod__383_comb;
  wire [15:0] p1_shifted_comb;
  wire [7:0] p1_smul_57326_TrailingBits__comb;
  wire [15:0] p1_shifted__1_comb;
  wire [7:0] p1_smul_57326_TrailingBits___1_comb;
  wire [15:0] p1_shifted__2_comb;
  wire [7:0] p1_smul_57326_TrailingBits___2_comb;
  wire [15:0] p1_shifted__3_comb;
  wire [7:0] p1_smul_57326_TrailingBits___3_comb;
  wire [15:0] p1_shifted__4_comb;
  wire [7:0] p1_smul_57326_TrailingBits___4_comb;
  wire [15:0] p1_shifted__5_comb;
  wire [7:0] p1_smul_57326_TrailingBits___5_comb;
  wire [15:0] p1_shifted__6_comb;
  wire [7:0] p1_smul_57326_TrailingBits___6_comb;
  wire [15:0] p1_shifted__7_comb;
  wire [7:0] p1_smul_57326_TrailingBits___7_comb;
  wire [15:0] p1_shifted__8_comb;
  wire [7:0] p1_smul_57326_TrailingBits___8_comb;
  wire [15:0] p1_shifted__9_comb;
  wire [7:0] p1_smul_57326_TrailingBits___9_comb;
  wire [15:0] p1_shifted__10_comb;
  wire [7:0] p1_smul_57326_TrailingBits___10_comb;
  wire [15:0] p1_shifted__11_comb;
  wire [7:0] p1_smul_57326_TrailingBits___11_comb;
  wire [15:0] p1_shifted__12_comb;
  wire [7:0] p1_smul_57326_TrailingBits___12_comb;
  wire [15:0] p1_shifted__13_comb;
  wire [7:0] p1_smul_57326_TrailingBits___13_comb;
  wire [15:0] p1_shifted__14_comb;
  wire [7:0] p1_smul_57326_TrailingBits___14_comb;
  wire [15:0] p1_shifted__15_comb;
  wire [7:0] p1_smul_57326_TrailingBits___15_comb;
  wire [15:0] p1_shifted__24_comb;
  wire [7:0] p1_smul_57326_TrailingBits___24_comb;
  wire [15:0] p1_shifted__25_comb;
  wire [7:0] p1_smul_57326_TrailingBits___25_comb;
  wire [15:0] p1_shifted__26_comb;
  wire [7:0] p1_smul_57326_TrailingBits___26_comb;
  wire [15:0] p1_shifted__27_comb;
  wire [7:0] p1_smul_57326_TrailingBits___27_comb;
  wire [15:0] p1_shifted__28_comb;
  wire [7:0] p1_smul_57326_TrailingBits___28_comb;
  wire [15:0] p1_shifted__29_comb;
  wire [7:0] p1_smul_57326_TrailingBits___29_comb;
  wire [15:0] p1_shifted__30_comb;
  wire [7:0] p1_smul_57326_TrailingBits___30_comb;
  wire [15:0] p1_shifted__31_comb;
  wire [7:0] p1_smul_57326_TrailingBits___31_comb;
  wire [15:0] p1_shifted__32_comb;
  wire [7:0] p1_smul_57326_TrailingBits___32_comb;
  wire [15:0] p1_shifted__33_comb;
  wire [7:0] p1_smul_57326_TrailingBits___33_comb;
  wire [15:0] p1_shifted__34_comb;
  wire [7:0] p1_smul_57326_TrailingBits___34_comb;
  wire [15:0] p1_shifted__35_comb;
  wire [7:0] p1_smul_57326_TrailingBits___35_comb;
  wire [15:0] p1_shifted__36_comb;
  wire [7:0] p1_smul_57326_TrailingBits___36_comb;
  wire [15:0] p1_shifted__37_comb;
  wire [7:0] p1_smul_57326_TrailingBits___37_comb;
  wire [15:0] p1_shifted__38_comb;
  wire [7:0] p1_smul_57326_TrailingBits___38_comb;
  wire [15:0] p1_shifted__39_comb;
  wire [7:0] p1_smul_57326_TrailingBits___39_comb;
  wire [15:0] p1_shifted__48_comb;
  wire [7:0] p1_smul_57326_TrailingBits___48_comb;
  wire [15:0] p1_shifted__49_comb;
  wire [7:0] p1_smul_57326_TrailingBits___49_comb;
  wire [15:0] p1_shifted__50_comb;
  wire [7:0] p1_smul_57326_TrailingBits___50_comb;
  wire [15:0] p1_shifted__51_comb;
  wire [7:0] p1_smul_57326_TrailingBits___51_comb;
  wire [15:0] p1_shifted__52_comb;
  wire [7:0] p1_smul_57326_TrailingBits___52_comb;
  wire [15:0] p1_shifted__53_comb;
  wire [7:0] p1_smul_57326_TrailingBits___53_comb;
  wire [15:0] p1_shifted__54_comb;
  wire [7:0] p1_smul_57326_TrailingBits___54_comb;
  wire [15:0] p1_shifted__55_comb;
  wire [7:0] p1_smul_57326_TrailingBits___55_comb;
  wire [15:0] p1_shifted__56_comb;
  wire [7:0] p1_smul_57326_TrailingBits___56_comb;
  wire [15:0] p1_shifted__57_comb;
  wire [7:0] p1_smul_57326_TrailingBits___57_comb;
  wire [15:0] p1_shifted__58_comb;
  wire [7:0] p1_smul_57326_TrailingBits___58_comb;
  wire [15:0] p1_shifted__59_comb;
  wire [7:0] p1_smul_57326_TrailingBits___59_comb;
  wire [15:0] p1_shifted__60_comb;
  wire [7:0] p1_smul_57326_TrailingBits___60_comb;
  wire [15:0] p1_shifted__61_comb;
  wire [7:0] p1_smul_57326_TrailingBits___61_comb;
  wire [15:0] p1_shifted__62_comb;
  wire [7:0] p1_smul_57326_TrailingBits___62_comb;
  wire [15:0] p1_shifted__63_comb;
  wire [7:0] p1_smul_57326_TrailingBits___63_comb;
  wire [31:0] p1_or_136311_comb;
  wire [31:0] p1_prod__11_comb;
  wire [31:0] p1_prod__12_comb;
  wire [31:0] p1_or_136318_comb;
  wire [31:0] p1_or_136325_comb;
  wire [31:0] p1_prod__75_comb;
  wire [31:0] p1_prod__80_comb;
  wire [31:0] p1_or_136332_comb;
  wire [31:0] p1_or_136339_comb;
  wire [31:0] p1_prod__203_comb;
  wire [31:0] p1_prod__208_comb;
  wire [31:0] p1_or_136346_comb;
  wire [31:0] p1_or_136353_comb;
  wire [31:0] p1_prod__267_comb;
  wire [31:0] p1_prod__272_comb;
  wire [31:0] p1_or_136360_comb;
  wire [31:0] p1_or_136367_comb;
  wire [31:0] p1_prod__395_comb;
  wire [31:0] p1_prod__400_comb;
  wire [31:0] p1_or_136374_comb;
  wire [31:0] p1_or_136381_comb;
  wire [31:0] p1_prod__459_comb;
  wire [31:0] p1_prod__464_comb;
  wire [31:0] p1_or_136388_comb;
  wire [31:0] p1_or_136393_comb;
  wire [31:0] p1_or_136400_comb;
  wire [31:0] p1_or_136403_comb;
  wire [31:0] p1_or_136410_comb;
  wire [31:0] p1_or_136413_comb;
  wire [31:0] p1_or_136420_comb;
  wire [31:0] p1_or_136423_comb;
  wire [31:0] p1_or_136430_comb;
  wire [31:0] p1_or_136433_comb;
  wire [31:0] p1_or_136440_comb;
  wire [31:0] p1_or_136443_comb;
  wire [31:0] p1_or_136450_comb;
  wire [31:0] p1_or_136453_comb;
  wire [31:0] p1_or_136460_comb;
  wire [31:0] p1_or_136463_comb;
  wire [31:0] p1_or_136470_comb;
  wire [31:0] p1_or_136473_comb;
  wire [31:0] p1_or_136480_comb;
  wire [31:0] p1_or_136483_comb;
  wire [31:0] p1_or_136490_comb;
  wire [31:0] p1_or_136493_comb;
  wire [31:0] p1_or_136500_comb;
  wire [31:0] p1_or_136503_comb;
  wire [31:0] p1_or_136510_comb;
  wire [31:0] p1_prod__25_comb;
  wire [31:0] p1_or_136517_comb;
  wire [31:0] p1_or_136520_comb;
  wire [31:0] p1_prod__30_comb;
  wire [31:0] p1_prod__77_comb;
  wire [31:0] p1_or_136531_comb;
  wire [31:0] p1_or_136534_comb;
  wire [31:0] p1_prod__108_comb;
  wire [31:0] p1_prod__205_comb;
  wire [31:0] p1_or_136545_comb;
  wire [31:0] p1_or_136548_comb;
  wire [31:0] p1_prod__236_comb;
  wire [31:0] p1_prod__269_comb;
  wire [31:0] p1_or_136559_comb;
  wire [31:0] p1_or_136562_comb;
  wire [31:0] p1_prod__300_comb;
  wire [31:0] p1_prod__397_comb;
  wire [31:0] p1_or_136573_comb;
  wire [31:0] p1_or_136576_comb;
  wire [31:0] p1_prod__428_comb;
  wire [31:0] p1_prod__461_comb;
  wire [31:0] p1_or_136587_comb;
  wire [31:0] p1_or_136590_comb;
  wire [31:0] p1_prod__492_comb;
  wire [31:0] p1_or_136645_comb;
  wire [31:0] p1_prod__42_comb;
  wire [31:0] p1_prod__45_comb;
  wire [31:0] p1_or_136656_comb;
  wire [31:0] p1_or_136659_comb;
  wire [31:0] p1_prod__97_comb;
  wire [31:0] p1_prod__115_comb;
  wire [31:0] p1_or_136670_comb;
  wire [31:0] p1_or_136673_comb;
  wire [31:0] p1_prod__225_comb;
  wire [31:0] p1_prod__243_comb;
  wire [31:0] p1_or_136684_comb;
  wire [31:0] p1_or_136687_comb;
  wire [31:0] p1_prod__289_comb;
  wire [31:0] p1_prod__307_comb;
  wire [31:0] p1_or_136698_comb;
  wire [31:0] p1_or_136701_comb;
  wire [31:0] p1_prod__417_comb;
  wire [31:0] p1_prod__435_comb;
  wire [31:0] p1_or_136712_comb;
  wire [31:0] p1_or_136715_comb;
  wire [31:0] p1_prod__481_comb;
  wire [31:0] p1_prod__499_comb;
  wire [31:0] p1_or_136726_comb;
  wire [31:0] p1_or_136731_comb;
  wire [31:0] p1_or_136736_comb;
  wire [31:0] p1_or_136739_comb;
  wire [31:0] p1_or_136744_comb;
  wire [31:0] p1_or_136751_comb;
  wire [31:0] p1_or_136756_comb;
  wire [31:0] p1_or_136759_comb;
  wire [31:0] p1_or_136764_comb;
  wire [31:0] p1_or_136771_comb;
  wire [31:0] p1_or_136776_comb;
  wire [31:0] p1_or_136779_comb;
  wire [31:0] p1_or_136784_comb;
  wire [31:0] p1_or_136791_comb;
  wire [31:0] p1_or_136796_comb;
  wire [31:0] p1_or_136799_comb;
  wire [31:0] p1_or_136804_comb;
  wire [31:0] p1_or_136811_comb;
  wire [31:0] p1_or_136816_comb;
  wire [31:0] p1_or_136819_comb;
  wire [31:0] p1_or_136824_comb;
  wire [31:0] p1_or_136831_comb;
  wire [31:0] p1_or_136836_comb;
  wire [31:0] p1_or_136839_comb;
  wire [31:0] p1_or_136844_comb;
  wire [31:0] p1_prod__56_comb;
  wire [31:0] p1_or_136851_comb;
  wire [31:0] p1_or_136858_comb;
  wire [31:0] p1_prod__63_comb;
  wire [31:0] p1_prod__99_comb;
  wire [31:0] p1_or_136865_comb;
  wire [31:0] p1_or_136872_comb;
  wire [31:0] p1_prod__127_comb;
  wire [31:0] p1_prod__227_comb;
  wire [31:0] p1_or_136879_comb;
  wire [31:0] p1_or_136886_comb;
  wire [31:0] p1_prod__255_comb;
  wire [31:0] p1_prod__291_comb;
  wire [31:0] p1_or_136893_comb;
  wire [31:0] p1_or_136900_comb;
  wire [31:0] p1_prod__319_comb;
  wire [31:0] p1_prod__419_comb;
  wire [31:0] p1_or_136907_comb;
  wire [31:0] p1_or_136914_comb;
  wire [31:0] p1_prod__447_comb;
  wire [31:0] p1_prod__483_comb;
  wire [31:0] p1_or_136921_comb;
  wire [31:0] p1_or_136928_comb;
  wire [31:0] p1_prod__511_comb;
  wire [16:0] p1_smul_57358_NarrowedMult__comb;
  wire [16:0] p1_smul_57360_NarrowedMult__comb;
  wire [31:0] p1_or_136986_comb;
  wire [31:0] p1_or_136987_comb;
  wire [16:0] p1_smul_57370_NarrowedMult__comb;
  wire [16:0] p1_smul_57372_NarrowedMult__comb;
  wire [16:0] p1_smul_57406_NarrowedMult__comb;
  wire [16:0] p1_smul_57408_NarrowedMult__comb;
  wire [31:0] p1_or_137002_comb;
  wire [31:0] p1_or_137003_comb;
  wire [16:0] p1_smul_57418_NarrowedMult__comb;
  wire [16:0] p1_smul_57420_NarrowedMult__comb;
  wire [16:0] p1_smul_57614_NarrowedMult__comb;
  wire [31:0] p1_or_137053_comb;
  wire [16:0] p1_smul_57618_NarrowedMult__comb;
  wire [16:0] p1_smul_57624_NarrowedMult__comb;
  wire [31:0] p1_or_137064_comb;
  wire [16:0] p1_smul_57628_NarrowedMult__comb;
  wire [16:0] p1_smul_57662_NarrowedMult__comb;
  wire [31:0] p1_or_137069_comb;
  wire [16:0] p1_smul_57666_NarrowedMult__comb;
  wire [16:0] p1_smul_57672_NarrowedMult__comb;
  wire [31:0] p1_or_137080_comb;
  wire [16:0] p1_smul_57676_NarrowedMult__comb;
  wire [16:0] p1_smul_57742_NarrowedMult__comb;
  wire [16:0] p1_smul_57744_NarrowedMult__comb;
  wire [16:0] p1_smul_57746_NarrowedMult__comb;
  wire [16:0] p1_smul_57748_NarrowedMult__comb;
  wire [16:0] p1_smul_57750_NarrowedMult__comb;
  wire [16:0] p1_smul_57752_NarrowedMult__comb;
  wire [16:0] p1_smul_57754_NarrowedMult__comb;
  wire [16:0] p1_smul_57756_NarrowedMult__comb;
  wire [16:0] p1_smul_57790_NarrowedMult__comb;
  wire [16:0] p1_smul_57792_NarrowedMult__comb;
  wire [16:0] p1_smul_57794_NarrowedMult__comb;
  wire [16:0] p1_smul_57796_NarrowedMult__comb;
  wire [16:0] p1_smul_57798_NarrowedMult__comb;
  wire [16:0] p1_smul_57800_NarrowedMult__comb;
  wire [16:0] p1_smul_57802_NarrowedMult__comb;
  wire [16:0] p1_smul_57804_NarrowedMult__comb;
  wire [16:0] p1_smul_57872_NarrowedMult__comb;
  wire [31:0] p1_or_137120_comb;
  wire [16:0] p1_smul_57876_NarrowedMult__comb;
  wire [16:0] p1_smul_57878_NarrowedMult__comb;
  wire [31:0] p1_or_137125_comb;
  wire [16:0] p1_smul_57882_NarrowedMult__comb;
  wire [16:0] p1_smul_57920_NarrowedMult__comb;
  wire [31:0] p1_or_137136_comb;
  wire [16:0] p1_smul_57924_NarrowedMult__comb;
  wire [16:0] p1_smul_57926_NarrowedMult__comb;
  wire [31:0] p1_or_137141_comb;
  wire [16:0] p1_smul_57930_NarrowedMult__comb;
  wire [31:0] p1_or_137187_comb;
  wire [16:0] p1_smul_58130_NarrowedMult__comb;
  wire [16:0] p1_smul_58132_NarrowedMult__comb;
  wire [16:0] p1_smul_58134_NarrowedMult__comb;
  wire [16:0] p1_smul_58136_NarrowedMult__comb;
  wire [31:0] p1_or_137202_comb;
  wire [31:0] p1_or_137203_comb;
  wire [16:0] p1_smul_58178_NarrowedMult__comb;
  wire [16:0] p1_smul_58180_NarrowedMult__comb;
  wire [16:0] p1_smul_58182_NarrowedMult__comb;
  wire [16:0] p1_smul_58184_NarrowedMult__comb;
  wire [31:0] p1_or_137218_comb;
  wire [16:0] p1_smul_57326_NarrowedMult__comb;
  wire [16:0] p1_smul_57328_NarrowedMult__comb;
  wire [31:0] p1_or_137370_comb;
  wire [31:0] p1_or_137371_comb;
  wire [16:0] p1_smul_57338_NarrowedMult__comb;
  wire [16:0] p1_smul_57340_NarrowedMult__comb;
  wire [16:0] p1_smul_57342_NarrowedMult__comb;
  wire [16:0] p1_smul_57344_NarrowedMult__comb;
  wire [31:0] p1_or_137386_comb;
  wire [31:0] p1_or_137387_comb;
  wire [16:0] p1_smul_57354_NarrowedMult__comb;
  wire [16:0] p1_smul_57356_NarrowedMult__comb;
  wire [16:0] p1_smul_57374_NarrowedMult__comb;
  wire [16:0] p1_smul_57376_NarrowedMult__comb;
  wire [31:0] p1_or_137402_comb;
  wire [31:0] p1_or_137403_comb;
  wire [16:0] p1_smul_57386_NarrowedMult__comb;
  wire [16:0] p1_smul_57388_NarrowedMult__comb;
  wire [16:0] p1_smul_57390_NarrowedMult__comb;
  wire [16:0] p1_smul_57392_NarrowedMult__comb;
  wire [31:0] p1_or_137418_comb;
  wire [31:0] p1_or_137419_comb;
  wire [16:0] p1_smul_57402_NarrowedMult__comb;
  wire [16:0] p1_smul_57404_NarrowedMult__comb;
  wire [16:0] p1_smul_57422_NarrowedMult__comb;
  wire [16:0] p1_smul_57424_NarrowedMult__comb;
  wire [31:0] p1_or_137434_comb;
  wire [31:0] p1_or_137435_comb;
  wire [16:0] p1_smul_57434_NarrowedMult__comb;
  wire [16:0] p1_smul_57436_NarrowedMult__comb;
  wire [16:0] p1_smul_57438_NarrowedMult__comb;
  wire [16:0] p1_smul_57440_NarrowedMult__comb;
  wire [31:0] p1_or_137450_comb;
  wire [31:0] p1_or_137451_comb;
  wire [16:0] p1_smul_57450_NarrowedMult__comb;
  wire [16:0] p1_smul_57452_NarrowedMult__comb;
  wire [16:0] p1_smul_57582_NarrowedMult__comb;
  wire [31:0] p1_or_137581_comb;
  wire [16:0] p1_smul_57586_NarrowedMult__comb;
  wire [16:0] p1_smul_57592_NarrowedMult__comb;
  wire [31:0] p1_or_137592_comb;
  wire [16:0] p1_smul_57596_NarrowedMult__comb;
  wire [16:0] p1_smul_57598_NarrowedMult__comb;
  wire [31:0] p1_or_137597_comb;
  wire [16:0] p1_smul_57602_NarrowedMult__comb;
  wire [16:0] p1_smul_57608_NarrowedMult__comb;
  wire [31:0] p1_or_137608_comb;
  wire [16:0] p1_smul_57612_NarrowedMult__comb;
  wire [16:0] p1_smul_57630_NarrowedMult__comb;
  wire [31:0] p1_or_137613_comb;
  wire [16:0] p1_smul_57634_NarrowedMult__comb;
  wire [16:0] p1_smul_57640_NarrowedMult__comb;
  wire [31:0] p1_or_137624_comb;
  wire [16:0] p1_smul_57644_NarrowedMult__comb;
  wire [16:0] p1_smul_57646_NarrowedMult__comb;
  wire [31:0] p1_or_137629_comb;
  wire [16:0] p1_smul_57650_NarrowedMult__comb;
  wire [16:0] p1_smul_57656_NarrowedMult__comb;
  wire [31:0] p1_or_137640_comb;
  wire [16:0] p1_smul_57660_NarrowedMult__comb;
  wire [16:0] p1_smul_57678_NarrowedMult__comb;
  wire [31:0] p1_or_137645_comb;
  wire [16:0] p1_smul_57682_NarrowedMult__comb;
  wire [16:0] p1_smul_57688_NarrowedMult__comb;
  wire [31:0] p1_or_137656_comb;
  wire [16:0] p1_smul_57692_NarrowedMult__comb;
  wire [16:0] p1_smul_57694_NarrowedMult__comb;
  wire [31:0] p1_or_137661_comb;
  wire [16:0] p1_smul_57698_NarrowedMult__comb;
  wire [16:0] p1_smul_57704_NarrowedMult__comb;
  wire [31:0] p1_or_137672_comb;
  wire [16:0] p1_smul_57708_NarrowedMult__comb;
  wire [16:0] p1_smul_57710_NarrowedMult__comb;
  wire [16:0] p1_smul_57712_NarrowedMult__comb;
  wire [16:0] p1_smul_57714_NarrowedMult__comb;
  wire [16:0] p1_smul_57716_NarrowedMult__comb;
  wire [16:0] p1_smul_57718_NarrowedMult__comb;
  wire [16:0] p1_smul_57720_NarrowedMult__comb;
  wire [16:0] p1_smul_57722_NarrowedMult__comb;
  wire [16:0] p1_smul_57724_NarrowedMult__comb;
  wire [16:0] p1_smul_57726_NarrowedMult__comb;
  wire [16:0] p1_smul_57728_NarrowedMult__comb;
  wire [16:0] p1_smul_57730_NarrowedMult__comb;
  wire [16:0] p1_smul_57732_NarrowedMult__comb;
  wire [16:0] p1_smul_57734_NarrowedMult__comb;
  wire [16:0] p1_smul_57736_NarrowedMult__comb;
  wire [16:0] p1_smul_57738_NarrowedMult__comb;
  wire [16:0] p1_smul_57740_NarrowedMult__comb;
  wire [16:0] p1_smul_57758_NarrowedMult__comb;
  wire [16:0] p1_smul_57760_NarrowedMult__comb;
  wire [16:0] p1_smul_57762_NarrowedMult__comb;
  wire [16:0] p1_smul_57764_NarrowedMult__comb;
  wire [16:0] p1_smul_57766_NarrowedMult__comb;
  wire [16:0] p1_smul_57768_NarrowedMult__comb;
  wire [16:0] p1_smul_57770_NarrowedMult__comb;
  wire [16:0] p1_smul_57772_NarrowedMult__comb;
  wire [16:0] p1_smul_57774_NarrowedMult__comb;
  wire [16:0] p1_smul_57776_NarrowedMult__comb;
  wire [16:0] p1_smul_57778_NarrowedMult__comb;
  wire [16:0] p1_smul_57780_NarrowedMult__comb;
  wire [16:0] p1_smul_57782_NarrowedMult__comb;
  wire [16:0] p1_smul_57784_NarrowedMult__comb;
  wire [16:0] p1_smul_57786_NarrowedMult__comb;
  wire [16:0] p1_smul_57788_NarrowedMult__comb;
  wire [16:0] p1_smul_57806_NarrowedMult__comb;
  wire [16:0] p1_smul_57808_NarrowedMult__comb;
  wire [16:0] p1_smul_57810_NarrowedMult__comb;
  wire [16:0] p1_smul_57812_NarrowedMult__comb;
  wire [16:0] p1_smul_57814_NarrowedMult__comb;
  wire [16:0] p1_smul_57816_NarrowedMult__comb;
  wire [16:0] p1_smul_57818_NarrowedMult__comb;
  wire [16:0] p1_smul_57820_NarrowedMult__comb;
  wire [16:0] p1_smul_57822_NarrowedMult__comb;
  wire [16:0] p1_smul_57824_NarrowedMult__comb;
  wire [16:0] p1_smul_57826_NarrowedMult__comb;
  wire [16:0] p1_smul_57828_NarrowedMult__comb;
  wire [16:0] p1_smul_57830_NarrowedMult__comb;
  wire [16:0] p1_smul_57832_NarrowedMult__comb;
  wire [16:0] p1_smul_57834_NarrowedMult__comb;
  wire [16:0] p1_smul_57836_NarrowedMult__comb;
  wire [16:0] p1_smul_57840_NarrowedMult__comb;
  wire [31:0] p1_or_137776_comb;
  wire [16:0] p1_smul_57844_NarrowedMult__comb;
  wire [16:0] p1_smul_57846_NarrowedMult__comb;
  wire [31:0] p1_or_137781_comb;
  wire [16:0] p1_smul_57850_NarrowedMult__comb;
  wire [16:0] p1_smul_57856_NarrowedMult__comb;
  wire [31:0] p1_or_137792_comb;
  wire [16:0] p1_smul_57860_NarrowedMult__comb;
  wire [16:0] p1_smul_57862_NarrowedMult__comb;
  wire [31:0] p1_or_137797_comb;
  wire [16:0] p1_smul_57866_NarrowedMult__comb;
  wire [16:0] p1_smul_57888_NarrowedMult__comb;
  wire [31:0] p1_or_137808_comb;
  wire [16:0] p1_smul_57892_NarrowedMult__comb;
  wire [16:0] p1_smul_57894_NarrowedMult__comb;
  wire [31:0] p1_or_137813_comb;
  wire [16:0] p1_smul_57898_NarrowedMult__comb;
  wire [16:0] p1_smul_57904_NarrowedMult__comb;
  wire [31:0] p1_or_137824_comb;
  wire [16:0] p1_smul_57908_NarrowedMult__comb;
  wire [16:0] p1_smul_57910_NarrowedMult__comb;
  wire [31:0] p1_or_137829_comb;
  wire [16:0] p1_smul_57914_NarrowedMult__comb;
  wire [16:0] p1_smul_57936_NarrowedMult__comb;
  wire [31:0] p1_or_137840_comb;
  wire [16:0] p1_smul_57940_NarrowedMult__comb;
  wire [16:0] p1_smul_57942_NarrowedMult__comb;
  wire [31:0] p1_or_137845_comb;
  wire [16:0] p1_smul_57946_NarrowedMult__comb;
  wire [16:0] p1_smul_57952_NarrowedMult__comb;
  wire [31:0] p1_or_137856_comb;
  wire [16:0] p1_smul_57956_NarrowedMult__comb;
  wire [16:0] p1_smul_57958_NarrowedMult__comb;
  wire [31:0] p1_or_137861_comb;
  wire [16:0] p1_smul_57962_NarrowedMult__comb;
  wire [31:0] p1_or_137987_comb;
  wire [16:0] p1_smul_58098_NarrowedMult__comb;
  wire [16:0] p1_smul_58100_NarrowedMult__comb;
  wire [16:0] p1_smul_58102_NarrowedMult__comb;
  wire [16:0] p1_smul_58104_NarrowedMult__comb;
  wire [31:0] p1_or_138002_comb;
  wire [31:0] p1_or_138003_comb;
  wire [16:0] p1_smul_58114_NarrowedMult__comb;
  wire [16:0] p1_smul_58116_NarrowedMult__comb;
  wire [16:0] p1_smul_58118_NarrowedMult__comb;
  wire [16:0] p1_smul_58120_NarrowedMult__comb;
  wire [31:0] p1_or_138018_comb;
  wire [31:0] p1_or_138019_comb;
  wire [16:0] p1_smul_58146_NarrowedMult__comb;
  wire [16:0] p1_smul_58148_NarrowedMult__comb;
  wire [16:0] p1_smul_58150_NarrowedMult__comb;
  wire [16:0] p1_smul_58152_NarrowedMult__comb;
  wire [31:0] p1_or_138034_comb;
  wire [31:0] p1_or_138035_comb;
  wire [16:0] p1_smul_58162_NarrowedMult__comb;
  wire [16:0] p1_smul_58164_NarrowedMult__comb;
  wire [16:0] p1_smul_58166_NarrowedMult__comb;
  wire [16:0] p1_smul_58168_NarrowedMult__comb;
  wire [31:0] p1_or_138050_comb;
  wire [31:0] p1_or_138051_comb;
  wire [16:0] p1_smul_58194_NarrowedMult__comb;
  wire [16:0] p1_smul_58196_NarrowedMult__comb;
  wire [16:0] p1_smul_58198_NarrowedMult__comb;
  wire [16:0] p1_smul_58200_NarrowedMult__comb;
  wire [31:0] p1_or_138066_comb;
  wire [31:0] p1_or_138067_comb;
  wire [16:0] p1_smul_58210_NarrowedMult__comb;
  wire [16:0] p1_smul_58212_NarrowedMult__comb;
  wire [16:0] p1_smul_58214_NarrowedMult__comb;
  wire [16:0] p1_smul_58216_NarrowedMult__comb;
  wire [31:0] p1_or_138082_comb;
  wire [15:0] p1_sel_138083_comb;
  wire [15:0] p1_sel_138084_comb;
  wire [15:0] p1_sel_138085_comb;
  wire [15:0] p1_sel_138086_comb;
  wire [15:0] p1_sel_138087_comb;
  wire [15:0] p1_sel_138088_comb;
  wire [15:0] p1_sel_138089_comb;
  wire [15:0] p1_sel_138090_comb;
  wire [15:0] p1_sel_138091_comb;
  wire [15:0] p1_sel_138092_comb;
  wire [15:0] p1_sel_138093_comb;
  wire [15:0] p1_sel_138094_comb;
  wire [15:0] p1_sel_138095_comb;
  wire [15:0] p1_sel_138096_comb;
  wire [15:0] p1_sel_138097_comb;
  wire [15:0] p1_sel_138098_comb;
  wire [15:0] p1_sel_138547_comb;
  wire [15:0] p1_sel_138548_comb;
  wire [15:0] p1_sel_138549_comb;
  wire [15:0] p1_sel_138550_comb;
  wire [15:0] p1_sel_138551_comb;
  wire [15:0] p1_sel_138552_comb;
  wire [15:0] p1_sel_138553_comb;
  wire [15:0] p1_sel_138554_comb;
  wire [15:0] p1_sel_138555_comb;
  wire [15:0] p1_sel_138556_comb;
  wire [15:0] p1_sel_138557_comb;
  wire [15:0] p1_sel_138558_comb;
  wire [15:0] p1_sel_138559_comb;
  wire [15:0] p1_sel_138560_comb;
  wire [15:0] p1_sel_138561_comb;
  wire [15:0] p1_sel_138562_comb;
  wire [15:0] p1_sel_138563_comb;
  wire [15:0] p1_sel_138564_comb;
  wire [15:0] p1_sel_138565_comb;
  wire [15:0] p1_sel_138566_comb;
  wire [15:0] p1_sel_138567_comb;
  wire [15:0] p1_sel_138568_comb;
  wire [15:0] p1_sel_138569_comb;
  wire [15:0] p1_sel_138570_comb;
  wire [15:0] p1_sel_138571_comb;
  wire [15:0] p1_sel_138572_comb;
  wire [15:0] p1_sel_138573_comb;
  wire [15:0] p1_sel_138574_comb;
  wire [15:0] p1_sel_138575_comb;
  wire [15:0] p1_sel_138576_comb;
  wire [15:0] p1_sel_138577_comb;
  wire [15:0] p1_sel_138578_comb;
  wire [15:0] p1_sel_138579_comb;
  wire [15:0] p1_sel_138580_comb;
  wire [15:0] p1_sel_138581_comb;
  wire [15:0] p1_sel_138582_comb;
  wire [15:0] p1_sel_138583_comb;
  wire [15:0] p1_sel_138584_comb;
  wire [15:0] p1_sel_138585_comb;
  wire [15:0] p1_sel_138586_comb;
  wire [15:0] p1_sel_138587_comb;
  wire [15:0] p1_sel_138588_comb;
  wire [15:0] p1_sel_138589_comb;
  wire [15:0] p1_sel_138590_comb;
  wire [15:0] p1_sel_138591_comb;
  wire [15:0] p1_sel_138592_comb;
  wire [15:0] p1_sel_138593_comb;
  wire [15:0] p1_sel_138594_comb;
  wire [16:0] p1_add_141347_comb;
  wire [16:0] p1_add_141348_comb;
  wire [16:0] p1_add_141349_comb;
  wire [16:0] p1_add_141350_comb;
  wire [16:0] p1_add_141351_comb;
  wire [16:0] p1_add_141352_comb;
  wire [16:0] p1_add_141353_comb;
  wire [16:0] p1_add_141354_comb;
  wire [15:0] p1_sel_141355_comb;
  wire [15:0] p1_sel_141356_comb;
  wire [15:0] p1_sel_141357_comb;
  wire [15:0] p1_sel_141358_comb;
  wire [15:0] p1_sel_141359_comb;
  wire [15:0] p1_sel_141360_comb;
  wire [15:0] p1_sel_141361_comb;
  wire [15:0] p1_sel_141362_comb;
  wire [15:0] p1_sel_141363_comb;
  wire [15:0] p1_sel_141364_comb;
  wire [15:0] p1_sel_141365_comb;
  wire [15:0] p1_sel_141366_comb;
  wire [15:0] p1_sel_141367_comb;
  wire [15:0] p1_sel_141368_comb;
  wire [15:0] p1_sel_141369_comb;
  wire [15:0] p1_sel_141370_comb;
  wire [15:0] p1_sel_141371_comb;
  wire [15:0] p1_sel_141372_comb;
  wire [15:0] p1_sel_141373_comb;
  wire [15:0] p1_sel_141374_comb;
  wire [15:0] p1_sel_141375_comb;
  wire [15:0] p1_sel_141376_comb;
  wire [15:0] p1_sel_141377_comb;
  wire [15:0] p1_sel_141378_comb;
  wire [15:0] p1_sel_141379_comb;
  wire [15:0] p1_sel_141380_comb;
  wire [15:0] p1_sel_141381_comb;
  wire [15:0] p1_sel_141382_comb;
  wire [15:0] p1_sel_141383_comb;
  wire [15:0] p1_sel_141384_comb;
  wire [15:0] p1_sel_141385_comb;
  wire [15:0] p1_sel_141386_comb;
  wire [15:0] p1_sel_141387_comb;
  wire [15:0] p1_sel_141388_comb;
  wire [15:0] p1_sel_141389_comb;
  wire [15:0] p1_sel_141390_comb;
  wire [15:0] p1_sel_141391_comb;
  wire [15:0] p1_sel_141392_comb;
  wire [15:0] p1_sel_141393_comb;
  wire [15:0] p1_sel_141394_comb;
  wire [15:0] p1_sel_141395_comb;
  wire [15:0] p1_sel_141396_comb;
  wire [15:0] p1_sel_141397_comb;
  wire [15:0] p1_sel_141398_comb;
  wire [15:0] p1_sel_141399_comb;
  wire [15:0] p1_sel_141400_comb;
  wire [15:0] p1_sel_141401_comb;
  wire [15:0] p1_sel_141402_comb;
  wire [15:0] p1_sel_141403_comb;
  wire [15:0] p1_sel_141404_comb;
  wire [15:0] p1_sel_141405_comb;
  wire [15:0] p1_sel_141406_comb;
  wire [15:0] p1_sel_141407_comb;
  wire [15:0] p1_sel_141408_comb;
  wire [15:0] p1_sel_141409_comb;
  wire [15:0] p1_sel_141410_comb;
  wire [15:0] p1_sel_141411_comb;
  wire [15:0] p1_sel_141412_comb;
  wire [15:0] p1_sel_141413_comb;
  wire [15:0] p1_sel_141414_comb;
  wire [15:0] p1_sel_141415_comb;
  wire [15:0] p1_sel_141416_comb;
  wire [15:0] p1_sel_141417_comb;
  wire [15:0] p1_sel_141418_comb;
  wire [15:0] p1_sel_141419_comb;
  wire [15:0] p1_sel_141420_comb;
  wire [15:0] p1_sel_141421_comb;
  wire [15:0] p1_sel_141422_comb;
  wire [15:0] p1_sel_141423_comb;
  wire [15:0] p1_sel_141424_comb;
  wire [15:0] p1_sel_141425_comb;
  wire [15:0] p1_sel_141426_comb;
  wire [15:0] p1_sel_141427_comb;
  wire [15:0] p1_sel_141428_comb;
  wire [15:0] p1_sel_141429_comb;
  wire [15:0] p1_sel_141430_comb;
  wire [15:0] p1_sel_141431_comb;
  wire [15:0] p1_sel_141432_comb;
  wire [15:0] p1_sel_141433_comb;
  wire [15:0] p1_sel_141434_comb;
  wire [15:0] p1_sel_141435_comb;
  wire [15:0] p1_sel_141436_comb;
  wire [15:0] p1_sel_141437_comb;
  wire [15:0] p1_sel_141438_comb;
  wire [15:0] p1_sel_141439_comb;
  wire [15:0] p1_sel_141440_comb;
  wire [15:0] p1_sel_141441_comb;
  wire [15:0] p1_sel_141442_comb;
  wire [15:0] p1_sel_141443_comb;
  wire [15:0] p1_sel_141444_comb;
  wire [15:0] p1_sel_141445_comb;
  wire [15:0] p1_sel_141446_comb;
  wire [15:0] p1_sel_141447_comb;
  wire [15:0] p1_sel_141448_comb;
  wire [15:0] p1_sel_141449_comb;
  wire [15:0] p1_sel_141450_comb;
  wire [15:0] p1_sel_141451_comb;
  wire [15:0] p1_sel_141452_comb;
  wire [15:0] p1_sel_141453_comb;
  wire [15:0] p1_sel_141454_comb;
  wire [15:0] p1_sel_141455_comb;
  wire [15:0] p1_sel_141456_comb;
  wire [15:0] p1_sel_141457_comb;
  wire [15:0] p1_sel_141458_comb;
  wire [15:0] p1_sel_141459_comb;
  wire [15:0] p1_sel_141460_comb;
  wire [15:0] p1_sel_141461_comb;
  wire [15:0] p1_sel_141462_comb;
  wire [15:0] p1_sel_141463_comb;
  wire [15:0] p1_sel_141464_comb;
  wire [15:0] p1_sel_141465_comb;
  wire [15:0] p1_sel_141466_comb;
  wire [16:0] p1_add_141467_comb;
  wire [16:0] p1_add_141468_comb;
  wire [16:0] p1_add_141469_comb;
  wire [16:0] p1_add_141470_comb;
  wire [16:0] p1_add_141471_comb;
  wire [16:0] p1_add_141472_comb;
  wire [16:0] p1_add_141473_comb;
  wire [16:0] p1_add_141474_comb;
  wire [16:0] p1_add_141475_comb;
  wire [16:0] p1_add_141476_comb;
  wire [16:0] p1_add_141477_comb;
  wire [16:0] p1_add_141478_comb;
  wire [16:0] p1_add_141479_comb;
  wire [16:0] p1_add_141480_comb;
  wire [16:0] p1_add_141481_comb;
  wire [16:0] p1_add_141482_comb;
  wire [16:0] p1_add_141483_comb;
  wire [16:0] p1_add_141484_comb;
  wire [16:0] p1_add_141485_comb;
  wire [16:0] p1_add_141486_comb;
  wire [16:0] p1_add_141487_comb;
  wire [16:0] p1_add_141488_comb;
  wire [16:0] p1_add_141489_comb;
  wire [16:0] p1_add_141490_comb;
  wire [15:0] p1_sel_141491_comb;
  wire [15:0] p1_sel_141492_comb;
  wire [15:0] p1_sel_141493_comb;
  wire [15:0] p1_sel_141494_comb;
  wire [15:0] p1_sel_141495_comb;
  wire [15:0] p1_sel_141496_comb;
  wire [15:0] p1_sel_141497_comb;
  wire [15:0] p1_sel_141498_comb;
  wire [15:0] p1_sel_141499_comb;
  wire [15:0] p1_sel_141500_comb;
  wire [15:0] p1_sel_141501_comb;
  wire [15:0] p1_sel_141502_comb;
  wire [15:0] p1_sel_141503_comb;
  wire [15:0] p1_sel_141504_comb;
  wire [15:0] p1_sel_141505_comb;
  wire [15:0] p1_sel_141506_comb;
  wire [15:0] p1_sel_141507_comb;
  wire [15:0] p1_sel_141508_comb;
  wire [15:0] p1_sel_141509_comb;
  wire [15:0] p1_sel_141510_comb;
  wire [15:0] p1_sel_141511_comb;
  wire [15:0] p1_sel_141512_comb;
  wire [15:0] p1_sel_141513_comb;
  wire [15:0] p1_sel_141514_comb;
  wire [15:0] p1_sel_141515_comb;
  wire [15:0] p1_sel_141516_comb;
  wire [15:0] p1_sel_141517_comb;
  wire [15:0] p1_sel_141518_comb;
  wire [15:0] p1_sel_141519_comb;
  wire [15:0] p1_sel_141520_comb;
  wire [15:0] p1_sel_141521_comb;
  wire [15:0] p1_sel_141522_comb;
  wire [15:0] p1_sel_141523_comb;
  wire [15:0] p1_sel_141524_comb;
  wire [15:0] p1_sel_141525_comb;
  wire [15:0] p1_sel_141526_comb;
  wire [15:0] p1_sel_141527_comb;
  wire [15:0] p1_sel_141528_comb;
  wire [15:0] p1_sel_141529_comb;
  wire [15:0] p1_sel_141530_comb;
  wire [15:0] p1_sel_141531_comb;
  wire [15:0] p1_sel_141532_comb;
  wire [15:0] p1_sel_141533_comb;
  wire [15:0] p1_sel_141534_comb;
  wire [15:0] p1_sel_141535_comb;
  wire [15:0] p1_sel_141536_comb;
  wire [15:0] p1_sel_141537_comb;
  wire [15:0] p1_sel_141538_comb;
  wire [15:0] p1_sel_141539_comb;
  wire [15:0] p1_sel_141540_comb;
  wire [15:0] p1_sel_141541_comb;
  wire [15:0] p1_sel_141542_comb;
  wire [15:0] p1_sel_141543_comb;
  wire [15:0] p1_sel_141544_comb;
  wire [15:0] p1_sel_141545_comb;
  wire [15:0] p1_sel_141546_comb;
  wire [15:0] p1_sel_141547_comb;
  wire [15:0] p1_sel_141548_comb;
  wire [15:0] p1_sel_141549_comb;
  wire [15:0] p1_sel_141550_comb;
  wire [15:0] p1_sel_141551_comb;
  wire [15:0] p1_sel_141552_comb;
  wire [15:0] p1_sel_141553_comb;
  wire [15:0] p1_sel_141554_comb;
  wire [15:0] p1_sel_141555_comb;
  wire [15:0] p1_sel_141556_comb;
  wire [15:0] p1_sel_141557_comb;
  wire [15:0] p1_sel_141558_comb;
  wire [15:0] p1_sel_141559_comb;
  wire [15:0] p1_sel_141560_comb;
  wire [15:0] p1_sel_141561_comb;
  wire [15:0] p1_sel_141562_comb;
  wire [15:0] p1_sel_141563_comb;
  wire [15:0] p1_sel_141564_comb;
  wire [15:0] p1_sel_141565_comb;
  wire [15:0] p1_sel_141566_comb;
  wire [15:0] p1_sel_141567_comb;
  wire [15:0] p1_sel_141568_comb;
  wire [15:0] p1_sel_141569_comb;
  wire [15:0] p1_sel_141570_comb;
  wire [15:0] p1_sel_141571_comb;
  wire [15:0] p1_sel_141572_comb;
  wire [15:0] p1_sel_141573_comb;
  wire [15:0] p1_sel_141574_comb;
  wire [15:0] p1_sel_141575_comb;
  wire [15:0] p1_sel_141576_comb;
  wire [15:0] p1_sel_141577_comb;
  wire [15:0] p1_sel_141578_comb;
  wire [15:0] p1_sel_141579_comb;
  wire [15:0] p1_sel_141580_comb;
  wire [15:0] p1_sel_141581_comb;
  wire [15:0] p1_sel_141582_comb;
  wire [15:0] p1_sel_141583_comb;
  wire [15:0] p1_sel_141584_comb;
  wire [15:0] p1_sel_141585_comb;
  wire [15:0] p1_sel_141586_comb;
  wire [15:0] p1_sel_141587_comb;
  wire [15:0] p1_sel_141588_comb;
  wire [15:0] p1_sel_141589_comb;
  wire [15:0] p1_sel_141590_comb;
  wire [15:0] p1_sel_141591_comb;
  wire [15:0] p1_sel_141592_comb;
  wire [15:0] p1_sel_141593_comb;
  wire [15:0] p1_sel_141594_comb;
  wire [15:0] p1_sel_141595_comb;
  wire [15:0] p1_sel_141596_comb;
  wire [15:0] p1_sel_141597_comb;
  wire [15:0] p1_sel_141598_comb;
  wire [15:0] p1_sel_141599_comb;
  wire [15:0] p1_sel_141600_comb;
  wire [15:0] p1_sel_141601_comb;
  wire [15:0] p1_sel_141602_comb;
  wire [15:0] p1_sel_141603_comb;
  wire [15:0] p1_sel_141604_comb;
  wire [15:0] p1_sel_141605_comb;
  wire [15:0] p1_sel_141606_comb;
  wire [15:0] p1_sel_141607_comb;
  wire [15:0] p1_sel_141608_comb;
  wire [15:0] p1_sel_141609_comb;
  wire [15:0] p1_sel_141610_comb;
  wire [15:0] p1_sel_141611_comb;
  wire [15:0] p1_sel_141612_comb;
  wire [15:0] p1_sel_141613_comb;
  wire [15:0] p1_sel_141614_comb;
  wire [15:0] p1_sel_141615_comb;
  wire [15:0] p1_sel_141616_comb;
  wire [15:0] p1_sel_141617_comb;
  wire [15:0] p1_sel_141618_comb;
  wire [15:0] p1_sel_141619_comb;
  wire [15:0] p1_sel_141620_comb;
  wire [15:0] p1_sel_141621_comb;
  wire [15:0] p1_sel_141622_comb;
  wire [15:0] p1_sel_141623_comb;
  wire [15:0] p1_sel_141624_comb;
  wire [15:0] p1_sel_141625_comb;
  wire [15:0] p1_sel_141626_comb;
  wire [15:0] p1_sel_141627_comb;
  wire [15:0] p1_sel_141628_comb;
  wire [15:0] p1_sel_141629_comb;
  wire [15:0] p1_sel_141630_comb;
  wire [15:0] p1_sel_141631_comb;
  wire [15:0] p1_sel_141632_comb;
  wire [15:0] p1_sel_141633_comb;
  wire [15:0] p1_sel_141634_comb;
  wire [15:0] p1_sel_141635_comb;
  wire [15:0] p1_sel_141636_comb;
  wire [15:0] p1_sel_141637_comb;
  wire [15:0] p1_sel_141638_comb;
  wire [15:0] p1_sel_141639_comb;
  wire [15:0] p1_sel_141640_comb;
  wire [15:0] p1_sel_141641_comb;
  wire [15:0] p1_sel_141642_comb;
  wire [15:0] p1_sel_141643_comb;
  wire [15:0] p1_sel_141644_comb;
  wire [15:0] p1_sel_141645_comb;
  wire [15:0] p1_sel_141646_comb;
  wire [15:0] p1_sel_141647_comb;
  wire [15:0] p1_sel_141648_comb;
  wire [15:0] p1_sel_141649_comb;
  wire [15:0] p1_sel_141650_comb;
  wire [15:0] p1_sel_141651_comb;
  wire [15:0] p1_sel_141652_comb;
  wire [15:0] p1_sel_141653_comb;
  wire [15:0] p1_sel_141654_comb;
  wire [15:0] p1_sel_141655_comb;
  wire [15:0] p1_sel_141656_comb;
  wire [15:0] p1_sel_141657_comb;
  wire [15:0] p1_sel_141658_comb;
  wire [15:0] p1_sel_141659_comb;
  wire [15:0] p1_sel_141660_comb;
  wire [15:0] p1_sel_141661_comb;
  wire [15:0] p1_sel_141662_comb;
  wire [15:0] p1_sel_141663_comb;
  wire [15:0] p1_sel_141664_comb;
  wire [15:0] p1_sel_141665_comb;
  wire [15:0] p1_sel_141666_comb;
  wire [15:0] p1_sel_141667_comb;
  wire [15:0] p1_sel_141668_comb;
  wire [15:0] p1_sel_141669_comb;
  wire [15:0] p1_sel_141670_comb;
  wire [15:0] p1_sel_141671_comb;
  wire [15:0] p1_sel_141672_comb;
  wire [15:0] p1_sel_141673_comb;
  wire [15:0] p1_sel_141674_comb;
  wire [15:0] p1_sel_141675_comb;
  wire [15:0] p1_sel_141676_comb;
  wire [15:0] p1_sel_141677_comb;
  wire [15:0] p1_sel_141678_comb;
  wire [15:0] p1_sel_141679_comb;
  wire [15:0] p1_sel_141680_comb;
  wire [15:0] p1_sel_141681_comb;
  wire [15:0] p1_sel_141682_comb;
  wire [15:0] p1_sel_141683_comb;
  wire [15:0] p1_sel_141684_comb;
  wire [15:0] p1_sel_141685_comb;
  wire [15:0] p1_sel_141686_comb;
  wire [15:0] p1_sel_141687_comb;
  wire [15:0] p1_sel_141688_comb;
  wire [15:0] p1_sel_141689_comb;
  wire [15:0] p1_sel_141690_comb;
  wire [15:0] p1_sel_141691_comb;
  wire [15:0] p1_sel_141692_comb;
  wire [15:0] p1_sel_141693_comb;
  wire [15:0] p1_sel_141694_comb;
  wire [15:0] p1_sel_141695_comb;
  wire [15:0] p1_sel_141696_comb;
  wire [15:0] p1_sel_141697_comb;
  wire [15:0] p1_sel_141698_comb;
  wire [15:0] p1_sel_141699_comb;
  wire [15:0] p1_sel_141700_comb;
  wire [15:0] p1_sel_141701_comb;
  wire [15:0] p1_sel_141702_comb;
  wire [15:0] p1_sel_141703_comb;
  wire [15:0] p1_sel_141704_comb;
  wire [15:0] p1_sel_141705_comb;
  wire [15:0] p1_sel_141706_comb;
  wire [15:0] p1_sel_141707_comb;
  wire [15:0] p1_sel_141708_comb;
  wire [15:0] p1_sel_141709_comb;
  wire [15:0] p1_sel_141710_comb;
  wire [15:0] p1_sel_141711_comb;
  wire [15:0] p1_sel_141712_comb;
  wire [15:0] p1_sel_141713_comb;
  wire [15:0] p1_sel_141714_comb;
  wire [15:0] p1_sel_141715_comb;
  wire [15:0] p1_sel_141716_comb;
  wire [15:0] p1_sel_141717_comb;
  wire [15:0] p1_sel_141718_comb;
  wire [15:0] p1_sel_141719_comb;
  wire [15:0] p1_sel_141720_comb;
  wire [15:0] p1_sel_141721_comb;
  wire [15:0] p1_sel_141722_comb;
  wire [15:0] p1_sel_141723_comb;
  wire [15:0] p1_sel_141724_comb;
  wire [15:0] p1_sel_141725_comb;
  wire [15:0] p1_sel_141726_comb;
  wire [15:0] p1_sel_141727_comb;
  wire [15:0] p1_sel_141728_comb;
  wire [15:0] p1_sel_141729_comb;
  wire [15:0] p1_sel_141730_comb;
  wire [15:0] p1_sel_141731_comb;
  wire [15:0] p1_sel_141732_comb;
  wire [15:0] p1_sel_141733_comb;
  wire [15:0] p1_sel_141734_comb;
  wire [15:0] p1_sel_141735_comb;
  wire [15:0] p1_sel_141736_comb;
  wire [15:0] p1_sel_141737_comb;
  wire [15:0] p1_sel_141738_comb;
  wire [15:0] p1_sel_141739_comb;
  wire [15:0] p1_sel_141740_comb;
  wire [15:0] p1_sel_141741_comb;
  wire [15:0] p1_sel_141742_comb;
  wire [15:0] p1_sel_141743_comb;
  wire [15:0] p1_sel_141744_comb;
  wire [15:0] p1_sel_141745_comb;
  wire [15:0] p1_sel_141746_comb;
  wire [15:0] p1_sel_141747_comb;
  wire [15:0] p1_sel_141748_comb;
  wire [15:0] p1_sel_141749_comb;
  wire [15:0] p1_sel_141750_comb;
  wire [15:0] p1_sel_141751_comb;
  wire [15:0] p1_sel_141752_comb;
  wire [15:0] p1_sel_141753_comb;
  wire [15:0] p1_sel_141754_comb;
  wire [15:0] p1_sel_141755_comb;
  wire [15:0] p1_sel_141756_comb;
  wire [15:0] p1_sel_141757_comb;
  wire [15:0] p1_sel_141758_comb;
  wire [15:0] p1_sel_141759_comb;
  wire [15:0] p1_sel_141760_comb;
  wire [15:0] p1_sel_141761_comb;
  wire [15:0] p1_sel_141762_comb;
  wire [15:0] p1_sel_141763_comb;
  wire [15:0] p1_sel_141764_comb;
  wire [15:0] p1_sel_141765_comb;
  wire [15:0] p1_sel_141766_comb;
  wire [15:0] p1_sel_141767_comb;
  wire [15:0] p1_sel_141768_comb;
  wire [15:0] p1_sel_141769_comb;
  wire [15:0] p1_sel_141770_comb;
  wire [15:0] p1_sel_141771_comb;
  wire [15:0] p1_sel_141772_comb;
  wire [15:0] p1_sel_141773_comb;
  wire [15:0] p1_sel_141774_comb;
  wire [15:0] p1_sel_141775_comb;
  wire [15:0] p1_sel_141776_comb;
  wire [15:0] p1_sel_141777_comb;
  wire [15:0] p1_sel_141778_comb;
  wire [15:0] p1_sel_141779_comb;
  wire [15:0] p1_sel_141780_comb;
  wire [15:0] p1_sel_141781_comb;
  wire [15:0] p1_sel_141782_comb;
  wire [15:0] p1_sel_141783_comb;
  wire [15:0] p1_sel_141784_comb;
  wire [15:0] p1_sel_141785_comb;
  wire [15:0] p1_sel_141786_comb;
  wire [15:0] p1_sel_141787_comb;
  wire [15:0] p1_sel_141788_comb;
  wire [15:0] p1_sel_141789_comb;
  wire [15:0] p1_sel_141790_comb;
  wire [15:0] p1_sel_141791_comb;
  wire [15:0] p1_sel_141792_comb;
  wire [15:0] p1_sel_141793_comb;
  wire [15:0] p1_sel_141794_comb;
  wire [15:0] p1_sel_141795_comb;
  wire [15:0] p1_sel_141796_comb;
  wire [15:0] p1_sel_141797_comb;
  wire [15:0] p1_sel_141798_comb;
  wire [15:0] p1_sel_141799_comb;
  wire [15:0] p1_sel_141800_comb;
  wire [15:0] p1_sel_141801_comb;
  wire [15:0] p1_sel_141802_comb;
  wire [15:0] p1_sel_141803_comb;
  wire [15:0] p1_sel_141804_comb;
  wire [15:0] p1_sel_141805_comb;
  wire [15:0] p1_sel_141806_comb;
  wire [15:0] p1_sel_141807_comb;
  wire [15:0] p1_sel_141808_comb;
  wire [15:0] p1_sel_141809_comb;
  wire [15:0] p1_sel_141810_comb;
  wire [15:0] p1_sel_141811_comb;
  wire [15:0] p1_sel_141812_comb;
  wire [15:0] p1_sel_141813_comb;
  wire [15:0] p1_sel_141814_comb;
  wire [15:0] p1_sel_141815_comb;
  wire [15:0] p1_sel_141816_comb;
  wire [15:0] p1_sel_141817_comb;
  wire [15:0] p1_sel_141818_comb;
  wire [15:0] p1_sel_141819_comb;
  wire [15:0] p1_sel_141820_comb;
  wire [15:0] p1_sel_141821_comb;
  wire [15:0] p1_sel_141822_comb;
  wire [15:0] p1_sel_141823_comb;
  wire [15:0] p1_sel_141824_comb;
  wire [15:0] p1_sel_141825_comb;
  wire [15:0] p1_sel_141826_comb;
  wire [31:0] p1_sum__989_comb;
  wire [31:0] p1_sum__990_comb;
  wire [31:0] p1_sum__991_comb;
  wire [31:0] p1_sum__992_comb;
  wire [31:0] p1_sum__884_comb;
  wire [31:0] p1_sum__885_comb;
  wire [31:0] p1_sum__886_comb;
  wire [31:0] p1_sum__887_comb;
  wire [31:0] p1_sum__1017_comb;
  wire [31:0] p1_sum__1018_comb;
  wire [31:0] p1_sum__1019_comb;
  wire [31:0] p1_sum__1020_comb;
  wire [31:0] p1_sum__1010_comb;
  wire [31:0] p1_sum__1011_comb;
  wire [31:0] p1_sum__1012_comb;
  wire [31:0] p1_sum__1013_comb;
  wire [31:0] p1_sum__961_comb;
  wire [31:0] p1_sum__962_comb;
  wire [31:0] p1_sum__963_comb;
  wire [31:0] p1_sum__964_comb;
  wire [31:0] p1_sum__926_comb;
  wire [31:0] p1_sum__927_comb;
  wire [31:0] p1_sum__928_comb;
  wire [31:0] p1_sum__929_comb;
  wire [31:0] p1_sum__835_comb;
  wire [31:0] p1_sum__836_comb;
  wire [31:0] p1_sum__837_comb;
  wire [31:0] p1_sum__838_comb;
  wire [31:0] p1_sum__779_comb;
  wire [31:0] p1_sum__780_comb;
  wire [31:0] p1_sum__781_comb;
  wire [31:0] p1_sum__782_comb;
  wire [31:0] p1_sum__993_comb;
  wire [31:0] p1_sum__994_comb;
  wire [31:0] p1_sum__888_comb;
  wire [31:0] p1_sum__889_comb;
  wire [16:0] p1_add_142311_comb;
  wire [16:0] p1_add_142312_comb;
  wire [16:0] p1_add_142313_comb;
  wire [16:0] p1_add_142314_comb;
  wire [16:0] p1_add_142315_comb;
  wire [16:0] p1_add_142316_comb;
  wire [16:0] p1_add_142317_comb;
  wire [16:0] p1_add_142318_comb;
  wire [16:0] p1_add_142319_comb;
  wire [16:0] p1_add_142320_comb;
  wire [16:0] p1_add_142321_comb;
  wire [16:0] p1_add_142322_comb;
  wire [16:0] p1_add_142323_comb;
  wire [16:0] p1_add_142324_comb;
  wire [16:0] p1_add_142325_comb;
  wire [16:0] p1_add_142326_comb;
  wire [16:0] p1_add_142327_comb;
  wire [16:0] p1_add_142328_comb;
  wire [16:0] p1_add_142329_comb;
  wire [16:0] p1_add_142330_comb;
  wire [16:0] p1_add_142331_comb;
  wire [16:0] p1_add_142332_comb;
  wire [16:0] p1_add_142333_comb;
  wire [16:0] p1_add_142334_comb;
  wire [16:0] p1_add_142335_comb;
  wire [16:0] p1_add_142336_comb;
  wire [16:0] p1_add_142337_comb;
  wire [16:0] p1_add_142338_comb;
  wire [16:0] p1_add_142339_comb;
  wire [16:0] p1_add_142340_comb;
  wire [16:0] p1_add_142341_comb;
  wire [16:0] p1_add_142342_comb;
  wire [16:0] p1_add_142343_comb;
  wire [16:0] p1_add_142344_comb;
  wire [16:0] p1_add_142345_comb;
  wire [16:0] p1_add_142346_comb;
  wire [16:0] p1_add_142347_comb;
  wire [16:0] p1_add_142348_comb;
  wire [16:0] p1_add_142349_comb;
  wire [16:0] p1_add_142350_comb;
  wire [16:0] p1_add_142351_comb;
  wire [16:0] p1_add_142352_comb;
  wire [16:0] p1_add_142353_comb;
  wire [16:0] p1_add_142354_comb;
  wire [16:0] p1_add_142355_comb;
  wire [16:0] p1_add_142356_comb;
  wire [16:0] p1_add_142357_comb;
  wire [16:0] p1_add_142358_comb;
  wire [16:0] p1_add_142359_comb;
  wire [16:0] p1_add_142360_comb;
  wire [16:0] p1_add_142361_comb;
  wire [16:0] p1_add_142362_comb;
  wire [16:0] p1_add_142363_comb;
  wire [16:0] p1_add_142364_comb;
  wire [16:0] p1_add_142365_comb;
  wire [16:0] p1_add_142366_comb;
  wire [31:0] p1_sum__1021_comb;
  wire [31:0] p1_sum__1022_comb;
  wire [31:0] p1_sum__1014_comb;
  wire [31:0] p1_sum__1015_comb;
  wire [31:0] p1_sum__965_comb;
  wire [31:0] p1_sum__966_comb;
  wire [31:0] p1_sum__930_comb;
  wire [31:0] p1_sum__931_comb;
  wire [31:0] p1_sum__839_comb;
  wire [31:0] p1_sum__840_comb;
  wire [31:0] p1_sum__783_comb;
  wire [31:0] p1_sum__784_comb;
  wire [16:0] p1_add_142379_comb;
  wire [16:0] p1_add_142380_comb;
  wire [16:0] p1_add_142381_comb;
  wire [16:0] p1_add_142382_comb;
  wire [16:0] p1_add_142383_comb;
  wire [16:0] p1_add_142384_comb;
  wire [16:0] p1_add_142385_comb;
  wire [16:0] p1_add_142386_comb;
  wire [16:0] p1_add_142387_comb;
  wire [16:0] p1_add_142388_comb;
  wire [16:0] p1_add_142389_comb;
  wire [16:0] p1_add_142390_comb;
  wire [16:0] p1_add_142391_comb;
  wire [16:0] p1_add_142392_comb;
  wire [16:0] p1_add_142393_comb;
  wire [16:0] p1_add_142394_comb;
  wire [16:0] p1_add_142395_comb;
  wire [16:0] p1_add_142396_comb;
  wire [16:0] p1_add_142397_comb;
  wire [16:0] p1_add_142398_comb;
  wire [16:0] p1_add_142399_comb;
  wire [16:0] p1_add_142400_comb;
  wire [16:0] p1_add_142401_comb;
  wire [16:0] p1_add_142402_comb;
  wire [16:0] p1_add_142403_comb;
  wire [16:0] p1_add_142404_comb;
  wire [16:0] p1_add_142405_comb;
  wire [16:0] p1_add_142406_comb;
  wire [16:0] p1_add_142407_comb;
  wire [16:0] p1_add_142408_comb;
  wire [16:0] p1_add_142409_comb;
  wire [16:0] p1_add_142410_comb;
  wire [16:0] p1_add_142411_comb;
  wire [16:0] p1_add_142412_comb;
  wire [16:0] p1_add_142413_comb;
  wire [16:0] p1_add_142414_comb;
  wire [16:0] p1_add_142415_comb;
  wire [16:0] p1_add_142416_comb;
  wire [16:0] p1_add_142417_comb;
  wire [16:0] p1_add_142418_comb;
  wire [16:0] p1_add_142419_comb;
  wire [16:0] p1_add_142420_comb;
  wire [16:0] p1_add_142421_comb;
  wire [16:0] p1_add_142422_comb;
  wire [16:0] p1_add_142423_comb;
  wire [16:0] p1_add_142424_comb;
  wire [16:0] p1_add_142425_comb;
  wire [16:0] p1_add_142426_comb;
  wire [16:0] p1_add_142427_comb;
  wire [16:0] p1_add_142428_comb;
  wire [16:0] p1_add_142429_comb;
  wire [16:0] p1_add_142430_comb;
  wire [16:0] p1_add_142431_comb;
  wire [16:0] p1_add_142432_comb;
  wire [16:0] p1_add_142433_comb;
  wire [16:0] p1_add_142434_comb;
  wire [16:0] p1_add_142435_comb;
  wire [16:0] p1_add_142436_comb;
  wire [16:0] p1_add_142437_comb;
  wire [16:0] p1_add_142438_comb;
  wire [16:0] p1_add_142439_comb;
  wire [16:0] p1_add_142440_comb;
  wire [16:0] p1_add_142441_comb;
  wire [16:0] p1_add_142442_comb;
  wire [16:0] p1_add_142443_comb;
  wire [16:0] p1_add_142444_comb;
  wire [16:0] p1_add_142445_comb;
  wire [16:0] p1_add_142446_comb;
  wire [16:0] p1_add_142447_comb;
  wire [16:0] p1_add_142448_comb;
  wire [16:0] p1_add_142449_comb;
  wire [16:0] p1_add_142450_comb;
  wire [16:0] p1_add_142451_comb;
  wire [16:0] p1_add_142452_comb;
  wire [16:0] p1_add_142453_comb;
  wire [16:0] p1_add_142454_comb;
  wire [16:0] p1_add_142455_comb;
  wire [16:0] p1_add_142456_comb;
  wire [16:0] p1_add_142457_comb;
  wire [16:0] p1_add_142458_comb;
  wire [16:0] p1_add_142459_comb;
  wire [16:0] p1_add_142460_comb;
  wire [16:0] p1_add_142461_comb;
  wire [16:0] p1_add_142462_comb;
  wire [16:0] p1_add_142463_comb;
  wire [16:0] p1_add_142464_comb;
  wire [16:0] p1_add_142465_comb;
  wire [16:0] p1_add_142466_comb;
  wire [16:0] p1_add_142467_comb;
  wire [16:0] p1_add_142468_comb;
  wire [16:0] p1_add_142469_comb;
  wire [16:0] p1_add_142470_comb;
  wire [16:0] p1_add_142471_comb;
  wire [16:0] p1_add_142472_comb;
  wire [16:0] p1_add_142473_comb;
  wire [16:0] p1_add_142474_comb;
  wire [16:0] p1_add_142475_comb;
  wire [16:0] p1_add_142476_comb;
  wire [16:0] p1_add_142477_comb;
  wire [16:0] p1_add_142478_comb;
  wire [16:0] p1_add_142479_comb;
  wire [16:0] p1_add_142480_comb;
  wire [16:0] p1_add_142481_comb;
  wire [16:0] p1_add_142482_comb;
  wire [16:0] p1_add_142483_comb;
  wire [16:0] p1_add_142484_comb;
  wire [16:0] p1_add_142485_comb;
  wire [16:0] p1_add_142486_comb;
  wire [16:0] p1_add_142487_comb;
  wire [16:0] p1_add_142488_comb;
  wire [16:0] p1_add_142489_comb;
  wire [16:0] p1_add_142490_comb;
  wire [16:0] p1_add_142491_comb;
  wire [16:0] p1_add_142492_comb;
  wire [16:0] p1_add_142493_comb;
  wire [16:0] p1_add_142494_comb;
  wire [16:0] p1_add_142495_comb;
  wire [16:0] p1_add_142496_comb;
  wire [16:0] p1_add_142497_comb;
  wire [16:0] p1_add_142498_comb;
  wire [16:0] p1_add_142499_comb;
  wire [16:0] p1_add_142500_comb;
  wire [16:0] p1_add_142501_comb;
  wire [16:0] p1_add_142502_comb;
  wire [16:0] p1_add_142503_comb;
  wire [16:0] p1_add_142504_comb;
  wire [16:0] p1_add_142505_comb;
  wire [16:0] p1_add_142506_comb;
  wire [16:0] p1_add_142507_comb;
  wire [16:0] p1_add_142508_comb;
  wire [16:0] p1_add_142509_comb;
  wire [16:0] p1_add_142510_comb;
  wire [16:0] p1_add_142511_comb;
  wire [16:0] p1_add_142512_comb;
  wire [16:0] p1_add_142513_comb;
  wire [16:0] p1_add_142514_comb;
  wire [16:0] p1_add_142515_comb;
  wire [16:0] p1_add_142516_comb;
  wire [16:0] p1_add_142517_comb;
  wire [16:0] p1_add_142518_comb;
  wire [16:0] p1_add_142519_comb;
  wire [16:0] p1_add_142520_comb;
  wire [16:0] p1_add_142521_comb;
  wire [16:0] p1_add_142522_comb;
  wire [16:0] p1_add_142523_comb;
  wire [16:0] p1_add_142524_comb;
  wire [16:0] p1_add_142525_comb;
  wire [16:0] p1_add_142526_comb;
  wire [16:0] p1_add_142527_comb;
  wire [16:0] p1_add_142528_comb;
  wire [16:0] p1_add_142529_comb;
  wire [16:0] p1_add_142530_comb;
  wire [16:0] p1_add_142531_comb;
  wire [16:0] p1_add_142532_comb;
  wire [16:0] p1_add_142533_comb;
  wire [16:0] p1_add_142534_comb;
  wire [16:0] p1_add_142535_comb;
  wire [16:0] p1_add_142536_comb;
  wire [16:0] p1_add_142537_comb;
  wire [16:0] p1_add_142538_comb;
  wire [16:0] p1_add_142539_comb;
  wire [16:0] p1_add_142540_comb;
  wire [16:0] p1_add_142541_comb;
  wire [16:0] p1_add_142542_comb;
  wire [16:0] p1_add_142543_comb;
  wire [16:0] p1_add_142544_comb;
  wire [16:0] p1_add_142545_comb;
  wire [16:0] p1_add_142546_comb;
  wire [31:0] p1_sum__995_comb;
  wire [31:0] p1_sum__890_comb;
  wire [24:0] p1_sum__1784_comb;
  wire [24:0] p1_sum__1785_comb;
  wire [24:0] p1_sum__1786_comb;
  wire [24:0] p1_sum__1787_comb;
  wire [24:0] p1_sum__1724_comb;
  wire [24:0] p1_sum__1725_comb;
  wire [24:0] p1_sum__1726_comb;
  wire [24:0] p1_sum__1727_comb;
  wire [24:0] p1_sum__1772_comb;
  wire [24:0] p1_sum__1773_comb;
  wire [24:0] p1_sum__1774_comb;
  wire [24:0] p1_sum__1775_comb;
  wire [24:0] p1_sum__1700_comb;
  wire [24:0] p1_sum__1701_comb;
  wire [24:0] p1_sum__1702_comb;
  wire [24:0] p1_sum__1703_comb;
  wire [24:0] p1_sum__1756_comb;
  wire [24:0] p1_sum__1757_comb;
  wire [24:0] p1_sum__1758_comb;
  wire [24:0] p1_sum__1759_comb;
  wire [24:0] p1_sum__1676_comb;
  wire [24:0] p1_sum__1677_comb;
  wire [24:0] p1_sum__1678_comb;
  wire [24:0] p1_sum__1679_comb;
  wire [24:0] p1_sum__1736_comb;
  wire [24:0] p1_sum__1737_comb;
  wire [24:0] p1_sum__1738_comb;
  wire [24:0] p1_sum__1739_comb;
  wire [24:0] p1_sum__1652_comb;
  wire [24:0] p1_sum__1653_comb;
  wire [24:0] p1_sum__1654_comb;
  wire [24:0] p1_sum__1655_comb;
  wire [24:0] p1_sum__1712_comb;
  wire [24:0] p1_sum__1713_comb;
  wire [24:0] p1_sum__1714_comb;
  wire [24:0] p1_sum__1715_comb;
  wire [24:0] p1_sum__1632_comb;
  wire [24:0] p1_sum__1633_comb;
  wire [24:0] p1_sum__1634_comb;
  wire [24:0] p1_sum__1635_comb;
  wire [24:0] p1_sum__1688_comb;
  wire [24:0] p1_sum__1689_comb;
  wire [24:0] p1_sum__1690_comb;
  wire [24:0] p1_sum__1691_comb;
  wire [24:0] p1_sum__1616_comb;
  wire [24:0] p1_sum__1617_comb;
  wire [24:0] p1_sum__1618_comb;
  wire [24:0] p1_sum__1619_comb;
  wire [24:0] p1_sum__1664_comb;
  wire [24:0] p1_sum__1665_comb;
  wire [24:0] p1_sum__1666_comb;
  wire [24:0] p1_sum__1667_comb;
  wire [24:0] p1_sum__1604_comb;
  wire [24:0] p1_sum__1605_comb;
  wire [24:0] p1_sum__1606_comb;
  wire [24:0] p1_sum__1607_comb;
  wire [31:0] p1_sum__1023_comb;
  wire [31:0] p1_sum__1016_comb;
  wire [31:0] p1_sum__967_comb;
  wire [31:0] p1_sum__932_comb;
  wire [31:0] p1_sum__841_comb;
  wire [31:0] p1_sum__785_comb;
  wire [24:0] p1_sum__1804_comb;
  wire [24:0] p1_sum__1805_comb;
  wire [24:0] p1_sum__1806_comb;
  wire [24:0] p1_sum__1807_comb;
  wire [24:0] p1_sum__1796_comb;
  wire [24:0] p1_sum__1797_comb;
  wire [24:0] p1_sum__1798_comb;
  wire [24:0] p1_sum__1799_comb;
  wire [24:0] p1_sum__1768_comb;
  wire [24:0] p1_sum__1769_comb;
  wire [24:0] p1_sum__1770_comb;
  wire [24:0] p1_sum__1771_comb;
  wire [24:0] p1_sum__1748_comb;
  wire [24:0] p1_sum__1749_comb;
  wire [24:0] p1_sum__1750_comb;
  wire [24:0] p1_sum__1751_comb;
  wire [24:0] p1_sum__1696_comb;
  wire [24:0] p1_sum__1697_comb;
  wire [24:0] p1_sum__1698_comb;
  wire [24:0] p1_sum__1699_comb;
  wire [24:0] p1_sum__1668_comb;
  wire [24:0] p1_sum__1669_comb;
  wire [24:0] p1_sum__1670_comb;
  wire [24:0] p1_sum__1671_comb;
  wire [24:0] p1_sum__1800_comb;
  wire [24:0] p1_sum__1801_comb;
  wire [24:0] p1_sum__1802_comb;
  wire [24:0] p1_sum__1803_comb;
  wire [24:0] p1_sum__1788_comb;
  wire [24:0] p1_sum__1789_comb;
  wire [24:0] p1_sum__1790_comb;
  wire [24:0] p1_sum__1791_comb;
  wire [24:0] p1_sum__1752_comb;
  wire [24:0] p1_sum__1753_comb;
  wire [24:0] p1_sum__1754_comb;
  wire [24:0] p1_sum__1755_comb;
  wire [24:0] p1_sum__1728_comb;
  wire [24:0] p1_sum__1729_comb;
  wire [24:0] p1_sum__1730_comb;
  wire [24:0] p1_sum__1731_comb;
  wire [24:0] p1_sum__1672_comb;
  wire [24:0] p1_sum__1673_comb;
  wire [24:0] p1_sum__1674_comb;
  wire [24:0] p1_sum__1675_comb;
  wire [24:0] p1_sum__1644_comb;
  wire [24:0] p1_sum__1645_comb;
  wire [24:0] p1_sum__1646_comb;
  wire [24:0] p1_sum__1647_comb;
  wire [24:0] p1_sum__1792_comb;
  wire [24:0] p1_sum__1793_comb;
  wire [24:0] p1_sum__1794_comb;
  wire [24:0] p1_sum__1795_comb;
  wire [24:0] p1_sum__1776_comb;
  wire [24:0] p1_sum__1777_comb;
  wire [24:0] p1_sum__1778_comb;
  wire [24:0] p1_sum__1779_comb;
  wire [24:0] p1_sum__1732_comb;
  wire [24:0] p1_sum__1733_comb;
  wire [24:0] p1_sum__1734_comb;
  wire [24:0] p1_sum__1735_comb;
  wire [24:0] p1_sum__1704_comb;
  wire [24:0] p1_sum__1705_comb;
  wire [24:0] p1_sum__1706_comb;
  wire [24:0] p1_sum__1707_comb;
  wire [24:0] p1_sum__1648_comb;
  wire [24:0] p1_sum__1649_comb;
  wire [24:0] p1_sum__1650_comb;
  wire [24:0] p1_sum__1651_comb;
  wire [24:0] p1_sum__1624_comb;
  wire [24:0] p1_sum__1625_comb;
  wire [24:0] p1_sum__1626_comb;
  wire [24:0] p1_sum__1627_comb;
  wire [24:0] p1_sum__1780_comb;
  wire [24:0] p1_sum__1781_comb;
  wire [24:0] p1_sum__1782_comb;
  wire [24:0] p1_sum__1783_comb;
  wire [24:0] p1_sum__1760_comb;
  wire [24:0] p1_sum__1761_comb;
  wire [24:0] p1_sum__1762_comb;
  wire [24:0] p1_sum__1763_comb;
  wire [24:0] p1_sum__1708_comb;
  wire [24:0] p1_sum__1709_comb;
  wire [24:0] p1_sum__1710_comb;
  wire [24:0] p1_sum__1711_comb;
  wire [24:0] p1_sum__1680_comb;
  wire [24:0] p1_sum__1681_comb;
  wire [24:0] p1_sum__1682_comb;
  wire [24:0] p1_sum__1683_comb;
  wire [24:0] p1_sum__1628_comb;
  wire [24:0] p1_sum__1629_comb;
  wire [24:0] p1_sum__1630_comb;
  wire [24:0] p1_sum__1631_comb;
  wire [24:0] p1_sum__1608_comb;
  wire [24:0] p1_sum__1609_comb;
  wire [24:0] p1_sum__1610_comb;
  wire [24:0] p1_sum__1611_comb;
  wire [24:0] p1_sum__1764_comb;
  wire [24:0] p1_sum__1765_comb;
  wire [24:0] p1_sum__1766_comb;
  wire [24:0] p1_sum__1767_comb;
  wire [24:0] p1_sum__1740_comb;
  wire [24:0] p1_sum__1741_comb;
  wire [24:0] p1_sum__1742_comb;
  wire [24:0] p1_sum__1743_comb;
  wire [24:0] p1_sum__1684_comb;
  wire [24:0] p1_sum__1685_comb;
  wire [24:0] p1_sum__1686_comb;
  wire [24:0] p1_sum__1687_comb;
  wire [24:0] p1_sum__1656_comb;
  wire [24:0] p1_sum__1657_comb;
  wire [24:0] p1_sum__1658_comb;
  wire [24:0] p1_sum__1659_comb;
  wire [24:0] p1_sum__1612_comb;
  wire [24:0] p1_sum__1613_comb;
  wire [24:0] p1_sum__1614_comb;
  wire [24:0] p1_sum__1615_comb;
  wire [24:0] p1_sum__1596_comb;
  wire [24:0] p1_sum__1597_comb;
  wire [24:0] p1_sum__1598_comb;
  wire [24:0] p1_sum__1599_comb;
  wire [24:0] p1_sum__1744_comb;
  wire [24:0] p1_sum__1745_comb;
  wire [24:0] p1_sum__1746_comb;
  wire [24:0] p1_sum__1747_comb;
  wire [24:0] p1_sum__1716_comb;
  wire [24:0] p1_sum__1717_comb;
  wire [24:0] p1_sum__1718_comb;
  wire [24:0] p1_sum__1719_comb;
  wire [24:0] p1_sum__1660_comb;
  wire [24:0] p1_sum__1661_comb;
  wire [24:0] p1_sum__1662_comb;
  wire [24:0] p1_sum__1663_comb;
  wire [24:0] p1_sum__1636_comb;
  wire [24:0] p1_sum__1637_comb;
  wire [24:0] p1_sum__1638_comb;
  wire [24:0] p1_sum__1639_comb;
  wire [24:0] p1_sum__1600_comb;
  wire [24:0] p1_sum__1601_comb;
  wire [24:0] p1_sum__1602_comb;
  wire [24:0] p1_sum__1603_comb;
  wire [24:0] p1_sum__1588_comb;
  wire [24:0] p1_sum__1589_comb;
  wire [24:0] p1_sum__1590_comb;
  wire [24:0] p1_sum__1591_comb;
  wire [24:0] p1_sum__1720_comb;
  wire [24:0] p1_sum__1721_comb;
  wire [24:0] p1_sum__1722_comb;
  wire [24:0] p1_sum__1723_comb;
  wire [24:0] p1_sum__1692_comb;
  wire [24:0] p1_sum__1693_comb;
  wire [24:0] p1_sum__1694_comb;
  wire [24:0] p1_sum__1695_comb;
  wire [24:0] p1_sum__1640_comb;
  wire [24:0] p1_sum__1641_comb;
  wire [24:0] p1_sum__1642_comb;
  wire [24:0] p1_sum__1643_comb;
  wire [24:0] p1_sum__1620_comb;
  wire [24:0] p1_sum__1621_comb;
  wire [24:0] p1_sum__1622_comb;
  wire [24:0] p1_sum__1623_comb;
  wire [24:0] p1_sum__1592_comb;
  wire [24:0] p1_sum__1593_comb;
  wire [24:0] p1_sum__1594_comb;
  wire [24:0] p1_sum__1595_comb;
  wire [24:0] p1_sum__1584_comb;
  wire [24:0] p1_sum__1585_comb;
  wire [24:0] p1_sum__1586_comb;
  wire [24:0] p1_sum__1587_comb;
  wire [31:0] p1_umul_142787_comb;
  wire [31:0] p1_umul_142788_comb;
  wire [24:0] p1_sum__1348_comb;
  wire [24:0] p1_sum__1349_comb;
  wire [24:0] p1_sum__1318_comb;
  wire [24:0] p1_sum__1319_comb;
  wire [24:0] p1_sum__1342_comb;
  wire [24:0] p1_sum__1343_comb;
  wire [24:0] p1_sum__1306_comb;
  wire [24:0] p1_sum__1307_comb;
  wire [24:0] p1_sum__1334_comb;
  wire [24:0] p1_sum__1335_comb;
  wire [24:0] p1_sum__1294_comb;
  wire [24:0] p1_sum__1295_comb;
  wire [24:0] p1_sum__1324_comb;
  wire [24:0] p1_sum__1325_comb;
  wire [24:0] p1_sum__1282_comb;
  wire [24:0] p1_sum__1283_comb;
  wire [24:0] p1_sum__1312_comb;
  wire [24:0] p1_sum__1313_comb;
  wire [24:0] p1_sum__1272_comb;
  wire [24:0] p1_sum__1273_comb;
  wire [24:0] p1_sum__1300_comb;
  wire [24:0] p1_sum__1301_comb;
  wire [24:0] p1_sum__1264_comb;
  wire [24:0] p1_sum__1265_comb;
  wire [24:0] p1_sum__1288_comb;
  wire [24:0] p1_sum__1289_comb;
  wire [24:0] p1_sum__1258_comb;
  wire [24:0] p1_sum__1259_comb;
  wire [31:0] p1_umul_142817_comb;
  wire [31:0] p1_umul_142818_comb;
  wire [31:0] p1_umul_142819_comb;
  wire [31:0] p1_umul_142820_comb;
  wire [31:0] p1_umul_142821_comb;
  wire [31:0] p1_umul_142822_comb;
  wire [24:0] p1_sum__1358_comb;
  wire [24:0] p1_sum__1359_comb;
  wire [24:0] p1_sum__1354_comb;
  wire [24:0] p1_sum__1355_comb;
  wire [24:0] p1_sum__1340_comb;
  wire [24:0] p1_sum__1341_comb;
  wire [24:0] p1_sum__1330_comb;
  wire [24:0] p1_sum__1331_comb;
  wire [24:0] p1_sum__1304_comb;
  wire [24:0] p1_sum__1305_comb;
  wire [24:0] p1_sum__1290_comb;
  wire [24:0] p1_sum__1291_comb;
  wire [24:0] p1_sum__1356_comb;
  wire [24:0] p1_sum__1357_comb;
  wire [24:0] p1_sum__1350_comb;
  wire [24:0] p1_sum__1351_comb;
  wire [24:0] p1_sum__1332_comb;
  wire [24:0] p1_sum__1333_comb;
  wire [24:0] p1_sum__1320_comb;
  wire [24:0] p1_sum__1321_comb;
  wire [24:0] p1_sum__1292_comb;
  wire [24:0] p1_sum__1293_comb;
  wire [24:0] p1_sum__1278_comb;
  wire [24:0] p1_sum__1279_comb;
  wire [24:0] p1_sum__1352_comb;
  wire [24:0] p1_sum__1353_comb;
  wire [24:0] p1_sum__1344_comb;
  wire [24:0] p1_sum__1345_comb;
  wire [24:0] p1_sum__1322_comb;
  wire [24:0] p1_sum__1323_comb;
  wire [24:0] p1_sum__1308_comb;
  wire [24:0] p1_sum__1309_comb;
  wire [24:0] p1_sum__1280_comb;
  wire [24:0] p1_sum__1281_comb;
  wire [24:0] p1_sum__1268_comb;
  wire [24:0] p1_sum__1269_comb;
  wire [24:0] p1_sum__1346_comb;
  wire [24:0] p1_sum__1347_comb;
  wire [24:0] p1_sum__1336_comb;
  wire [24:0] p1_sum__1337_comb;
  wire [24:0] p1_sum__1310_comb;
  wire [24:0] p1_sum__1311_comb;
  wire [24:0] p1_sum__1296_comb;
  wire [24:0] p1_sum__1297_comb;
  wire [24:0] p1_sum__1270_comb;
  wire [24:0] p1_sum__1271_comb;
  wire [24:0] p1_sum__1260_comb;
  wire [24:0] p1_sum__1261_comb;
  wire [24:0] p1_sum__1338_comb;
  wire [24:0] p1_sum__1339_comb;
  wire [24:0] p1_sum__1326_comb;
  wire [24:0] p1_sum__1327_comb;
  wire [24:0] p1_sum__1298_comb;
  wire [24:0] p1_sum__1299_comb;
  wire [24:0] p1_sum__1284_comb;
  wire [24:0] p1_sum__1285_comb;
  wire [24:0] p1_sum__1262_comb;
  wire [24:0] p1_sum__1263_comb;
  wire [24:0] p1_sum__1254_comb;
  wire [24:0] p1_sum__1255_comb;
  wire [24:0] p1_sum__1328_comb;
  wire [24:0] p1_sum__1329_comb;
  wire [24:0] p1_sum__1314_comb;
  wire [24:0] p1_sum__1315_comb;
  wire [24:0] p1_sum__1286_comb;
  wire [24:0] p1_sum__1287_comb;
  wire [24:0] p1_sum__1274_comb;
  wire [24:0] p1_sum__1275_comb;
  wire [24:0] p1_sum__1256_comb;
  wire [24:0] p1_sum__1257_comb;
  wire [24:0] p1_sum__1250_comb;
  wire [24:0] p1_sum__1251_comb;
  wire [24:0] p1_sum__1316_comb;
  wire [24:0] p1_sum__1317_comb;
  wire [24:0] p1_sum__1302_comb;
  wire [24:0] p1_sum__1303_comb;
  wire [24:0] p1_sum__1276_comb;
  wire [24:0] p1_sum__1277_comb;
  wire [24:0] p1_sum__1266_comb;
  wire [24:0] p1_sum__1267_comb;
  wire [24:0] p1_sum__1252_comb;
  wire [24:0] p1_sum__1253_comb;
  wire [24:0] p1_sum__1248_comb;
  wire [24:0] p1_sum__1249_comb;
  wire [24:0] p1_sum__1130_comb;
  wire [24:0] p1_sum__1115_comb;
  wire [24:0] p1_sum__1127_comb;
  wire [24:0] p1_sum__1109_comb;
  wire [24:0] p1_sum__1123_comb;
  wire [24:0] p1_sum__1103_comb;
  wire [24:0] p1_sum__1118_comb;
  wire [24:0] p1_sum__1097_comb;
  wire [24:0] p1_sum__1112_comb;
  wire [24:0] p1_sum__1092_comb;
  wire [24:0] p1_sum__1106_comb;
  wire [24:0] p1_sum__1088_comb;
  wire [24:0] p1_sum__1100_comb;
  wire [24:0] p1_sum__1085_comb;
  wire [24:0] p1_sum__1135_comb;
  wire [24:0] p1_sum__1133_comb;
  wire [24:0] p1_sum__1126_comb;
  wire [24:0] p1_sum__1121_comb;
  wire [24:0] p1_sum__1108_comb;
  wire [24:0] p1_sum__1101_comb;
  wire [24:0] p1_sum__1134_comb;
  wire [24:0] p1_sum__1131_comb;
  wire [24:0] p1_sum__1122_comb;
  wire [24:0] p1_sum__1116_comb;
  wire [24:0] p1_sum__1102_comb;
  wire [24:0] p1_sum__1095_comb;
  wire [24:0] p1_sum__1132_comb;
  wire [24:0] p1_sum__1128_comb;
  wire [24:0] p1_sum__1117_comb;
  wire [24:0] p1_sum__1110_comb;
  wire [24:0] p1_sum__1096_comb;
  wire [24:0] p1_sum__1090_comb;
  wire [24:0] p1_sum__1129_comb;
  wire [24:0] p1_sum__1124_comb;
  wire [24:0] p1_sum__1111_comb;
  wire [24:0] p1_sum__1104_comb;
  wire [24:0] p1_sum__1091_comb;
  wire [24:0] p1_sum__1086_comb;
  wire [24:0] p1_sum__1125_comb;
  wire [24:0] p1_sum__1119_comb;
  wire [24:0] p1_sum__1105_comb;
  wire [24:0] p1_sum__1098_comb;
  wire [24:0] p1_sum__1087_comb;
  wire [24:0] p1_sum__1083_comb;
  wire [24:0] p1_sum__1120_comb;
  wire [24:0] p1_sum__1113_comb;
  wire [24:0] p1_sum__1099_comb;
  wire [24:0] p1_sum__1093_comb;
  wire [24:0] p1_sum__1084_comb;
  wire [24:0] p1_sum__1081_comb;
  wire [24:0] p1_sum__1114_comb;
  wire [24:0] p1_sum__1107_comb;
  wire [24:0] p1_sum__1094_comb;
  wire [24:0] p1_sum__1089_comb;
  wire [24:0] p1_sum__1082_comb;
  wire [24:0] p1_sum__1080_comb;
  wire [24:0] p1_add_143035_comb;
  wire [24:0] p1_add_143036_comb;
  wire [24:0] p1_add_143037_comb;
  wire [24:0] p1_add_143038_comb;
  wire [24:0] p1_add_143039_comb;
  wire [24:0] p1_add_143040_comb;
  wire [24:0] p1_add_143041_comb;
  wire [24:0] p1_add_143042_comb;
  wire [24:0] p1_add_143043_comb;
  wire [24:0] p1_add_143044_comb;
  wire [24:0] p1_add_143045_comb;
  wire [24:0] p1_add_143046_comb;
  wire [24:0] p1_add_143047_comb;
  wire [24:0] p1_add_143048_comb;
  wire [24:0] p1_add_143049_comb;
  wire [24:0] p1_add_143050_comb;
  wire [24:0] p1_add_143051_comb;
  wire [24:0] p1_add_143052_comb;
  wire [24:0] p1_add_143053_comb;
  wire [24:0] p1_add_143054_comb;
  wire [24:0] p1_add_143055_comb;
  wire [24:0] p1_add_143056_comb;
  wire [24:0] p1_add_143057_comb;
  wire [24:0] p1_add_143058_comb;
  wire [24:0] p1_add_143059_comb;
  wire [24:0] p1_add_143060_comb;
  wire [24:0] p1_add_143061_comb;
  wire [24:0] p1_add_143062_comb;
  wire [24:0] p1_add_143063_comb;
  wire [24:0] p1_add_143064_comb;
  wire [24:0] p1_add_143065_comb;
  wire [24:0] p1_add_143066_comb;
  wire [24:0] p1_add_143067_comb;
  wire [24:0] p1_add_143068_comb;
  wire [24:0] p1_add_143069_comb;
  wire [24:0] p1_add_143070_comb;
  wire [24:0] p1_add_143071_comb;
  wire [24:0] p1_add_143072_comb;
  wire [24:0] p1_add_143073_comb;
  wire [24:0] p1_add_143074_comb;
  wire [24:0] p1_add_143075_comb;
  wire [24:0] p1_add_143076_comb;
  wire [24:0] p1_add_143077_comb;
  wire [24:0] p1_add_143078_comb;
  wire [24:0] p1_add_143079_comb;
  wire [24:0] p1_add_143080_comb;
  wire [24:0] p1_add_143081_comb;
  wire [24:0] p1_add_143082_comb;
  wire [24:0] p1_add_143083_comb;
  wire [24:0] p1_add_143084_comb;
  wire [24:0] p1_add_143085_comb;
  wire [24:0] p1_add_143086_comb;
  wire [24:0] p1_add_143087_comb;
  wire [24:0] p1_add_143088_comb;
  wire [24:0] p1_add_143089_comb;
  wire [24:0] p1_add_143090_comb;
  wire [24:0] p1_add_143091_comb;
  wire [24:0] p1_add_143092_comb;
  wire [24:0] p1_add_143093_comb;
  wire [24:0] p1_add_143094_comb;
  wire [24:0] p1_add_143095_comb;
  wire [24:0] p1_add_143096_comb;
  wire [24:0] p1_add_143097_comb;
  wire [24:0] p1_add_143098_comb;
  wire [8:0] p1_clipped__256_comb;
  wire [8:0] p1_clipped__259_comb;
  wire [8:0] p1_clipped__260_comb;
  wire [8:0] p1_clipped__263_comb;
  wire [8:0] p1_clipped__264_comb;
  wire [8:0] p1_clipped__267_comb;
  wire [8:0] p1_clipped__268_comb;
  wire [8:0] p1_clipped__271_comb;
  wire [8:0] p1_clipped__272_comb;
  wire [8:0] p1_clipped__275_comb;
  wire [8:0] p1_clipped__276_comb;
  wire [8:0] p1_clipped__279_comb;
  wire [8:0] p1_clipped__280_comb;
  wire [8:0] p1_clipped__283_comb;
  wire [8:0] p1_clipped__284_comb;
  wire [8:0] p1_clipped__287_comb;
  wire [8:0] p1_clipped__288_comb;
  wire [8:0] p1_clipped__289_comb;
  wire [8:0] p1_clipped__257_comb;
  wire [8:0] p1_clipped__258_comb;
  wire [8:0] p1_clipped__290_comb;
  wire [8:0] p1_clipped__291_comb;
  wire [8:0] p1_clipped__292_comb;
  wire [8:0] p1_clipped__293_comb;
  wire [8:0] p1_clipped__261_comb;
  wire [8:0] p1_clipped__262_comb;
  wire [8:0] p1_clipped__294_comb;
  wire [8:0] p1_clipped__295_comb;
  wire [8:0] p1_clipped__296_comb;
  wire [8:0] p1_clipped__297_comb;
  wire [8:0] p1_clipped__265_comb;
  wire [8:0] p1_clipped__266_comb;
  wire [8:0] p1_clipped__298_comb;
  wire [8:0] p1_clipped__299_comb;
  wire [8:0] p1_clipped__300_comb;
  wire [8:0] p1_clipped__301_comb;
  wire [8:0] p1_clipped__269_comb;
  wire [8:0] p1_clipped__270_comb;
  wire [8:0] p1_clipped__302_comb;
  wire [8:0] p1_clipped__303_comb;
  wire [8:0] p1_clipped__304_comb;
  wire [8:0] p1_clipped__305_comb;
  wire [8:0] p1_clipped__273_comb;
  wire [8:0] p1_clipped__274_comb;
  wire [8:0] p1_clipped__306_comb;
  wire [8:0] p1_clipped__307_comb;
  wire [8:0] p1_clipped__308_comb;
  wire [8:0] p1_clipped__309_comb;
  wire [8:0] p1_clipped__277_comb;
  wire [8:0] p1_clipped__278_comb;
  wire [8:0] p1_clipped__310_comb;
  wire [8:0] p1_clipped__311_comb;
  wire [8:0] p1_clipped__312_comb;
  wire [8:0] p1_clipped__313_comb;
  wire [8:0] p1_clipped__281_comb;
  wire [8:0] p1_clipped__282_comb;
  wire [8:0] p1_clipped__314_comb;
  wire [8:0] p1_clipped__315_comb;
  wire [8:0] p1_clipped__316_comb;
  wire [8:0] p1_clipped__317_comb;
  wire [8:0] p1_clipped__285_comb;
  wire [8:0] p1_clipped__286_comb;
  wire [8:0] p1_clipped__318_comb;
  wire [8:0] p1_clipped__319_comb;
  wire [9:0] p1_add_143867_comb;
  wire [9:0] p1_add_143868_comb;
  wire [9:0] p1_add_143869_comb;
  wire [9:0] p1_add_143870_comb;
  wire [9:0] p1_add_143871_comb;
  wire [9:0] p1_add_143872_comb;
  wire [9:0] p1_add_143873_comb;
  wire [9:0] p1_add_143874_comb;
  wire [9:0] p1_add_143875_comb;
  wire [9:0] p1_add_143876_comb;
  wire [9:0] p1_add_143877_comb;
  wire [9:0] p1_add_143878_comb;
  wire [9:0] p1_add_143879_comb;
  wire [9:0] p1_add_143880_comb;
  wire [9:0] p1_add_143881_comb;
  wire [9:0] p1_add_143882_comb;
  wire [9:0] p1_add_143883_comb;
  wire [9:0] p1_add_143884_comb;
  wire [9:0] p1_add_143885_comb;
  wire [9:0] p1_add_143886_comb;
  wire [9:0] p1_add_143887_comb;
  wire [9:0] p1_add_143888_comb;
  wire [9:0] p1_add_143889_comb;
  wire [9:0] p1_add_143890_comb;
  wire [9:0] p1_add_143891_comb;
  wire [9:0] p1_add_143892_comb;
  wire [9:0] p1_add_143893_comb;
  wire [9:0] p1_add_143894_comb;
  wire [9:0] p1_add_143895_comb;
  wire [9:0] p1_add_143896_comb;
  wire [9:0] p1_add_143897_comb;
  wire [9:0] p1_add_143898_comb;
  wire [9:0] p1_add_143899_comb;
  wire [9:0] p1_add_143900_comb;
  wire [9:0] p1_add_143901_comb;
  wire [9:0] p1_add_143902_comb;
  wire [9:0] p1_add_143903_comb;
  wire [9:0] p1_add_143904_comb;
  wire [9:0] p1_add_143905_comb;
  wire [9:0] p1_add_143906_comb;
  wire [9:0] p1_add_143907_comb;
  wire [9:0] p1_add_143908_comb;
  wire [9:0] p1_add_143909_comb;
  wire [9:0] p1_add_143910_comb;
  wire [9:0] p1_add_143911_comb;
  wire [9:0] p1_add_143912_comb;
  wire [9:0] p1_add_143913_comb;
  wire [9:0] p1_add_143914_comb;
  wire [9:0] p1_add_143915_comb;
  wire [9:0] p1_add_143916_comb;
  wire [9:0] p1_add_143917_comb;
  wire [9:0] p1_add_143918_comb;
  wire [9:0] p1_add_143919_comb;
  wire [9:0] p1_add_143920_comb;
  wire [9:0] p1_add_143921_comb;
  wire [9:0] p1_add_143922_comb;
  wire [9:0] p1_add_143923_comb;
  wire [9:0] p1_add_143924_comb;
  wire [9:0] p1_add_143925_comb;
  wire [9:0] p1_add_143926_comb;
  wire [9:0] p1_add_143927_comb;
  wire [9:0] p1_add_143928_comb;
  wire [9:0] p1_add_143929_comb;
  wire [9:0] p1_add_143930_comb;
  wire [1:0] p1_bit_slice_143931_comb;
  wire [1:0] p1_bit_slice_143932_comb;
  wire [1:0] p1_bit_slice_143933_comb;
  wire [1:0] p1_bit_slice_143934_comb;
  wire [1:0] p1_bit_slice_143935_comb;
  wire [1:0] p1_bit_slice_143936_comb;
  wire [1:0] p1_bit_slice_143937_comb;
  wire [1:0] p1_bit_slice_143938_comb;
  wire [1:0] p1_bit_slice_143939_comb;
  wire [1:0] p1_bit_slice_143940_comb;
  wire [1:0] p1_bit_slice_143941_comb;
  wire [1:0] p1_bit_slice_143942_comb;
  wire [1:0] p1_bit_slice_143943_comb;
  wire [1:0] p1_bit_slice_143944_comb;
  wire [1:0] p1_bit_slice_143945_comb;
  wire [1:0] p1_bit_slice_143946_comb;
  wire [1:0] p1_bit_slice_143947_comb;
  wire [1:0] p1_bit_slice_143948_comb;
  wire [1:0] p1_bit_slice_143949_comb;
  wire [1:0] p1_bit_slice_143950_comb;
  wire [1:0] p1_bit_slice_143951_comb;
  wire [1:0] p1_bit_slice_143952_comb;
  wire [1:0] p1_bit_slice_143953_comb;
  wire [1:0] p1_bit_slice_143954_comb;
  wire [1:0] p1_bit_slice_143955_comb;
  wire [1:0] p1_bit_slice_143956_comb;
  wire [1:0] p1_bit_slice_143957_comb;
  wire [1:0] p1_bit_slice_143958_comb;
  wire [1:0] p1_bit_slice_143959_comb;
  wire [1:0] p1_bit_slice_143960_comb;
  wire [1:0] p1_bit_slice_143961_comb;
  wire [1:0] p1_bit_slice_143962_comb;
  wire [1:0] p1_bit_slice_143963_comb;
  wire [1:0] p1_bit_slice_143964_comb;
  wire [1:0] p1_bit_slice_143965_comb;
  wire [1:0] p1_bit_slice_143966_comb;
  wire [1:0] p1_bit_slice_143967_comb;
  wire [1:0] p1_bit_slice_143968_comb;
  wire [1:0] p1_bit_slice_143969_comb;
  wire [1:0] p1_bit_slice_143970_comb;
  wire [1:0] p1_bit_slice_143971_comb;
  wire [1:0] p1_bit_slice_143972_comb;
  wire [1:0] p1_bit_slice_143973_comb;
  wire [1:0] p1_bit_slice_143974_comb;
  wire [1:0] p1_bit_slice_143975_comb;
  wire [1:0] p1_bit_slice_143976_comb;
  wire [1:0] p1_bit_slice_143977_comb;
  wire [1:0] p1_bit_slice_143978_comb;
  wire [1:0] p1_bit_slice_143979_comb;
  wire [1:0] p1_bit_slice_143980_comb;
  wire [1:0] p1_bit_slice_143981_comb;
  wire [1:0] p1_bit_slice_143982_comb;
  wire [1:0] p1_bit_slice_143983_comb;
  wire [1:0] p1_bit_slice_143984_comb;
  wire [1:0] p1_bit_slice_143985_comb;
  wire [1:0] p1_bit_slice_143986_comb;
  wire [1:0] p1_bit_slice_143987_comb;
  wire [1:0] p1_bit_slice_143988_comb;
  wire [1:0] p1_bit_slice_143989_comb;
  wire [1:0] p1_bit_slice_143990_comb;
  wire [1:0] p1_bit_slice_143991_comb;
  wire [1:0] p1_bit_slice_143992_comb;
  wire [1:0] p1_bit_slice_143993_comb;
  wire [1:0] p1_bit_slice_143994_comb;
  wire [2:0] p1_add_144123_comb;
  wire [2:0] p1_add_144124_comb;
  wire [2:0] p1_add_144125_comb;
  wire [2:0] p1_add_144126_comb;
  wire [2:0] p1_add_144127_comb;
  wire [2:0] p1_add_144128_comb;
  wire [2:0] p1_add_144129_comb;
  wire [2:0] p1_add_144130_comb;
  wire [2:0] p1_add_144131_comb;
  wire [2:0] p1_add_144132_comb;
  wire [2:0] p1_add_144133_comb;
  wire [2:0] p1_add_144134_comb;
  wire [2:0] p1_add_144135_comb;
  wire [2:0] p1_add_144136_comb;
  wire [2:0] p1_add_144137_comb;
  wire [2:0] p1_add_144138_comb;
  wire [2:0] p1_add_144139_comb;
  wire [2:0] p1_add_144140_comb;
  wire [2:0] p1_add_144141_comb;
  wire [2:0] p1_add_144142_comb;
  wire [2:0] p1_add_144143_comb;
  wire [2:0] p1_add_144144_comb;
  wire [2:0] p1_add_144145_comb;
  wire [2:0] p1_add_144146_comb;
  wire [2:0] p1_add_144147_comb;
  wire [2:0] p1_add_144148_comb;
  wire [2:0] p1_add_144149_comb;
  wire [2:0] p1_add_144150_comb;
  wire [2:0] p1_add_144151_comb;
  wire [2:0] p1_add_144152_comb;
  wire [2:0] p1_add_144153_comb;
  wire [2:0] p1_add_144154_comb;
  wire [2:0] p1_add_144155_comb;
  wire [2:0] p1_add_144156_comb;
  wire [2:0] p1_add_144157_comb;
  wire [2:0] p1_add_144158_comb;
  wire [2:0] p1_add_144159_comb;
  wire [2:0] p1_add_144160_comb;
  wire [2:0] p1_add_144161_comb;
  wire [2:0] p1_add_144162_comb;
  wire [2:0] p1_add_144163_comb;
  wire [2:0] p1_add_144164_comb;
  wire [2:0] p1_add_144165_comb;
  wire [2:0] p1_add_144166_comb;
  wire [2:0] p1_add_144167_comb;
  wire [2:0] p1_add_144168_comb;
  wire [2:0] p1_add_144169_comb;
  wire [2:0] p1_add_144170_comb;
  wire [2:0] p1_add_144171_comb;
  wire [2:0] p1_add_144172_comb;
  wire [2:0] p1_add_144173_comb;
  wire [2:0] p1_add_144174_comb;
  wire [2:0] p1_add_144175_comb;
  wire [2:0] p1_add_144176_comb;
  wire [2:0] p1_add_144177_comb;
  wire [2:0] p1_add_144178_comb;
  wire [2:0] p1_add_144179_comb;
  wire [2:0] p1_add_144180_comb;
  wire [2:0] p1_add_144181_comb;
  wire [2:0] p1_add_144182_comb;
  wire [2:0] p1_add_144183_comb;
  wire [2:0] p1_add_144184_comb;
  wire [2:0] p1_add_144185_comb;
  wire [2:0] p1_add_144186_comb;
  wire [7:0] p1_clipped__40_comb;
  wire [7:0] p1_clipped__88_comb;
  wire [7:0] p1_clipped__41_comb;
  wire [7:0] p1_clipped__89_comb;
  wire [7:0] p1_clipped__42_comb;
  wire [7:0] p1_clipped__90_comb;
  wire [7:0] p1_clipped__43_comb;
  wire [7:0] p1_clipped__91_comb;
  wire [7:0] p1_clipped__44_comb;
  wire [7:0] p1_clipped__92_comb;
  wire [7:0] p1_clipped__45_comb;
  wire [7:0] p1_clipped__93_comb;
  wire [7:0] p1_clipped__46_comb;
  wire [7:0] p1_clipped__94_comb;
  wire [7:0] p1_clipped__47_comb;
  wire [7:0] p1_clipped__95_comb;
  wire [7:0] p1_clipped__8_comb;
  wire [7:0] p1_clipped__24_comb;
  wire [7:0] p1_clipped__56_comb;
  wire [7:0] p1_clipped__72_comb;
  wire [7:0] p1_clipped__104_comb;
  wire [7:0] p1_clipped__120_comb;
  wire [7:0] p1_clipped__9_comb;
  wire [7:0] p1_clipped__25_comb;
  wire [7:0] p1_clipped__57_comb;
  wire [7:0] p1_clipped__73_comb;
  wire [7:0] p1_clipped__105_comb;
  wire [7:0] p1_clipped__121_comb;
  wire [7:0] p1_clipped__10_comb;
  wire [7:0] p1_clipped__26_comb;
  wire [7:0] p1_clipped__58_comb;
  wire [7:0] p1_clipped__74_comb;
  wire [7:0] p1_clipped__106_comb;
  wire [7:0] p1_clipped__122_comb;
  wire [7:0] p1_clipped__11_comb;
  wire [7:0] p1_clipped__27_comb;
  wire [7:0] p1_clipped__59_comb;
  wire [7:0] p1_clipped__75_comb;
  wire [7:0] p1_clipped__107_comb;
  wire [7:0] p1_clipped__123_comb;
  wire [7:0] p1_clipped__12_comb;
  wire [7:0] p1_clipped__28_comb;
  wire [7:0] p1_clipped__60_comb;
  wire [7:0] p1_clipped__76_comb;
  wire [7:0] p1_clipped__108_comb;
  wire [7:0] p1_clipped__124_comb;
  wire [7:0] p1_clipped__13_comb;
  wire [7:0] p1_clipped__29_comb;
  wire [7:0] p1_clipped__61_comb;
  wire [7:0] p1_clipped__77_comb;
  wire [7:0] p1_clipped__109_comb;
  wire [7:0] p1_clipped__125_comb;
  wire [7:0] p1_clipped__14_comb;
  wire [7:0] p1_clipped__30_comb;
  wire [7:0] p1_clipped__62_comb;
  wire [7:0] p1_clipped__78_comb;
  wire [7:0] p1_clipped__110_comb;
  wire [7:0] p1_clipped__126_comb;
  wire [7:0] p1_clipped__15_comb;
  wire [7:0] p1_clipped__31_comb;
  wire [7:0] p1_clipped__63_comb;
  wire [7:0] p1_clipped__79_comb;
  wire [7:0] p1_clipped__111_comb;
  wire [7:0] p1_clipped__127_comb;
  wire [7:0] p1_shifted__66_squeezed_comb;
  wire [7:0] p1_shifted__69_squeezed_comb;
  wire [7:0] p1_shifted__74_squeezed_comb;
  wire [7:0] p1_shifted__77_squeezed_comb;
  wire [7:0] p1_shifted__82_squeezed_comb;
  wire [7:0] p1_shifted__85_squeezed_comb;
  wire [7:0] p1_shifted__90_squeezed_comb;
  wire [7:0] p1_shifted__93_squeezed_comb;
  wire [7:0] p1_shifted__98_squeezed_comb;
  wire [7:0] p1_shifted__101_squeezed_comb;
  wire [7:0] p1_shifted__106_squeezed_comb;
  wire [7:0] p1_shifted__109_squeezed_comb;
  wire [7:0] p1_shifted__114_squeezed_comb;
  wire [7:0] p1_shifted__117_squeezed_comb;
  wire [7:0] p1_shifted__122_squeezed_comb;
  wire [7:0] p1_shifted__125_squeezed_comb;
  wire [7:0] p1_shifted__64_squeezed_comb;
  wire [7:0] p1_shifted__65_squeezed_comb;
  wire [7:0] p1_shifted__67_squeezed_comb;
  wire [7:0] p1_shifted__68_squeezed_comb;
  wire [7:0] p1_shifted__70_squeezed_comb;
  wire [7:0] p1_shifted__71_squeezed_comb;
  wire [7:0] p1_shifted__72_squeezed_comb;
  wire [7:0] p1_shifted__73_squeezed_comb;
  wire [7:0] p1_shifted__75_squeezed_comb;
  wire [7:0] p1_shifted__76_squeezed_comb;
  wire [7:0] p1_shifted__78_squeezed_comb;
  wire [7:0] p1_shifted__79_squeezed_comb;
  wire [7:0] p1_shifted__80_squeezed_comb;
  wire [7:0] p1_shifted__81_squeezed_comb;
  wire [7:0] p1_shifted__83_squeezed_comb;
  wire [7:0] p1_shifted__84_squeezed_comb;
  wire [7:0] p1_shifted__86_squeezed_comb;
  wire [7:0] p1_shifted__87_squeezed_comb;
  wire [7:0] p1_shifted__88_squeezed_comb;
  wire [7:0] p1_shifted__89_squeezed_comb;
  wire [7:0] p1_shifted__91_squeezed_comb;
  wire [7:0] p1_shifted__92_squeezed_comb;
  wire [7:0] p1_shifted__94_squeezed_comb;
  wire [7:0] p1_shifted__95_squeezed_comb;
  wire [7:0] p1_shifted__96_squeezed_comb;
  wire [7:0] p1_shifted__97_squeezed_comb;
  wire [7:0] p1_shifted__99_squeezed_comb;
  wire [7:0] p1_shifted__100_squeezed_comb;
  wire [7:0] p1_shifted__102_squeezed_comb;
  wire [7:0] p1_shifted__103_squeezed_comb;
  wire [7:0] p1_shifted__104_squeezed_comb;
  wire [7:0] p1_shifted__105_squeezed_comb;
  wire [7:0] p1_shifted__107_squeezed_comb;
  wire [7:0] p1_shifted__108_squeezed_comb;
  wire [7:0] p1_shifted__110_squeezed_comb;
  wire [7:0] p1_shifted__111_squeezed_comb;
  wire [7:0] p1_shifted__112_squeezed_comb;
  wire [7:0] p1_shifted__113_squeezed_comb;
  wire [7:0] p1_shifted__115_squeezed_comb;
  wire [7:0] p1_shifted__116_squeezed_comb;
  wire [7:0] p1_shifted__118_squeezed_comb;
  wire [7:0] p1_shifted__119_squeezed_comb;
  wire [7:0] p1_shifted__120_squeezed_comb;
  wire [7:0] p1_shifted__121_squeezed_comb;
  wire [7:0] p1_shifted__123_squeezed_comb;
  wire [7:0] p1_shifted__124_squeezed_comb;
  wire [7:0] p1_shifted__126_squeezed_comb;
  wire [7:0] p1_shifted__127_squeezed_comb;
  wire [15:0] p1_smul_58226_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___192_comb;
  wire [15:0] p1_smul_58232_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___195_comb;
  wire [15:0] p1_smul_58242_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___196_comb;
  wire [15:0] p1_smul_58248_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___199_comb;
  wire [15:0] p1_smul_58258_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___200_comb;
  wire [15:0] p1_smul_58264_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___203_comb;
  wire [15:0] p1_smul_58274_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___204_comb;
  wire [15:0] p1_smul_58280_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___207_comb;
  wire [15:0] p1_smul_58290_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___208_comb;
  wire [15:0] p1_smul_58296_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___211_comb;
  wire [15:0] p1_smul_58306_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___212_comb;
  wire [15:0] p1_smul_58312_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___215_comb;
  wire [15:0] p1_smul_58322_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___216_comb;
  wire [15:0] p1_smul_58328_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___219_comb;
  wire [15:0] p1_smul_58338_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___220_comb;
  wire [15:0] p1_smul_58344_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___223_comb;
  wire [14:0] p1_smul_58350_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___64_comb;
  wire [14:0] p1_smul_58352_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___224_comb;
  wire [14:0] p1_smul_58354_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___225_comb;
  wire [14:0] p1_smul_58356_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___65_comb;
  wire [14:0] p1_smul_58358_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___66_comb;
  wire [14:0] p1_smul_58360_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___226_comb;
  wire [14:0] p1_smul_58362_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___227_comb;
  wire [14:0] p1_smul_58364_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___67_comb;
  wire [14:0] p1_smul_58366_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___68_comb;
  wire [14:0] p1_smul_58368_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___228_comb;
  wire [14:0] p1_smul_58370_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___229_comb;
  wire [14:0] p1_smul_58372_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___69_comb;
  wire [14:0] p1_smul_58374_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___70_comb;
  wire [14:0] p1_smul_58376_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___230_comb;
  wire [14:0] p1_smul_58378_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___231_comb;
  wire [14:0] p1_smul_58380_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___71_comb;
  wire [14:0] p1_smul_58382_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___72_comb;
  wire [14:0] p1_smul_58384_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___232_comb;
  wire [14:0] p1_smul_58386_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___233_comb;
  wire [14:0] p1_smul_58388_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___73_comb;
  wire [14:0] p1_smul_58390_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___74_comb;
  wire [14:0] p1_smul_58392_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___234_comb;
  wire [14:0] p1_smul_58394_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___235_comb;
  wire [14:0] p1_smul_58396_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___75_comb;
  wire [14:0] p1_smul_58398_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___76_comb;
  wire [14:0] p1_smul_58400_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___236_comb;
  wire [14:0] p1_smul_58402_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___237_comb;
  wire [14:0] p1_smul_58404_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___77_comb;
  wire [14:0] p1_smul_58406_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___78_comb;
  wire [14:0] p1_smul_58408_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___238_comb;
  wire [14:0] p1_smul_58410_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___239_comb;
  wire [14:0] p1_smul_58412_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___79_comb;
  wire [14:0] p1_smul_58414_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___80_comb;
  wire [14:0] p1_smul_58416_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___240_comb;
  wire [14:0] p1_smul_58418_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___241_comb;
  wire [14:0] p1_smul_58420_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___81_comb;
  wire [14:0] p1_smul_58422_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___82_comb;
  wire [14:0] p1_smul_58424_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___242_comb;
  wire [14:0] p1_smul_58426_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___243_comb;
  wire [14:0] p1_smul_58428_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___83_comb;
  wire [14:0] p1_smul_58430_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___84_comb;
  wire [14:0] p1_smul_58432_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___244_comb;
  wire [14:0] p1_smul_58434_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___245_comb;
  wire [14:0] p1_smul_58436_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___85_comb;
  wire [14:0] p1_smul_58438_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___86_comb;
  wire [14:0] p1_smul_58440_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___246_comb;
  wire [14:0] p1_smul_58442_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___247_comb;
  wire [14:0] p1_smul_58444_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___87_comb;
  wire [14:0] p1_smul_58446_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___88_comb;
  wire [14:0] p1_smul_58448_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___248_comb;
  wire [14:0] p1_smul_58450_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___249_comb;
  wire [14:0] p1_smul_58452_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___89_comb;
  wire [14:0] p1_smul_58454_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___90_comb;
  wire [14:0] p1_smul_58456_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___250_comb;
  wire [14:0] p1_smul_58458_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___251_comb;
  wire [14:0] p1_smul_58460_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___91_comb;
  wire [14:0] p1_smul_58462_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___92_comb;
  wire [14:0] p1_smul_58464_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___252_comb;
  wire [14:0] p1_smul_58466_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___253_comb;
  wire [14:0] p1_smul_58468_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___93_comb;
  wire [14:0] p1_smul_58470_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___94_comb;
  wire [14:0] p1_smul_58472_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___254_comb;
  wire [14:0] p1_smul_58474_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___255_comb;
  wire [14:0] p1_smul_58476_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___95_comb;
  wire [15:0] p1_smul_58484_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___257_comb;
  wire [15:0] p1_smul_58486_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___258_comb;
  wire [15:0] p1_smul_58500_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___261_comb;
  wire [15:0] p1_smul_58502_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___262_comb;
  wire [15:0] p1_smul_58516_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___265_comb;
  wire [15:0] p1_smul_58518_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___266_comb;
  wire [15:0] p1_smul_58532_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___269_comb;
  wire [15:0] p1_smul_58534_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___270_comb;
  wire [15:0] p1_smul_58548_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___273_comb;
  wire [15:0] p1_smul_58550_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___274_comb;
  wire [15:0] p1_smul_58564_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___277_comb;
  wire [15:0] p1_smul_58566_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___278_comb;
  wire [15:0] p1_smul_58580_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___281_comb;
  wire [15:0] p1_smul_58582_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___282_comb;
  wire [15:0] p1_smul_58596_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___285_comb;
  wire [15:0] p1_smul_58598_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___286_comb;
  wire [15:0] p1_smul_58734_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___288_comb;
  wire [15:0] p1_smul_58748_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___291_comb;
  wire [15:0] p1_smul_58750_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___292_comb;
  wire [15:0] p1_smul_58764_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___295_comb;
  wire [15:0] p1_smul_58766_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___296_comb;
  wire [15:0] p1_smul_58780_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___299_comb;
  wire [15:0] p1_smul_58782_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___300_comb;
  wire [15:0] p1_smul_58796_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___303_comb;
  wire [15:0] p1_smul_58798_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___304_comb;
  wire [15:0] p1_smul_58812_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___307_comb;
  wire [15:0] p1_smul_58814_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___308_comb;
  wire [15:0] p1_smul_58828_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___311_comb;
  wire [15:0] p1_smul_58830_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___312_comb;
  wire [15:0] p1_smul_58844_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___315_comb;
  wire [15:0] p1_smul_58846_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___316_comb;
  wire [15:0] p1_smul_58860_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___319_comb;
  wire [14:0] p1_smul_58862_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___320_comb;
  wire [14:0] p1_smul_58864_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___96_comb;
  wire [14:0] p1_smul_58866_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___321_comb;
  wire [14:0] p1_smul_58868_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___97_comb;
  wire [14:0] p1_smul_58870_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___98_comb;
  wire [14:0] p1_smul_58872_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___322_comb;
  wire [14:0] p1_smul_58874_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___99_comb;
  wire [14:0] p1_smul_58876_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___323_comb;
  wire [14:0] p1_smul_58878_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___324_comb;
  wire [14:0] p1_smul_58880_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___100_comb;
  wire [14:0] p1_smul_58882_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___325_comb;
  wire [14:0] p1_smul_58884_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___101_comb;
  wire [14:0] p1_smul_58886_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___102_comb;
  wire [14:0] p1_smul_58888_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___326_comb;
  wire [14:0] p1_smul_58890_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___103_comb;
  wire [14:0] p1_smul_58892_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___327_comb;
  wire [14:0] p1_smul_58894_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___328_comb;
  wire [14:0] p1_smul_58896_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___104_comb;
  wire [14:0] p1_smul_58898_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___329_comb;
  wire [14:0] p1_smul_58900_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___105_comb;
  wire [14:0] p1_smul_58902_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___106_comb;
  wire [14:0] p1_smul_58904_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___330_comb;
  wire [14:0] p1_smul_58906_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___107_comb;
  wire [14:0] p1_smul_58908_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___331_comb;
  wire [14:0] p1_smul_58910_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___332_comb;
  wire [14:0] p1_smul_58912_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___108_comb;
  wire [14:0] p1_smul_58914_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___333_comb;
  wire [14:0] p1_smul_58916_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___109_comb;
  wire [14:0] p1_smul_58918_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___110_comb;
  wire [14:0] p1_smul_58920_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___334_comb;
  wire [14:0] p1_smul_58922_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___111_comb;
  wire [14:0] p1_smul_58924_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___335_comb;
  wire [14:0] p1_smul_58926_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___336_comb;
  wire [14:0] p1_smul_58928_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___112_comb;
  wire [14:0] p1_smul_58930_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___337_comb;
  wire [14:0] p1_smul_58932_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___113_comb;
  wire [14:0] p1_smul_58934_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___114_comb;
  wire [14:0] p1_smul_58936_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___338_comb;
  wire [14:0] p1_smul_58938_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___115_comb;
  wire [14:0] p1_smul_58940_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___339_comb;
  wire [14:0] p1_smul_58942_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___340_comb;
  wire [14:0] p1_smul_58944_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___116_comb;
  wire [14:0] p1_smul_58946_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___341_comb;
  wire [14:0] p1_smul_58948_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___117_comb;
  wire [14:0] p1_smul_58950_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___118_comb;
  wire [14:0] p1_smul_58952_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___342_comb;
  wire [14:0] p1_smul_58954_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___119_comb;
  wire [14:0] p1_smul_58956_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___343_comb;
  wire [14:0] p1_smul_58958_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___344_comb;
  wire [14:0] p1_smul_58960_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___120_comb;
  wire [14:0] p1_smul_58962_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___345_comb;
  wire [14:0] p1_smul_58964_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___121_comb;
  wire [14:0] p1_smul_58966_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___122_comb;
  wire [14:0] p1_smul_58968_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___346_comb;
  wire [14:0] p1_smul_58970_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___123_comb;
  wire [14:0] p1_smul_58972_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___347_comb;
  wire [14:0] p1_smul_58974_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___348_comb;
  wire [14:0] p1_smul_58976_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___124_comb;
  wire [14:0] p1_smul_58978_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___349_comb;
  wire [14:0] p1_smul_58980_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___125_comb;
  wire [14:0] p1_smul_58982_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___126_comb;
  wire [14:0] p1_smul_58984_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___350_comb;
  wire [14:0] p1_smul_58986_NarrowedMult__comb;
  wire [9:0] p1_smul_57454_TrailingBits___127_comb;
  wire [14:0] p1_smul_58988_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___351_comb;
  wire [15:0] p1_smul_58992_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___353_comb;
  wire [15:0] p1_smul_59002_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___354_comb;
  wire [15:0] p1_smul_59008_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___357_comb;
  wire [15:0] p1_smul_59018_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___358_comb;
  wire [15:0] p1_smul_59024_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___361_comb;
  wire [15:0] p1_smul_59034_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___362_comb;
  wire [15:0] p1_smul_59040_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___365_comb;
  wire [15:0] p1_smul_59050_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___366_comb;
  wire [15:0] p1_smul_59056_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___369_comb;
  wire [15:0] p1_smul_59066_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___370_comb;
  wire [15:0] p1_smul_59072_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___373_comb;
  wire [15:0] p1_smul_59082_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___374_comb;
  wire [15:0] p1_smul_59088_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___377_comb;
  wire [15:0] p1_smul_59098_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___378_comb;
  wire [15:0] p1_smul_59104_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___381_comb;
  wire [15:0] p1_smul_59114_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___382_comb;
  wire [24:0] p1_concat_145531_comb;
  wire [13:0] p1_smul_58228_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___193_comb;
  wire [13:0] p1_smul_58230_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___194_comb;
  wire [24:0] p1_concat_145536_comb;
  wire [24:0] p1_concat_145537_comb;
  wire [13:0] p1_smul_58244_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___197_comb;
  wire [13:0] p1_smul_58246_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___198_comb;
  wire [24:0] p1_concat_145542_comb;
  wire [24:0] p1_concat_145543_comb;
  wire [13:0] p1_smul_58260_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___201_comb;
  wire [13:0] p1_smul_58262_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___202_comb;
  wire [24:0] p1_concat_145548_comb;
  wire [24:0] p1_concat_145549_comb;
  wire [13:0] p1_smul_58276_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___205_comb;
  wire [13:0] p1_smul_58278_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___206_comb;
  wire [24:0] p1_concat_145554_comb;
  wire [24:0] p1_concat_145555_comb;
  wire [13:0] p1_smul_58292_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___209_comb;
  wire [13:0] p1_smul_58294_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___210_comb;
  wire [24:0] p1_concat_145560_comb;
  wire [24:0] p1_concat_145561_comb;
  wire [13:0] p1_smul_58308_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___213_comb;
  wire [13:0] p1_smul_58310_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___214_comb;
  wire [24:0] p1_concat_145566_comb;
  wire [24:0] p1_concat_145567_comb;
  wire [13:0] p1_smul_58324_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___217_comb;
  wire [13:0] p1_smul_58326_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___218_comb;
  wire [24:0] p1_concat_145572_comb;
  wire [24:0] p1_concat_145573_comb;
  wire [13:0] p1_smul_58340_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___221_comb;
  wire [13:0] p1_smul_58342_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___222_comb;
  wire [24:0] p1_concat_145578_comb;
  wire [24:0] p1_concat_145579_comb;
  wire [23:0] p1_concat_145580_comb;
  wire [23:0] p1_concat_145581_comb;
  wire [24:0] p1_concat_145582_comb;
  wire [24:0] p1_concat_145583_comb;
  wire [23:0] p1_concat_145584_comb;
  wire [23:0] p1_concat_145585_comb;
  wire [24:0] p1_concat_145586_comb;
  wire [24:0] p1_concat_145587_comb;
  wire [23:0] p1_concat_145588_comb;
  wire [23:0] p1_concat_145589_comb;
  wire [24:0] p1_concat_145590_comb;
  wire [24:0] p1_concat_145591_comb;
  wire [23:0] p1_concat_145592_comb;
  wire [23:0] p1_concat_145593_comb;
  wire [24:0] p1_concat_145594_comb;
  wire [24:0] p1_concat_145595_comb;
  wire [23:0] p1_concat_145596_comb;
  wire [23:0] p1_concat_145597_comb;
  wire [24:0] p1_concat_145598_comb;
  wire [24:0] p1_concat_145599_comb;
  wire [23:0] p1_concat_145600_comb;
  wire [23:0] p1_concat_145601_comb;
  wire [24:0] p1_concat_145602_comb;
  wire [24:0] p1_concat_145603_comb;
  wire [23:0] p1_concat_145604_comb;
  wire [23:0] p1_concat_145605_comb;
  wire [24:0] p1_concat_145606_comb;
  wire [24:0] p1_concat_145607_comb;
  wire [23:0] p1_concat_145608_comb;
  wire [23:0] p1_concat_145609_comb;
  wire [24:0] p1_concat_145610_comb;
  wire [24:0] p1_concat_145611_comb;
  wire [23:0] p1_concat_145612_comb;
  wire [23:0] p1_concat_145613_comb;
  wire [24:0] p1_concat_145614_comb;
  wire [24:0] p1_concat_145615_comb;
  wire [23:0] p1_concat_145616_comb;
  wire [23:0] p1_concat_145617_comb;
  wire [24:0] p1_concat_145618_comb;
  wire [24:0] p1_concat_145619_comb;
  wire [23:0] p1_concat_145620_comb;
  wire [23:0] p1_concat_145621_comb;
  wire [24:0] p1_concat_145622_comb;
  wire [24:0] p1_concat_145623_comb;
  wire [23:0] p1_concat_145624_comb;
  wire [23:0] p1_concat_145625_comb;
  wire [24:0] p1_concat_145626_comb;
  wire [24:0] p1_concat_145627_comb;
  wire [23:0] p1_concat_145628_comb;
  wire [23:0] p1_concat_145629_comb;
  wire [24:0] p1_concat_145630_comb;
  wire [24:0] p1_concat_145631_comb;
  wire [23:0] p1_concat_145632_comb;
  wire [23:0] p1_concat_145633_comb;
  wire [24:0] p1_concat_145634_comb;
  wire [24:0] p1_concat_145635_comb;
  wire [23:0] p1_concat_145636_comb;
  wire [23:0] p1_concat_145637_comb;
  wire [24:0] p1_concat_145638_comb;
  wire [24:0] p1_concat_145639_comb;
  wire [23:0] p1_concat_145640_comb;
  wire [23:0] p1_concat_145641_comb;
  wire [24:0] p1_concat_145642_comb;
  wire [13:0] p1_smul_58480_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___256_comb;
  wire [24:0] p1_concat_145645_comb;
  wire [24:0] p1_concat_145646_comb;
  wire [13:0] p1_smul_58490_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___259_comb;
  wire [13:0] p1_smul_58496_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___260_comb;
  wire [24:0] p1_concat_145651_comb;
  wire [24:0] p1_concat_145652_comb;
  wire [13:0] p1_smul_58506_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___263_comb;
  wire [13:0] p1_smul_58512_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___264_comb;
  wire [24:0] p1_concat_145657_comb;
  wire [24:0] p1_concat_145658_comb;
  wire [13:0] p1_smul_58522_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___267_comb;
  wire [13:0] p1_smul_58528_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___268_comb;
  wire [24:0] p1_concat_145663_comb;
  wire [24:0] p1_concat_145664_comb;
  wire [13:0] p1_smul_58538_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___271_comb;
  wire [13:0] p1_smul_58544_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___272_comb;
  wire [24:0] p1_concat_145669_comb;
  wire [24:0] p1_concat_145670_comb;
  wire [13:0] p1_smul_58554_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___275_comb;
  wire [13:0] p1_smul_58560_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___276_comb;
  wire [24:0] p1_concat_145675_comb;
  wire [24:0] p1_concat_145676_comb;
  wire [13:0] p1_smul_58570_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___279_comb;
  wire [13:0] p1_smul_58576_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___280_comb;
  wire [24:0] p1_concat_145681_comb;
  wire [24:0] p1_concat_145682_comb;
  wire [13:0] p1_smul_58586_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___283_comb;
  wire [13:0] p1_smul_58592_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___284_comb;
  wire [24:0] p1_concat_145687_comb;
  wire [24:0] p1_concat_145688_comb;
  wire [13:0] p1_smul_58602_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___287_comb;
  wire [24:0] p1_concat_145691_comb;
  wire [13:0] p1_smul_58738_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___289_comb;
  wire [13:0] p1_smul_58744_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___290_comb;
  wire [24:0] p1_concat_145696_comb;
  wire [24:0] p1_concat_145697_comb;
  wire [13:0] p1_smul_58754_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___293_comb;
  wire [13:0] p1_smul_58760_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___294_comb;
  wire [24:0] p1_concat_145702_comb;
  wire [24:0] p1_concat_145703_comb;
  wire [13:0] p1_smul_58770_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___297_comb;
  wire [13:0] p1_smul_58776_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___298_comb;
  wire [24:0] p1_concat_145708_comb;
  wire [24:0] p1_concat_145709_comb;
  wire [13:0] p1_smul_58786_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___301_comb;
  wire [13:0] p1_smul_58792_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___302_comb;
  wire [24:0] p1_concat_145714_comb;
  wire [24:0] p1_concat_145715_comb;
  wire [13:0] p1_smul_58802_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___305_comb;
  wire [13:0] p1_smul_58808_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___306_comb;
  wire [24:0] p1_concat_145720_comb;
  wire [24:0] p1_concat_145721_comb;
  wire [13:0] p1_smul_58818_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___309_comb;
  wire [13:0] p1_smul_58824_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___310_comb;
  wire [24:0] p1_concat_145726_comb;
  wire [24:0] p1_concat_145727_comb;
  wire [13:0] p1_smul_58834_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___313_comb;
  wire [13:0] p1_smul_58840_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___314_comb;
  wire [24:0] p1_concat_145732_comb;
  wire [24:0] p1_concat_145733_comb;
  wire [13:0] p1_smul_58850_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___317_comb;
  wire [13:0] p1_smul_58856_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___318_comb;
  wire [24:0] p1_concat_145738_comb;
  wire [23:0] p1_concat_145739_comb;
  wire [24:0] p1_concat_145740_comb;
  wire [23:0] p1_concat_145741_comb;
  wire [24:0] p1_concat_145742_comb;
  wire [24:0] p1_concat_145743_comb;
  wire [23:0] p1_concat_145744_comb;
  wire [24:0] p1_concat_145745_comb;
  wire [23:0] p1_concat_145746_comb;
  wire [23:0] p1_concat_145747_comb;
  wire [24:0] p1_concat_145748_comb;
  wire [23:0] p1_concat_145749_comb;
  wire [24:0] p1_concat_145750_comb;
  wire [24:0] p1_concat_145751_comb;
  wire [23:0] p1_concat_145752_comb;
  wire [24:0] p1_concat_145753_comb;
  wire [23:0] p1_concat_145754_comb;
  wire [23:0] p1_concat_145755_comb;
  wire [24:0] p1_concat_145756_comb;
  wire [23:0] p1_concat_145757_comb;
  wire [24:0] p1_concat_145758_comb;
  wire [24:0] p1_concat_145759_comb;
  wire [23:0] p1_concat_145760_comb;
  wire [24:0] p1_concat_145761_comb;
  wire [23:0] p1_concat_145762_comb;
  wire [23:0] p1_concat_145763_comb;
  wire [24:0] p1_concat_145764_comb;
  wire [23:0] p1_concat_145765_comb;
  wire [24:0] p1_concat_145766_comb;
  wire [24:0] p1_concat_145767_comb;
  wire [23:0] p1_concat_145768_comb;
  wire [24:0] p1_concat_145769_comb;
  wire [23:0] p1_concat_145770_comb;
  wire [23:0] p1_concat_145771_comb;
  wire [24:0] p1_concat_145772_comb;
  wire [23:0] p1_concat_145773_comb;
  wire [24:0] p1_concat_145774_comb;
  wire [24:0] p1_concat_145775_comb;
  wire [23:0] p1_concat_145776_comb;
  wire [24:0] p1_concat_145777_comb;
  wire [23:0] p1_concat_145778_comb;
  wire [23:0] p1_concat_145779_comb;
  wire [24:0] p1_concat_145780_comb;
  wire [23:0] p1_concat_145781_comb;
  wire [24:0] p1_concat_145782_comb;
  wire [24:0] p1_concat_145783_comb;
  wire [23:0] p1_concat_145784_comb;
  wire [24:0] p1_concat_145785_comb;
  wire [23:0] p1_concat_145786_comb;
  wire [23:0] p1_concat_145787_comb;
  wire [24:0] p1_concat_145788_comb;
  wire [23:0] p1_concat_145789_comb;
  wire [24:0] p1_concat_145790_comb;
  wire [24:0] p1_concat_145791_comb;
  wire [23:0] p1_concat_145792_comb;
  wire [24:0] p1_concat_145793_comb;
  wire [23:0] p1_concat_145794_comb;
  wire [23:0] p1_concat_145795_comb;
  wire [24:0] p1_concat_145796_comb;
  wire [23:0] p1_concat_145797_comb;
  wire [24:0] p1_concat_145798_comb;
  wire [24:0] p1_concat_145799_comb;
  wire [23:0] p1_concat_145800_comb;
  wire [24:0] p1_concat_145801_comb;
  wire [23:0] p1_concat_145802_comb;
  wire [13:0] p1_smul_58990_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___352_comb;
  wire [24:0] p1_concat_145805_comb;
  wire [24:0] p1_concat_145806_comb;
  wire [13:0] p1_smul_59004_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___355_comb;
  wire [13:0] p1_smul_59006_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___356_comb;
  wire [24:0] p1_concat_145811_comb;
  wire [24:0] p1_concat_145812_comb;
  wire [13:0] p1_smul_59020_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___359_comb;
  wire [13:0] p1_smul_59022_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___360_comb;
  wire [24:0] p1_concat_145817_comb;
  wire [24:0] p1_concat_145818_comb;
  wire [13:0] p1_smul_59036_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___363_comb;
  wire [13:0] p1_smul_59038_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___364_comb;
  wire [24:0] p1_concat_145823_comb;
  wire [24:0] p1_concat_145824_comb;
  wire [13:0] p1_smul_59052_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___367_comb;
  wire [13:0] p1_smul_59054_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___368_comb;
  wire [24:0] p1_concat_145829_comb;
  wire [24:0] p1_concat_145830_comb;
  wire [13:0] p1_smul_59068_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___371_comb;
  wire [13:0] p1_smul_59070_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___372_comb;
  wire [24:0] p1_concat_145835_comb;
  wire [24:0] p1_concat_145836_comb;
  wire [13:0] p1_smul_59084_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___375_comb;
  wire [13:0] p1_smul_59086_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___376_comb;
  wire [24:0] p1_concat_145841_comb;
  wire [24:0] p1_concat_145842_comb;
  wire [13:0] p1_smul_59100_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___379_comb;
  wire [13:0] p1_smul_59102_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___380_comb;
  wire [24:0] p1_concat_145847_comb;
  wire [24:0] p1_concat_145848_comb;
  wire [13:0] p1_smul_59116_NarrowedMult__comb;
  wire [8:0] p1_smul_57330_TrailingBits___383_comb;
  wire [7:0] p1_smul_57326_TrailingBits___192_comb;
  wire [7:0] p1_smul_57326_TrailingBits___193_comb;
  wire [7:0] p1_smul_57326_TrailingBits___194_comb;
  wire [7:0] p1_smul_57326_TrailingBits___195_comb;
  wire [7:0] p1_smul_57326_TrailingBits___196_comb;
  wire [7:0] p1_smul_57326_TrailingBits___197_comb;
  wire [7:0] p1_smul_57326_TrailingBits___198_comb;
  wire [7:0] p1_smul_57326_TrailingBits___199_comb;
  wire [7:0] p1_smul_57326_TrailingBits___200_comb;
  wire [7:0] p1_smul_57326_TrailingBits___201_comb;
  wire [7:0] p1_smul_57326_TrailingBits___202_comb;
  wire [7:0] p1_smul_57326_TrailingBits___203_comb;
  wire [7:0] p1_smul_57326_TrailingBits___204_comb;
  wire [7:0] p1_smul_57326_TrailingBits___205_comb;
  wire [7:0] p1_smul_57326_TrailingBits___206_comb;
  wire [7:0] p1_smul_57326_TrailingBits___207_comb;
  wire [7:0] p1_smul_57326_TrailingBits___208_comb;
  wire [7:0] p1_smul_57326_TrailingBits___209_comb;
  wire [7:0] p1_smul_57326_TrailingBits___210_comb;
  wire [7:0] p1_smul_57326_TrailingBits___211_comb;
  wire [7:0] p1_smul_57326_TrailingBits___212_comb;
  wire [7:0] p1_smul_57326_TrailingBits___213_comb;
  wire [7:0] p1_smul_57326_TrailingBits___214_comb;
  wire [7:0] p1_smul_57326_TrailingBits___215_comb;
  wire [7:0] p1_smul_57326_TrailingBits___216_comb;
  wire [7:0] p1_smul_57326_TrailingBits___217_comb;
  wire [7:0] p1_smul_57326_TrailingBits___218_comb;
  wire [7:0] p1_smul_57326_TrailingBits___219_comb;
  wire [7:0] p1_smul_57326_TrailingBits___220_comb;
  wire [7:0] p1_smul_57326_TrailingBits___221_comb;
  wire [7:0] p1_smul_57326_TrailingBits___222_comb;
  wire [7:0] p1_smul_57326_TrailingBits___223_comb;
  wire [7:0] p1_smul_57326_TrailingBits___224_comb;
  wire [7:0] p1_smul_57326_TrailingBits___225_comb;
  wire [7:0] p1_smul_57326_TrailingBits___226_comb;
  wire [7:0] p1_smul_57326_TrailingBits___227_comb;
  wire [7:0] p1_smul_57326_TrailingBits___228_comb;
  wire [7:0] p1_smul_57326_TrailingBits___229_comb;
  wire [7:0] p1_smul_57326_TrailingBits___230_comb;
  wire [7:0] p1_smul_57326_TrailingBits___231_comb;
  wire [7:0] p1_smul_57326_TrailingBits___232_comb;
  wire [7:0] p1_smul_57326_TrailingBits___233_comb;
  wire [7:0] p1_smul_57326_TrailingBits___234_comb;
  wire [7:0] p1_smul_57326_TrailingBits___235_comb;
  wire [7:0] p1_smul_57326_TrailingBits___236_comb;
  wire [7:0] p1_smul_57326_TrailingBits___237_comb;
  wire [7:0] p1_smul_57326_TrailingBits___238_comb;
  wire [7:0] p1_smul_57326_TrailingBits___239_comb;
  wire [7:0] p1_smul_57326_TrailingBits___240_comb;
  wire [7:0] p1_smul_57326_TrailingBits___241_comb;
  wire [7:0] p1_smul_57326_TrailingBits___242_comb;
  wire [7:0] p1_smul_57326_TrailingBits___243_comb;
  wire [7:0] p1_smul_57326_TrailingBits___244_comb;
  wire [7:0] p1_smul_57326_TrailingBits___245_comb;
  wire [7:0] p1_smul_57326_TrailingBits___246_comb;
  wire [7:0] p1_smul_57326_TrailingBits___247_comb;
  wire [7:0] p1_smul_57326_TrailingBits___248_comb;
  wire [7:0] p1_smul_57326_TrailingBits___249_comb;
  wire [7:0] p1_smul_57326_TrailingBits___250_comb;
  wire [7:0] p1_smul_57326_TrailingBits___251_comb;
  wire [7:0] p1_smul_57326_TrailingBits___252_comb;
  wire [7:0] p1_smul_57326_TrailingBits___253_comb;
  wire [7:0] p1_smul_57326_TrailingBits___254_comb;
  wire [7:0] p1_smul_57326_TrailingBits___255_comb;
  wire [31:0] p1_prod__519_comb;
  wire [22:0] p1_concat_146045_comb;
  wire [22:0] p1_concat_146046_comb;
  wire [31:0] p1_prod__534_comb;
  wire [31:0] p1_prod__583_comb;
  wire [22:0] p1_concat_146051_comb;
  wire [22:0] p1_concat_146052_comb;
  wire [31:0] p1_prod__598_comb;
  wire [31:0] p1_prod__647_comb;
  wire [22:0] p1_concat_146057_comb;
  wire [22:0] p1_concat_146058_comb;
  wire [31:0] p1_prod__662_comb;
  wire [31:0] p1_prod__711_comb;
  wire [22:0] p1_concat_146063_comb;
  wire [22:0] p1_concat_146064_comb;
  wire [31:0] p1_prod__726_comb;
  wire [31:0] p1_prod__775_comb;
  wire [22:0] p1_concat_146069_comb;
  wire [22:0] p1_concat_146070_comb;
  wire [31:0] p1_prod__790_comb;
  wire [31:0] p1_prod__839_comb;
  wire [22:0] p1_concat_146075_comb;
  wire [22:0] p1_concat_146076_comb;
  wire [31:0] p1_prod__854_comb;
  wire [31:0] p1_prod__903_comb;
  wire [22:0] p1_concat_146081_comb;
  wire [22:0] p1_concat_146082_comb;
  wire [31:0] p1_prod__918_comb;
  wire [31:0] p1_prod__967_comb;
  wire [22:0] p1_concat_146087_comb;
  wire [22:0] p1_concat_146088_comb;
  wire [31:0] p1_prod__982_comb;
  wire [31:0] p1_prod__517_comb;
  wire [31:0] p1_prod__520_comb;
  wire [31:0] p1_prod__524_comb;
  wire [31:0] p1_prod__529_comb;
  wire [31:0] p1_prod__535_comb;
  wire [31:0] p1_prod__542_comb;
  wire [31:0] p1_prod__549_comb;
  wire [31:0] p1_prod__555_comb;
  wire [31:0] p1_prod__581_comb;
  wire [31:0] p1_prod__584_comb;
  wire [31:0] p1_prod__588_comb;
  wire [31:0] p1_prod__593_comb;
  wire [31:0] p1_prod__599_comb;
  wire [31:0] p1_prod__606_comb;
  wire [31:0] p1_prod__613_comb;
  wire [31:0] p1_prod__619_comb;
  wire [31:0] p1_prod__645_comb;
  wire [31:0] p1_prod__648_comb;
  wire [31:0] p1_prod__652_comb;
  wire [31:0] p1_prod__657_comb;
  wire [31:0] p1_prod__663_comb;
  wire [31:0] p1_prod__670_comb;
  wire [31:0] p1_prod__677_comb;
  wire [31:0] p1_prod__683_comb;
  wire [31:0] p1_prod__709_comb;
  wire [31:0] p1_prod__712_comb;
  wire [31:0] p1_prod__716_comb;
  wire [31:0] p1_prod__721_comb;
  wire [31:0] p1_prod__727_comb;
  wire [31:0] p1_prod__734_comb;
  wire [31:0] p1_prod__741_comb;
  wire [31:0] p1_prod__747_comb;
  wire [31:0] p1_prod__773_comb;
  wire [31:0] p1_prod__776_comb;
  wire [31:0] p1_prod__780_comb;
  wire [31:0] p1_prod__785_comb;
  wire [31:0] p1_prod__791_comb;
  wire [31:0] p1_prod__798_comb;
  wire [31:0] p1_prod__805_comb;
  wire [31:0] p1_prod__811_comb;
  wire [31:0] p1_prod__837_comb;
  wire [31:0] p1_prod__840_comb;
  wire [31:0] p1_prod__844_comb;
  wire [31:0] p1_prod__849_comb;
  wire [31:0] p1_prod__855_comb;
  wire [31:0] p1_prod__862_comb;
  wire [31:0] p1_prod__869_comb;
  wire [31:0] p1_prod__875_comb;
  wire [31:0] p1_prod__901_comb;
  wire [31:0] p1_prod__904_comb;
  wire [31:0] p1_prod__908_comb;
  wire [31:0] p1_prod__913_comb;
  wire [31:0] p1_prod__919_comb;
  wire [31:0] p1_prod__926_comb;
  wire [31:0] p1_prod__933_comb;
  wire [31:0] p1_prod__939_comb;
  wire [31:0] p1_prod__965_comb;
  wire [31:0] p1_prod__968_comb;
  wire [31:0] p1_prod__972_comb;
  wire [31:0] p1_prod__977_comb;
  wire [31:0] p1_prod__983_comb;
  wire [31:0] p1_prod__990_comb;
  wire [31:0] p1_prod__997_comb;
  wire [31:0] p1_prod__1003_comb;
  wire [22:0] p1_concat_146187_comb;
  wire [31:0] p1_prod__536_comb;
  wire [31:0] p1_prod__543_comb;
  wire [22:0] p1_concat_146192_comb;
  wire [22:0] p1_concat_146193_comb;
  wire [31:0] p1_prod__600_comb;
  wire [31:0] p1_prod__607_comb;
  wire [22:0] p1_concat_146198_comb;
  wire [22:0] p1_concat_146199_comb;
  wire [31:0] p1_prod__664_comb;
  wire [31:0] p1_prod__671_comb;
  wire [22:0] p1_concat_146204_comb;
  wire [22:0] p1_concat_146205_comb;
  wire [31:0] p1_prod__728_comb;
  wire [31:0] p1_prod__735_comb;
  wire [22:0] p1_concat_146210_comb;
  wire [22:0] p1_concat_146211_comb;
  wire [31:0] p1_prod__792_comb;
  wire [31:0] p1_prod__799_comb;
  wire [22:0] p1_concat_146216_comb;
  wire [22:0] p1_concat_146217_comb;
  wire [31:0] p1_prod__856_comb;
  wire [31:0] p1_prod__863_comb;
  wire [22:0] p1_concat_146222_comb;
  wire [22:0] p1_concat_146223_comb;
  wire [31:0] p1_prod__920_comb;
  wire [31:0] p1_prod__927_comb;
  wire [22:0] p1_concat_146228_comb;
  wire [22:0] p1_concat_146229_comb;
  wire [31:0] p1_prod__984_comb;
  wire [31:0] p1_prod__991_comb;
  wire [22:0] p1_concat_146234_comb;
  wire [31:0] p1_prod__532_comb;
  wire [22:0] p1_concat_146237_comb;
  wire [22:0] p1_concat_146238_comb;
  wire [31:0] p1_prod__570_comb;
  wire [31:0] p1_prod__596_comb;
  wire [22:0] p1_concat_146243_comb;
  wire [22:0] p1_concat_146244_comb;
  wire [31:0] p1_prod__634_comb;
  wire [31:0] p1_prod__660_comb;
  wire [22:0] p1_concat_146249_comb;
  wire [22:0] p1_concat_146250_comb;
  wire [31:0] p1_prod__698_comb;
  wire [31:0] p1_prod__724_comb;
  wire [22:0] p1_concat_146255_comb;
  wire [22:0] p1_concat_146256_comb;
  wire [31:0] p1_prod__762_comb;
  wire [31:0] p1_prod__788_comb;
  wire [22:0] p1_concat_146261_comb;
  wire [22:0] p1_concat_146262_comb;
  wire [31:0] p1_prod__826_comb;
  wire [31:0] p1_prod__852_comb;
  wire [22:0] p1_concat_146267_comb;
  wire [22:0] p1_concat_146268_comb;
  wire [31:0] p1_prod__890_comb;
  wire [31:0] p1_prod__916_comb;
  wire [22:0] p1_concat_146273_comb;
  wire [22:0] p1_concat_146274_comb;
  wire [31:0] p1_prod__954_comb;
  wire [31:0] p1_prod__980_comb;
  wire [22:0] p1_concat_146279_comb;
  wire [22:0] p1_concat_146280_comb;
  wire [31:0] p1_prod__1018_comb;
  wire [31:0] p1_prod__539_comb;
  wire [31:0] p1_prod__546_comb;
  wire [31:0] p1_prod__553_comb;
  wire [31:0] p1_prod__559_comb;
  wire [31:0] p1_prod__564_comb;
  wire [31:0] p1_prod__568_comb;
  wire [31:0] p1_prod__571_comb;
  wire [31:0] p1_prod__573_comb;
  wire [31:0] p1_prod__603_comb;
  wire [31:0] p1_prod__610_comb;
  wire [31:0] p1_prod__617_comb;
  wire [31:0] p1_prod__623_comb;
  wire [31:0] p1_prod__628_comb;
  wire [31:0] p1_prod__632_comb;
  wire [31:0] p1_prod__635_comb;
  wire [31:0] p1_prod__637_comb;
  wire [31:0] p1_prod__667_comb;
  wire [31:0] p1_prod__674_comb;
  wire [31:0] p1_prod__681_comb;
  wire [31:0] p1_prod__687_comb;
  wire [31:0] p1_prod__692_comb;
  wire [31:0] p1_prod__696_comb;
  wire [31:0] p1_prod__699_comb;
  wire [31:0] p1_prod__701_comb;
  wire [31:0] p1_prod__731_comb;
  wire [31:0] p1_prod__738_comb;
  wire [31:0] p1_prod__745_comb;
  wire [31:0] p1_prod__751_comb;
  wire [31:0] p1_prod__756_comb;
  wire [31:0] p1_prod__760_comb;
  wire [31:0] p1_prod__763_comb;
  wire [31:0] p1_prod__765_comb;
  wire [31:0] p1_prod__795_comb;
  wire [31:0] p1_prod__802_comb;
  wire [31:0] p1_prod__809_comb;
  wire [31:0] p1_prod__815_comb;
  wire [31:0] p1_prod__820_comb;
  wire [31:0] p1_prod__824_comb;
  wire [31:0] p1_prod__827_comb;
  wire [31:0] p1_prod__829_comb;
  wire [31:0] p1_prod__859_comb;
  wire [31:0] p1_prod__866_comb;
  wire [31:0] p1_prod__873_comb;
  wire [31:0] p1_prod__879_comb;
  wire [31:0] p1_prod__884_comb;
  wire [31:0] p1_prod__888_comb;
  wire [31:0] p1_prod__891_comb;
  wire [31:0] p1_prod__893_comb;
  wire [31:0] p1_prod__923_comb;
  wire [31:0] p1_prod__930_comb;
  wire [31:0] p1_prod__937_comb;
  wire [31:0] p1_prod__943_comb;
  wire [31:0] p1_prod__948_comb;
  wire [31:0] p1_prod__952_comb;
  wire [31:0] p1_prod__955_comb;
  wire [31:0] p1_prod__957_comb;
  wire [31:0] p1_prod__987_comb;
  wire [31:0] p1_prod__994_comb;
  wire [31:0] p1_prod__1001_comb;
  wire [31:0] p1_prod__1007_comb;
  wire [31:0] p1_prod__1012_comb;
  wire [31:0] p1_prod__1016_comb;
  wire [31:0] p1_prod__1019_comb;
  wire [31:0] p1_prod__1021_comb;
  wire [22:0] p1_concat_146379_comb;
  wire [31:0] p1_prod__554_comb;
  wire [31:0] p1_prod__574_comb;
  wire [22:0] p1_concat_146384_comb;
  wire [22:0] p1_concat_146385_comb;
  wire [31:0] p1_prod__618_comb;
  wire [31:0] p1_prod__638_comb;
  wire [22:0] p1_concat_146390_comb;
  wire [22:0] p1_concat_146391_comb;
  wire [31:0] p1_prod__682_comb;
  wire [31:0] p1_prod__702_comb;
  wire [22:0] p1_concat_146396_comb;
  wire [22:0] p1_concat_146397_comb;
  wire [31:0] p1_prod__746_comb;
  wire [31:0] p1_prod__766_comb;
  wire [22:0] p1_concat_146402_comb;
  wire [22:0] p1_concat_146403_comb;
  wire [31:0] p1_prod__810_comb;
  wire [31:0] p1_prod__830_comb;
  wire [22:0] p1_concat_146408_comb;
  wire [22:0] p1_concat_146409_comb;
  wire [31:0] p1_prod__874_comb;
  wire [31:0] p1_prod__894_comb;
  wire [22:0] p1_concat_146414_comb;
  wire [22:0] p1_concat_146415_comb;
  wire [31:0] p1_prod__938_comb;
  wire [31:0] p1_prod__958_comb;
  wire [22:0] p1_concat_146420_comb;
  wire [22:0] p1_concat_146421_comb;
  wire [31:0] p1_prod__1002_comb;
  wire [31:0] p1_prod__1022_comb;
  wire [22:0] p1_concat_146426_comb;
  wire [15:0] p1_shifted__64_comb;
  wire [7:0] p1_smul_57326_TrailingBits___64_comb;
  wire [15:0] p1_shifted__65_comb;
  wire [7:0] p1_smul_57326_TrailingBits___65_comb;
  wire [15:0] p1_shifted__66_comb;
  wire [7:0] p1_smul_57326_TrailingBits___66_comb;
  wire [15:0] p1_shifted__67_comb;
  wire [7:0] p1_smul_57326_TrailingBits___67_comb;
  wire [15:0] p1_shifted__68_comb;
  wire [7:0] p1_smul_57326_TrailingBits___68_comb;
  wire [15:0] p1_shifted__69_comb;
  wire [7:0] p1_smul_57326_TrailingBits___69_comb;
  wire [15:0] p1_shifted__70_comb;
  wire [7:0] p1_smul_57326_TrailingBits___70_comb;
  wire [15:0] p1_shifted__71_comb;
  wire [7:0] p1_smul_57326_TrailingBits___71_comb;
  wire [15:0] p1_shifted__72_comb;
  wire [7:0] p1_smul_57326_TrailingBits___72_comb;
  wire [15:0] p1_shifted__73_comb;
  wire [7:0] p1_smul_57326_TrailingBits___73_comb;
  wire [15:0] p1_shifted__74_comb;
  wire [7:0] p1_smul_57326_TrailingBits___74_comb;
  wire [15:0] p1_shifted__75_comb;
  wire [7:0] p1_smul_57326_TrailingBits___75_comb;
  wire [15:0] p1_shifted__76_comb;
  wire [7:0] p1_smul_57326_TrailingBits___76_comb;
  wire [15:0] p1_shifted__77_comb;
  wire [7:0] p1_smul_57326_TrailingBits___77_comb;
  wire [15:0] p1_shifted__78_comb;
  wire [7:0] p1_smul_57326_TrailingBits___78_comb;
  wire [15:0] p1_shifted__79_comb;
  wire [7:0] p1_smul_57326_TrailingBits___79_comb;
  wire [15:0] p1_shifted__80_comb;
  wire [7:0] p1_smul_57326_TrailingBits___80_comb;
  wire [15:0] p1_shifted__81_comb;
  wire [7:0] p1_smul_57326_TrailingBits___81_comb;
  wire [15:0] p1_shifted__82_comb;
  wire [7:0] p1_smul_57326_TrailingBits___82_comb;
  wire [15:0] p1_shifted__83_comb;
  wire [7:0] p1_smul_57326_TrailingBits___83_comb;
  wire [15:0] p1_shifted__84_comb;
  wire [7:0] p1_smul_57326_TrailingBits___84_comb;
  wire [15:0] p1_shifted__85_comb;
  wire [7:0] p1_smul_57326_TrailingBits___85_comb;
  wire [15:0] p1_shifted__86_comb;
  wire [7:0] p1_smul_57326_TrailingBits___86_comb;
  wire [15:0] p1_shifted__87_comb;
  wire [7:0] p1_smul_57326_TrailingBits___87_comb;
  wire [15:0] p1_shifted__88_comb;
  wire [7:0] p1_smul_57326_TrailingBits___88_comb;
  wire [15:0] p1_shifted__89_comb;
  wire [7:0] p1_smul_57326_TrailingBits___89_comb;
  wire [15:0] p1_shifted__90_comb;
  wire [7:0] p1_smul_57326_TrailingBits___90_comb;
  wire [15:0] p1_shifted__91_comb;
  wire [7:0] p1_smul_57326_TrailingBits___91_comb;
  wire [15:0] p1_shifted__92_comb;
  wire [7:0] p1_smul_57326_TrailingBits___92_comb;
  wire [15:0] p1_shifted__93_comb;
  wire [7:0] p1_smul_57326_TrailingBits___93_comb;
  wire [15:0] p1_shifted__94_comb;
  wire [7:0] p1_smul_57326_TrailingBits___94_comb;
  wire [15:0] p1_shifted__95_comb;
  wire [7:0] p1_smul_57326_TrailingBits___95_comb;
  wire [15:0] p1_shifted__96_comb;
  wire [7:0] p1_smul_57326_TrailingBits___96_comb;
  wire [15:0] p1_shifted__97_comb;
  wire [7:0] p1_smul_57326_TrailingBits___97_comb;
  wire [15:0] p1_shifted__98_comb;
  wire [7:0] p1_smul_57326_TrailingBits___98_comb;
  wire [15:0] p1_shifted__99_comb;
  wire [7:0] p1_smul_57326_TrailingBits___99_comb;
  wire [15:0] p1_shifted__100_comb;
  wire [7:0] p1_smul_57326_TrailingBits___100_comb;
  wire [15:0] p1_shifted__101_comb;
  wire [7:0] p1_smul_57326_TrailingBits___101_comb;
  wire [15:0] p1_shifted__102_comb;
  wire [7:0] p1_smul_57326_TrailingBits___102_comb;
  wire [15:0] p1_shifted__103_comb;
  wire [7:0] p1_smul_57326_TrailingBits___103_comb;
  wire [15:0] p1_shifted__104_comb;
  wire [7:0] p1_smul_57326_TrailingBits___104_comb;
  wire [15:0] p1_shifted__105_comb;
  wire [7:0] p1_smul_57326_TrailingBits___105_comb;
  wire [15:0] p1_shifted__106_comb;
  wire [7:0] p1_smul_57326_TrailingBits___106_comb;
  wire [15:0] p1_shifted__107_comb;
  wire [7:0] p1_smul_57326_TrailingBits___107_comb;
  wire [15:0] p1_shifted__108_comb;
  wire [7:0] p1_smul_57326_TrailingBits___108_comb;
  wire [15:0] p1_shifted__109_comb;
  wire [7:0] p1_smul_57326_TrailingBits___109_comb;
  wire [15:0] p1_shifted__110_comb;
  wire [7:0] p1_smul_57326_TrailingBits___110_comb;
  wire [15:0] p1_shifted__111_comb;
  wire [7:0] p1_smul_57326_TrailingBits___111_comb;
  wire [15:0] p1_shifted__112_comb;
  wire [7:0] p1_smul_57326_TrailingBits___112_comb;
  wire [15:0] p1_shifted__113_comb;
  wire [7:0] p1_smul_57326_TrailingBits___113_comb;
  wire [15:0] p1_shifted__114_comb;
  wire [7:0] p1_smul_57326_TrailingBits___114_comb;
  wire [15:0] p1_shifted__115_comb;
  wire [7:0] p1_smul_57326_TrailingBits___115_comb;
  wire [15:0] p1_shifted__116_comb;
  wire [7:0] p1_smul_57326_TrailingBits___116_comb;
  wire [15:0] p1_shifted__117_comb;
  wire [7:0] p1_smul_57326_TrailingBits___117_comb;
  wire [15:0] p1_shifted__118_comb;
  wire [7:0] p1_smul_57326_TrailingBits___118_comb;
  wire [15:0] p1_shifted__119_comb;
  wire [7:0] p1_smul_57326_TrailingBits___119_comb;
  wire [15:0] p1_shifted__120_comb;
  wire [7:0] p1_smul_57326_TrailingBits___120_comb;
  wire [15:0] p1_shifted__121_comb;
  wire [7:0] p1_smul_57326_TrailingBits___121_comb;
  wire [15:0] p1_shifted__122_comb;
  wire [7:0] p1_smul_57326_TrailingBits___122_comb;
  wire [15:0] p1_shifted__123_comb;
  wire [7:0] p1_smul_57326_TrailingBits___123_comb;
  wire [15:0] p1_shifted__124_comb;
  wire [7:0] p1_smul_57326_TrailingBits___124_comb;
  wire [15:0] p1_shifted__125_comb;
  wire [7:0] p1_smul_57326_TrailingBits___125_comb;
  wire [15:0] p1_shifted__126_comb;
  wire [7:0] p1_smul_57326_TrailingBits___126_comb;
  wire [15:0] p1_shifted__127_comb;
  wire [7:0] p1_smul_57326_TrailingBits___127_comb;
  wire [31:0] p1_or_146687_comb;
  wire [31:0] p1_prod__523_comb;
  wire [31:0] p1_prod__528_comb;
  wire [31:0] p1_or_146694_comb;
  wire [31:0] p1_or_146701_comb;
  wire [31:0] p1_prod__587_comb;
  wire [31:0] p1_prod__592_comb;
  wire [31:0] p1_or_146708_comb;
  wire [31:0] p1_or_146715_comb;
  wire [31:0] p1_prod__651_comb;
  wire [31:0] p1_prod__656_comb;
  wire [31:0] p1_or_146722_comb;
  wire [31:0] p1_or_146729_comb;
  wire [31:0] p1_prod__715_comb;
  wire [31:0] p1_prod__720_comb;
  wire [31:0] p1_or_146736_comb;
  wire [31:0] p1_or_146743_comb;
  wire [31:0] p1_prod__779_comb;
  wire [31:0] p1_prod__784_comb;
  wire [31:0] p1_or_146750_comb;
  wire [31:0] p1_or_146757_comb;
  wire [31:0] p1_prod__843_comb;
  wire [31:0] p1_prod__848_comb;
  wire [31:0] p1_or_146764_comb;
  wire [31:0] p1_or_146771_comb;
  wire [31:0] p1_prod__907_comb;
  wire [31:0] p1_prod__912_comb;
  wire [31:0] p1_or_146778_comb;
  wire [31:0] p1_or_146785_comb;
  wire [31:0] p1_prod__971_comb;
  wire [31:0] p1_prod__976_comb;
  wire [31:0] p1_or_146792_comb;
  wire [31:0] p1_or_146797_comb;
  wire [31:0] p1_or_146804_comb;
  wire [31:0] p1_or_146807_comb;
  wire [31:0] p1_or_146814_comb;
  wire [31:0] p1_or_146817_comb;
  wire [31:0] p1_or_146824_comb;
  wire [31:0] p1_or_146827_comb;
  wire [31:0] p1_or_146834_comb;
  wire [31:0] p1_or_146837_comb;
  wire [31:0] p1_or_146844_comb;
  wire [31:0] p1_or_146847_comb;
  wire [31:0] p1_or_146854_comb;
  wire [31:0] p1_or_146857_comb;
  wire [31:0] p1_or_146864_comb;
  wire [31:0] p1_or_146867_comb;
  wire [31:0] p1_or_146874_comb;
  wire [31:0] p1_or_146877_comb;
  wire [31:0] p1_or_146884_comb;
  wire [31:0] p1_or_146887_comb;
  wire [31:0] p1_or_146894_comb;
  wire [31:0] p1_or_146897_comb;
  wire [31:0] p1_or_146904_comb;
  wire [31:0] p1_or_146907_comb;
  wire [31:0] p1_or_146914_comb;
  wire [31:0] p1_or_146917_comb;
  wire [31:0] p1_or_146924_comb;
  wire [31:0] p1_or_146927_comb;
  wire [31:0] p1_or_146934_comb;
  wire [31:0] p1_or_146937_comb;
  wire [31:0] p1_or_146944_comb;
  wire [31:0] p1_or_146947_comb;
  wire [31:0] p1_or_146954_comb;
  wire [31:0] p1_prod__525_comb;
  wire [31:0] p1_or_146961_comb;
  wire [31:0] p1_or_146964_comb;
  wire [31:0] p1_prod__556_comb;
  wire [31:0] p1_prod__589_comb;
  wire [31:0] p1_or_146975_comb;
  wire [31:0] p1_or_146978_comb;
  wire [31:0] p1_prod__620_comb;
  wire [31:0] p1_prod__653_comb;
  wire [31:0] p1_or_146989_comb;
  wire [31:0] p1_or_146992_comb;
  wire [31:0] p1_prod__684_comb;
  wire [31:0] p1_prod__717_comb;
  wire [31:0] p1_or_147003_comb;
  wire [31:0] p1_or_147006_comb;
  wire [31:0] p1_prod__748_comb;
  wire [31:0] p1_prod__781_comb;
  wire [31:0] p1_or_147017_comb;
  wire [31:0] p1_or_147020_comb;
  wire [31:0] p1_prod__812_comb;
  wire [31:0] p1_prod__845_comb;
  wire [31:0] p1_or_147031_comb;
  wire [31:0] p1_or_147034_comb;
  wire [31:0] p1_prod__876_comb;
  wire [31:0] p1_prod__909_comb;
  wire [31:0] p1_or_147045_comb;
  wire [31:0] p1_or_147048_comb;
  wire [31:0] p1_prod__940_comb;
  wire [31:0] p1_prod__973_comb;
  wire [31:0] p1_or_147059_comb;
  wire [31:0] p1_or_147062_comb;
  wire [31:0] p1_prod__1004_comb;
  wire [31:0] p1_or_147133_comb;
  wire [31:0] p1_prod__545_comb;
  wire [31:0] p1_prod__563_comb;
  wire [31:0] p1_or_147144_comb;
  wire [31:0] p1_or_147147_comb;
  wire [31:0] p1_prod__609_comb;
  wire [31:0] p1_prod__627_comb;
  wire [31:0] p1_or_147158_comb;
  wire [31:0] p1_or_147161_comb;
  wire [31:0] p1_prod__673_comb;
  wire [31:0] p1_prod__691_comb;
  wire [31:0] p1_or_147172_comb;
  wire [31:0] p1_or_147175_comb;
  wire [31:0] p1_prod__737_comb;
  wire [31:0] p1_prod__755_comb;
  wire [31:0] p1_or_147186_comb;
  wire [31:0] p1_or_147189_comb;
  wire [31:0] p1_prod__801_comb;
  wire [31:0] p1_prod__819_comb;
  wire [31:0] p1_or_147200_comb;
  wire [31:0] p1_or_147203_comb;
  wire [31:0] p1_prod__865_comb;
  wire [31:0] p1_prod__883_comb;
  wire [31:0] p1_or_147214_comb;
  wire [31:0] p1_or_147217_comb;
  wire [31:0] p1_prod__929_comb;
  wire [31:0] p1_prod__947_comb;
  wire [31:0] p1_or_147228_comb;
  wire [31:0] p1_or_147231_comb;
  wire [31:0] p1_prod__993_comb;
  wire [31:0] p1_prod__1011_comb;
  wire [31:0] p1_or_147242_comb;
  wire [31:0] p1_or_147247_comb;
  wire [31:0] p1_or_147252_comb;
  wire [31:0] p1_or_147255_comb;
  wire [31:0] p1_or_147260_comb;
  wire [31:0] p1_or_147267_comb;
  wire [31:0] p1_or_147272_comb;
  wire [31:0] p1_or_147275_comb;
  wire [31:0] p1_or_147280_comb;
  wire [31:0] p1_or_147287_comb;
  wire [31:0] p1_or_147292_comb;
  wire [31:0] p1_or_147295_comb;
  wire [31:0] p1_or_147300_comb;
  wire [31:0] p1_or_147307_comb;
  wire [31:0] p1_or_147312_comb;
  wire [31:0] p1_or_147315_comb;
  wire [31:0] p1_or_147320_comb;
  wire [31:0] p1_or_147327_comb;
  wire [31:0] p1_or_147332_comb;
  wire [31:0] p1_or_147335_comb;
  wire [31:0] p1_or_147340_comb;
  wire [31:0] p1_or_147347_comb;
  wire [31:0] p1_or_147352_comb;
  wire [31:0] p1_or_147355_comb;
  wire [31:0] p1_or_147360_comb;
  wire [31:0] p1_or_147367_comb;
  wire [31:0] p1_or_147372_comb;
  wire [31:0] p1_or_147375_comb;
  wire [31:0] p1_or_147380_comb;
  wire [31:0] p1_or_147387_comb;
  wire [31:0] p1_or_147392_comb;
  wire [31:0] p1_or_147395_comb;
  wire [31:0] p1_or_147400_comb;
  wire [31:0] p1_prod__547_comb;
  wire [31:0] p1_or_147407_comb;
  wire [31:0] p1_or_147414_comb;
  wire [31:0] p1_prod__575_comb;
  wire [31:0] p1_prod__611_comb;
  wire [31:0] p1_or_147421_comb;
  wire [31:0] p1_or_147428_comb;
  wire [31:0] p1_prod__639_comb;
  wire [31:0] p1_prod__675_comb;
  wire [31:0] p1_or_147435_comb;
  wire [31:0] p1_or_147442_comb;
  wire [31:0] p1_prod__703_comb;
  wire [31:0] p1_prod__739_comb;
  wire [31:0] p1_or_147449_comb;
  wire [31:0] p1_or_147456_comb;
  wire [31:0] p1_prod__767_comb;
  wire [31:0] p1_prod__803_comb;
  wire [31:0] p1_or_147463_comb;
  wire [31:0] p1_or_147470_comb;
  wire [31:0] p1_prod__831_comb;
  wire [31:0] p1_prod__867_comb;
  wire [31:0] p1_or_147477_comb;
  wire [31:0] p1_or_147484_comb;
  wire [31:0] p1_prod__895_comb;
  wire [31:0] p1_prod__931_comb;
  wire [31:0] p1_or_147491_comb;
  wire [31:0] p1_or_147498_comb;
  wire [31:0] p1_prod__959_comb;
  wire [31:0] p1_prod__995_comb;
  wire [31:0] p1_or_147505_comb;
  wire [31:0] p1_or_147512_comb;
  wire [31:0] p1_prod__1023_comb;
  wire [16:0] p1_smul_58222_NarrowedMult__comb;
  wire [16:0] p1_smul_58224_NarrowedMult__comb;
  wire [31:0] p1_or_147714_comb;
  wire [31:0] p1_or_147715_comb;
  wire [16:0] p1_smul_58234_NarrowedMult__comb;
  wire [16:0] p1_smul_58236_NarrowedMult__comb;
  wire [16:0] p1_smul_58238_NarrowedMult__comb;
  wire [16:0] p1_smul_58240_NarrowedMult__comb;
  wire [31:0] p1_or_147730_comb;
  wire [31:0] p1_or_147731_comb;
  wire [16:0] p1_smul_58250_NarrowedMult__comb;
  wire [16:0] p1_smul_58252_NarrowedMult__comb;
  wire [16:0] p1_smul_58254_NarrowedMult__comb;
  wire [16:0] p1_smul_58256_NarrowedMult__comb;
  wire [31:0] p1_or_147746_comb;
  wire [31:0] p1_or_147747_comb;
  wire [16:0] p1_smul_58266_NarrowedMult__comb;
  wire [16:0] p1_smul_58268_NarrowedMult__comb;
  wire [16:0] p1_smul_58270_NarrowedMult__comb;
  wire [16:0] p1_smul_58272_NarrowedMult__comb;
  wire [31:0] p1_or_147762_comb;
  wire [31:0] p1_or_147763_comb;
  wire [16:0] p1_smul_58282_NarrowedMult__comb;
  wire [16:0] p1_smul_58284_NarrowedMult__comb;
  wire [16:0] p1_smul_58286_NarrowedMult__comb;
  wire [16:0] p1_smul_58288_NarrowedMult__comb;
  wire [31:0] p1_or_147778_comb;
  wire [31:0] p1_or_147779_comb;
  wire [16:0] p1_smul_58298_NarrowedMult__comb;
  wire [16:0] p1_smul_58300_NarrowedMult__comb;
  wire [16:0] p1_smul_58302_NarrowedMult__comb;
  wire [16:0] p1_smul_58304_NarrowedMult__comb;
  wire [31:0] p1_or_147794_comb;
  wire [31:0] p1_or_147795_comb;
  wire [16:0] p1_smul_58314_NarrowedMult__comb;
  wire [16:0] p1_smul_58316_NarrowedMult__comb;
  wire [16:0] p1_smul_58318_NarrowedMult__comb;
  wire [16:0] p1_smul_58320_NarrowedMult__comb;
  wire [31:0] p1_or_147810_comb;
  wire [31:0] p1_or_147811_comb;
  wire [16:0] p1_smul_58330_NarrowedMult__comb;
  wire [16:0] p1_smul_58332_NarrowedMult__comb;
  wire [16:0] p1_smul_58334_NarrowedMult__comb;
  wire [16:0] p1_smul_58336_NarrowedMult__comb;
  wire [31:0] p1_or_147826_comb;
  wire [31:0] p1_or_147827_comb;
  wire [16:0] p1_smul_58346_NarrowedMult__comb;
  wire [16:0] p1_smul_58348_NarrowedMult__comb;
  wire [16:0] p1_smul_58478_NarrowedMult__comb;
  wire [31:0] p1_or_147997_comb;
  wire [16:0] p1_smul_58482_NarrowedMult__comb;
  wire [16:0] p1_smul_58488_NarrowedMult__comb;
  wire [31:0] p1_or_148008_comb;
  wire [16:0] p1_smul_58492_NarrowedMult__comb;
  wire [16:0] p1_smul_58494_NarrowedMult__comb;
  wire [31:0] p1_or_148013_comb;
  wire [16:0] p1_smul_58498_NarrowedMult__comb;
  wire [16:0] p1_smul_58504_NarrowedMult__comb;
  wire [31:0] p1_or_148024_comb;
  wire [16:0] p1_smul_58508_NarrowedMult__comb;
  wire [16:0] p1_smul_58510_NarrowedMult__comb;
  wire [31:0] p1_or_148029_comb;
  wire [16:0] p1_smul_58514_NarrowedMult__comb;
  wire [16:0] p1_smul_58520_NarrowedMult__comb;
  wire [31:0] p1_or_148040_comb;
  wire [16:0] p1_smul_58524_NarrowedMult__comb;
  wire [16:0] p1_smul_58526_NarrowedMult__comb;
  wire [31:0] p1_or_148045_comb;
  wire [16:0] p1_smul_58530_NarrowedMult__comb;
  wire [16:0] p1_smul_58536_NarrowedMult__comb;
  wire [31:0] p1_or_148056_comb;
  wire [16:0] p1_smul_58540_NarrowedMult__comb;
  wire [16:0] p1_smul_58542_NarrowedMult__comb;
  wire [31:0] p1_or_148061_comb;
  wire [16:0] p1_smul_58546_NarrowedMult__comb;
  wire [16:0] p1_smul_58552_NarrowedMult__comb;
  wire [31:0] p1_or_148072_comb;
  wire [16:0] p1_smul_58556_NarrowedMult__comb;
  wire [16:0] p1_smul_58558_NarrowedMult__comb;
  wire [31:0] p1_or_148077_comb;
  wire [16:0] p1_smul_58562_NarrowedMult__comb;
  wire [16:0] p1_smul_58568_NarrowedMult__comb;
  wire [31:0] p1_or_148088_comb;
  wire [16:0] p1_smul_58572_NarrowedMult__comb;
  wire [16:0] p1_smul_58574_NarrowedMult__comb;
  wire [31:0] p1_or_148093_comb;
  wire [16:0] p1_smul_58578_NarrowedMult__comb;
  wire [16:0] p1_smul_58584_NarrowedMult__comb;
  wire [31:0] p1_or_148104_comb;
  wire [16:0] p1_smul_58588_NarrowedMult__comb;
  wire [16:0] p1_smul_58590_NarrowedMult__comb;
  wire [31:0] p1_or_148109_comb;
  wire [16:0] p1_smul_58594_NarrowedMult__comb;
  wire [16:0] p1_smul_58600_NarrowedMult__comb;
  wire [31:0] p1_or_148120_comb;
  wire [16:0] p1_smul_58604_NarrowedMult__comb;
  wire [16:0] p1_smul_58606_NarrowedMult__comb;
  wire [16:0] p1_smul_58608_NarrowedMult__comb;
  wire [16:0] p1_smul_58610_NarrowedMult__comb;
  wire [16:0] p1_smul_58612_NarrowedMult__comb;
  wire [16:0] p1_smul_58614_NarrowedMult__comb;
  wire [16:0] p1_smul_58616_NarrowedMult__comb;
  wire [16:0] p1_smul_58618_NarrowedMult__comb;
  wire [16:0] p1_smul_58620_NarrowedMult__comb;
  wire [16:0] p1_smul_58622_NarrowedMult__comb;
  wire [16:0] p1_smul_58624_NarrowedMult__comb;
  wire [16:0] p1_smul_58626_NarrowedMult__comb;
  wire [16:0] p1_smul_58628_NarrowedMult__comb;
  wire [16:0] p1_smul_58630_NarrowedMult__comb;
  wire [16:0] p1_smul_58632_NarrowedMult__comb;
  wire [16:0] p1_smul_58634_NarrowedMult__comb;
  wire [16:0] p1_smul_58636_NarrowedMult__comb;
  wire [16:0] p1_smul_58638_NarrowedMult__comb;
  wire [16:0] p1_smul_58640_NarrowedMult__comb;
  wire [16:0] p1_smul_58642_NarrowedMult__comb;
  wire [16:0] p1_smul_58644_NarrowedMult__comb;
  wire [16:0] p1_smul_58646_NarrowedMult__comb;
  wire [16:0] p1_smul_58648_NarrowedMult__comb;
  wire [16:0] p1_smul_58650_NarrowedMult__comb;
  wire [16:0] p1_smul_58652_NarrowedMult__comb;
  wire [16:0] p1_smul_58654_NarrowedMult__comb;
  wire [16:0] p1_smul_58656_NarrowedMult__comb;
  wire [16:0] p1_smul_58658_NarrowedMult__comb;
  wire [16:0] p1_smul_58660_NarrowedMult__comb;
  wire [16:0] p1_smul_58662_NarrowedMult__comb;
  wire [16:0] p1_smul_58664_NarrowedMult__comb;
  wire [16:0] p1_smul_58666_NarrowedMult__comb;
  wire [16:0] p1_smul_58668_NarrowedMult__comb;
  wire [16:0] p1_smul_58670_NarrowedMult__comb;
  wire [16:0] p1_smul_58672_NarrowedMult__comb;
  wire [16:0] p1_smul_58674_NarrowedMult__comb;
  wire [16:0] p1_smul_58676_NarrowedMult__comb;
  wire [16:0] p1_smul_58678_NarrowedMult__comb;
  wire [16:0] p1_smul_58680_NarrowedMult__comb;
  wire [16:0] p1_smul_58682_NarrowedMult__comb;
  wire [16:0] p1_smul_58684_NarrowedMult__comb;
  wire [16:0] p1_smul_58686_NarrowedMult__comb;
  wire [16:0] p1_smul_58688_NarrowedMult__comb;
  wire [16:0] p1_smul_58690_NarrowedMult__comb;
  wire [16:0] p1_smul_58692_NarrowedMult__comb;
  wire [16:0] p1_smul_58694_NarrowedMult__comb;
  wire [16:0] p1_smul_58696_NarrowedMult__comb;
  wire [16:0] p1_smul_58698_NarrowedMult__comb;
  wire [16:0] p1_smul_58700_NarrowedMult__comb;
  wire [16:0] p1_smul_58702_NarrowedMult__comb;
  wire [16:0] p1_smul_58704_NarrowedMult__comb;
  wire [16:0] p1_smul_58706_NarrowedMult__comb;
  wire [16:0] p1_smul_58708_NarrowedMult__comb;
  wire [16:0] p1_smul_58710_NarrowedMult__comb;
  wire [16:0] p1_smul_58712_NarrowedMult__comb;
  wire [16:0] p1_smul_58714_NarrowedMult__comb;
  wire [16:0] p1_smul_58716_NarrowedMult__comb;
  wire [16:0] p1_smul_58718_NarrowedMult__comb;
  wire [16:0] p1_smul_58720_NarrowedMult__comb;
  wire [16:0] p1_smul_58722_NarrowedMult__comb;
  wire [16:0] p1_smul_58724_NarrowedMult__comb;
  wire [16:0] p1_smul_58726_NarrowedMult__comb;
  wire [16:0] p1_smul_58728_NarrowedMult__comb;
  wire [16:0] p1_smul_58730_NarrowedMult__comb;
  wire [16:0] p1_smul_58732_NarrowedMult__comb;
  wire [16:0] p1_smul_58736_NarrowedMult__comb;
  wire [31:0] p1_or_148256_comb;
  wire [16:0] p1_smul_58740_NarrowedMult__comb;
  wire [16:0] p1_smul_58742_NarrowedMult__comb;
  wire [31:0] p1_or_148261_comb;
  wire [16:0] p1_smul_58746_NarrowedMult__comb;
  wire [16:0] p1_smul_58752_NarrowedMult__comb;
  wire [31:0] p1_or_148272_comb;
  wire [16:0] p1_smul_58756_NarrowedMult__comb;
  wire [16:0] p1_smul_58758_NarrowedMult__comb;
  wire [31:0] p1_or_148277_comb;
  wire [16:0] p1_smul_58762_NarrowedMult__comb;
  wire [16:0] p1_smul_58768_NarrowedMult__comb;
  wire [31:0] p1_or_148288_comb;
  wire [16:0] p1_smul_58772_NarrowedMult__comb;
  wire [16:0] p1_smul_58774_NarrowedMult__comb;
  wire [31:0] p1_or_148293_comb;
  wire [16:0] p1_smul_58778_NarrowedMult__comb;
  wire [16:0] p1_smul_58784_NarrowedMult__comb;
  wire [31:0] p1_or_148304_comb;
  wire [16:0] p1_smul_58788_NarrowedMult__comb;
  wire [16:0] p1_smul_58790_NarrowedMult__comb;
  wire [31:0] p1_or_148309_comb;
  wire [16:0] p1_smul_58794_NarrowedMult__comb;
  wire [16:0] p1_smul_58800_NarrowedMult__comb;
  wire [31:0] p1_or_148320_comb;
  wire [16:0] p1_smul_58804_NarrowedMult__comb;
  wire [16:0] p1_smul_58806_NarrowedMult__comb;
  wire [31:0] p1_or_148325_comb;
  wire [16:0] p1_smul_58810_NarrowedMult__comb;
  wire [16:0] p1_smul_58816_NarrowedMult__comb;
  wire [31:0] p1_or_148336_comb;
  wire [16:0] p1_smul_58820_NarrowedMult__comb;
  wire [16:0] p1_smul_58822_NarrowedMult__comb;
  wire [31:0] p1_or_148341_comb;
  wire [16:0] p1_smul_58826_NarrowedMult__comb;
  wire [16:0] p1_smul_58832_NarrowedMult__comb;
  wire [31:0] p1_or_148352_comb;
  wire [16:0] p1_smul_58836_NarrowedMult__comb;
  wire [16:0] p1_smul_58838_NarrowedMult__comb;
  wire [31:0] p1_or_148357_comb;
  wire [16:0] p1_smul_58842_NarrowedMult__comb;
  wire [16:0] p1_smul_58848_NarrowedMult__comb;
  wire [31:0] p1_or_148368_comb;
  wire [16:0] p1_smul_58852_NarrowedMult__comb;
  wire [16:0] p1_smul_58854_NarrowedMult__comb;
  wire [31:0] p1_or_148373_comb;
  wire [16:0] p1_smul_58858_NarrowedMult__comb;
  wire [31:0] p1_or_148539_comb;
  wire [16:0] p1_smul_58994_NarrowedMult__comb;
  wire [16:0] p1_smul_58996_NarrowedMult__comb;
  wire [16:0] p1_smul_58998_NarrowedMult__comb;
  wire [16:0] p1_smul_59000_NarrowedMult__comb;
  wire [31:0] p1_or_148554_comb;
  wire [31:0] p1_or_148555_comb;
  wire [16:0] p1_smul_59010_NarrowedMult__comb;
  wire [16:0] p1_smul_59012_NarrowedMult__comb;
  wire [16:0] p1_smul_59014_NarrowedMult__comb;
  wire [16:0] p1_smul_59016_NarrowedMult__comb;
  wire [31:0] p1_or_148570_comb;
  wire [31:0] p1_or_148571_comb;
  wire [16:0] p1_smul_59026_NarrowedMult__comb;
  wire [16:0] p1_smul_59028_NarrowedMult__comb;
  wire [16:0] p1_smul_59030_NarrowedMult__comb;
  wire [16:0] p1_smul_59032_NarrowedMult__comb;
  wire [31:0] p1_or_148586_comb;
  wire [31:0] p1_or_148587_comb;
  wire [16:0] p1_smul_59042_NarrowedMult__comb;
  wire [16:0] p1_smul_59044_NarrowedMult__comb;
  wire [16:0] p1_smul_59046_NarrowedMult__comb;
  wire [16:0] p1_smul_59048_NarrowedMult__comb;
  wire [31:0] p1_or_148602_comb;
  wire [31:0] p1_or_148603_comb;
  wire [16:0] p1_smul_59058_NarrowedMult__comb;
  wire [16:0] p1_smul_59060_NarrowedMult__comb;
  wire [16:0] p1_smul_59062_NarrowedMult__comb;
  wire [16:0] p1_smul_59064_NarrowedMult__comb;
  wire [31:0] p1_or_148618_comb;
  wire [31:0] p1_or_148619_comb;
  wire [16:0] p1_smul_59074_NarrowedMult__comb;
  wire [16:0] p1_smul_59076_NarrowedMult__comb;
  wire [16:0] p1_smul_59078_NarrowedMult__comb;
  wire [16:0] p1_smul_59080_NarrowedMult__comb;
  wire [31:0] p1_or_148634_comb;
  wire [31:0] p1_or_148635_comb;
  wire [16:0] p1_smul_59090_NarrowedMult__comb;
  wire [16:0] p1_smul_59092_NarrowedMult__comb;
  wire [16:0] p1_smul_59094_NarrowedMult__comb;
  wire [16:0] p1_smul_59096_NarrowedMult__comb;
  wire [31:0] p1_or_148650_comb;
  wire [31:0] p1_or_148651_comb;
  wire [16:0] p1_smul_59106_NarrowedMult__comb;
  wire [16:0] p1_smul_59108_NarrowedMult__comb;
  wire [16:0] p1_smul_59110_NarrowedMult__comb;
  wire [16:0] p1_smul_59112_NarrowedMult__comb;
  wire [31:0] p1_or_148666_comb;
  wire [15:0] p1_sel_148667_comb;
  wire [15:0] p1_sel_148668_comb;
  wire [15:0] p1_sel_148669_comb;
  wire [15:0] p1_sel_148670_comb;
  wire [15:0] p1_sel_148671_comb;
  wire [15:0] p1_sel_148672_comb;
  wire [15:0] p1_sel_148673_comb;
  wire [15:0] p1_sel_148674_comb;
  wire [15:0] p1_sel_148675_comb;
  wire [15:0] p1_sel_148676_comb;
  wire [15:0] p1_sel_148677_comb;
  wire [15:0] p1_sel_148678_comb;
  wire [15:0] p1_sel_148679_comb;
  wire [15:0] p1_sel_148680_comb;
  wire [15:0] p1_sel_148681_comb;
  wire [15:0] p1_sel_148682_comb;
  wire [15:0] p1_sel_148683_comb;
  wire [15:0] p1_sel_148684_comb;
  wire [15:0] p1_sel_148685_comb;
  wire [15:0] p1_sel_148686_comb;
  wire [15:0] p1_sel_148687_comb;
  wire [15:0] p1_sel_148688_comb;
  wire [15:0] p1_sel_148689_comb;
  wire [15:0] p1_sel_148690_comb;
  wire [15:0] p1_sel_148691_comb;
  wire [15:0] p1_sel_148692_comb;
  wire [15:0] p1_sel_148693_comb;
  wire [15:0] p1_sel_148694_comb;
  wire [15:0] p1_sel_148695_comb;
  wire [15:0] p1_sel_148696_comb;
  wire [15:0] p1_sel_148697_comb;
  wire [15:0] p1_sel_148698_comb;
  wire [15:0] p1_sel_148699_comb;
  wire [15:0] p1_sel_148700_comb;
  wire [15:0] p1_sel_148701_comb;
  wire [15:0] p1_sel_148702_comb;
  wire [15:0] p1_sel_148703_comb;
  wire [15:0] p1_sel_148704_comb;
  wire [15:0] p1_sel_148705_comb;
  wire [15:0] p1_sel_148706_comb;
  wire [15:0] p1_sel_148707_comb;
  wire [15:0] p1_sel_148708_comb;
  wire [15:0] p1_sel_148709_comb;
  wire [15:0] p1_sel_148710_comb;
  wire [15:0] p1_sel_148711_comb;
  wire [15:0] p1_sel_148712_comb;
  wire [15:0] p1_sel_148713_comb;
  wire [15:0] p1_sel_148714_comb;
  wire [15:0] p1_sel_148715_comb;
  wire [15:0] p1_sel_148716_comb;
  wire [15:0] p1_sel_148717_comb;
  wire [15:0] p1_sel_148718_comb;
  wire [15:0] p1_sel_148719_comb;
  wire [15:0] p1_sel_148720_comb;
  wire [15:0] p1_sel_148721_comb;
  wire [15:0] p1_sel_148722_comb;
  wire [15:0] p1_sel_148723_comb;
  wire [15:0] p1_sel_148724_comb;
  wire [15:0] p1_sel_148725_comb;
  wire [15:0] p1_sel_148726_comb;
  wire [15:0] p1_sel_148727_comb;
  wire [15:0] p1_sel_148728_comb;
  wire [15:0] p1_sel_148729_comb;
  wire [15:0] p1_sel_148730_comb;
  wire [16:0] p1_add_151931_comb;
  wire [16:0] p1_add_151932_comb;
  wire [16:0] p1_add_151933_comb;
  wire [16:0] p1_add_151934_comb;
  wire [16:0] p1_add_151935_comb;
  wire [16:0] p1_add_151936_comb;
  wire [16:0] p1_add_151937_comb;
  wire [16:0] p1_add_151938_comb;
  wire [16:0] p1_add_151939_comb;
  wire [16:0] p1_add_151940_comb;
  wire [16:0] p1_add_151941_comb;
  wire [16:0] p1_add_151942_comb;
  wire [16:0] p1_add_151943_comb;
  wire [16:0] p1_add_151944_comb;
  wire [16:0] p1_add_151945_comb;
  wire [16:0] p1_add_151946_comb;
  wire [16:0] p1_add_151947_comb;
  wire [16:0] p1_add_151948_comb;
  wire [16:0] p1_add_151949_comb;
  wire [16:0] p1_add_151950_comb;
  wire [16:0] p1_add_151951_comb;
  wire [16:0] p1_add_151952_comb;
  wire [16:0] p1_add_151953_comb;
  wire [16:0] p1_add_151954_comb;
  wire [16:0] p1_add_151955_comb;
  wire [16:0] p1_add_151956_comb;
  wire [16:0] p1_add_151957_comb;
  wire [16:0] p1_add_151958_comb;
  wire [16:0] p1_add_151959_comb;
  wire [16:0] p1_add_151960_comb;
  wire [16:0] p1_add_151961_comb;
  wire [16:0] p1_add_151962_comb;
  wire [15:0] p1_sel_151963_comb;
  wire [15:0] p1_sel_151964_comb;
  wire [15:0] p1_sel_151965_comb;
  wire [15:0] p1_sel_151966_comb;
  wire [15:0] p1_sel_151967_comb;
  wire [15:0] p1_sel_151968_comb;
  wire [15:0] p1_sel_151969_comb;
  wire [15:0] p1_sel_151970_comb;
  wire [15:0] p1_sel_151971_comb;
  wire [15:0] p1_sel_151972_comb;
  wire [15:0] p1_sel_151973_comb;
  wire [15:0] p1_sel_151974_comb;
  wire [15:0] p1_sel_151975_comb;
  wire [15:0] p1_sel_151976_comb;
  wire [15:0] p1_sel_151977_comb;
  wire [15:0] p1_sel_151978_comb;
  wire [15:0] p1_sel_151979_comb;
  wire [15:0] p1_sel_151980_comb;
  wire [15:0] p1_sel_151981_comb;
  wire [15:0] p1_sel_151982_comb;
  wire [15:0] p1_sel_151983_comb;
  wire [15:0] p1_sel_151984_comb;
  wire [15:0] p1_sel_151985_comb;
  wire [15:0] p1_sel_151986_comb;
  wire [15:0] p1_sel_151987_comb;
  wire [15:0] p1_sel_151988_comb;
  wire [15:0] p1_sel_151989_comb;
  wire [15:0] p1_sel_151990_comb;
  wire [15:0] p1_sel_151991_comb;
  wire [15:0] p1_sel_151992_comb;
  wire [15:0] p1_sel_151993_comb;
  wire [15:0] p1_sel_151994_comb;
  wire [15:0] p1_sel_151995_comb;
  wire [15:0] p1_sel_151996_comb;
  wire [15:0] p1_sel_151997_comb;
  wire [15:0] p1_sel_151998_comb;
  wire [15:0] p1_sel_151999_comb;
  wire [15:0] p1_sel_152000_comb;
  wire [15:0] p1_sel_152001_comb;
  wire [15:0] p1_sel_152002_comb;
  wire [15:0] p1_sel_152003_comb;
  wire [15:0] p1_sel_152004_comb;
  wire [15:0] p1_sel_152005_comb;
  wire [15:0] p1_sel_152006_comb;
  wire [15:0] p1_sel_152007_comb;
  wire [15:0] p1_sel_152008_comb;
  wire [15:0] p1_sel_152009_comb;
  wire [15:0] p1_sel_152010_comb;
  wire [15:0] p1_sel_152011_comb;
  wire [15:0] p1_sel_152012_comb;
  wire [15:0] p1_sel_152013_comb;
  wire [15:0] p1_sel_152014_comb;
  wire [15:0] p1_sel_152015_comb;
  wire [15:0] p1_sel_152016_comb;
  wire [15:0] p1_sel_152017_comb;
  wire [15:0] p1_sel_152018_comb;
  wire [15:0] p1_sel_152019_comb;
  wire [15:0] p1_sel_152020_comb;
  wire [15:0] p1_sel_152021_comb;
  wire [15:0] p1_sel_152022_comb;
  wire [15:0] p1_sel_152023_comb;
  wire [15:0] p1_sel_152024_comb;
  wire [15:0] p1_sel_152025_comb;
  wire [15:0] p1_sel_152026_comb;
  wire [15:0] p1_sel_152027_comb;
  wire [15:0] p1_sel_152028_comb;
  wire [15:0] p1_sel_152029_comb;
  wire [15:0] p1_sel_152030_comb;
  wire [15:0] p1_sel_152031_comb;
  wire [15:0] p1_sel_152032_comb;
  wire [15:0] p1_sel_152033_comb;
  wire [15:0] p1_sel_152034_comb;
  wire [15:0] p1_sel_152035_comb;
  wire [15:0] p1_sel_152036_comb;
  wire [15:0] p1_sel_152037_comb;
  wire [15:0] p1_sel_152038_comb;
  wire [15:0] p1_sel_152039_comb;
  wire [15:0] p1_sel_152040_comb;
  wire [15:0] p1_sel_152041_comb;
  wire [15:0] p1_sel_152042_comb;
  wire [15:0] p1_sel_152043_comb;
  wire [15:0] p1_sel_152044_comb;
  wire [15:0] p1_sel_152045_comb;
  wire [15:0] p1_sel_152046_comb;
  wire [15:0] p1_sel_152047_comb;
  wire [15:0] p1_sel_152048_comb;
  wire [15:0] p1_sel_152049_comb;
  wire [15:0] p1_sel_152050_comb;
  wire [15:0] p1_sel_152051_comb;
  wire [15:0] p1_sel_152052_comb;
  wire [15:0] p1_sel_152053_comb;
  wire [15:0] p1_sel_152054_comb;
  wire [15:0] p1_sel_152055_comb;
  wire [15:0] p1_sel_152056_comb;
  wire [15:0] p1_sel_152057_comb;
  wire [15:0] p1_sel_152058_comb;
  wire [15:0] p1_sel_152059_comb;
  wire [15:0] p1_sel_152060_comb;
  wire [15:0] p1_sel_152061_comb;
  wire [15:0] p1_sel_152062_comb;
  wire [15:0] p1_sel_152063_comb;
  wire [15:0] p1_sel_152064_comb;
  wire [15:0] p1_sel_152065_comb;
  wire [15:0] p1_sel_152066_comb;
  wire [15:0] p1_sel_152067_comb;
  wire [15:0] p1_sel_152068_comb;
  wire [15:0] p1_sel_152069_comb;
  wire [15:0] p1_sel_152070_comb;
  wire [15:0] p1_sel_152071_comb;
  wire [15:0] p1_sel_152072_comb;
  wire [15:0] p1_sel_152073_comb;
  wire [15:0] p1_sel_152074_comb;
  wire [15:0] p1_sel_152075_comb;
  wire [15:0] p1_sel_152076_comb;
  wire [15:0] p1_sel_152077_comb;
  wire [15:0] p1_sel_152078_comb;
  wire [15:0] p1_sel_152079_comb;
  wire [15:0] p1_sel_152080_comb;
  wire [15:0] p1_sel_152081_comb;
  wire [15:0] p1_sel_152082_comb;
  wire [15:0] p1_sel_152083_comb;
  wire [15:0] p1_sel_152084_comb;
  wire [15:0] p1_sel_152085_comb;
  wire [15:0] p1_sel_152086_comb;
  wire [15:0] p1_sel_152087_comb;
  wire [15:0] p1_sel_152088_comb;
  wire [15:0] p1_sel_152089_comb;
  wire [15:0] p1_sel_152090_comb;
  wire [15:0] p1_sel_152091_comb;
  wire [15:0] p1_sel_152092_comb;
  wire [15:0] p1_sel_152093_comb;
  wire [15:0] p1_sel_152094_comb;
  wire [15:0] p1_sel_152095_comb;
  wire [15:0] p1_sel_152096_comb;
  wire [15:0] p1_sel_152097_comb;
  wire [15:0] p1_sel_152098_comb;
  wire [15:0] p1_sel_152099_comb;
  wire [15:0] p1_sel_152100_comb;
  wire [15:0] p1_sel_152101_comb;
  wire [15:0] p1_sel_152102_comb;
  wire [15:0] p1_sel_152103_comb;
  wire [15:0] p1_sel_152104_comb;
  wire [15:0] p1_sel_152105_comb;
  wire [15:0] p1_sel_152106_comb;
  wire [15:0] p1_sel_152107_comb;
  wire [15:0] p1_sel_152108_comb;
  wire [15:0] p1_sel_152109_comb;
  wire [15:0] p1_sel_152110_comb;
  wire [15:0] p1_sel_152111_comb;
  wire [15:0] p1_sel_152112_comb;
  wire [15:0] p1_sel_152113_comb;
  wire [15:0] p1_sel_152114_comb;
  wire [15:0] p1_sel_152115_comb;
  wire [15:0] p1_sel_152116_comb;
  wire [15:0] p1_sel_152117_comb;
  wire [15:0] p1_sel_152118_comb;
  wire [15:0] p1_sel_152119_comb;
  wire [15:0] p1_sel_152120_comb;
  wire [15:0] p1_sel_152121_comb;
  wire [15:0] p1_sel_152122_comb;
  wire [15:0] p1_sel_152123_comb;
  wire [15:0] p1_sel_152124_comb;
  wire [15:0] p1_sel_152125_comb;
  wire [15:0] p1_sel_152126_comb;
  wire [15:0] p1_sel_152127_comb;
  wire [15:0] p1_sel_152128_comb;
  wire [15:0] p1_sel_152129_comb;
  wire [15:0] p1_sel_152130_comb;
  wire [15:0] p1_sel_152131_comb;
  wire [15:0] p1_sel_152132_comb;
  wire [15:0] p1_sel_152133_comb;
  wire [15:0] p1_sel_152134_comb;
  wire [15:0] p1_sel_152135_comb;
  wire [15:0] p1_sel_152136_comb;
  wire [15:0] p1_sel_152137_comb;
  wire [15:0] p1_sel_152138_comb;
  wire [15:0] p1_sel_152139_comb;
  wire [15:0] p1_sel_152140_comb;
  wire [15:0] p1_sel_152141_comb;
  wire [15:0] p1_sel_152142_comb;
  wire [15:0] p1_sel_152143_comb;
  wire [15:0] p1_sel_152144_comb;
  wire [15:0] p1_sel_152145_comb;
  wire [15:0] p1_sel_152146_comb;
  wire [15:0] p1_sel_152147_comb;
  wire [15:0] p1_sel_152148_comb;
  wire [15:0] p1_sel_152149_comb;
  wire [15:0] p1_sel_152150_comb;
  wire [15:0] p1_sel_152151_comb;
  wire [15:0] p1_sel_152152_comb;
  wire [15:0] p1_sel_152153_comb;
  wire [15:0] p1_sel_152154_comb;
  wire [15:0] p1_sel_152155_comb;
  wire [15:0] p1_sel_152156_comb;
  wire [15:0] p1_sel_152157_comb;
  wire [15:0] p1_sel_152158_comb;
  wire [15:0] p1_sel_152159_comb;
  wire [15:0] p1_sel_152160_comb;
  wire [15:0] p1_sel_152161_comb;
  wire [15:0] p1_sel_152162_comb;
  wire [15:0] p1_sel_152163_comb;
  wire [15:0] p1_sel_152164_comb;
  wire [15:0] p1_sel_152165_comb;
  wire [15:0] p1_sel_152166_comb;
  wire [15:0] p1_sel_152167_comb;
  wire [15:0] p1_sel_152168_comb;
  wire [15:0] p1_sel_152169_comb;
  wire [15:0] p1_sel_152170_comb;
  wire [15:0] p1_sel_152171_comb;
  wire [15:0] p1_sel_152172_comb;
  wire [15:0] p1_sel_152173_comb;
  wire [15:0] p1_sel_152174_comb;
  wire [15:0] p1_sel_152175_comb;
  wire [15:0] p1_sel_152176_comb;
  wire [15:0] p1_sel_152177_comb;
  wire [15:0] p1_sel_152178_comb;
  wire [15:0] p1_sel_152179_comb;
  wire [15:0] p1_sel_152180_comb;
  wire [15:0] p1_sel_152181_comb;
  wire [15:0] p1_sel_152182_comb;
  wire [15:0] p1_sel_152183_comb;
  wire [15:0] p1_sel_152184_comb;
  wire [15:0] p1_sel_152185_comb;
  wire [15:0] p1_sel_152186_comb;
  wire [15:0] p1_sel_152187_comb;
  wire [15:0] p1_sel_152188_comb;
  wire [15:0] p1_sel_152189_comb;
  wire [15:0] p1_sel_152190_comb;
  wire [15:0] p1_sel_152191_comb;
  wire [15:0] p1_sel_152192_comb;
  wire [15:0] p1_sel_152193_comb;
  wire [15:0] p1_sel_152194_comb;
  wire [15:0] p1_sel_152195_comb;
  wire [15:0] p1_sel_152196_comb;
  wire [15:0] p1_sel_152197_comb;
  wire [15:0] p1_sel_152198_comb;
  wire [15:0] p1_sel_152199_comb;
  wire [15:0] p1_sel_152200_comb;
  wire [15:0] p1_sel_152201_comb;
  wire [15:0] p1_sel_152202_comb;
  wire [15:0] p1_sel_152203_comb;
  wire [15:0] p1_sel_152204_comb;
  wire [15:0] p1_sel_152205_comb;
  wire [15:0] p1_sel_152206_comb;
  wire [15:0] p1_sel_152207_comb;
  wire [15:0] p1_sel_152208_comb;
  wire [15:0] p1_sel_152209_comb;
  wire [15:0] p1_sel_152210_comb;
  wire [15:0] p1_sel_152211_comb;
  wire [15:0] p1_sel_152212_comb;
  wire [15:0] p1_sel_152213_comb;
  wire [15:0] p1_sel_152214_comb;
  wire [15:0] p1_sel_152215_comb;
  wire [15:0] p1_sel_152216_comb;
  wire [15:0] p1_sel_152217_comb;
  wire [15:0] p1_sel_152218_comb;
  wire [15:0] p1_sel_152219_comb;
  wire [15:0] p1_sel_152220_comb;
  wire [15:0] p1_sel_152221_comb;
  wire [15:0] p1_sel_152222_comb;
  wire [15:0] p1_sel_152223_comb;
  wire [15:0] p1_sel_152224_comb;
  wire [15:0] p1_sel_152225_comb;
  wire [15:0] p1_sel_152226_comb;
  wire [15:0] p1_sel_152227_comb;
  wire [15:0] p1_sel_152228_comb;
  wire [15:0] p1_sel_152229_comb;
  wire [15:0] p1_sel_152230_comb;
  wire [15:0] p1_sel_152231_comb;
  wire [15:0] p1_sel_152232_comb;
  wire [15:0] p1_sel_152233_comb;
  wire [15:0] p1_sel_152234_comb;
  wire [15:0] p1_sel_152235_comb;
  wire [15:0] p1_sel_152236_comb;
  wire [15:0] p1_sel_152237_comb;
  wire [15:0] p1_sel_152238_comb;
  wire [15:0] p1_sel_152239_comb;
  wire [15:0] p1_sel_152240_comb;
  wire [15:0] p1_sel_152241_comb;
  wire [15:0] p1_sel_152242_comb;
  wire [15:0] p1_sel_152243_comb;
  wire [15:0] p1_sel_152244_comb;
  wire [15:0] p1_sel_152245_comb;
  wire [15:0] p1_sel_152246_comb;
  wire [15:0] p1_sel_152247_comb;
  wire [15:0] p1_sel_152248_comb;
  wire [15:0] p1_sel_152249_comb;
  wire [15:0] p1_sel_152250_comb;
  wire [15:0] p1_sel_152251_comb;
  wire [15:0] p1_sel_152252_comb;
  wire [15:0] p1_sel_152253_comb;
  wire [15:0] p1_sel_152254_comb;
  wire [15:0] p1_sel_152255_comb;
  wire [15:0] p1_sel_152256_comb;
  wire [15:0] p1_sel_152257_comb;
  wire [15:0] p1_sel_152258_comb;
  wire [15:0] p1_sel_152259_comb;
  wire [15:0] p1_sel_152260_comb;
  wire [15:0] p1_sel_152261_comb;
  wire [15:0] p1_sel_152262_comb;
  wire [15:0] p1_sel_152263_comb;
  wire [15:0] p1_sel_152264_comb;
  wire [15:0] p1_sel_152265_comb;
  wire [15:0] p1_sel_152266_comb;
  wire [15:0] p1_sel_152267_comb;
  wire [15:0] p1_sel_152268_comb;
  wire [15:0] p1_sel_152269_comb;
  wire [15:0] p1_sel_152270_comb;
  wire [15:0] p1_sel_152271_comb;
  wire [15:0] p1_sel_152272_comb;
  wire [15:0] p1_sel_152273_comb;
  wire [15:0] p1_sel_152274_comb;
  wire [15:0] p1_sel_152275_comb;
  wire [15:0] p1_sel_152276_comb;
  wire [15:0] p1_sel_152277_comb;
  wire [15:0] p1_sel_152278_comb;
  wire [15:0] p1_sel_152279_comb;
  wire [15:0] p1_sel_152280_comb;
  wire [15:0] p1_sel_152281_comb;
  wire [15:0] p1_sel_152282_comb;
  wire [15:0] p1_sel_152283_comb;
  wire [15:0] p1_sel_152284_comb;
  wire [15:0] p1_sel_152285_comb;
  wire [15:0] p1_sel_152286_comb;
  wire [15:0] p1_sel_152287_comb;
  wire [15:0] p1_sel_152288_comb;
  wire [15:0] p1_sel_152289_comb;
  wire [15:0] p1_sel_152290_comb;
  wire [15:0] p1_sel_152291_comb;
  wire [15:0] p1_sel_152292_comb;
  wire [15:0] p1_sel_152293_comb;
  wire [15:0] p1_sel_152294_comb;
  wire [15:0] p1_sel_152295_comb;
  wire [15:0] p1_sel_152296_comb;
  wire [15:0] p1_sel_152297_comb;
  wire [15:0] p1_sel_152298_comb;
  wire [15:0] p1_sel_152299_comb;
  wire [15:0] p1_sel_152300_comb;
  wire [15:0] p1_sel_152301_comb;
  wire [15:0] p1_sel_152302_comb;
  wire [15:0] p1_sel_152303_comb;
  wire [15:0] p1_sel_152304_comb;
  wire [15:0] p1_sel_152305_comb;
  wire [15:0] p1_sel_152306_comb;
  wire [15:0] p1_sel_152307_comb;
  wire [15:0] p1_sel_152308_comb;
  wire [15:0] p1_sel_152309_comb;
  wire [15:0] p1_sel_152310_comb;
  wire [15:0] p1_sel_152311_comb;
  wire [15:0] p1_sel_152312_comb;
  wire [15:0] p1_sel_152313_comb;
  wire [15:0] p1_sel_152314_comb;
  wire [15:0] p1_sel_152315_comb;
  wire [15:0] p1_sel_152316_comb;
  wire [15:0] p1_sel_152317_comb;
  wire [15:0] p1_sel_152318_comb;
  wire [15:0] p1_sel_152319_comb;
  wire [15:0] p1_sel_152320_comb;
  wire [15:0] p1_sel_152321_comb;
  wire [15:0] p1_sel_152322_comb;
  wire [15:0] p1_sel_152323_comb;
  wire [15:0] p1_sel_152324_comb;
  wire [15:0] p1_sel_152325_comb;
  wire [15:0] p1_sel_152326_comb;
  wire [15:0] p1_sel_152327_comb;
  wire [15:0] p1_sel_152328_comb;
  wire [15:0] p1_sel_152329_comb;
  wire [15:0] p1_sel_152330_comb;
  wire [15:0] p1_sel_152331_comb;
  wire [15:0] p1_sel_152332_comb;
  wire [15:0] p1_sel_152333_comb;
  wire [15:0] p1_sel_152334_comb;
  wire [15:0] p1_sel_152335_comb;
  wire [15:0] p1_sel_152336_comb;
  wire [15:0] p1_sel_152337_comb;
  wire [15:0] p1_sel_152338_comb;
  wire [15:0] p1_sel_152339_comb;
  wire [15:0] p1_sel_152340_comb;
  wire [15:0] p1_sel_152341_comb;
  wire [15:0] p1_sel_152342_comb;
  wire [15:0] p1_sel_152343_comb;
  wire [15:0] p1_sel_152344_comb;
  wire [15:0] p1_sel_152345_comb;
  wire [15:0] p1_sel_152346_comb;
  wire [15:0] p1_sel_152347_comb;
  wire [15:0] p1_sel_152348_comb;
  wire [15:0] p1_sel_152349_comb;
  wire [15:0] p1_sel_152350_comb;
  wire [15:0] p1_sel_152351_comb;
  wire [15:0] p1_sel_152352_comb;
  wire [15:0] p1_sel_152353_comb;
  wire [15:0] p1_sel_152354_comb;
  wire [15:0] p1_sel_152355_comb;
  wire [15:0] p1_sel_152356_comb;
  wire [15:0] p1_sel_152357_comb;
  wire [15:0] p1_sel_152358_comb;
  wire [15:0] p1_sel_152359_comb;
  wire [15:0] p1_sel_152360_comb;
  wire [15:0] p1_sel_152361_comb;
  wire [15:0] p1_sel_152362_comb;
  wire [15:0] p1_sel_152363_comb;
  wire [15:0] p1_sel_152364_comb;
  wire [15:0] p1_sel_152365_comb;
  wire [15:0] p1_sel_152366_comb;
  wire [15:0] p1_sel_152367_comb;
  wire [15:0] p1_sel_152368_comb;
  wire [15:0] p1_sel_152369_comb;
  wire [15:0] p1_sel_152370_comb;
  wire [15:0] p1_sel_152371_comb;
  wire [15:0] p1_sel_152372_comb;
  wire [15:0] p1_sel_152373_comb;
  wire [15:0] p1_sel_152374_comb;
  wire [15:0] p1_sel_152375_comb;
  wire [15:0] p1_sel_152376_comb;
  wire [15:0] p1_sel_152377_comb;
  wire [15:0] p1_sel_152378_comb;
  wire [15:0] p1_sel_152379_comb;
  wire [15:0] p1_sel_152380_comb;
  wire [15:0] p1_sel_152381_comb;
  wire [15:0] p1_sel_152382_comb;
  wire [15:0] p1_sel_152383_comb;
  wire [15:0] p1_sel_152384_comb;
  wire [15:0] p1_sel_152385_comb;
  wire [15:0] p1_sel_152386_comb;
  wire [15:0] p1_sel_152387_comb;
  wire [15:0] p1_sel_152388_comb;
  wire [15:0] p1_sel_152389_comb;
  wire [15:0] p1_sel_152390_comb;
  wire [15:0] p1_sel_152391_comb;
  wire [15:0] p1_sel_152392_comb;
  wire [15:0] p1_sel_152393_comb;
  wire [15:0] p1_sel_152394_comb;
  wire [15:0] p1_sel_152395_comb;
  wire [15:0] p1_sel_152396_comb;
  wire [15:0] p1_sel_152397_comb;
  wire [15:0] p1_sel_152398_comb;
  wire [15:0] p1_sel_152399_comb;
  wire [15:0] p1_sel_152400_comb;
  wire [15:0] p1_sel_152401_comb;
  wire [15:0] p1_sel_152402_comb;
  wire [15:0] p1_sel_152403_comb;
  wire [15:0] p1_sel_152404_comb;
  wire [15:0] p1_sel_152405_comb;
  wire [15:0] p1_sel_152406_comb;
  wire [15:0] p1_sel_152407_comb;
  wire [15:0] p1_sel_152408_comb;
  wire [15:0] p1_sel_152409_comb;
  wire [15:0] p1_sel_152410_comb;
  wire [31:0] p1_sum__520_comb;
  wire [31:0] p1_sum__521_comb;
  wire [31:0] p1_sum__522_comb;
  wire [31:0] p1_sum__523_comb;
  wire [31:0] p1_sum__464_comb;
  wire [31:0] p1_sum__465_comb;
  wire [31:0] p1_sum__466_comb;
  wire [31:0] p1_sum__467_comb;
  wire [31:0] p1_sum__408_comb;
  wire [31:0] p1_sum__409_comb;
  wire [31:0] p1_sum__410_comb;
  wire [31:0] p1_sum__411_comb;
  wire [31:0] p1_sum__352_comb;
  wire [31:0] p1_sum__353_comb;
  wire [31:0] p1_sum__354_comb;
  wire [31:0] p1_sum__355_comb;
  wire [31:0] p1_sum__296_comb;
  wire [31:0] p1_sum__297_comb;
  wire [31:0] p1_sum__298_comb;
  wire [31:0] p1_sum__299_comb;
  wire [31:0] p1_sum__240_comb;
  wire [31:0] p1_sum__241_comb;
  wire [31:0] p1_sum__242_comb;
  wire [31:0] p1_sum__243_comb;
  wire [31:0] p1_sum__184_comb;
  wire [31:0] p1_sum__185_comb;
  wire [31:0] p1_sum__186_comb;
  wire [31:0] p1_sum__187_comb;
  wire [31:0] p1_sum__128_comb;
  wire [31:0] p1_sum__129_comb;
  wire [31:0] p1_sum__130_comb;
  wire [31:0] p1_sum__131_comb;
  wire [31:0] p1_sum__524_comb;
  wire [31:0] p1_sum__525_comb;
  wire [31:0] p1_sum__468_comb;
  wire [31:0] p1_sum__469_comb;
  wire [31:0] p1_sum__412_comb;
  wire [31:0] p1_sum__413_comb;
  wire [31:0] p1_sum__356_comb;
  wire [31:0] p1_sum__357_comb;
  wire [31:0] p1_sum__300_comb;
  wire [31:0] p1_sum__301_comb;
  wire [31:0] p1_sum__244_comb;
  wire [31:0] p1_sum__245_comb;
  wire [31:0] p1_sum__188_comb;
  wire [31:0] p1_sum__189_comb;
  wire [31:0] p1_sum__132_comb;
  wire [31:0] p1_sum__133_comb;
  wire [16:0] p1_add_152907_comb;
  wire [16:0] p1_add_152908_comb;
  wire [16:0] p1_add_152909_comb;
  wire [16:0] p1_add_152910_comb;
  wire [16:0] p1_add_152911_comb;
  wire [16:0] p1_add_152912_comb;
  wire [16:0] p1_add_152913_comb;
  wire [16:0] p1_add_152914_comb;
  wire [16:0] p1_add_152915_comb;
  wire [16:0] p1_add_152916_comb;
  wire [16:0] p1_add_152917_comb;
  wire [16:0] p1_add_152918_comb;
  wire [16:0] p1_add_152919_comb;
  wire [16:0] p1_add_152920_comb;
  wire [16:0] p1_add_152921_comb;
  wire [16:0] p1_add_152922_comb;
  wire [16:0] p1_add_152923_comb;
  wire [16:0] p1_add_152924_comb;
  wire [16:0] p1_add_152925_comb;
  wire [16:0] p1_add_152926_comb;
  wire [16:0] p1_add_152927_comb;
  wire [16:0] p1_add_152928_comb;
  wire [16:0] p1_add_152929_comb;
  wire [16:0] p1_add_152930_comb;
  wire [16:0] p1_add_152931_comb;
  wire [16:0] p1_add_152932_comb;
  wire [16:0] p1_add_152933_comb;
  wire [16:0] p1_add_152934_comb;
  wire [16:0] p1_add_152935_comb;
  wire [16:0] p1_add_152936_comb;
  wire [16:0] p1_add_152937_comb;
  wire [16:0] p1_add_152938_comb;
  wire [16:0] p1_add_152939_comb;
  wire [16:0] p1_add_152940_comb;
  wire [16:0] p1_add_152941_comb;
  wire [16:0] p1_add_152942_comb;
  wire [16:0] p1_add_152943_comb;
  wire [16:0] p1_add_152944_comb;
  wire [16:0] p1_add_152945_comb;
  wire [16:0] p1_add_152946_comb;
  wire [16:0] p1_add_152947_comb;
  wire [16:0] p1_add_152948_comb;
  wire [16:0] p1_add_152949_comb;
  wire [16:0] p1_add_152950_comb;
  wire [16:0] p1_add_152951_comb;
  wire [16:0] p1_add_152952_comb;
  wire [16:0] p1_add_152953_comb;
  wire [16:0] p1_add_152954_comb;
  wire [16:0] p1_add_152955_comb;
  wire [16:0] p1_add_152956_comb;
  wire [16:0] p1_add_152957_comb;
  wire [16:0] p1_add_152958_comb;
  wire [16:0] p1_add_152959_comb;
  wire [16:0] p1_add_152960_comb;
  wire [16:0] p1_add_152961_comb;
  wire [16:0] p1_add_152962_comb;
  wire [16:0] p1_add_152963_comb;
  wire [16:0] p1_add_152964_comb;
  wire [16:0] p1_add_152965_comb;
  wire [16:0] p1_add_152966_comb;
  wire [16:0] p1_add_152967_comb;
  wire [16:0] p1_add_152968_comb;
  wire [16:0] p1_add_152969_comb;
  wire [16:0] p1_add_152970_comb;
  wire [16:0] p1_add_152971_comb;
  wire [16:0] p1_add_152972_comb;
  wire [16:0] p1_add_152973_comb;
  wire [16:0] p1_add_152974_comb;
  wire [16:0] p1_add_152975_comb;
  wire [16:0] p1_add_152976_comb;
  wire [16:0] p1_add_152977_comb;
  wire [16:0] p1_add_152978_comb;
  wire [16:0] p1_add_152979_comb;
  wire [16:0] p1_add_152980_comb;
  wire [16:0] p1_add_152981_comb;
  wire [16:0] p1_add_152982_comb;
  wire [16:0] p1_add_152983_comb;
  wire [16:0] p1_add_152984_comb;
  wire [16:0] p1_add_152985_comb;
  wire [16:0] p1_add_152986_comb;
  wire [16:0] p1_add_152987_comb;
  wire [16:0] p1_add_152988_comb;
  wire [16:0] p1_add_152989_comb;
  wire [16:0] p1_add_152990_comb;
  wire [16:0] p1_add_152991_comb;
  wire [16:0] p1_add_152992_comb;
  wire [16:0] p1_add_152993_comb;
  wire [16:0] p1_add_152994_comb;
  wire [16:0] p1_add_152995_comb;
  wire [16:0] p1_add_152996_comb;
  wire [16:0] p1_add_152997_comb;
  wire [16:0] p1_add_152998_comb;
  wire [16:0] p1_add_152999_comb;
  wire [16:0] p1_add_153000_comb;
  wire [16:0] p1_add_153001_comb;
  wire [16:0] p1_add_153002_comb;
  wire [16:0] p1_add_153003_comb;
  wire [16:0] p1_add_153004_comb;
  wire [16:0] p1_add_153005_comb;
  wire [16:0] p1_add_153006_comb;
  wire [16:0] p1_add_153007_comb;
  wire [16:0] p1_add_153008_comb;
  wire [16:0] p1_add_153009_comb;
  wire [16:0] p1_add_153010_comb;
  wire [16:0] p1_add_153011_comb;
  wire [16:0] p1_add_153012_comb;
  wire [16:0] p1_add_153013_comb;
  wire [16:0] p1_add_153014_comb;
  wire [16:0] p1_add_153015_comb;
  wire [16:0] p1_add_153016_comb;
  wire [16:0] p1_add_153017_comb;
  wire [16:0] p1_add_153018_comb;
  wire [16:0] p1_add_153019_comb;
  wire [16:0] p1_add_153020_comb;
  wire [16:0] p1_add_153021_comb;
  wire [16:0] p1_add_153022_comb;
  wire [16:0] p1_add_153023_comb;
  wire [16:0] p1_add_153024_comb;
  wire [16:0] p1_add_153025_comb;
  wire [16:0] p1_add_153026_comb;
  wire [16:0] p1_add_153027_comb;
  wire [16:0] p1_add_153028_comb;
  wire [16:0] p1_add_153029_comb;
  wire [16:0] p1_add_153030_comb;
  wire [16:0] p1_add_153031_comb;
  wire [16:0] p1_add_153032_comb;
  wire [16:0] p1_add_153033_comb;
  wire [16:0] p1_add_153034_comb;
  wire [16:0] p1_add_153035_comb;
  wire [16:0] p1_add_153036_comb;
  wire [16:0] p1_add_153037_comb;
  wire [16:0] p1_add_153038_comb;
  wire [16:0] p1_add_153039_comb;
  wire [16:0] p1_add_153040_comb;
  wire [16:0] p1_add_153041_comb;
  wire [16:0] p1_add_153042_comb;
  wire [16:0] p1_add_153043_comb;
  wire [16:0] p1_add_153044_comb;
  wire [16:0] p1_add_153045_comb;
  wire [16:0] p1_add_153046_comb;
  wire [16:0] p1_add_153047_comb;
  wire [16:0] p1_add_153048_comb;
  wire [16:0] p1_add_153049_comb;
  wire [16:0] p1_add_153050_comb;
  wire [16:0] p1_add_153051_comb;
  wire [16:0] p1_add_153052_comb;
  wire [16:0] p1_add_153053_comb;
  wire [16:0] p1_add_153054_comb;
  wire [16:0] p1_add_153055_comb;
  wire [16:0] p1_add_153056_comb;
  wire [16:0] p1_add_153057_comb;
  wire [16:0] p1_add_153058_comb;
  wire [16:0] p1_add_153059_comb;
  wire [16:0] p1_add_153060_comb;
  wire [16:0] p1_add_153061_comb;
  wire [16:0] p1_add_153062_comb;
  wire [16:0] p1_add_153063_comb;
  wire [16:0] p1_add_153064_comb;
  wire [16:0] p1_add_153065_comb;
  wire [16:0] p1_add_153066_comb;
  wire [16:0] p1_add_153067_comb;
  wire [16:0] p1_add_153068_comb;
  wire [16:0] p1_add_153069_comb;
  wire [16:0] p1_add_153070_comb;
  wire [16:0] p1_add_153071_comb;
  wire [16:0] p1_add_153072_comb;
  wire [16:0] p1_add_153073_comb;
  wire [16:0] p1_add_153074_comb;
  wire [16:0] p1_add_153075_comb;
  wire [16:0] p1_add_153076_comb;
  wire [16:0] p1_add_153077_comb;
  wire [16:0] p1_add_153078_comb;
  wire [16:0] p1_add_153079_comb;
  wire [16:0] p1_add_153080_comb;
  wire [16:0] p1_add_153081_comb;
  wire [16:0] p1_add_153082_comb;
  wire [16:0] p1_add_153083_comb;
  wire [16:0] p1_add_153084_comb;
  wire [16:0] p1_add_153085_comb;
  wire [16:0] p1_add_153086_comb;
  wire [16:0] p1_add_153087_comb;
  wire [16:0] p1_add_153088_comb;
  wire [16:0] p1_add_153089_comb;
  wire [16:0] p1_add_153090_comb;
  wire [16:0] p1_add_153091_comb;
  wire [16:0] p1_add_153092_comb;
  wire [16:0] p1_add_153093_comb;
  wire [16:0] p1_add_153094_comb;
  wire [16:0] p1_add_153095_comb;
  wire [16:0] p1_add_153096_comb;
  wire [16:0] p1_add_153097_comb;
  wire [16:0] p1_add_153098_comb;
  wire [16:0] p1_add_153099_comb;
  wire [16:0] p1_add_153100_comb;
  wire [16:0] p1_add_153101_comb;
  wire [16:0] p1_add_153102_comb;
  wire [16:0] p1_add_153103_comb;
  wire [16:0] p1_add_153104_comb;
  wire [16:0] p1_add_153105_comb;
  wire [16:0] p1_add_153106_comb;
  wire [16:0] p1_add_153107_comb;
  wire [16:0] p1_add_153108_comb;
  wire [16:0] p1_add_153109_comb;
  wire [16:0] p1_add_153110_comb;
  wire [16:0] p1_add_153111_comb;
  wire [16:0] p1_add_153112_comb;
  wire [16:0] p1_add_153113_comb;
  wire [16:0] p1_add_153114_comb;
  wire [16:0] p1_add_153115_comb;
  wire [16:0] p1_add_153116_comb;
  wire [16:0] p1_add_153117_comb;
  wire [16:0] p1_add_153118_comb;
  wire [16:0] p1_add_153119_comb;
  wire [16:0] p1_add_153120_comb;
  wire [16:0] p1_add_153121_comb;
  wire [16:0] p1_add_153122_comb;
  wire [16:0] p1_add_153123_comb;
  wire [16:0] p1_add_153124_comb;
  wire [16:0] p1_add_153125_comb;
  wire [16:0] p1_add_153126_comb;
  wire [16:0] p1_add_153127_comb;
  wire [16:0] p1_add_153128_comb;
  wire [16:0] p1_add_153129_comb;
  wire [16:0] p1_add_153130_comb;
  wire [31:0] p1_sum__526_comb;
  wire [31:0] p1_sum__470_comb;
  wire [31:0] p1_sum__414_comb;
  wire [31:0] p1_sum__358_comb;
  wire [31:0] p1_sum__302_comb;
  wire [31:0] p1_sum__246_comb;
  wire [31:0] p1_sum__190_comb;
  wire [31:0] p1_sum__134_comb;
  wire [24:0] p1_sum__1580_comb;
  wire [24:0] p1_sum__1581_comb;
  wire [24:0] p1_sum__1582_comb;
  wire [24:0] p1_sum__1583_comb;
  wire [24:0] p1_sum__1552_comb;
  wire [24:0] p1_sum__1553_comb;
  wire [24:0] p1_sum__1554_comb;
  wire [24:0] p1_sum__1555_comb;
  wire [24:0] p1_sum__1524_comb;
  wire [24:0] p1_sum__1525_comb;
  wire [24:0] p1_sum__1526_comb;
  wire [24:0] p1_sum__1527_comb;
  wire [24:0] p1_sum__1496_comb;
  wire [24:0] p1_sum__1497_comb;
  wire [24:0] p1_sum__1498_comb;
  wire [24:0] p1_sum__1499_comb;
  wire [24:0] p1_sum__1468_comb;
  wire [24:0] p1_sum__1469_comb;
  wire [24:0] p1_sum__1470_comb;
  wire [24:0] p1_sum__1471_comb;
  wire [24:0] p1_sum__1440_comb;
  wire [24:0] p1_sum__1441_comb;
  wire [24:0] p1_sum__1442_comb;
  wire [24:0] p1_sum__1443_comb;
  wire [24:0] p1_sum__1412_comb;
  wire [24:0] p1_sum__1413_comb;
  wire [24:0] p1_sum__1414_comb;
  wire [24:0] p1_sum__1415_comb;
  wire [24:0] p1_sum__1384_comb;
  wire [24:0] p1_sum__1385_comb;
  wire [24:0] p1_sum__1386_comb;
  wire [24:0] p1_sum__1387_comb;
  wire [24:0] p1_sum__1576_comb;
  wire [24:0] p1_sum__1577_comb;
  wire [24:0] p1_sum__1578_comb;
  wire [24:0] p1_sum__1579_comb;
  wire [24:0] p1_sum__1548_comb;
  wire [24:0] p1_sum__1549_comb;
  wire [24:0] p1_sum__1550_comb;
  wire [24:0] p1_sum__1551_comb;
  wire [24:0] p1_sum__1520_comb;
  wire [24:0] p1_sum__1521_comb;
  wire [24:0] p1_sum__1522_comb;
  wire [24:0] p1_sum__1523_comb;
  wire [24:0] p1_sum__1492_comb;
  wire [24:0] p1_sum__1493_comb;
  wire [24:0] p1_sum__1494_comb;
  wire [24:0] p1_sum__1495_comb;
  wire [24:0] p1_sum__1464_comb;
  wire [24:0] p1_sum__1465_comb;
  wire [24:0] p1_sum__1466_comb;
  wire [24:0] p1_sum__1467_comb;
  wire [24:0] p1_sum__1436_comb;
  wire [24:0] p1_sum__1437_comb;
  wire [24:0] p1_sum__1438_comb;
  wire [24:0] p1_sum__1439_comb;
  wire [24:0] p1_sum__1408_comb;
  wire [24:0] p1_sum__1409_comb;
  wire [24:0] p1_sum__1410_comb;
  wire [24:0] p1_sum__1411_comb;
  wire [24:0] p1_sum__1380_comb;
  wire [24:0] p1_sum__1381_comb;
  wire [24:0] p1_sum__1382_comb;
  wire [24:0] p1_sum__1383_comb;
  wire [24:0] p1_sum__1572_comb;
  wire [24:0] p1_sum__1573_comb;
  wire [24:0] p1_sum__1574_comb;
  wire [24:0] p1_sum__1575_comb;
  wire [24:0] p1_sum__1544_comb;
  wire [24:0] p1_sum__1545_comb;
  wire [24:0] p1_sum__1546_comb;
  wire [24:0] p1_sum__1547_comb;
  wire [24:0] p1_sum__1516_comb;
  wire [24:0] p1_sum__1517_comb;
  wire [24:0] p1_sum__1518_comb;
  wire [24:0] p1_sum__1519_comb;
  wire [24:0] p1_sum__1488_comb;
  wire [24:0] p1_sum__1489_comb;
  wire [24:0] p1_sum__1490_comb;
  wire [24:0] p1_sum__1491_comb;
  wire [24:0] p1_sum__1460_comb;
  wire [24:0] p1_sum__1461_comb;
  wire [24:0] p1_sum__1462_comb;
  wire [24:0] p1_sum__1463_comb;
  wire [24:0] p1_sum__1432_comb;
  wire [24:0] p1_sum__1433_comb;
  wire [24:0] p1_sum__1434_comb;
  wire [24:0] p1_sum__1435_comb;
  wire [24:0] p1_sum__1404_comb;
  wire [24:0] p1_sum__1405_comb;
  wire [24:0] p1_sum__1406_comb;
  wire [24:0] p1_sum__1407_comb;
  wire [24:0] p1_sum__1376_comb;
  wire [24:0] p1_sum__1377_comb;
  wire [24:0] p1_sum__1378_comb;
  wire [24:0] p1_sum__1379_comb;
  wire [24:0] p1_sum__1568_comb;
  wire [24:0] p1_sum__1569_comb;
  wire [24:0] p1_sum__1570_comb;
  wire [24:0] p1_sum__1571_comb;
  wire [24:0] p1_sum__1540_comb;
  wire [24:0] p1_sum__1541_comb;
  wire [24:0] p1_sum__1542_comb;
  wire [24:0] p1_sum__1543_comb;
  wire [24:0] p1_sum__1512_comb;
  wire [24:0] p1_sum__1513_comb;
  wire [24:0] p1_sum__1514_comb;
  wire [24:0] p1_sum__1515_comb;
  wire [24:0] p1_sum__1484_comb;
  wire [24:0] p1_sum__1485_comb;
  wire [24:0] p1_sum__1486_comb;
  wire [24:0] p1_sum__1487_comb;
  wire [24:0] p1_sum__1456_comb;
  wire [24:0] p1_sum__1457_comb;
  wire [24:0] p1_sum__1458_comb;
  wire [24:0] p1_sum__1459_comb;
  wire [24:0] p1_sum__1428_comb;
  wire [24:0] p1_sum__1429_comb;
  wire [24:0] p1_sum__1430_comb;
  wire [24:0] p1_sum__1431_comb;
  wire [24:0] p1_sum__1400_comb;
  wire [24:0] p1_sum__1401_comb;
  wire [24:0] p1_sum__1402_comb;
  wire [24:0] p1_sum__1403_comb;
  wire [24:0] p1_sum__1372_comb;
  wire [24:0] p1_sum__1373_comb;
  wire [24:0] p1_sum__1374_comb;
  wire [24:0] p1_sum__1375_comb;
  wire [24:0] p1_sum__1564_comb;
  wire [24:0] p1_sum__1565_comb;
  wire [24:0] p1_sum__1566_comb;
  wire [24:0] p1_sum__1567_comb;
  wire [24:0] p1_sum__1536_comb;
  wire [24:0] p1_sum__1537_comb;
  wire [24:0] p1_sum__1538_comb;
  wire [24:0] p1_sum__1539_comb;
  wire [24:0] p1_sum__1508_comb;
  wire [24:0] p1_sum__1509_comb;
  wire [24:0] p1_sum__1510_comb;
  wire [24:0] p1_sum__1511_comb;
  wire [24:0] p1_sum__1480_comb;
  wire [24:0] p1_sum__1481_comb;
  wire [24:0] p1_sum__1482_comb;
  wire [24:0] p1_sum__1483_comb;
  wire [24:0] p1_sum__1452_comb;
  wire [24:0] p1_sum__1453_comb;
  wire [24:0] p1_sum__1454_comb;
  wire [24:0] p1_sum__1455_comb;
  wire [24:0] p1_sum__1424_comb;
  wire [24:0] p1_sum__1425_comb;
  wire [24:0] p1_sum__1426_comb;
  wire [24:0] p1_sum__1427_comb;
  wire [24:0] p1_sum__1396_comb;
  wire [24:0] p1_sum__1397_comb;
  wire [24:0] p1_sum__1398_comb;
  wire [24:0] p1_sum__1399_comb;
  wire [24:0] p1_sum__1368_comb;
  wire [24:0] p1_sum__1369_comb;
  wire [24:0] p1_sum__1370_comb;
  wire [24:0] p1_sum__1371_comb;
  wire [24:0] p1_sum__1560_comb;
  wire [24:0] p1_sum__1561_comb;
  wire [24:0] p1_sum__1562_comb;
  wire [24:0] p1_sum__1563_comb;
  wire [24:0] p1_sum__1532_comb;
  wire [24:0] p1_sum__1533_comb;
  wire [24:0] p1_sum__1534_comb;
  wire [24:0] p1_sum__1535_comb;
  wire [24:0] p1_sum__1504_comb;
  wire [24:0] p1_sum__1505_comb;
  wire [24:0] p1_sum__1506_comb;
  wire [24:0] p1_sum__1507_comb;
  wire [24:0] p1_sum__1476_comb;
  wire [24:0] p1_sum__1477_comb;
  wire [24:0] p1_sum__1478_comb;
  wire [24:0] p1_sum__1479_comb;
  wire [24:0] p1_sum__1448_comb;
  wire [24:0] p1_sum__1449_comb;
  wire [24:0] p1_sum__1450_comb;
  wire [24:0] p1_sum__1451_comb;
  wire [24:0] p1_sum__1420_comb;
  wire [24:0] p1_sum__1421_comb;
  wire [24:0] p1_sum__1422_comb;
  wire [24:0] p1_sum__1423_comb;
  wire [24:0] p1_sum__1392_comb;
  wire [24:0] p1_sum__1393_comb;
  wire [24:0] p1_sum__1394_comb;
  wire [24:0] p1_sum__1395_comb;
  wire [24:0] p1_sum__1364_comb;
  wire [24:0] p1_sum__1365_comb;
  wire [24:0] p1_sum__1366_comb;
  wire [24:0] p1_sum__1367_comb;
  wire [24:0] p1_sum__1556_comb;
  wire [24:0] p1_sum__1557_comb;
  wire [24:0] p1_sum__1558_comb;
  wire [24:0] p1_sum__1559_comb;
  wire [24:0] p1_sum__1528_comb;
  wire [24:0] p1_sum__1529_comb;
  wire [24:0] p1_sum__1530_comb;
  wire [24:0] p1_sum__1531_comb;
  wire [24:0] p1_sum__1500_comb;
  wire [24:0] p1_sum__1501_comb;
  wire [24:0] p1_sum__1502_comb;
  wire [24:0] p1_sum__1503_comb;
  wire [24:0] p1_sum__1472_comb;
  wire [24:0] p1_sum__1473_comb;
  wire [24:0] p1_sum__1474_comb;
  wire [24:0] p1_sum__1475_comb;
  wire [24:0] p1_sum__1444_comb;
  wire [24:0] p1_sum__1445_comb;
  wire [24:0] p1_sum__1446_comb;
  wire [24:0] p1_sum__1447_comb;
  wire [24:0] p1_sum__1416_comb;
  wire [24:0] p1_sum__1417_comb;
  wire [24:0] p1_sum__1418_comb;
  wire [24:0] p1_sum__1419_comb;
  wire [24:0] p1_sum__1388_comb;
  wire [24:0] p1_sum__1389_comb;
  wire [24:0] p1_sum__1390_comb;
  wire [24:0] p1_sum__1391_comb;
  wire [24:0] p1_sum__1360_comb;
  wire [24:0] p1_sum__1361_comb;
  wire [24:0] p1_sum__1362_comb;
  wire [24:0] p1_sum__1363_comb;
  wire [31:0] p1_umul_153371_comb;
  wire [31:0] p1_umul_153372_comb;
  wire [31:0] p1_umul_153373_comb;
  wire [31:0] p1_umul_153374_comb;
  wire [31:0] p1_umul_153375_comb;
  wire [31:0] p1_umul_153376_comb;
  wire [31:0] p1_umul_153377_comb;
  wire [31:0] p1_umul_153378_comb;
  wire [24:0] p1_sum__1246_comb;
  wire [24:0] p1_sum__1247_comb;
  wire [24:0] p1_sum__1232_comb;
  wire [24:0] p1_sum__1233_comb;
  wire [24:0] p1_sum__1218_comb;
  wire [24:0] p1_sum__1219_comb;
  wire [24:0] p1_sum__1204_comb;
  wire [24:0] p1_sum__1205_comb;
  wire [24:0] p1_sum__1190_comb;
  wire [24:0] p1_sum__1191_comb;
  wire [24:0] p1_sum__1176_comb;
  wire [24:0] p1_sum__1177_comb;
  wire [24:0] p1_sum__1162_comb;
  wire [24:0] p1_sum__1163_comb;
  wire [24:0] p1_sum__1148_comb;
  wire [24:0] p1_sum__1149_comb;
  wire [24:0] p1_sum__1244_comb;
  wire [24:0] p1_sum__1245_comb;
  wire [24:0] p1_sum__1230_comb;
  wire [24:0] p1_sum__1231_comb;
  wire [24:0] p1_sum__1216_comb;
  wire [24:0] p1_sum__1217_comb;
  wire [24:0] p1_sum__1202_comb;
  wire [24:0] p1_sum__1203_comb;
  wire [24:0] p1_sum__1188_comb;
  wire [24:0] p1_sum__1189_comb;
  wire [24:0] p1_sum__1174_comb;
  wire [24:0] p1_sum__1175_comb;
  wire [24:0] p1_sum__1160_comb;
  wire [24:0] p1_sum__1161_comb;
  wire [24:0] p1_sum__1146_comb;
  wire [24:0] p1_sum__1147_comb;
  wire [24:0] p1_sum__1242_comb;
  wire [24:0] p1_sum__1243_comb;
  wire [24:0] p1_sum__1228_comb;
  wire [24:0] p1_sum__1229_comb;
  wire [24:0] p1_sum__1214_comb;
  wire [24:0] p1_sum__1215_comb;
  wire [24:0] p1_sum__1200_comb;
  wire [24:0] p1_sum__1201_comb;
  wire [24:0] p1_sum__1186_comb;
  wire [24:0] p1_sum__1187_comb;
  wire [24:0] p1_sum__1172_comb;
  wire [24:0] p1_sum__1173_comb;
  wire [24:0] p1_sum__1158_comb;
  wire [24:0] p1_sum__1159_comb;
  wire [24:0] p1_sum__1144_comb;
  wire [24:0] p1_sum__1145_comb;
  wire [24:0] p1_sum__1240_comb;
  wire [24:0] p1_sum__1241_comb;
  wire [24:0] p1_sum__1226_comb;
  wire [24:0] p1_sum__1227_comb;
  wire [24:0] p1_sum__1212_comb;
  wire [24:0] p1_sum__1213_comb;
  wire [24:0] p1_sum__1198_comb;
  wire [24:0] p1_sum__1199_comb;
  wire [24:0] p1_sum__1184_comb;
  wire [24:0] p1_sum__1185_comb;
  wire [24:0] p1_sum__1170_comb;
  wire [24:0] p1_sum__1171_comb;
  wire [24:0] p1_sum__1156_comb;
  wire [24:0] p1_sum__1157_comb;
  wire [24:0] p1_sum__1142_comb;
  wire [24:0] p1_sum__1143_comb;
  wire [24:0] p1_sum__1238_comb;
  wire [24:0] p1_sum__1239_comb;
  wire [24:0] p1_sum__1224_comb;
  wire [24:0] p1_sum__1225_comb;
  wire [24:0] p1_sum__1210_comb;
  wire [24:0] p1_sum__1211_comb;
  wire [24:0] p1_sum__1196_comb;
  wire [24:0] p1_sum__1197_comb;
  wire [24:0] p1_sum__1182_comb;
  wire [24:0] p1_sum__1183_comb;
  wire [24:0] p1_sum__1168_comb;
  wire [24:0] p1_sum__1169_comb;
  wire [24:0] p1_sum__1154_comb;
  wire [24:0] p1_sum__1155_comb;
  wire [24:0] p1_sum__1140_comb;
  wire [24:0] p1_sum__1141_comb;
  wire [24:0] p1_sum__1236_comb;
  wire [24:0] p1_sum__1237_comb;
  wire [24:0] p1_sum__1222_comb;
  wire [24:0] p1_sum__1223_comb;
  wire [24:0] p1_sum__1208_comb;
  wire [24:0] p1_sum__1209_comb;
  wire [24:0] p1_sum__1194_comb;
  wire [24:0] p1_sum__1195_comb;
  wire [24:0] p1_sum__1180_comb;
  wire [24:0] p1_sum__1181_comb;
  wire [24:0] p1_sum__1166_comb;
  wire [24:0] p1_sum__1167_comb;
  wire [24:0] p1_sum__1152_comb;
  wire [24:0] p1_sum__1153_comb;
  wire [24:0] p1_sum__1138_comb;
  wire [24:0] p1_sum__1139_comb;
  wire [24:0] p1_sum__1234_comb;
  wire [24:0] p1_sum__1235_comb;
  wire [24:0] p1_sum__1220_comb;
  wire [24:0] p1_sum__1221_comb;
  wire [24:0] p1_sum__1206_comb;
  wire [24:0] p1_sum__1207_comb;
  wire [24:0] p1_sum__1192_comb;
  wire [24:0] p1_sum__1193_comb;
  wire [24:0] p1_sum__1178_comb;
  wire [24:0] p1_sum__1179_comb;
  wire [24:0] p1_sum__1164_comb;
  wire [24:0] p1_sum__1165_comb;
  wire [24:0] p1_sum__1150_comb;
  wire [24:0] p1_sum__1151_comb;
  wire [24:0] p1_sum__1136_comb;
  wire [24:0] p1_sum__1137_comb;
  wire [24:0] p1_sum__1079_comb;
  wire [24:0] p1_sum__1072_comb;
  wire [24:0] p1_sum__1065_comb;
  wire [24:0] p1_sum__1058_comb;
  wire [24:0] p1_sum__1051_comb;
  wire [24:0] p1_sum__1044_comb;
  wire [24:0] p1_sum__1037_comb;
  wire [24:0] p1_sum__1030_comb;
  wire [24:0] p1_sum__1078_comb;
  wire [24:0] p1_sum__1071_comb;
  wire [24:0] p1_sum__1064_comb;
  wire [24:0] p1_sum__1057_comb;
  wire [24:0] p1_sum__1050_comb;
  wire [24:0] p1_sum__1043_comb;
  wire [24:0] p1_sum__1036_comb;
  wire [24:0] p1_sum__1029_comb;
  wire [24:0] p1_sum__1077_comb;
  wire [24:0] p1_sum__1070_comb;
  wire [24:0] p1_sum__1063_comb;
  wire [24:0] p1_sum__1056_comb;
  wire [24:0] p1_sum__1049_comb;
  wire [24:0] p1_sum__1042_comb;
  wire [24:0] p1_sum__1035_comb;
  wire [24:0] p1_sum__1028_comb;
  wire [24:0] p1_sum__1076_comb;
  wire [24:0] p1_sum__1069_comb;
  wire [24:0] p1_sum__1062_comb;
  wire [24:0] p1_sum__1055_comb;
  wire [24:0] p1_sum__1048_comb;
  wire [24:0] p1_sum__1041_comb;
  wire [24:0] p1_sum__1034_comb;
  wire [24:0] p1_sum__1027_comb;
  wire [24:0] p1_sum__1075_comb;
  wire [24:0] p1_sum__1068_comb;
  wire [24:0] p1_sum__1061_comb;
  wire [24:0] p1_sum__1054_comb;
  wire [24:0] p1_sum__1047_comb;
  wire [24:0] p1_sum__1040_comb;
  wire [24:0] p1_sum__1033_comb;
  wire [24:0] p1_sum__1026_comb;
  wire [24:0] p1_sum__1074_comb;
  wire [24:0] p1_sum__1067_comb;
  wire [24:0] p1_sum__1060_comb;
  wire [24:0] p1_sum__1053_comb;
  wire [24:0] p1_sum__1046_comb;
  wire [24:0] p1_sum__1039_comb;
  wire [24:0] p1_sum__1032_comb;
  wire [24:0] p1_sum__1025_comb;
  wire [24:0] p1_sum__1073_comb;
  wire [24:0] p1_sum__1066_comb;
  wire [24:0] p1_sum__1059_comb;
  wire [24:0] p1_sum__1052_comb;
  wire [24:0] p1_sum__1045_comb;
  wire [24:0] p1_sum__1038_comb;
  wire [24:0] p1_sum__1031_comb;
  wire [24:0] p1_sum__1024_comb;
  wire [24:0] p1_add_153619_comb;
  wire [24:0] p1_add_153620_comb;
  wire [24:0] p1_add_153621_comb;
  wire [24:0] p1_add_153622_comb;
  wire [24:0] p1_add_153623_comb;
  wire [24:0] p1_add_153624_comb;
  wire [24:0] p1_add_153625_comb;
  wire [24:0] p1_add_153626_comb;
  wire [24:0] p1_add_153627_comb;
  wire [24:0] p1_add_153628_comb;
  wire [24:0] p1_add_153629_comb;
  wire [24:0] p1_add_153630_comb;
  wire [24:0] p1_add_153631_comb;
  wire [24:0] p1_add_153632_comb;
  wire [24:0] p1_add_153633_comb;
  wire [24:0] p1_add_153634_comb;
  wire [24:0] p1_add_153635_comb;
  wire [24:0] p1_add_153636_comb;
  wire [24:0] p1_add_153637_comb;
  wire [24:0] p1_add_153638_comb;
  wire [24:0] p1_add_153639_comb;
  wire [24:0] p1_add_153640_comb;
  wire [24:0] p1_add_153641_comb;
  wire [24:0] p1_add_153642_comb;
  wire [24:0] p1_add_153643_comb;
  wire [24:0] p1_add_153644_comb;
  wire [24:0] p1_add_153645_comb;
  wire [24:0] p1_add_153646_comb;
  wire [24:0] p1_add_153647_comb;
  wire [24:0] p1_add_153648_comb;
  wire [24:0] p1_add_153649_comb;
  wire [24:0] p1_add_153650_comb;
  wire [24:0] p1_add_153651_comb;
  wire [24:0] p1_add_153652_comb;
  wire [24:0] p1_add_153653_comb;
  wire [24:0] p1_add_153654_comb;
  wire [24:0] p1_add_153655_comb;
  wire [24:0] p1_add_153656_comb;
  wire [24:0] p1_add_153657_comb;
  wire [24:0] p1_add_153658_comb;
  wire [24:0] p1_add_153659_comb;
  wire [24:0] p1_add_153660_comb;
  wire [24:0] p1_add_153661_comb;
  wire [24:0] p1_add_153662_comb;
  wire [24:0] p1_add_153663_comb;
  wire [24:0] p1_add_153664_comb;
  wire [24:0] p1_add_153665_comb;
  wire [24:0] p1_add_153666_comb;
  wire [24:0] p1_add_153667_comb;
  wire [24:0] p1_add_153668_comb;
  wire [24:0] p1_add_153669_comb;
  wire [24:0] p1_add_153670_comb;
  wire [24:0] p1_add_153671_comb;
  wire [24:0] p1_add_153672_comb;
  wire [24:0] p1_add_153673_comb;
  wire [24:0] p1_add_153674_comb;
  wire [24:0] p1_add_153675_comb;
  wire [24:0] p1_add_153676_comb;
  wire [24:0] p1_add_153677_comb;
  wire [24:0] p1_add_153678_comb;
  wire [24:0] p1_add_153679_comb;
  wire [24:0] p1_add_153680_comb;
  wire [24:0] p1_add_153681_comb;
  wire [24:0] p1_add_153682_comb;
  wire [8:0] p1_clipped__320_comb;
  wire [8:0] p1_clipped__321_comb;
  wire [8:0] p1_clipped__322_comb;
  wire [8:0] p1_clipped__323_comb;
  wire [8:0] p1_clipped__324_comb;
  wire [8:0] p1_clipped__325_comb;
  wire [8:0] p1_clipped__326_comb;
  wire [8:0] p1_clipped__327_comb;
  wire [8:0] p1_clipped__328_comb;
  wire [8:0] p1_clipped__329_comb;
  wire [8:0] p1_clipped__330_comb;
  wire [8:0] p1_clipped__331_comb;
  wire [8:0] p1_clipped__332_comb;
  wire [8:0] p1_clipped__333_comb;
  wire [8:0] p1_clipped__334_comb;
  wire [8:0] p1_clipped__335_comb;
  wire [8:0] p1_clipped__336_comb;
  wire [8:0] p1_clipped__337_comb;
  wire [8:0] p1_clipped__338_comb;
  wire [8:0] p1_clipped__339_comb;
  wire [8:0] p1_clipped__340_comb;
  wire [8:0] p1_clipped__341_comb;
  wire [8:0] p1_clipped__342_comb;
  wire [8:0] p1_clipped__343_comb;
  wire [8:0] p1_clipped__344_comb;
  wire [8:0] p1_clipped__345_comb;
  wire [8:0] p1_clipped__346_comb;
  wire [8:0] p1_clipped__347_comb;
  wire [8:0] p1_clipped__348_comb;
  wire [8:0] p1_clipped__349_comb;
  wire [8:0] p1_clipped__350_comb;
  wire [8:0] p1_clipped__351_comb;
  wire [8:0] p1_clipped__352_comb;
  wire [8:0] p1_clipped__353_comb;
  wire [8:0] p1_clipped__354_comb;
  wire [8:0] p1_clipped__355_comb;
  wire [8:0] p1_clipped__356_comb;
  wire [8:0] p1_clipped__357_comb;
  wire [8:0] p1_clipped__358_comb;
  wire [8:0] p1_clipped__359_comb;
  wire [8:0] p1_clipped__360_comb;
  wire [8:0] p1_clipped__361_comb;
  wire [8:0] p1_clipped__362_comb;
  wire [8:0] p1_clipped__363_comb;
  wire [8:0] p1_clipped__364_comb;
  wire [8:0] p1_clipped__365_comb;
  wire [8:0] p1_clipped__366_comb;
  wire [8:0] p1_clipped__367_comb;
  wire [8:0] p1_clipped__368_comb;
  wire [8:0] p1_clipped__369_comb;
  wire [8:0] p1_clipped__370_comb;
  wire [8:0] p1_clipped__371_comb;
  wire [8:0] p1_clipped__372_comb;
  wire [8:0] p1_clipped__373_comb;
  wire [8:0] p1_clipped__374_comb;
  wire [8:0] p1_clipped__375_comb;
  wire [8:0] p1_clipped__376_comb;
  wire [8:0] p1_clipped__377_comb;
  wire [8:0] p1_clipped__378_comb;
  wire [8:0] p1_clipped__379_comb;
  wire [8:0] p1_clipped__380_comb;
  wire [8:0] p1_clipped__381_comb;
  wire [8:0] p1_clipped__382_comb;
  wire [8:0] p1_clipped__383_comb;
  wire [9:0] p1_add_154451_comb;
  wire [9:0] p1_add_154452_comb;
  wire [9:0] p1_add_154453_comb;
  wire [9:0] p1_add_154454_comb;
  wire [9:0] p1_add_154455_comb;
  wire [9:0] p1_add_154456_comb;
  wire [9:0] p1_add_154457_comb;
  wire [9:0] p1_add_154458_comb;
  wire [9:0] p1_add_154459_comb;
  wire [9:0] p1_add_154460_comb;
  wire [9:0] p1_add_154461_comb;
  wire [9:0] p1_add_154462_comb;
  wire [9:0] p1_add_154463_comb;
  wire [9:0] p1_add_154464_comb;
  wire [9:0] p1_add_154465_comb;
  wire [9:0] p1_add_154466_comb;
  wire [9:0] p1_add_154467_comb;
  wire [9:0] p1_add_154468_comb;
  wire [9:0] p1_add_154469_comb;
  wire [9:0] p1_add_154470_comb;
  wire [9:0] p1_add_154471_comb;
  wire [9:0] p1_add_154472_comb;
  wire [9:0] p1_add_154473_comb;
  wire [9:0] p1_add_154474_comb;
  wire [9:0] p1_add_154475_comb;
  wire [9:0] p1_add_154476_comb;
  wire [9:0] p1_add_154477_comb;
  wire [9:0] p1_add_154478_comb;
  wire [9:0] p1_add_154479_comb;
  wire [9:0] p1_add_154480_comb;
  wire [9:0] p1_add_154481_comb;
  wire [9:0] p1_add_154482_comb;
  wire [9:0] p1_add_154483_comb;
  wire [9:0] p1_add_154484_comb;
  wire [9:0] p1_add_154485_comb;
  wire [9:0] p1_add_154486_comb;
  wire [9:0] p1_add_154487_comb;
  wire [9:0] p1_add_154488_comb;
  wire [9:0] p1_add_154489_comb;
  wire [9:0] p1_add_154490_comb;
  wire [9:0] p1_add_154491_comb;
  wire [9:0] p1_add_154492_comb;
  wire [9:0] p1_add_154493_comb;
  wire [9:0] p1_add_154494_comb;
  wire [9:0] p1_add_154495_comb;
  wire [9:0] p1_add_154496_comb;
  wire [9:0] p1_add_154497_comb;
  wire [9:0] p1_add_154498_comb;
  wire [9:0] p1_add_154499_comb;
  wire [9:0] p1_add_154500_comb;
  wire [9:0] p1_add_154501_comb;
  wire [9:0] p1_add_154502_comb;
  wire [9:0] p1_add_154503_comb;
  wire [9:0] p1_add_154504_comb;
  wire [9:0] p1_add_154505_comb;
  wire [9:0] p1_add_154506_comb;
  wire [9:0] p1_add_154507_comb;
  wire [9:0] p1_add_154508_comb;
  wire [9:0] p1_add_154509_comb;
  wire [9:0] p1_add_154510_comb;
  wire [9:0] p1_add_154511_comb;
  wire [9:0] p1_add_154512_comb;
  wire [9:0] p1_add_154513_comb;
  wire [9:0] p1_add_154514_comb;
  wire [1:0] p1_bit_slice_154515_comb;
  wire [1:0] p1_bit_slice_154516_comb;
  wire [1:0] p1_bit_slice_154517_comb;
  wire [1:0] p1_bit_slice_154518_comb;
  wire [1:0] p1_bit_slice_154519_comb;
  wire [1:0] p1_bit_slice_154520_comb;
  wire [1:0] p1_bit_slice_154521_comb;
  wire [1:0] p1_bit_slice_154522_comb;
  wire [1:0] p1_bit_slice_154523_comb;
  wire [1:0] p1_bit_slice_154524_comb;
  wire [1:0] p1_bit_slice_154525_comb;
  wire [1:0] p1_bit_slice_154526_comb;
  wire [1:0] p1_bit_slice_154527_comb;
  wire [1:0] p1_bit_slice_154528_comb;
  wire [1:0] p1_bit_slice_154529_comb;
  wire [1:0] p1_bit_slice_154530_comb;
  wire [1:0] p1_bit_slice_154531_comb;
  wire [1:0] p1_bit_slice_154532_comb;
  wire [1:0] p1_bit_slice_154533_comb;
  wire [1:0] p1_bit_slice_154534_comb;
  wire [1:0] p1_bit_slice_154535_comb;
  wire [1:0] p1_bit_slice_154536_comb;
  wire [1:0] p1_bit_slice_154537_comb;
  wire [1:0] p1_bit_slice_154538_comb;
  wire [1:0] p1_bit_slice_154539_comb;
  wire [1:0] p1_bit_slice_154540_comb;
  wire [1:0] p1_bit_slice_154541_comb;
  wire [1:0] p1_bit_slice_154542_comb;
  wire [1:0] p1_bit_slice_154543_comb;
  wire [1:0] p1_bit_slice_154544_comb;
  wire [1:0] p1_bit_slice_154545_comb;
  wire [1:0] p1_bit_slice_154546_comb;
  wire [1:0] p1_bit_slice_154547_comb;
  wire [1:0] p1_bit_slice_154548_comb;
  wire [1:0] p1_bit_slice_154549_comb;
  wire [1:0] p1_bit_slice_154550_comb;
  wire [1:0] p1_bit_slice_154551_comb;
  wire [1:0] p1_bit_slice_154552_comb;
  wire [1:0] p1_bit_slice_154553_comb;
  wire [1:0] p1_bit_slice_154554_comb;
  wire [1:0] p1_bit_slice_154555_comb;
  wire [1:0] p1_bit_slice_154556_comb;
  wire [1:0] p1_bit_slice_154557_comb;
  wire [1:0] p1_bit_slice_154558_comb;
  wire [1:0] p1_bit_slice_154559_comb;
  wire [1:0] p1_bit_slice_154560_comb;
  wire [1:0] p1_bit_slice_154561_comb;
  wire [1:0] p1_bit_slice_154562_comb;
  wire [1:0] p1_bit_slice_154563_comb;
  wire [1:0] p1_bit_slice_154564_comb;
  wire [1:0] p1_bit_slice_154565_comb;
  wire [1:0] p1_bit_slice_154566_comb;
  wire [1:0] p1_bit_slice_154567_comb;
  wire [1:0] p1_bit_slice_154568_comb;
  wire [1:0] p1_bit_slice_154569_comb;
  wire [1:0] p1_bit_slice_154570_comb;
  wire [1:0] p1_bit_slice_154571_comb;
  wire [1:0] p1_bit_slice_154572_comb;
  wire [1:0] p1_bit_slice_154573_comb;
  wire [1:0] p1_bit_slice_154574_comb;
  wire [1:0] p1_bit_slice_154575_comb;
  wire [1:0] p1_bit_slice_154576_comb;
  wire [1:0] p1_bit_slice_154577_comb;
  wire [1:0] p1_bit_slice_154578_comb;
  wire [2:0] p1_add_154707_comb;
  wire [2:0] p1_add_154708_comb;
  wire [2:0] p1_add_154709_comb;
  wire [2:0] p1_add_154710_comb;
  wire [2:0] p1_add_154711_comb;
  wire [2:0] p1_add_154712_comb;
  wire [2:0] p1_add_154713_comb;
  wire [2:0] p1_add_154714_comb;
  wire [2:0] p1_add_154715_comb;
  wire [2:0] p1_add_154716_comb;
  wire [2:0] p1_add_154717_comb;
  wire [2:0] p1_add_154718_comb;
  wire [2:0] p1_add_154719_comb;
  wire [2:0] p1_add_154720_comb;
  wire [2:0] p1_add_154721_comb;
  wire [2:0] p1_add_154722_comb;
  wire [2:0] p1_add_154723_comb;
  wire [2:0] p1_add_154724_comb;
  wire [2:0] p1_add_154725_comb;
  wire [2:0] p1_add_154726_comb;
  wire [2:0] p1_add_154727_comb;
  wire [2:0] p1_add_154728_comb;
  wire [2:0] p1_add_154729_comb;
  wire [2:0] p1_add_154730_comb;
  wire [2:0] p1_add_154731_comb;
  wire [2:0] p1_add_154732_comb;
  wire [2:0] p1_add_154733_comb;
  wire [2:0] p1_add_154734_comb;
  wire [2:0] p1_add_154735_comb;
  wire [2:0] p1_add_154736_comb;
  wire [2:0] p1_add_154737_comb;
  wire [2:0] p1_add_154738_comb;
  wire [2:0] p1_add_154739_comb;
  wire [2:0] p1_add_154740_comb;
  wire [2:0] p1_add_154741_comb;
  wire [2:0] p1_add_154742_comb;
  wire [2:0] p1_add_154743_comb;
  wire [2:0] p1_add_154744_comb;
  wire [2:0] p1_add_154745_comb;
  wire [2:0] p1_add_154746_comb;
  wire [2:0] p1_add_154747_comb;
  wire [2:0] p1_add_154748_comb;
  wire [2:0] p1_add_154749_comb;
  wire [2:0] p1_add_154750_comb;
  wire [2:0] p1_add_154751_comb;
  wire [2:0] p1_add_154752_comb;
  wire [2:0] p1_add_154753_comb;
  wire [2:0] p1_add_154754_comb;
  wire [2:0] p1_add_154755_comb;
  wire [2:0] p1_add_154756_comb;
  wire [2:0] p1_add_154757_comb;
  wire [2:0] p1_add_154758_comb;
  wire [2:0] p1_add_154759_comb;
  wire [2:0] p1_add_154760_comb;
  wire [2:0] p1_add_154761_comb;
  wire [2:0] p1_add_154762_comb;
  wire [2:0] p1_add_154763_comb;
  wire [2:0] p1_add_154764_comb;
  wire [2:0] p1_add_154765_comb;
  wire [2:0] p1_add_154766_comb;
  wire [2:0] p1_add_154767_comb;
  wire [2:0] p1_add_154768_comb;
  wire [2:0] p1_add_154769_comb;
  wire [2:0] p1_add_154770_comb;
  wire [7:0] p1_clipped__136_comb;
  wire [7:0] p1_clipped__152_comb;
  wire [7:0] p1_clipped__168_comb;
  wire [7:0] p1_clipped__184_comb;
  wire [7:0] p1_clipped__200_comb;
  wire [7:0] p1_clipped__216_comb;
  wire [7:0] p1_clipped__232_comb;
  wire [7:0] p1_clipped__248_comb;
  wire [7:0] p1_clipped__137_comb;
  wire [7:0] p1_clipped__153_comb;
  wire [7:0] p1_clipped__169_comb;
  wire [7:0] p1_clipped__185_comb;
  wire [7:0] p1_clipped__201_comb;
  wire [7:0] p1_clipped__217_comb;
  wire [7:0] p1_clipped__233_comb;
  wire [7:0] p1_clipped__249_comb;
  wire [7:0] p1_clipped__138_comb;
  wire [7:0] p1_clipped__154_comb;
  wire [7:0] p1_clipped__170_comb;
  wire [7:0] p1_clipped__186_comb;
  wire [7:0] p1_clipped__202_comb;
  wire [7:0] p1_clipped__218_comb;
  wire [7:0] p1_clipped__234_comb;
  wire [7:0] p1_clipped__250_comb;
  wire [7:0] p1_clipped__139_comb;
  wire [7:0] p1_clipped__155_comb;
  wire [7:0] p1_clipped__171_comb;
  wire [7:0] p1_clipped__187_comb;
  wire [7:0] p1_clipped__203_comb;
  wire [7:0] p1_clipped__219_comb;
  wire [7:0] p1_clipped__235_comb;
  wire [7:0] p1_clipped__251_comb;
  wire [7:0] p1_clipped__140_comb;
  wire [7:0] p1_clipped__156_comb;
  wire [7:0] p1_clipped__172_comb;
  wire [7:0] p1_clipped__188_comb;
  wire [7:0] p1_clipped__204_comb;
  wire [7:0] p1_clipped__220_comb;
  wire [7:0] p1_clipped__236_comb;
  wire [7:0] p1_clipped__252_comb;
  wire [7:0] p1_clipped__141_comb;
  wire [7:0] p1_clipped__157_comb;
  wire [7:0] p1_clipped__173_comb;
  wire [7:0] p1_clipped__189_comb;
  wire [7:0] p1_clipped__205_comb;
  wire [7:0] p1_clipped__221_comb;
  wire [7:0] p1_clipped__237_comb;
  wire [7:0] p1_clipped__253_comb;
  wire [7:0] p1_clipped__142_comb;
  wire [7:0] p1_clipped__158_comb;
  wire [7:0] p1_clipped__174_comb;
  wire [7:0] p1_clipped__190_comb;
  wire [7:0] p1_clipped__206_comb;
  wire [7:0] p1_clipped__222_comb;
  wire [7:0] p1_clipped__238_comb;
  wire [7:0] p1_clipped__254_comb;
  wire [7:0] p1_clipped__143_comb;
  wire [7:0] p1_clipped__159_comb;
  wire [7:0] p1_clipped__175_comb;
  wire [7:0] p1_clipped__191_comb;
  wire [7:0] p1_clipped__207_comb;
  wire [7:0] p1_clipped__223_comb;
  wire [7:0] p1_clipped__239_comb;
  wire [7:0] p1_clipped__255_comb;
  wire [7:0] p1_array_155155_comb[0:7];
  wire [7:0] p1_array_155156_comb[0:7];
  wire [7:0] p1_array_155157_comb[0:7];
  wire [7:0] p1_array_155158_comb[0:7];
  wire [7:0] p1_array_155159_comb[0:7];
  wire [7:0] p1_array_155160_comb[0:7];
  wire [7:0] p1_array_155161_comb[0:7];
  wire [7:0] p1_array_155162_comb[0:7];
  wire [7:0] p1_col_transformed_comb[0:7][0:7];
  assign p1_array_index_133923_comb = p0_x[3'h2][3'h2];
  assign p1_array_index_133924_comb = p0_x[3'h2][3'h5];
  assign p1_array_index_133925_comb = p0_x[3'h5][3'h2];
  assign p1_array_index_133926_comb = p0_x[3'h5][3'h5];
  assign p1_array_index_133927_comb = p0_x[3'h2][3'h0];
  assign p1_array_index_133928_comb = p0_x[3'h2][3'h1];
  assign p1_array_index_133929_comb = p0_x[3'h2][3'h3];
  assign p1_array_index_133930_comb = p0_x[3'h2][3'h4];
  assign p1_array_index_133931_comb = p0_x[3'h2][3'h6];
  assign p1_array_index_133932_comb = p0_x[3'h2][3'h7];
  assign p1_array_index_133933_comb = p0_x[3'h5][3'h0];
  assign p1_array_index_133934_comb = p0_x[3'h5][3'h1];
  assign p1_array_index_133935_comb = p0_x[3'h5][3'h3];
  assign p1_array_index_133936_comb = p0_x[3'h5][3'h4];
  assign p1_array_index_133937_comb = p0_x[3'h5][3'h6];
  assign p1_array_index_133938_comb = p0_x[3'h5][3'h7];
  assign p1_array_index_133939_comb = p0_x[3'h0][3'h2];
  assign p1_array_index_133940_comb = p0_x[3'h0][3'h5];
  assign p1_array_index_133941_comb = p0_x[3'h1][3'h2];
  assign p1_array_index_133942_comb = p0_x[3'h1][3'h5];
  assign p1_array_index_133943_comb = p0_x[3'h3][3'h2];
  assign p1_array_index_133944_comb = p0_x[3'h3][3'h5];
  assign p1_array_index_133945_comb = p0_x[3'h4][3'h2];
  assign p1_array_index_133946_comb = p0_x[3'h4][3'h5];
  assign p1_array_index_133947_comb = p0_x[3'h6][3'h2];
  assign p1_array_index_133948_comb = p0_x[3'h6][3'h5];
  assign p1_array_index_133949_comb = p0_x[3'h7][3'h2];
  assign p1_array_index_133950_comb = p0_x[3'h7][3'h5];
  assign p1_array_index_133951_comb = p0_x[3'h0][3'h0];
  assign p1_array_index_133952_comb = p0_x[3'h0][3'h1];
  assign p1_array_index_133953_comb = p0_x[3'h0][3'h3];
  assign p1_array_index_133954_comb = p0_x[3'h0][3'h4];
  assign p1_array_index_133955_comb = p0_x[3'h0][3'h6];
  assign p1_array_index_133956_comb = p0_x[3'h0][3'h7];
  assign p1_array_index_133957_comb = p0_x[3'h1][3'h0];
  assign p1_array_index_133958_comb = p0_x[3'h1][3'h1];
  assign p1_array_index_133959_comb = p0_x[3'h1][3'h3];
  assign p1_array_index_133960_comb = p0_x[3'h1][3'h4];
  assign p1_array_index_133961_comb = p0_x[3'h1][3'h6];
  assign p1_array_index_133962_comb = p0_x[3'h1][3'h7];
  assign p1_array_index_133963_comb = p0_x[3'h3][3'h0];
  assign p1_array_index_133964_comb = p0_x[3'h3][3'h1];
  assign p1_array_index_133965_comb = p0_x[3'h3][3'h3];
  assign p1_array_index_133966_comb = p0_x[3'h3][3'h4];
  assign p1_array_index_133967_comb = p0_x[3'h3][3'h6];
  assign p1_array_index_133968_comb = p0_x[3'h3][3'h7];
  assign p1_array_index_133969_comb = p0_x[3'h4][3'h0];
  assign p1_array_index_133970_comb = p0_x[3'h4][3'h1];
  assign p1_array_index_133971_comb = p0_x[3'h4][3'h3];
  assign p1_array_index_133972_comb = p0_x[3'h4][3'h4];
  assign p1_array_index_133973_comb = p0_x[3'h4][3'h6];
  assign p1_array_index_133974_comb = p0_x[3'h4][3'h7];
  assign p1_array_index_133975_comb = p0_x[3'h6][3'h0];
  assign p1_array_index_133976_comb = p0_x[3'h6][3'h1];
  assign p1_array_index_133977_comb = p0_x[3'h6][3'h3];
  assign p1_array_index_133978_comb = p0_x[3'h6][3'h4];
  assign p1_array_index_133979_comb = p0_x[3'h6][3'h6];
  assign p1_array_index_133980_comb = p0_x[3'h6][3'h7];
  assign p1_array_index_133981_comb = p0_x[3'h7][3'h0];
  assign p1_array_index_133982_comb = p0_x[3'h7][3'h1];
  assign p1_array_index_133983_comb = p0_x[3'h7][3'h3];
  assign p1_array_index_133984_comb = p0_x[3'h7][3'h4];
  assign p1_array_index_133985_comb = p0_x[3'h7][3'h6];
  assign p1_array_index_133986_comb = p0_x[3'h7][3'h7];
  assign p1_shifted__18_squeezed_comb = {~p1_array_index_133923_comb[7], p1_array_index_133923_comb[6:0]};
  assign p1_shifted__21_squeezed_comb = {~p1_array_index_133924_comb[7], p1_array_index_133924_comb[6:0]};
  assign p1_shifted__42_squeezed_comb = {~p1_array_index_133925_comb[7], p1_array_index_133925_comb[6:0]};
  assign p1_shifted__45_squeezed_comb = {~p1_array_index_133926_comb[7], p1_array_index_133926_comb[6:0]};
  assign p1_shifted__16_squeezed_comb = {~p1_array_index_133927_comb[7], p1_array_index_133927_comb[6:0]};
  assign p1_shifted__17_squeezed_comb = {~p1_array_index_133928_comb[7], p1_array_index_133928_comb[6:0]};
  assign p1_shifted__19_squeezed_comb = {~p1_array_index_133929_comb[7], p1_array_index_133929_comb[6:0]};
  assign p1_shifted__20_squeezed_comb = {~p1_array_index_133930_comb[7], p1_array_index_133930_comb[6:0]};
  assign p1_shifted__22_squeezed_comb = {~p1_array_index_133931_comb[7], p1_array_index_133931_comb[6:0]};
  assign p1_shifted__23_squeezed_comb = {~p1_array_index_133932_comb[7], p1_array_index_133932_comb[6:0]};
  assign p1_shifted__40_squeezed_comb = {~p1_array_index_133933_comb[7], p1_array_index_133933_comb[6:0]};
  assign p1_shifted__41_squeezed_comb = {~p1_array_index_133934_comb[7], p1_array_index_133934_comb[6:0]};
  assign p1_shifted__43_squeezed_comb = {~p1_array_index_133935_comb[7], p1_array_index_133935_comb[6:0]};
  assign p1_shifted__44_squeezed_comb = {~p1_array_index_133936_comb[7], p1_array_index_133936_comb[6:0]};
  assign p1_shifted__46_squeezed_comb = {~p1_array_index_133937_comb[7], p1_array_index_133937_comb[6:0]};
  assign p1_shifted__47_squeezed_comb = {~p1_array_index_133938_comb[7], p1_array_index_133938_comb[6:0]};
  assign p1_shifted__2_squeezed_comb = {~p1_array_index_133939_comb[7], p1_array_index_133939_comb[6:0]};
  assign p1_shifted__5_squeezed_comb = {~p1_array_index_133940_comb[7], p1_array_index_133940_comb[6:0]};
  assign p1_shifted__10_squeezed_comb = {~p1_array_index_133941_comb[7], p1_array_index_133941_comb[6:0]};
  assign p1_shifted__13_squeezed_comb = {~p1_array_index_133942_comb[7], p1_array_index_133942_comb[6:0]};
  assign p1_shifted__26_squeezed_comb = {~p1_array_index_133943_comb[7], p1_array_index_133943_comb[6:0]};
  assign p1_shifted__29_squeezed_comb = {~p1_array_index_133944_comb[7], p1_array_index_133944_comb[6:0]};
  assign p1_shifted__34_squeezed_comb = {~p1_array_index_133945_comb[7], p1_array_index_133945_comb[6:0]};
  assign p1_shifted__37_squeezed_comb = {~p1_array_index_133946_comb[7], p1_array_index_133946_comb[6:0]};
  assign p1_shifted__50_squeezed_comb = {~p1_array_index_133947_comb[7], p1_array_index_133947_comb[6:0]};
  assign p1_shifted__53_squeezed_comb = {~p1_array_index_133948_comb[7], p1_array_index_133948_comb[6:0]};
  assign p1_shifted__58_squeezed_comb = {~p1_array_index_133949_comb[7], p1_array_index_133949_comb[6:0]};
  assign p1_shifted__61_squeezed_comb = {~p1_array_index_133950_comb[7], p1_array_index_133950_comb[6:0]};
  assign p1_shifted_squeezed_comb = {~p1_array_index_133951_comb[7], p1_array_index_133951_comb[6:0]};
  assign p1_shifted__1_squeezed_comb = {~p1_array_index_133952_comb[7], p1_array_index_133952_comb[6:0]};
  assign p1_shifted__3_squeezed_comb = {~p1_array_index_133953_comb[7], p1_array_index_133953_comb[6:0]};
  assign p1_shifted__4_squeezed_comb = {~p1_array_index_133954_comb[7], p1_array_index_133954_comb[6:0]};
  assign p1_shifted__6_squeezed_comb = {~p1_array_index_133955_comb[7], p1_array_index_133955_comb[6:0]};
  assign p1_shifted__7_squeezed_comb = {~p1_array_index_133956_comb[7], p1_array_index_133956_comb[6:0]};
  assign p1_shifted__8_squeezed_comb = {~p1_array_index_133957_comb[7], p1_array_index_133957_comb[6:0]};
  assign p1_shifted__9_squeezed_comb = {~p1_array_index_133958_comb[7], p1_array_index_133958_comb[6:0]};
  assign p1_shifted__11_squeezed_comb = {~p1_array_index_133959_comb[7], p1_array_index_133959_comb[6:0]};
  assign p1_shifted__12_squeezed_comb = {~p1_array_index_133960_comb[7], p1_array_index_133960_comb[6:0]};
  assign p1_shifted__14_squeezed_comb = {~p1_array_index_133961_comb[7], p1_array_index_133961_comb[6:0]};
  assign p1_shifted__15_squeezed_comb = {~p1_array_index_133962_comb[7], p1_array_index_133962_comb[6:0]};
  assign p1_shifted__24_squeezed_comb = {~p1_array_index_133963_comb[7], p1_array_index_133963_comb[6:0]};
  assign p1_shifted__25_squeezed_comb = {~p1_array_index_133964_comb[7], p1_array_index_133964_comb[6:0]};
  assign p1_shifted__27_squeezed_comb = {~p1_array_index_133965_comb[7], p1_array_index_133965_comb[6:0]};
  assign p1_shifted__28_squeezed_comb = {~p1_array_index_133966_comb[7], p1_array_index_133966_comb[6:0]};
  assign p1_shifted__30_squeezed_comb = {~p1_array_index_133967_comb[7], p1_array_index_133967_comb[6:0]};
  assign p1_shifted__31_squeezed_comb = {~p1_array_index_133968_comb[7], p1_array_index_133968_comb[6:0]};
  assign p1_shifted__32_squeezed_comb = {~p1_array_index_133969_comb[7], p1_array_index_133969_comb[6:0]};
  assign p1_shifted__33_squeezed_comb = {~p1_array_index_133970_comb[7], p1_array_index_133970_comb[6:0]};
  assign p1_shifted__35_squeezed_comb = {~p1_array_index_133971_comb[7], p1_array_index_133971_comb[6:0]};
  assign p1_shifted__36_squeezed_comb = {~p1_array_index_133972_comb[7], p1_array_index_133972_comb[6:0]};
  assign p1_shifted__38_squeezed_comb = {~p1_array_index_133973_comb[7], p1_array_index_133973_comb[6:0]};
  assign p1_shifted__39_squeezed_comb = {~p1_array_index_133974_comb[7], p1_array_index_133974_comb[6:0]};
  assign p1_shifted__48_squeezed_comb = {~p1_array_index_133975_comb[7], p1_array_index_133975_comb[6:0]};
  assign p1_shifted__49_squeezed_comb = {~p1_array_index_133976_comb[7], p1_array_index_133976_comb[6:0]};
  assign p1_shifted__51_squeezed_comb = {~p1_array_index_133977_comb[7], p1_array_index_133977_comb[6:0]};
  assign p1_shifted__52_squeezed_comb = {~p1_array_index_133978_comb[7], p1_array_index_133978_comb[6:0]};
  assign p1_shifted__54_squeezed_comb = {~p1_array_index_133979_comb[7], p1_array_index_133979_comb[6:0]};
  assign p1_shifted__55_squeezed_comb = {~p1_array_index_133980_comb[7], p1_array_index_133980_comb[6:0]};
  assign p1_shifted__56_squeezed_comb = {~p1_array_index_133981_comb[7], p1_array_index_133981_comb[6:0]};
  assign p1_shifted__57_squeezed_comb = {~p1_array_index_133982_comb[7], p1_array_index_133982_comb[6:0]};
  assign p1_shifted__59_squeezed_comb = {~p1_array_index_133983_comb[7], p1_array_index_133983_comb[6:0]};
  assign p1_shifted__60_squeezed_comb = {~p1_array_index_133984_comb[7], p1_array_index_133984_comb[6:0]};
  assign p1_shifted__62_squeezed_comb = {~p1_array_index_133985_comb[7], p1_array_index_133985_comb[6:0]};
  assign p1_shifted__63_squeezed_comb = {~p1_array_index_133986_comb[7], p1_array_index_133986_comb[6:0]};
  assign p1_smul_57362_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__18_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___8_comb = 9'h000;
  assign p1_smul_57368_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__21_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___11_comb = 9'h000;
  assign p1_smul_57410_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__42_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___20_comb = 9'h000;
  assign p1_smul_57416_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__45_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___23_comb = 9'h000;
  assign p1_smul_57486_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__16_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___8_comb = 10'h000;
  assign p1_smul_57488_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__17_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___40_comb = 9'h000;
  assign p1_smul_57490_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__18_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___41_comb = 9'h000;
  assign p1_smul_57492_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__19_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___9_comb = 10'h000;
  assign p1_smul_57494_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__20_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___10_comb = 10'h000;
  assign p1_smul_57496_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__21_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___42_comb = 9'h000;
  assign p1_smul_57498_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__22_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___43_comb = 9'h000;
  assign p1_smul_57500_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__23_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___11_comb = 10'h000;
  assign p1_smul_57534_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__40_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___20_comb = 10'h000;
  assign p1_smul_57536_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__41_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___52_comb = 9'h000;
  assign p1_smul_57538_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__42_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___53_comb = 9'h000;
  assign p1_smul_57540_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__43_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___21_comb = 10'h000;
  assign p1_smul_57542_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__44_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___22_comb = 10'h000;
  assign p1_smul_57544_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__45_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___54_comb = 9'h000;
  assign p1_smul_57546_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__46_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___55_comb = 9'h000;
  assign p1_smul_57548_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__47_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___23_comb = 10'h000;
  assign p1_smul_57620_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__19_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___73_comb = 9'h000;
  assign p1_smul_57622_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__20_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___74_comb = 9'h000;
  assign p1_smul_57668_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__43_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___85_comb = 9'h000;
  assign p1_smul_57670_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__44_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___86_comb = 9'h000;
  assign p1_smul_57870_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__16_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___104_comb = 9'h000;
  assign p1_smul_57884_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__23_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___107_comb = 9'h000;
  assign p1_smul_57918_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__40_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___116_comb = 9'h000;
  assign p1_smul_57932_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__47_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___119_comb = 9'h000;
  assign p1_smul_57998_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__16_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___136_comb = 9'h000;
  assign p1_smul_58000_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__17_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___40_comb = 10'h000;
  assign p1_smul_58002_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__18_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___137_comb = 9'h000;
  assign p1_smul_58004_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__19_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___41_comb = 10'h000;
  assign p1_smul_58006_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__20_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___42_comb = 10'h000;
  assign p1_smul_58008_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__21_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___138_comb = 9'h000;
  assign p1_smul_58010_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__22_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___43_comb = 10'h000;
  assign p1_smul_58012_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__23_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___139_comb = 9'h000;
  assign p1_smul_58046_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__40_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___148_comb = 9'h000;
  assign p1_smul_58048_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__41_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___52_comb = 10'h000;
  assign p1_smul_58050_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__42_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___149_comb = 9'h000;
  assign p1_smul_58052_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__43_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___53_comb = 10'h000;
  assign p1_smul_58054_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__44_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___54_comb = 10'h000;
  assign p1_smul_58056_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__45_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___150_comb = 9'h000;
  assign p1_smul_58058_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__46_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___55_comb = 10'h000;
  assign p1_smul_58060_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__47_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___151_comb = 9'h000;
  assign p1_smul_58128_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__17_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___169_comb = 9'h000;
  assign p1_smul_58138_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__22_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___170_comb = 9'h000;
  assign p1_smul_58176_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__41_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___181_comb = 9'h000;
  assign p1_smul_58186_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__46_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___182_comb = 9'h000;
  assign p1_smul_57330_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__2_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits__comb = 9'h000;
  assign p1_smul_57336_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__5_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___3_comb = 9'h000;
  assign p1_smul_57346_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__10_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___4_comb = 9'h000;
  assign p1_smul_57352_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__13_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___7_comb = 9'h000;
  assign p1_smul_57378_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__26_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___12_comb = 9'h000;
  assign p1_smul_57384_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__29_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___15_comb = 9'h000;
  assign p1_smul_57394_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__34_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___16_comb = 9'h000;
  assign p1_smul_57400_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__37_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___19_comb = 9'h000;
  assign p1_smul_57426_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__50_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___24_comb = 9'h000;
  assign p1_smul_57432_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__53_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___27_comb = 9'h000;
  assign p1_smul_57442_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__58_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___28_comb = 9'h000;
  assign p1_smul_57448_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__61_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___31_comb = 9'h000;
  assign p1_smul_57454_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits__comb = 10'h000;
  assign p1_smul_57456_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__1_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___32_comb = 9'h000;
  assign p1_smul_57458_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__2_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___33_comb = 9'h000;
  assign p1_smul_57460_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__3_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___1_comb = 10'h000;
  assign p1_smul_57462_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__4_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___2_comb = 10'h000;
  assign p1_smul_57464_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__5_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___34_comb = 9'h000;
  assign p1_smul_57466_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__6_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___35_comb = 9'h000;
  assign p1_smul_57468_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__7_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___3_comb = 10'h000;
  assign p1_smul_57470_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__8_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___4_comb = 10'h000;
  assign p1_smul_57472_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__9_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___36_comb = 9'h000;
  assign p1_smul_57474_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__10_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___37_comb = 9'h000;
  assign p1_smul_57476_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__11_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___5_comb = 10'h000;
  assign p1_smul_57478_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__12_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___6_comb = 10'h000;
  assign p1_smul_57480_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__13_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___38_comb = 9'h000;
  assign p1_smul_57482_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__14_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___39_comb = 9'h000;
  assign p1_smul_57484_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__15_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___7_comb = 10'h000;
  assign p1_smul_57502_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__24_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___12_comb = 10'h000;
  assign p1_smul_57504_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__25_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___44_comb = 9'h000;
  assign p1_smul_57506_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__26_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___45_comb = 9'h000;
  assign p1_smul_57508_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__27_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___13_comb = 10'h000;
  assign p1_smul_57510_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__28_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___14_comb = 10'h000;
  assign p1_smul_57512_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__29_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___46_comb = 9'h000;
  assign p1_smul_57514_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__30_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___47_comb = 9'h000;
  assign p1_smul_57516_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__31_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___15_comb = 10'h000;
  assign p1_smul_57518_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__32_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___16_comb = 10'h000;
  assign p1_smul_57520_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__33_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___48_comb = 9'h000;
  assign p1_smul_57522_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__34_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___49_comb = 9'h000;
  assign p1_smul_57524_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__35_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___17_comb = 10'h000;
  assign p1_smul_57526_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__36_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___18_comb = 10'h000;
  assign p1_smul_57528_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__37_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___50_comb = 9'h000;
  assign p1_smul_57530_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__38_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___51_comb = 9'h000;
  assign p1_smul_57532_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__39_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___19_comb = 10'h000;
  assign p1_smul_57550_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__48_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___24_comb = 10'h000;
  assign p1_smul_57552_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__49_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___56_comb = 9'h000;
  assign p1_smul_57554_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__50_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___57_comb = 9'h000;
  assign p1_smul_57556_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__51_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___25_comb = 10'h000;
  assign p1_smul_57558_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__52_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___26_comb = 10'h000;
  assign p1_smul_57560_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__53_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___58_comb = 9'h000;
  assign p1_smul_57562_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__54_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___59_comb = 9'h000;
  assign p1_smul_57564_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__55_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___27_comb = 10'h000;
  assign p1_smul_57566_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__56_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___28_comb = 10'h000;
  assign p1_smul_57568_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__57_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___60_comb = 9'h000;
  assign p1_smul_57570_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__58_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___61_comb = 9'h000;
  assign p1_smul_57572_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__59_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___29_comb = 10'h000;
  assign p1_smul_57574_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__60_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___30_comb = 10'h000;
  assign p1_smul_57576_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__61_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___62_comb = 9'h000;
  assign p1_smul_57578_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__62_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___63_comb = 9'h000;
  assign p1_smul_57580_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__63_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___31_comb = 10'h000;
  assign p1_smul_57588_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__3_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___65_comb = 9'h000;
  assign p1_smul_57590_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__4_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___66_comb = 9'h000;
  assign p1_smul_57604_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__11_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___69_comb = 9'h000;
  assign p1_smul_57606_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__12_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___70_comb = 9'h000;
  assign p1_smul_57636_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__27_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___77_comb = 9'h000;
  assign p1_smul_57638_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__28_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___78_comb = 9'h000;
  assign p1_smul_57652_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__35_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___81_comb = 9'h000;
  assign p1_smul_57654_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__36_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___82_comb = 9'h000;
  assign p1_smul_57684_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__51_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___89_comb = 9'h000;
  assign p1_smul_57686_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__52_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___90_comb = 9'h000;
  assign p1_smul_57700_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__59_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___93_comb = 9'h000;
  assign p1_smul_57702_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__60_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___94_comb = 9'h000;
  assign p1_smul_57838_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___96_comb = 9'h000;
  assign p1_smul_57852_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__7_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___99_comb = 9'h000;
  assign p1_smul_57854_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__8_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___100_comb = 9'h000;
  assign p1_smul_57868_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__15_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___103_comb = 9'h000;
  assign p1_smul_57886_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__24_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___108_comb = 9'h000;
  assign p1_smul_57900_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__31_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___111_comb = 9'h000;
  assign p1_smul_57902_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__32_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___112_comb = 9'h000;
  assign p1_smul_57916_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__39_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___115_comb = 9'h000;
  assign p1_smul_57934_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__48_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___120_comb = 9'h000;
  assign p1_smul_57948_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__55_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___123_comb = 9'h000;
  assign p1_smul_57950_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__56_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___124_comb = 9'h000;
  assign p1_smul_57964_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__63_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___127_comb = 9'h000;
  assign p1_smul_57966_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___128_comb = 9'h000;
  assign p1_smul_57968_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__1_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___32_comb = 10'h000;
  assign p1_smul_57970_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__2_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___129_comb = 9'h000;
  assign p1_smul_57972_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__3_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___33_comb = 10'h000;
  assign p1_smul_57974_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__4_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___34_comb = 10'h000;
  assign p1_smul_57976_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__5_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___130_comb = 9'h000;
  assign p1_smul_57978_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__6_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___35_comb = 10'h000;
  assign p1_smul_57980_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__7_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___131_comb = 9'h000;
  assign p1_smul_57982_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__8_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___132_comb = 9'h000;
  assign p1_smul_57984_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__9_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___36_comb = 10'h000;
  assign p1_smul_57986_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__10_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___133_comb = 9'h000;
  assign p1_smul_57988_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__11_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___37_comb = 10'h000;
  assign p1_smul_57990_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__12_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___38_comb = 10'h000;
  assign p1_smul_57992_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__13_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___134_comb = 9'h000;
  assign p1_smul_57994_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__14_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___39_comb = 10'h000;
  assign p1_smul_57996_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__15_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___135_comb = 9'h000;
  assign p1_smul_58014_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__24_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___140_comb = 9'h000;
  assign p1_smul_58016_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__25_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___44_comb = 10'h000;
  assign p1_smul_58018_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__26_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___141_comb = 9'h000;
  assign p1_smul_58020_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__27_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___45_comb = 10'h000;
  assign p1_smul_58022_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__28_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___46_comb = 10'h000;
  assign p1_smul_58024_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__29_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___142_comb = 9'h000;
  assign p1_smul_58026_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__30_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___47_comb = 10'h000;
  assign p1_smul_58028_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__31_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___143_comb = 9'h000;
  assign p1_smul_58030_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__32_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___144_comb = 9'h000;
  assign p1_smul_58032_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__33_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___48_comb = 10'h000;
  assign p1_smul_58034_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__34_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___145_comb = 9'h000;
  assign p1_smul_58036_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__35_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___49_comb = 10'h000;
  assign p1_smul_58038_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__36_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___50_comb = 10'h000;
  assign p1_smul_58040_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__37_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___146_comb = 9'h000;
  assign p1_smul_58042_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__38_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___51_comb = 10'h000;
  assign p1_smul_58044_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__39_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___147_comb = 9'h000;
  assign p1_smul_58062_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__48_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___152_comb = 9'h000;
  assign p1_smul_58064_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__49_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___56_comb = 10'h000;
  assign p1_smul_58066_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__50_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___153_comb = 9'h000;
  assign p1_smul_58068_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__51_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___57_comb = 10'h000;
  assign p1_smul_58070_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__52_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___58_comb = 10'h000;
  assign p1_smul_58072_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__53_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___154_comb = 9'h000;
  assign p1_smul_58074_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__54_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___59_comb = 10'h000;
  assign p1_smul_58076_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__55_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___155_comb = 9'h000;
  assign p1_smul_58078_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__56_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___156_comb = 9'h000;
  assign p1_smul_58080_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__57_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___60_comb = 10'h000;
  assign p1_smul_58082_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__58_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___157_comb = 9'h000;
  assign p1_smul_58084_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__59_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___61_comb = 10'h000;
  assign p1_smul_58086_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__60_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___62_comb = 10'h000;
  assign p1_smul_58088_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__61_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___158_comb = 9'h000;
  assign p1_smul_58090_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__62_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___63_comb = 10'h000;
  assign p1_smul_58092_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__63_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___159_comb = 9'h000;
  assign p1_smul_58096_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__1_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___161_comb = 9'h000;
  assign p1_smul_58106_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__6_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___162_comb = 9'h000;
  assign p1_smul_58112_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__9_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___165_comb = 9'h000;
  assign p1_smul_58122_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__14_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___166_comb = 9'h000;
  assign p1_smul_58144_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__25_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___173_comb = 9'h000;
  assign p1_smul_58154_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__30_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___174_comb = 9'h000;
  assign p1_smul_58160_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__33_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___177_comb = 9'h000;
  assign p1_smul_58170_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__38_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___178_comb = 9'h000;
  assign p1_smul_58192_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__49_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___185_comb = 9'h000;
  assign p1_smul_58202_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__54_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___186_comb = 9'h000;
  assign p1_smul_58208_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__57_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___189_comb = 9'h000;
  assign p1_smul_58218_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__62_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___190_comb = 9'h000;
  assign p1_concat_134899_comb = {p1_smul_57362_NarrowedMult__comb, p1_smul_57330_TrailingBits___8_comb};
  assign p1_smul_57364_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__19_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___9_comb = 9'h000;
  assign p1_smul_57366_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__20_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___10_comb = 9'h000;
  assign p1_concat_134904_comb = {p1_smul_57368_NarrowedMult__comb, p1_smul_57330_TrailingBits___11_comb};
  assign p1_concat_134905_comb = {p1_smul_57410_NarrowedMult__comb, p1_smul_57330_TrailingBits___20_comb};
  assign p1_smul_57412_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__43_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___21_comb = 9'h000;
  assign p1_smul_57414_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__44_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___22_comb = 9'h000;
  assign p1_concat_134910_comb = {p1_smul_57416_NarrowedMult__comb, p1_smul_57330_TrailingBits___23_comb};
  assign p1_concat_134911_comb = {p1_smul_57486_NarrowedMult__comb, p1_smul_57454_TrailingBits___8_comb};
  assign p1_concat_134912_comb = {p1_smul_57488_NarrowedMult__comb, p1_smul_57330_TrailingBits___40_comb};
  assign p1_concat_134913_comb = {p1_smul_57490_NarrowedMult__comb, p1_smul_57330_TrailingBits___41_comb};
  assign p1_concat_134914_comb = {p1_smul_57492_NarrowedMult__comb, p1_smul_57454_TrailingBits___9_comb};
  assign p1_concat_134915_comb = {p1_smul_57494_NarrowedMult__comb, p1_smul_57454_TrailingBits___10_comb};
  assign p1_concat_134916_comb = {p1_smul_57496_NarrowedMult__comb, p1_smul_57330_TrailingBits___42_comb};
  assign p1_concat_134917_comb = {p1_smul_57498_NarrowedMult__comb, p1_smul_57330_TrailingBits___43_comb};
  assign p1_concat_134918_comb = {p1_smul_57500_NarrowedMult__comb, p1_smul_57454_TrailingBits___11_comb};
  assign p1_concat_134919_comb = {p1_smul_57534_NarrowedMult__comb, p1_smul_57454_TrailingBits___20_comb};
  assign p1_concat_134920_comb = {p1_smul_57536_NarrowedMult__comb, p1_smul_57330_TrailingBits___52_comb};
  assign p1_concat_134921_comb = {p1_smul_57538_NarrowedMult__comb, p1_smul_57330_TrailingBits___53_comb};
  assign p1_concat_134922_comb = {p1_smul_57540_NarrowedMult__comb, p1_smul_57454_TrailingBits___21_comb};
  assign p1_concat_134923_comb = {p1_smul_57542_NarrowedMult__comb, p1_smul_57454_TrailingBits___22_comb};
  assign p1_concat_134924_comb = {p1_smul_57544_NarrowedMult__comb, p1_smul_57330_TrailingBits___54_comb};
  assign p1_concat_134925_comb = {p1_smul_57546_NarrowedMult__comb, p1_smul_57330_TrailingBits___55_comb};
  assign p1_concat_134926_comb = {p1_smul_57548_NarrowedMult__comb, p1_smul_57454_TrailingBits___23_comb};
  assign p1_smul_57616_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__17_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___72_comb = 9'h000;
  assign p1_concat_134929_comb = {p1_smul_57620_NarrowedMult__comb, p1_smul_57330_TrailingBits___73_comb};
  assign p1_concat_134930_comb = {p1_smul_57622_NarrowedMult__comb, p1_smul_57330_TrailingBits___74_comb};
  assign p1_smul_57626_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__22_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___75_comb = 9'h000;
  assign p1_smul_57664_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__41_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___84_comb = 9'h000;
  assign p1_concat_134935_comb = {p1_smul_57668_NarrowedMult__comb, p1_smul_57330_TrailingBits___85_comb};
  assign p1_concat_134936_comb = {p1_smul_57670_NarrowedMult__comb, p1_smul_57330_TrailingBits___86_comb};
  assign p1_smul_57674_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__46_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___87_comb = 9'h000;
  assign p1_concat_134939_comb = {p1_smul_57870_NarrowedMult__comb, p1_smul_57330_TrailingBits___104_comb};
  assign p1_smul_57874_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__18_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___105_comb = 9'h000;
  assign p1_smul_57880_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__21_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___106_comb = 9'h000;
  assign p1_concat_134944_comb = {p1_smul_57884_NarrowedMult__comb, p1_smul_57330_TrailingBits___107_comb};
  assign p1_concat_134945_comb = {p1_smul_57918_NarrowedMult__comb, p1_smul_57330_TrailingBits___116_comb};
  assign p1_smul_57922_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__42_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___117_comb = 9'h000;
  assign p1_smul_57928_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__45_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___118_comb = 9'h000;
  assign p1_concat_134950_comb = {p1_smul_57932_NarrowedMult__comb, p1_smul_57330_TrailingBits___119_comb};
  assign p1_concat_134951_comb = {p1_smul_57998_NarrowedMult__comb, p1_smul_57330_TrailingBits___136_comb};
  assign p1_concat_134952_comb = {p1_smul_58000_NarrowedMult__comb, p1_smul_57454_TrailingBits___40_comb};
  assign p1_concat_134953_comb = {p1_smul_58002_NarrowedMult__comb, p1_smul_57330_TrailingBits___137_comb};
  assign p1_concat_134954_comb = {p1_smul_58004_NarrowedMult__comb, p1_smul_57454_TrailingBits___41_comb};
  assign p1_concat_134955_comb = {p1_smul_58006_NarrowedMult__comb, p1_smul_57454_TrailingBits___42_comb};
  assign p1_concat_134956_comb = {p1_smul_58008_NarrowedMult__comb, p1_smul_57330_TrailingBits___138_comb};
  assign p1_concat_134957_comb = {p1_smul_58010_NarrowedMult__comb, p1_smul_57454_TrailingBits___43_comb};
  assign p1_concat_134958_comb = {p1_smul_58012_NarrowedMult__comb, p1_smul_57330_TrailingBits___139_comb};
  assign p1_concat_134959_comb = {p1_smul_58046_NarrowedMult__comb, p1_smul_57330_TrailingBits___148_comb};
  assign p1_concat_134960_comb = {p1_smul_58048_NarrowedMult__comb, p1_smul_57454_TrailingBits___52_comb};
  assign p1_concat_134961_comb = {p1_smul_58050_NarrowedMult__comb, p1_smul_57330_TrailingBits___149_comb};
  assign p1_concat_134962_comb = {p1_smul_58052_NarrowedMult__comb, p1_smul_57454_TrailingBits___53_comb};
  assign p1_concat_134963_comb = {p1_smul_58054_NarrowedMult__comb, p1_smul_57454_TrailingBits___54_comb};
  assign p1_concat_134964_comb = {p1_smul_58056_NarrowedMult__comb, p1_smul_57330_TrailingBits___150_comb};
  assign p1_concat_134965_comb = {p1_smul_58058_NarrowedMult__comb, p1_smul_57454_TrailingBits___55_comb};
  assign p1_concat_134966_comb = {p1_smul_58060_NarrowedMult__comb, p1_smul_57330_TrailingBits___151_comb};
  assign p1_smul_58126_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__16_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___168_comb = 9'h000;
  assign p1_concat_134969_comb = {p1_smul_58128_NarrowedMult__comb, p1_smul_57330_TrailingBits___169_comb};
  assign p1_concat_134970_comb = {p1_smul_58138_NarrowedMult__comb, p1_smul_57330_TrailingBits___170_comb};
  assign p1_smul_58140_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__23_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___171_comb = 9'h000;
  assign p1_smul_58174_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__40_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___180_comb = 9'h000;
  assign p1_concat_134975_comb = {p1_smul_58176_NarrowedMult__comb, p1_smul_57330_TrailingBits___181_comb};
  assign p1_concat_134976_comb = {p1_smul_58186_NarrowedMult__comb, p1_smul_57330_TrailingBits___182_comb};
  assign p1_smul_58188_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__47_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___183_comb = 9'h000;
  assign p1_concat_135027_comb = {p1_smul_57330_NarrowedMult__comb, p1_smul_57330_TrailingBits__comb};
  assign p1_smul_57332_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__3_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___1_comb = 9'h000;
  assign p1_smul_57334_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__4_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___2_comb = 9'h000;
  assign p1_concat_135032_comb = {p1_smul_57336_NarrowedMult__comb, p1_smul_57330_TrailingBits___3_comb};
  assign p1_concat_135033_comb = {p1_smul_57346_NarrowedMult__comb, p1_smul_57330_TrailingBits___4_comb};
  assign p1_smul_57348_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__11_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___5_comb = 9'h000;
  assign p1_smul_57350_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__12_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___6_comb = 9'h000;
  assign p1_concat_135038_comb = {p1_smul_57352_NarrowedMult__comb, p1_smul_57330_TrailingBits___7_comb};
  assign p1_concat_135039_comb = {p1_smul_57378_NarrowedMult__comb, p1_smul_57330_TrailingBits___12_comb};
  assign p1_smul_57380_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__27_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___13_comb = 9'h000;
  assign p1_smul_57382_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__28_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___14_comb = 9'h000;
  assign p1_concat_135044_comb = {p1_smul_57384_NarrowedMult__comb, p1_smul_57330_TrailingBits___15_comb};
  assign p1_concat_135045_comb = {p1_smul_57394_NarrowedMult__comb, p1_smul_57330_TrailingBits___16_comb};
  assign p1_smul_57396_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__35_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___17_comb = 9'h000;
  assign p1_smul_57398_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__36_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___18_comb = 9'h000;
  assign p1_concat_135050_comb = {p1_smul_57400_NarrowedMult__comb, p1_smul_57330_TrailingBits___19_comb};
  assign p1_concat_135051_comb = {p1_smul_57426_NarrowedMult__comb, p1_smul_57330_TrailingBits___24_comb};
  assign p1_smul_57428_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__51_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___25_comb = 9'h000;
  assign p1_smul_57430_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__52_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___26_comb = 9'h000;
  assign p1_concat_135056_comb = {p1_smul_57432_NarrowedMult__comb, p1_smul_57330_TrailingBits___27_comb};
  assign p1_concat_135057_comb = {p1_smul_57442_NarrowedMult__comb, p1_smul_57330_TrailingBits___28_comb};
  assign p1_smul_57444_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__59_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___29_comb = 9'h000;
  assign p1_smul_57446_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__60_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___30_comb = 9'h000;
  assign p1_concat_135062_comb = {p1_smul_57448_NarrowedMult__comb, p1_smul_57330_TrailingBits___31_comb};
  assign p1_concat_135063_comb = {p1_smul_57454_NarrowedMult__comb, p1_smul_57454_TrailingBits__comb};
  assign p1_concat_135064_comb = {p1_smul_57456_NarrowedMult__comb, p1_smul_57330_TrailingBits___32_comb};
  assign p1_concat_135065_comb = {p1_smul_57458_NarrowedMult__comb, p1_smul_57330_TrailingBits___33_comb};
  assign p1_concat_135066_comb = {p1_smul_57460_NarrowedMult__comb, p1_smul_57454_TrailingBits___1_comb};
  assign p1_concat_135067_comb = {p1_smul_57462_NarrowedMult__comb, p1_smul_57454_TrailingBits___2_comb};
  assign p1_concat_135068_comb = {p1_smul_57464_NarrowedMult__comb, p1_smul_57330_TrailingBits___34_comb};
  assign p1_concat_135069_comb = {p1_smul_57466_NarrowedMult__comb, p1_smul_57330_TrailingBits___35_comb};
  assign p1_concat_135070_comb = {p1_smul_57468_NarrowedMult__comb, p1_smul_57454_TrailingBits___3_comb};
  assign p1_concat_135071_comb = {p1_smul_57470_NarrowedMult__comb, p1_smul_57454_TrailingBits___4_comb};
  assign p1_concat_135072_comb = {p1_smul_57472_NarrowedMult__comb, p1_smul_57330_TrailingBits___36_comb};
  assign p1_concat_135073_comb = {p1_smul_57474_NarrowedMult__comb, p1_smul_57330_TrailingBits___37_comb};
  assign p1_concat_135074_comb = {p1_smul_57476_NarrowedMult__comb, p1_smul_57454_TrailingBits___5_comb};
  assign p1_concat_135075_comb = {p1_smul_57478_NarrowedMult__comb, p1_smul_57454_TrailingBits___6_comb};
  assign p1_concat_135076_comb = {p1_smul_57480_NarrowedMult__comb, p1_smul_57330_TrailingBits___38_comb};
  assign p1_concat_135077_comb = {p1_smul_57482_NarrowedMult__comb, p1_smul_57330_TrailingBits___39_comb};
  assign p1_concat_135078_comb = {p1_smul_57484_NarrowedMult__comb, p1_smul_57454_TrailingBits___7_comb};
  assign p1_concat_135079_comb = {p1_smul_57502_NarrowedMult__comb, p1_smul_57454_TrailingBits___12_comb};
  assign p1_concat_135080_comb = {p1_smul_57504_NarrowedMult__comb, p1_smul_57330_TrailingBits___44_comb};
  assign p1_concat_135081_comb = {p1_smul_57506_NarrowedMult__comb, p1_smul_57330_TrailingBits___45_comb};
  assign p1_concat_135082_comb = {p1_smul_57508_NarrowedMult__comb, p1_smul_57454_TrailingBits___13_comb};
  assign p1_concat_135083_comb = {p1_smul_57510_NarrowedMult__comb, p1_smul_57454_TrailingBits___14_comb};
  assign p1_concat_135084_comb = {p1_smul_57512_NarrowedMult__comb, p1_smul_57330_TrailingBits___46_comb};
  assign p1_concat_135085_comb = {p1_smul_57514_NarrowedMult__comb, p1_smul_57330_TrailingBits___47_comb};
  assign p1_concat_135086_comb = {p1_smul_57516_NarrowedMult__comb, p1_smul_57454_TrailingBits___15_comb};
  assign p1_concat_135087_comb = {p1_smul_57518_NarrowedMult__comb, p1_smul_57454_TrailingBits___16_comb};
  assign p1_concat_135088_comb = {p1_smul_57520_NarrowedMult__comb, p1_smul_57330_TrailingBits___48_comb};
  assign p1_concat_135089_comb = {p1_smul_57522_NarrowedMult__comb, p1_smul_57330_TrailingBits___49_comb};
  assign p1_concat_135090_comb = {p1_smul_57524_NarrowedMult__comb, p1_smul_57454_TrailingBits___17_comb};
  assign p1_concat_135091_comb = {p1_smul_57526_NarrowedMult__comb, p1_smul_57454_TrailingBits___18_comb};
  assign p1_concat_135092_comb = {p1_smul_57528_NarrowedMult__comb, p1_smul_57330_TrailingBits___50_comb};
  assign p1_concat_135093_comb = {p1_smul_57530_NarrowedMult__comb, p1_smul_57330_TrailingBits___51_comb};
  assign p1_concat_135094_comb = {p1_smul_57532_NarrowedMult__comb, p1_smul_57454_TrailingBits___19_comb};
  assign p1_concat_135095_comb = {p1_smul_57550_NarrowedMult__comb, p1_smul_57454_TrailingBits___24_comb};
  assign p1_concat_135096_comb = {p1_smul_57552_NarrowedMult__comb, p1_smul_57330_TrailingBits___56_comb};
  assign p1_concat_135097_comb = {p1_smul_57554_NarrowedMult__comb, p1_smul_57330_TrailingBits___57_comb};
  assign p1_concat_135098_comb = {p1_smul_57556_NarrowedMult__comb, p1_smul_57454_TrailingBits___25_comb};
  assign p1_concat_135099_comb = {p1_smul_57558_NarrowedMult__comb, p1_smul_57454_TrailingBits___26_comb};
  assign p1_concat_135100_comb = {p1_smul_57560_NarrowedMult__comb, p1_smul_57330_TrailingBits___58_comb};
  assign p1_concat_135101_comb = {p1_smul_57562_NarrowedMult__comb, p1_smul_57330_TrailingBits___59_comb};
  assign p1_concat_135102_comb = {p1_smul_57564_NarrowedMult__comb, p1_smul_57454_TrailingBits___27_comb};
  assign p1_concat_135103_comb = {p1_smul_57566_NarrowedMult__comb, p1_smul_57454_TrailingBits___28_comb};
  assign p1_concat_135104_comb = {p1_smul_57568_NarrowedMult__comb, p1_smul_57330_TrailingBits___60_comb};
  assign p1_concat_135105_comb = {p1_smul_57570_NarrowedMult__comb, p1_smul_57330_TrailingBits___61_comb};
  assign p1_concat_135106_comb = {p1_smul_57572_NarrowedMult__comb, p1_smul_57454_TrailingBits___29_comb};
  assign p1_concat_135107_comb = {p1_smul_57574_NarrowedMult__comb, p1_smul_57454_TrailingBits___30_comb};
  assign p1_concat_135108_comb = {p1_smul_57576_NarrowedMult__comb, p1_smul_57330_TrailingBits___62_comb};
  assign p1_concat_135109_comb = {p1_smul_57578_NarrowedMult__comb, p1_smul_57330_TrailingBits___63_comb};
  assign p1_concat_135110_comb = {p1_smul_57580_NarrowedMult__comb, p1_smul_57454_TrailingBits___31_comb};
  assign p1_smul_57584_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__1_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___64_comb = 9'h000;
  assign p1_concat_135113_comb = {p1_smul_57588_NarrowedMult__comb, p1_smul_57330_TrailingBits___65_comb};
  assign p1_concat_135114_comb = {p1_smul_57590_NarrowedMult__comb, p1_smul_57330_TrailingBits___66_comb};
  assign p1_smul_57594_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__6_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___67_comb = 9'h000;
  assign p1_smul_57600_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__9_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___68_comb = 9'h000;
  assign p1_concat_135119_comb = {p1_smul_57604_NarrowedMult__comb, p1_smul_57330_TrailingBits___69_comb};
  assign p1_concat_135120_comb = {p1_smul_57606_NarrowedMult__comb, p1_smul_57330_TrailingBits___70_comb};
  assign p1_smul_57610_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__14_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___71_comb = 9'h000;
  assign p1_smul_57632_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__25_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___76_comb = 9'h000;
  assign p1_concat_135125_comb = {p1_smul_57636_NarrowedMult__comb, p1_smul_57330_TrailingBits___77_comb};
  assign p1_concat_135126_comb = {p1_smul_57638_NarrowedMult__comb, p1_smul_57330_TrailingBits___78_comb};
  assign p1_smul_57642_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__30_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___79_comb = 9'h000;
  assign p1_smul_57648_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__33_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___80_comb = 9'h000;
  assign p1_concat_135131_comb = {p1_smul_57652_NarrowedMult__comb, p1_smul_57330_TrailingBits___81_comb};
  assign p1_concat_135132_comb = {p1_smul_57654_NarrowedMult__comb, p1_smul_57330_TrailingBits___82_comb};
  assign p1_smul_57658_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__38_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___83_comb = 9'h000;
  assign p1_smul_57680_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__49_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___88_comb = 9'h000;
  assign p1_concat_135137_comb = {p1_smul_57684_NarrowedMult__comb, p1_smul_57330_TrailingBits___89_comb};
  assign p1_concat_135138_comb = {p1_smul_57686_NarrowedMult__comb, p1_smul_57330_TrailingBits___90_comb};
  assign p1_smul_57690_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__54_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___91_comb = 9'h000;
  assign p1_smul_57696_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__57_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___92_comb = 9'h000;
  assign p1_concat_135143_comb = {p1_smul_57700_NarrowedMult__comb, p1_smul_57330_TrailingBits___93_comb};
  assign p1_concat_135144_comb = {p1_smul_57702_NarrowedMult__comb, p1_smul_57330_TrailingBits___94_comb};
  assign p1_smul_57706_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__62_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___95_comb = 9'h000;
  assign p1_concat_135147_comb = {p1_smul_57838_NarrowedMult__comb, p1_smul_57330_TrailingBits___96_comb};
  assign p1_smul_57842_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__2_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___97_comb = 9'h000;
  assign p1_smul_57848_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__5_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___98_comb = 9'h000;
  assign p1_concat_135152_comb = {p1_smul_57852_NarrowedMult__comb, p1_smul_57330_TrailingBits___99_comb};
  assign p1_concat_135153_comb = {p1_smul_57854_NarrowedMult__comb, p1_smul_57330_TrailingBits___100_comb};
  assign p1_smul_57858_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__10_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___101_comb = 9'h000;
  assign p1_smul_57864_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__13_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___102_comb = 9'h000;
  assign p1_concat_135158_comb = {p1_smul_57868_NarrowedMult__comb, p1_smul_57330_TrailingBits___103_comb};
  assign p1_concat_135159_comb = {p1_smul_57886_NarrowedMult__comb, p1_smul_57330_TrailingBits___108_comb};
  assign p1_smul_57890_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__26_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___109_comb = 9'h000;
  assign p1_smul_57896_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__29_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___110_comb = 9'h000;
  assign p1_concat_135164_comb = {p1_smul_57900_NarrowedMult__comb, p1_smul_57330_TrailingBits___111_comb};
  assign p1_concat_135165_comb = {p1_smul_57902_NarrowedMult__comb, p1_smul_57330_TrailingBits___112_comb};
  assign p1_smul_57906_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__34_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___113_comb = 9'h000;
  assign p1_smul_57912_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__37_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___114_comb = 9'h000;
  assign p1_concat_135170_comb = {p1_smul_57916_NarrowedMult__comb, p1_smul_57330_TrailingBits___115_comb};
  assign p1_concat_135171_comb = {p1_smul_57934_NarrowedMult__comb, p1_smul_57330_TrailingBits___120_comb};
  assign p1_smul_57938_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__50_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___121_comb = 9'h000;
  assign p1_smul_57944_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__53_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___122_comb = 9'h000;
  assign p1_concat_135176_comb = {p1_smul_57948_NarrowedMult__comb, p1_smul_57330_TrailingBits___123_comb};
  assign p1_concat_135177_comb = {p1_smul_57950_NarrowedMult__comb, p1_smul_57330_TrailingBits___124_comb};
  assign p1_smul_57954_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__58_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___125_comb = 9'h000;
  assign p1_smul_57960_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__61_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___126_comb = 9'h000;
  assign p1_concat_135182_comb = {p1_smul_57964_NarrowedMult__comb, p1_smul_57330_TrailingBits___127_comb};
  assign p1_concat_135183_comb = {p1_smul_57966_NarrowedMult__comb, p1_smul_57330_TrailingBits___128_comb};
  assign p1_concat_135184_comb = {p1_smul_57968_NarrowedMult__comb, p1_smul_57454_TrailingBits___32_comb};
  assign p1_concat_135185_comb = {p1_smul_57970_NarrowedMult__comb, p1_smul_57330_TrailingBits___129_comb};
  assign p1_concat_135186_comb = {p1_smul_57972_NarrowedMult__comb, p1_smul_57454_TrailingBits___33_comb};
  assign p1_concat_135187_comb = {p1_smul_57974_NarrowedMult__comb, p1_smul_57454_TrailingBits___34_comb};
  assign p1_concat_135188_comb = {p1_smul_57976_NarrowedMult__comb, p1_smul_57330_TrailingBits___130_comb};
  assign p1_concat_135189_comb = {p1_smul_57978_NarrowedMult__comb, p1_smul_57454_TrailingBits___35_comb};
  assign p1_concat_135190_comb = {p1_smul_57980_NarrowedMult__comb, p1_smul_57330_TrailingBits___131_comb};
  assign p1_concat_135191_comb = {p1_smul_57982_NarrowedMult__comb, p1_smul_57330_TrailingBits___132_comb};
  assign p1_concat_135192_comb = {p1_smul_57984_NarrowedMult__comb, p1_smul_57454_TrailingBits___36_comb};
  assign p1_concat_135193_comb = {p1_smul_57986_NarrowedMult__comb, p1_smul_57330_TrailingBits___133_comb};
  assign p1_concat_135194_comb = {p1_smul_57988_NarrowedMult__comb, p1_smul_57454_TrailingBits___37_comb};
  assign p1_concat_135195_comb = {p1_smul_57990_NarrowedMult__comb, p1_smul_57454_TrailingBits___38_comb};
  assign p1_concat_135196_comb = {p1_smul_57992_NarrowedMult__comb, p1_smul_57330_TrailingBits___134_comb};
  assign p1_concat_135197_comb = {p1_smul_57994_NarrowedMult__comb, p1_smul_57454_TrailingBits___39_comb};
  assign p1_concat_135198_comb = {p1_smul_57996_NarrowedMult__comb, p1_smul_57330_TrailingBits___135_comb};
  assign p1_concat_135199_comb = {p1_smul_58014_NarrowedMult__comb, p1_smul_57330_TrailingBits___140_comb};
  assign p1_concat_135200_comb = {p1_smul_58016_NarrowedMult__comb, p1_smul_57454_TrailingBits___44_comb};
  assign p1_concat_135201_comb = {p1_smul_58018_NarrowedMult__comb, p1_smul_57330_TrailingBits___141_comb};
  assign p1_concat_135202_comb = {p1_smul_58020_NarrowedMult__comb, p1_smul_57454_TrailingBits___45_comb};
  assign p1_concat_135203_comb = {p1_smul_58022_NarrowedMult__comb, p1_smul_57454_TrailingBits___46_comb};
  assign p1_concat_135204_comb = {p1_smul_58024_NarrowedMult__comb, p1_smul_57330_TrailingBits___142_comb};
  assign p1_concat_135205_comb = {p1_smul_58026_NarrowedMult__comb, p1_smul_57454_TrailingBits___47_comb};
  assign p1_concat_135206_comb = {p1_smul_58028_NarrowedMult__comb, p1_smul_57330_TrailingBits___143_comb};
  assign p1_concat_135207_comb = {p1_smul_58030_NarrowedMult__comb, p1_smul_57330_TrailingBits___144_comb};
  assign p1_concat_135208_comb = {p1_smul_58032_NarrowedMult__comb, p1_smul_57454_TrailingBits___48_comb};
  assign p1_concat_135209_comb = {p1_smul_58034_NarrowedMult__comb, p1_smul_57330_TrailingBits___145_comb};
  assign p1_concat_135210_comb = {p1_smul_58036_NarrowedMult__comb, p1_smul_57454_TrailingBits___49_comb};
  assign p1_concat_135211_comb = {p1_smul_58038_NarrowedMult__comb, p1_smul_57454_TrailingBits___50_comb};
  assign p1_concat_135212_comb = {p1_smul_58040_NarrowedMult__comb, p1_smul_57330_TrailingBits___146_comb};
  assign p1_concat_135213_comb = {p1_smul_58042_NarrowedMult__comb, p1_smul_57454_TrailingBits___51_comb};
  assign p1_concat_135214_comb = {p1_smul_58044_NarrowedMult__comb, p1_smul_57330_TrailingBits___147_comb};
  assign p1_concat_135215_comb = {p1_smul_58062_NarrowedMult__comb, p1_smul_57330_TrailingBits___152_comb};
  assign p1_concat_135216_comb = {p1_smul_58064_NarrowedMult__comb, p1_smul_57454_TrailingBits___56_comb};
  assign p1_concat_135217_comb = {p1_smul_58066_NarrowedMult__comb, p1_smul_57330_TrailingBits___153_comb};
  assign p1_concat_135218_comb = {p1_smul_58068_NarrowedMult__comb, p1_smul_57454_TrailingBits___57_comb};
  assign p1_concat_135219_comb = {p1_smul_58070_NarrowedMult__comb, p1_smul_57454_TrailingBits___58_comb};
  assign p1_concat_135220_comb = {p1_smul_58072_NarrowedMult__comb, p1_smul_57330_TrailingBits___154_comb};
  assign p1_concat_135221_comb = {p1_smul_58074_NarrowedMult__comb, p1_smul_57454_TrailingBits___59_comb};
  assign p1_concat_135222_comb = {p1_smul_58076_NarrowedMult__comb, p1_smul_57330_TrailingBits___155_comb};
  assign p1_concat_135223_comb = {p1_smul_58078_NarrowedMult__comb, p1_smul_57330_TrailingBits___156_comb};
  assign p1_concat_135224_comb = {p1_smul_58080_NarrowedMult__comb, p1_smul_57454_TrailingBits___60_comb};
  assign p1_concat_135225_comb = {p1_smul_58082_NarrowedMult__comb, p1_smul_57330_TrailingBits___157_comb};
  assign p1_concat_135226_comb = {p1_smul_58084_NarrowedMult__comb, p1_smul_57454_TrailingBits___61_comb};
  assign p1_concat_135227_comb = {p1_smul_58086_NarrowedMult__comb, p1_smul_57454_TrailingBits___62_comb};
  assign p1_concat_135228_comb = {p1_smul_58088_NarrowedMult__comb, p1_smul_57330_TrailingBits___158_comb};
  assign p1_concat_135229_comb = {p1_smul_58090_NarrowedMult__comb, p1_smul_57454_TrailingBits___63_comb};
  assign p1_concat_135230_comb = {p1_smul_58092_NarrowedMult__comb, p1_smul_57330_TrailingBits___159_comb};
  assign p1_smul_58094_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___160_comb = 9'h000;
  assign p1_concat_135233_comb = {p1_smul_58096_NarrowedMult__comb, p1_smul_57330_TrailingBits___161_comb};
  assign p1_concat_135234_comb = {p1_smul_58106_NarrowedMult__comb, p1_smul_57330_TrailingBits___162_comb};
  assign p1_smul_58108_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__7_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___163_comb = 9'h000;
  assign p1_smul_58110_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__8_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___164_comb = 9'h000;
  assign p1_concat_135239_comb = {p1_smul_58112_NarrowedMult__comb, p1_smul_57330_TrailingBits___165_comb};
  assign p1_concat_135240_comb = {p1_smul_58122_NarrowedMult__comb, p1_smul_57330_TrailingBits___166_comb};
  assign p1_smul_58124_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__15_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___167_comb = 9'h000;
  assign p1_smul_58142_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__24_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___172_comb = 9'h000;
  assign p1_concat_135245_comb = {p1_smul_58144_NarrowedMult__comb, p1_smul_57330_TrailingBits___173_comb};
  assign p1_concat_135246_comb = {p1_smul_58154_NarrowedMult__comb, p1_smul_57330_TrailingBits___174_comb};
  assign p1_smul_58156_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__31_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___175_comb = 9'h000;
  assign p1_smul_58158_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__32_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___176_comb = 9'h000;
  assign p1_concat_135251_comb = {p1_smul_58160_NarrowedMult__comb, p1_smul_57330_TrailingBits___177_comb};
  assign p1_concat_135252_comb = {p1_smul_58170_NarrowedMult__comb, p1_smul_57330_TrailingBits___178_comb};
  assign p1_smul_58172_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__39_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___179_comb = 9'h000;
  assign p1_smul_58190_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__48_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___184_comb = 9'h000;
  assign p1_concat_135257_comb = {p1_smul_58192_NarrowedMult__comb, p1_smul_57330_TrailingBits___185_comb};
  assign p1_concat_135258_comb = {p1_smul_58202_NarrowedMult__comb, p1_smul_57330_TrailingBits___186_comb};
  assign p1_smul_58204_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__55_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___187_comb = 9'h000;
  assign p1_smul_58206_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__56_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___188_comb = 9'h000;
  assign p1_concat_135263_comb = {p1_smul_58208_NarrowedMult__comb, p1_smul_57330_TrailingBits___189_comb};
  assign p1_concat_135264_comb = {p1_smul_58218_NarrowedMult__comb, p1_smul_57330_TrailingBits___190_comb};
  assign p1_smul_58220_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__63_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___191_comb = 9'h000;
  assign p1_smul_57326_TrailingBits___144_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___145_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___146_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___147_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___148_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___149_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___150_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___151_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___168_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___169_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___170_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___171_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___172_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___173_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___174_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___175_comb = 8'h00;
  assign p1_prod__135_comb = {{7{p1_concat_134899_comb[24]}}, p1_concat_134899_comb};
  assign p1_concat_135317_comb = {p1_smul_57364_NarrowedMult__comb, p1_smul_57330_TrailingBits___9_comb};
  assign p1_concat_135318_comb = {p1_smul_57366_NarrowedMult__comb, p1_smul_57330_TrailingBits___10_comb};
  assign p1_prod__150_comb = {{7{p1_concat_134904_comb[24]}}, p1_concat_134904_comb};
  assign p1_prod__327_comb = {{7{p1_concat_134905_comb[24]}}, p1_concat_134905_comb};
  assign p1_concat_135323_comb = {p1_smul_57412_NarrowedMult__comb, p1_smul_57330_TrailingBits___21_comb};
  assign p1_concat_135324_comb = {p1_smul_57414_NarrowedMult__comb, p1_smul_57330_TrailingBits___22_comb};
  assign p1_prod__342_comb = {{7{p1_concat_134910_comb[24]}}, p1_concat_134910_comb};
  assign p1_prod__133_comb = {{7{p1_concat_134911_comb[24]}}, p1_concat_134911_comb};
  assign p1_prod__136_comb = {{8{p1_concat_134912_comb[23]}}, p1_concat_134912_comb};
  assign p1_prod__140_comb = {{8{p1_concat_134913_comb[23]}}, p1_concat_134913_comb};
  assign p1_prod__145_comb = {{7{p1_concat_134914_comb[24]}}, p1_concat_134914_comb};
  assign p1_prod__151_comb = {{7{p1_concat_134915_comb[24]}}, p1_concat_134915_comb};
  assign p1_prod__158_comb = {{8{p1_concat_134916_comb[23]}}, p1_concat_134916_comb};
  assign p1_prod__165_comb = {{8{p1_concat_134917_comb[23]}}, p1_concat_134917_comb};
  assign p1_prod__171_comb = {{7{p1_concat_134918_comb[24]}}, p1_concat_134918_comb};
  assign p1_prod__325_comb = {{7{p1_concat_134919_comb[24]}}, p1_concat_134919_comb};
  assign p1_prod__328_comb = {{8{p1_concat_134920_comb[23]}}, p1_concat_134920_comb};
  assign p1_prod__332_comb = {{8{p1_concat_134921_comb[23]}}, p1_concat_134921_comb};
  assign p1_prod__337_comb = {{7{p1_concat_134922_comb[24]}}, p1_concat_134922_comb};
  assign p1_prod__343_comb = {{7{p1_concat_134923_comb[24]}}, p1_concat_134923_comb};
  assign p1_prod__350_comb = {{8{p1_concat_134924_comb[23]}}, p1_concat_134924_comb};
  assign p1_prod__357_comb = {{8{p1_concat_134925_comb[23]}}, p1_concat_134925_comb};
  assign p1_prod__363_comb = {{7{p1_concat_134926_comb[24]}}, p1_concat_134926_comb};
  assign p1_concat_135351_comb = {p1_smul_57616_NarrowedMult__comb, p1_smul_57330_TrailingBits___72_comb};
  assign p1_prod__152_comb = {{7{p1_concat_134929_comb[24]}}, p1_concat_134929_comb};
  assign p1_prod__159_comb = {{7{p1_concat_134930_comb[24]}}, p1_concat_134930_comb};
  assign p1_concat_135356_comb = {p1_smul_57626_NarrowedMult__comb, p1_smul_57330_TrailingBits___75_comb};
  assign p1_concat_135357_comb = {p1_smul_57664_NarrowedMult__comb, p1_smul_57330_TrailingBits___84_comb};
  assign p1_prod__344_comb = {{7{p1_concat_134935_comb[24]}}, p1_concat_134935_comb};
  assign p1_prod__351_comb = {{7{p1_concat_134936_comb[24]}}, p1_concat_134936_comb};
  assign p1_concat_135362_comb = {p1_smul_57674_NarrowedMult__comb, p1_smul_57330_TrailingBits___87_comb};
  assign p1_prod__148_comb = {{7{p1_concat_134939_comb[24]}}, p1_concat_134939_comb};
  assign p1_concat_135365_comb = {p1_smul_57874_NarrowedMult__comb, p1_smul_57330_TrailingBits___105_comb};
  assign p1_concat_135366_comb = {p1_smul_57880_NarrowedMult__comb, p1_smul_57330_TrailingBits___106_comb};
  assign p1_prod__186_comb = {{7{p1_concat_134944_comb[24]}}, p1_concat_134944_comb};
  assign p1_prod__340_comb = {{7{p1_concat_134945_comb[24]}}, p1_concat_134945_comb};
  assign p1_concat_135371_comb = {p1_smul_57922_NarrowedMult__comb, p1_smul_57330_TrailingBits___117_comb};
  assign p1_concat_135372_comb = {p1_smul_57928_NarrowedMult__comb, p1_smul_57330_TrailingBits___118_comb};
  assign p1_prod__378_comb = {{7{p1_concat_134950_comb[24]}}, p1_concat_134950_comb};
  assign p1_prod__155_comb = {{8{p1_concat_134951_comb[23]}}, p1_concat_134951_comb};
  assign p1_prod__162_comb = {{7{p1_concat_134952_comb[24]}}, p1_concat_134952_comb};
  assign p1_prod__169_comb = {{8{p1_concat_134953_comb[23]}}, p1_concat_134953_comb};
  assign p1_prod__175_comb = {{7{p1_concat_134954_comb[24]}}, p1_concat_134954_comb};
  assign p1_prod__180_comb = {{7{p1_concat_134955_comb[24]}}, p1_concat_134955_comb};
  assign p1_prod__184_comb = {{8{p1_concat_134956_comb[23]}}, p1_concat_134956_comb};
  assign p1_prod__187_comb = {{7{p1_concat_134957_comb[24]}}, p1_concat_134957_comb};
  assign p1_prod__189_comb = {{8{p1_concat_134958_comb[23]}}, p1_concat_134958_comb};
  assign p1_prod__347_comb = {{8{p1_concat_134959_comb[23]}}, p1_concat_134959_comb};
  assign p1_prod__354_comb = {{7{p1_concat_134960_comb[24]}}, p1_concat_134960_comb};
  assign p1_prod__361_comb = {{8{p1_concat_134961_comb[23]}}, p1_concat_134961_comb};
  assign p1_prod__367_comb = {{7{p1_concat_134962_comb[24]}}, p1_concat_134962_comb};
  assign p1_prod__372_comb = {{7{p1_concat_134963_comb[24]}}, p1_concat_134963_comb};
  assign p1_prod__376_comb = {{8{p1_concat_134964_comb[23]}}, p1_concat_134964_comb};
  assign p1_prod__379_comb = {{7{p1_concat_134965_comb[24]}}, p1_concat_134965_comb};
  assign p1_prod__381_comb = {{8{p1_concat_134966_comb[23]}}, p1_concat_134966_comb};
  assign p1_concat_135399_comb = {p1_smul_58126_NarrowedMult__comb, p1_smul_57330_TrailingBits___168_comb};
  assign p1_prod__170_comb = {{7{p1_concat_134969_comb[24]}}, p1_concat_134969_comb};
  assign p1_prod__190_comb = {{7{p1_concat_134970_comb[24]}}, p1_concat_134970_comb};
  assign p1_concat_135404_comb = {p1_smul_58140_NarrowedMult__comb, p1_smul_57330_TrailingBits___171_comb};
  assign p1_concat_135405_comb = {p1_smul_58174_NarrowedMult__comb, p1_smul_57330_TrailingBits___180_comb};
  assign p1_prod__362_comb = {{7{p1_concat_134975_comb[24]}}, p1_concat_134975_comb};
  assign p1_prod__382_comb = {{7{p1_concat_134976_comb[24]}}, p1_concat_134976_comb};
  assign p1_concat_135410_comb = {p1_smul_58188_NarrowedMult__comb, p1_smul_57330_TrailingBits___183_comb};
  assign p1_smul_57326_TrailingBits___128_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___129_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___130_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___131_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___132_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___133_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___134_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___135_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___136_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___137_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___138_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___139_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___140_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___141_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___142_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___143_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___152_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___153_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___154_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___155_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___156_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___157_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___158_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___159_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___160_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___161_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___162_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___163_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___164_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___165_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___166_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___167_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___176_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___177_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___178_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___179_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___180_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___181_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___182_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___183_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___184_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___185_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___186_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___187_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___188_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___189_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___190_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___191_comb = 8'h00;
  assign p1_prod__10_comb = {{7{p1_concat_135027_comb[24]}}, p1_concat_135027_comb};
  assign p1_concat_135557_comb = {p1_smul_57332_NarrowedMult__comb, p1_smul_57330_TrailingBits___1_comb};
  assign p1_concat_135558_comb = {p1_smul_57334_NarrowedMult__comb, p1_smul_57330_TrailingBits___2_comb};
  assign p1_prod__13_comb = {{7{p1_concat_135032_comb[24]}}, p1_concat_135032_comb};
  assign p1_prod__71_comb = {{7{p1_concat_135033_comb[24]}}, p1_concat_135033_comb};
  assign p1_concat_135563_comb = {p1_smul_57348_NarrowedMult__comb, p1_smul_57330_TrailingBits___5_comb};
  assign p1_concat_135564_comb = {p1_smul_57350_NarrowedMult__comb, p1_smul_57330_TrailingBits___6_comb};
  assign p1_prod__86_comb = {{7{p1_concat_135038_comb[24]}}, p1_concat_135038_comb};
  assign p1_prod__199_comb = {{7{p1_concat_135039_comb[24]}}, p1_concat_135039_comb};
  assign p1_concat_135569_comb = {p1_smul_57380_NarrowedMult__comb, p1_smul_57330_TrailingBits___13_comb};
  assign p1_concat_135570_comb = {p1_smul_57382_NarrowedMult__comb, p1_smul_57330_TrailingBits___14_comb};
  assign p1_prod__214_comb = {{7{p1_concat_135044_comb[24]}}, p1_concat_135044_comb};
  assign p1_prod__263_comb = {{7{p1_concat_135045_comb[24]}}, p1_concat_135045_comb};
  assign p1_concat_135575_comb = {p1_smul_57396_NarrowedMult__comb, p1_smul_57330_TrailingBits___17_comb};
  assign p1_concat_135576_comb = {p1_smul_57398_NarrowedMult__comb, p1_smul_57330_TrailingBits___18_comb};
  assign p1_prod__278_comb = {{7{p1_concat_135050_comb[24]}}, p1_concat_135050_comb};
  assign p1_prod__391_comb = {{7{p1_concat_135051_comb[24]}}, p1_concat_135051_comb};
  assign p1_concat_135581_comb = {p1_smul_57428_NarrowedMult__comb, p1_smul_57330_TrailingBits___25_comb};
  assign p1_concat_135582_comb = {p1_smul_57430_NarrowedMult__comb, p1_smul_57330_TrailingBits___26_comb};
  assign p1_prod__406_comb = {{7{p1_concat_135056_comb[24]}}, p1_concat_135056_comb};
  assign p1_prod__455_comb = {{7{p1_concat_135057_comb[24]}}, p1_concat_135057_comb};
  assign p1_concat_135587_comb = {p1_smul_57444_NarrowedMult__comb, p1_smul_57330_TrailingBits___29_comb};
  assign p1_concat_135588_comb = {p1_smul_57446_NarrowedMult__comb, p1_smul_57330_TrailingBits___30_comb};
  assign p1_prod__470_comb = {{7{p1_concat_135062_comb[24]}}, p1_concat_135062_comb};
  assign p1_prod__16_comb = {{7{p1_concat_135063_comb[24]}}, p1_concat_135063_comb};
  assign p1_prod__17_comb = {{8{p1_concat_135064_comb[23]}}, p1_concat_135064_comb};
  assign p1_prod__18_comb = {{8{p1_concat_135065_comb[23]}}, p1_concat_135065_comb};
  assign p1_prod__19_comb = {{7{p1_concat_135066_comb[24]}}, p1_concat_135066_comb};
  assign p1_prod__20_comb = {{7{p1_concat_135067_comb[24]}}, p1_concat_135067_comb};
  assign p1_prod__21_comb = {{8{p1_concat_135068_comb[23]}}, p1_concat_135068_comb};
  assign p1_prod__22_comb = {{8{p1_concat_135069_comb[23]}}, p1_concat_135069_comb};
  assign p1_prod__23_comb = {{7{p1_concat_135070_comb[24]}}, p1_concat_135070_comb};
  assign p1_prod__69_comb = {{7{p1_concat_135071_comb[24]}}, p1_concat_135071_comb};
  assign p1_prod__72_comb = {{8{p1_concat_135072_comb[23]}}, p1_concat_135072_comb};
  assign p1_prod__76_comb = {{8{p1_concat_135073_comb[23]}}, p1_concat_135073_comb};
  assign p1_prod__81_comb = {{7{p1_concat_135074_comb[24]}}, p1_concat_135074_comb};
  assign p1_prod__87_comb = {{7{p1_concat_135075_comb[24]}}, p1_concat_135075_comb};
  assign p1_prod__94_comb = {{8{p1_concat_135076_comb[23]}}, p1_concat_135076_comb};
  assign p1_prod__101_comb = {{8{p1_concat_135077_comb[23]}}, p1_concat_135077_comb};
  assign p1_prod__107_comb = {{7{p1_concat_135078_comb[24]}}, p1_concat_135078_comb};
  assign p1_prod__197_comb = {{7{p1_concat_135079_comb[24]}}, p1_concat_135079_comb};
  assign p1_prod__200_comb = {{8{p1_concat_135080_comb[23]}}, p1_concat_135080_comb};
  assign p1_prod__204_comb = {{8{p1_concat_135081_comb[23]}}, p1_concat_135081_comb};
  assign p1_prod__209_comb = {{7{p1_concat_135082_comb[24]}}, p1_concat_135082_comb};
  assign p1_prod__215_comb = {{7{p1_concat_135083_comb[24]}}, p1_concat_135083_comb};
  assign p1_prod__222_comb = {{8{p1_concat_135084_comb[23]}}, p1_concat_135084_comb};
  assign p1_prod__229_comb = {{8{p1_concat_135085_comb[23]}}, p1_concat_135085_comb};
  assign p1_prod__235_comb = {{7{p1_concat_135086_comb[24]}}, p1_concat_135086_comb};
  assign p1_prod__261_comb = {{7{p1_concat_135087_comb[24]}}, p1_concat_135087_comb};
  assign p1_prod__264_comb = {{8{p1_concat_135088_comb[23]}}, p1_concat_135088_comb};
  assign p1_prod__268_comb = {{8{p1_concat_135089_comb[23]}}, p1_concat_135089_comb};
  assign p1_prod__273_comb = {{7{p1_concat_135090_comb[24]}}, p1_concat_135090_comb};
  assign p1_prod__279_comb = {{7{p1_concat_135091_comb[24]}}, p1_concat_135091_comb};
  assign p1_prod__286_comb = {{8{p1_concat_135092_comb[23]}}, p1_concat_135092_comb};
  assign p1_prod__293_comb = {{8{p1_concat_135093_comb[23]}}, p1_concat_135093_comb};
  assign p1_prod__299_comb = {{7{p1_concat_135094_comb[24]}}, p1_concat_135094_comb};
  assign p1_prod__389_comb = {{7{p1_concat_135095_comb[24]}}, p1_concat_135095_comb};
  assign p1_prod__392_comb = {{8{p1_concat_135096_comb[23]}}, p1_concat_135096_comb};
  assign p1_prod__396_comb = {{8{p1_concat_135097_comb[23]}}, p1_concat_135097_comb};
  assign p1_prod__401_comb = {{7{p1_concat_135098_comb[24]}}, p1_concat_135098_comb};
  assign p1_prod__407_comb = {{7{p1_concat_135099_comb[24]}}, p1_concat_135099_comb};
  assign p1_prod__414_comb = {{8{p1_concat_135100_comb[23]}}, p1_concat_135100_comb};
  assign p1_prod__421_comb = {{8{p1_concat_135101_comb[23]}}, p1_concat_135101_comb};
  assign p1_prod__427_comb = {{7{p1_concat_135102_comb[24]}}, p1_concat_135102_comb};
  assign p1_prod__453_comb = {{7{p1_concat_135103_comb[24]}}, p1_concat_135103_comb};
  assign p1_prod__456_comb = {{8{p1_concat_135104_comb[23]}}, p1_concat_135104_comb};
  assign p1_prod__460_comb = {{8{p1_concat_135105_comb[23]}}, p1_concat_135105_comb};
  assign p1_prod__465_comb = {{7{p1_concat_135106_comb[24]}}, p1_concat_135106_comb};
  assign p1_prod__471_comb = {{7{p1_concat_135107_comb[24]}}, p1_concat_135107_comb};
  assign p1_prod__478_comb = {{8{p1_concat_135108_comb[23]}}, p1_concat_135108_comb};
  assign p1_prod__485_comb = {{8{p1_concat_135109_comb[23]}}, p1_concat_135109_comb};
  assign p1_prod__491_comb = {{7{p1_concat_135110_comb[24]}}, p1_concat_135110_comb};
  assign p1_concat_135663_comb = {p1_smul_57584_NarrowedMult__comb, p1_smul_57330_TrailingBits___64_comb};
  assign p1_prod__27_comb = {{7{p1_concat_135113_comb[24]}}, p1_concat_135113_comb};
  assign p1_prod__28_comb = {{7{p1_concat_135114_comb[24]}}, p1_concat_135114_comb};
  assign p1_concat_135668_comb = {p1_smul_57594_NarrowedMult__comb, p1_smul_57330_TrailingBits___67_comb};
  assign p1_concat_135669_comb = {p1_smul_57600_NarrowedMult__comb, p1_smul_57330_TrailingBits___68_comb};
  assign p1_prod__88_comb = {{7{p1_concat_135119_comb[24]}}, p1_concat_135119_comb};
  assign p1_prod__95_comb = {{7{p1_concat_135120_comb[24]}}, p1_concat_135120_comb};
  assign p1_concat_135674_comb = {p1_smul_57610_NarrowedMult__comb, p1_smul_57330_TrailingBits___71_comb};
  assign p1_concat_135675_comb = {p1_smul_57632_NarrowedMult__comb, p1_smul_57330_TrailingBits___76_comb};
  assign p1_prod__216_comb = {{7{p1_concat_135125_comb[24]}}, p1_concat_135125_comb};
  assign p1_prod__223_comb = {{7{p1_concat_135126_comb[24]}}, p1_concat_135126_comb};
  assign p1_concat_135680_comb = {p1_smul_57642_NarrowedMult__comb, p1_smul_57330_TrailingBits___79_comb};
  assign p1_concat_135681_comb = {p1_smul_57648_NarrowedMult__comb, p1_smul_57330_TrailingBits___80_comb};
  assign p1_prod__280_comb = {{7{p1_concat_135131_comb[24]}}, p1_concat_135131_comb};
  assign p1_prod__287_comb = {{7{p1_concat_135132_comb[24]}}, p1_concat_135132_comb};
  assign p1_concat_135686_comb = {p1_smul_57658_NarrowedMult__comb, p1_smul_57330_TrailingBits___83_comb};
  assign p1_concat_135687_comb = {p1_smul_57680_NarrowedMult__comb, p1_smul_57330_TrailingBits___88_comb};
  assign p1_prod__408_comb = {{7{p1_concat_135137_comb[24]}}, p1_concat_135137_comb};
  assign p1_prod__415_comb = {{7{p1_concat_135138_comb[24]}}, p1_concat_135138_comb};
  assign p1_concat_135692_comb = {p1_smul_57690_NarrowedMult__comb, p1_smul_57330_TrailingBits___91_comb};
  assign p1_concat_135693_comb = {p1_smul_57696_NarrowedMult__comb, p1_smul_57330_TrailingBits___92_comb};
  assign p1_prod__472_comb = {{7{p1_concat_135143_comb[24]}}, p1_concat_135143_comb};
  assign p1_prod__479_comb = {{7{p1_concat_135144_comb[24]}}, p1_concat_135144_comb};
  assign p1_concat_135698_comb = {p1_smul_57706_NarrowedMult__comb, p1_smul_57330_TrailingBits___95_comb};
  assign p1_prod__40_comb = {{7{p1_concat_135147_comb[24]}}, p1_concat_135147_comb};
  assign p1_concat_135701_comb = {p1_smul_57842_NarrowedMult__comb, p1_smul_57330_TrailingBits___97_comb};
  assign p1_concat_135702_comb = {p1_smul_57848_NarrowedMult__comb, p1_smul_57330_TrailingBits___98_comb};
  assign p1_prod__47_comb = {{7{p1_concat_135152_comb[24]}}, p1_concat_135152_comb};
  assign p1_prod__84_comb = {{7{p1_concat_135153_comb[24]}}, p1_concat_135153_comb};
  assign p1_concat_135707_comb = {p1_smul_57858_NarrowedMult__comb, p1_smul_57330_TrailingBits___101_comb};
  assign p1_concat_135708_comb = {p1_smul_57864_NarrowedMult__comb, p1_smul_57330_TrailingBits___102_comb};
  assign p1_prod__122_comb = {{7{p1_concat_135158_comb[24]}}, p1_concat_135158_comb};
  assign p1_prod__212_comb = {{7{p1_concat_135159_comb[24]}}, p1_concat_135159_comb};
  assign p1_concat_135713_comb = {p1_smul_57890_NarrowedMult__comb, p1_smul_57330_TrailingBits___109_comb};
  assign p1_concat_135714_comb = {p1_smul_57896_NarrowedMult__comb, p1_smul_57330_TrailingBits___110_comb};
  assign p1_prod__250_comb = {{7{p1_concat_135164_comb[24]}}, p1_concat_135164_comb};
  assign p1_prod__276_comb = {{7{p1_concat_135165_comb[24]}}, p1_concat_135165_comb};
  assign p1_concat_135719_comb = {p1_smul_57906_NarrowedMult__comb, p1_smul_57330_TrailingBits___113_comb};
  assign p1_concat_135720_comb = {p1_smul_57912_NarrowedMult__comb, p1_smul_57330_TrailingBits___114_comb};
  assign p1_prod__314_comb = {{7{p1_concat_135170_comb[24]}}, p1_concat_135170_comb};
  assign p1_prod__404_comb = {{7{p1_concat_135171_comb[24]}}, p1_concat_135171_comb};
  assign p1_concat_135725_comb = {p1_smul_57938_NarrowedMult__comb, p1_smul_57330_TrailingBits___121_comb};
  assign p1_concat_135726_comb = {p1_smul_57944_NarrowedMult__comb, p1_smul_57330_TrailingBits___122_comb};
  assign p1_prod__442_comb = {{7{p1_concat_135176_comb[24]}}, p1_concat_135176_comb};
  assign p1_prod__468_comb = {{7{p1_concat_135177_comb[24]}}, p1_concat_135177_comb};
  assign p1_concat_135731_comb = {p1_smul_57954_NarrowedMult__comb, p1_smul_57330_TrailingBits___125_comb};
  assign p1_concat_135732_comb = {p1_smul_57960_NarrowedMult__comb, p1_smul_57330_TrailingBits___126_comb};
  assign p1_prod__506_comb = {{7{p1_concat_135182_comb[24]}}, p1_concat_135182_comb};
  assign p1_prod__48_comb = {{8{p1_concat_135183_comb[23]}}, p1_concat_135183_comb};
  assign p1_prod__49_comb = {{7{p1_concat_135184_comb[24]}}, p1_concat_135184_comb};
  assign p1_prod__50_comb = {{8{p1_concat_135185_comb[23]}}, p1_concat_135185_comb};
  assign p1_prod__51_comb = {{7{p1_concat_135186_comb[24]}}, p1_concat_135186_comb};
  assign p1_prod__52_comb = {{7{p1_concat_135187_comb[24]}}, p1_concat_135187_comb};
  assign p1_prod__53_comb = {{8{p1_concat_135188_comb[23]}}, p1_concat_135188_comb};
  assign p1_prod__54_comb = {{7{p1_concat_135189_comb[24]}}, p1_concat_135189_comb};
  assign p1_prod__55_comb = {{8{p1_concat_135190_comb[23]}}, p1_concat_135190_comb};
  assign p1_prod__91_comb = {{8{p1_concat_135191_comb[23]}}, p1_concat_135191_comb};
  assign p1_prod__98_comb = {{7{p1_concat_135192_comb[24]}}, p1_concat_135192_comb};
  assign p1_prod__105_comb = {{8{p1_concat_135193_comb[23]}}, p1_concat_135193_comb};
  assign p1_prod__111_comb = {{7{p1_concat_135194_comb[24]}}, p1_concat_135194_comb};
  assign p1_prod__116_comb = {{7{p1_concat_135195_comb[24]}}, p1_concat_135195_comb};
  assign p1_prod__120_comb = {{8{p1_concat_135196_comb[23]}}, p1_concat_135196_comb};
  assign p1_prod__123_comb = {{7{p1_concat_135197_comb[24]}}, p1_concat_135197_comb};
  assign p1_prod__125_comb = {{8{p1_concat_135198_comb[23]}}, p1_concat_135198_comb};
  assign p1_prod__219_comb = {{8{p1_concat_135199_comb[23]}}, p1_concat_135199_comb};
  assign p1_prod__226_comb = {{7{p1_concat_135200_comb[24]}}, p1_concat_135200_comb};
  assign p1_prod__233_comb = {{8{p1_concat_135201_comb[23]}}, p1_concat_135201_comb};
  assign p1_prod__239_comb = {{7{p1_concat_135202_comb[24]}}, p1_concat_135202_comb};
  assign p1_prod__244_comb = {{7{p1_concat_135203_comb[24]}}, p1_concat_135203_comb};
  assign p1_prod__248_comb = {{8{p1_concat_135204_comb[23]}}, p1_concat_135204_comb};
  assign p1_prod__251_comb = {{7{p1_concat_135205_comb[24]}}, p1_concat_135205_comb};
  assign p1_prod__253_comb = {{8{p1_concat_135206_comb[23]}}, p1_concat_135206_comb};
  assign p1_prod__283_comb = {{8{p1_concat_135207_comb[23]}}, p1_concat_135207_comb};
  assign p1_prod__290_comb = {{7{p1_concat_135208_comb[24]}}, p1_concat_135208_comb};
  assign p1_prod__297_comb = {{8{p1_concat_135209_comb[23]}}, p1_concat_135209_comb};
  assign p1_prod__303_comb = {{7{p1_concat_135210_comb[24]}}, p1_concat_135210_comb};
  assign p1_prod__308_comb = {{7{p1_concat_135211_comb[24]}}, p1_concat_135211_comb};
  assign p1_prod__312_comb = {{8{p1_concat_135212_comb[23]}}, p1_concat_135212_comb};
  assign p1_prod__315_comb = {{7{p1_concat_135213_comb[24]}}, p1_concat_135213_comb};
  assign p1_prod__317_comb = {{8{p1_concat_135214_comb[23]}}, p1_concat_135214_comb};
  assign p1_prod__411_comb = {{8{p1_concat_135215_comb[23]}}, p1_concat_135215_comb};
  assign p1_prod__418_comb = {{7{p1_concat_135216_comb[24]}}, p1_concat_135216_comb};
  assign p1_prod__425_comb = {{8{p1_concat_135217_comb[23]}}, p1_concat_135217_comb};
  assign p1_prod__431_comb = {{7{p1_concat_135218_comb[24]}}, p1_concat_135218_comb};
  assign p1_prod__436_comb = {{7{p1_concat_135219_comb[24]}}, p1_concat_135219_comb};
  assign p1_prod__440_comb = {{8{p1_concat_135220_comb[23]}}, p1_concat_135220_comb};
  assign p1_prod__443_comb = {{7{p1_concat_135221_comb[24]}}, p1_concat_135221_comb};
  assign p1_prod__445_comb = {{8{p1_concat_135222_comb[23]}}, p1_concat_135222_comb};
  assign p1_prod__475_comb = {{8{p1_concat_135223_comb[23]}}, p1_concat_135223_comb};
  assign p1_prod__482_comb = {{7{p1_concat_135224_comb[24]}}, p1_concat_135224_comb};
  assign p1_prod__489_comb = {{8{p1_concat_135225_comb[23]}}, p1_concat_135225_comb};
  assign p1_prod__495_comb = {{7{p1_concat_135226_comb[24]}}, p1_concat_135226_comb};
  assign p1_prod__500_comb = {{7{p1_concat_135227_comb[24]}}, p1_concat_135227_comb};
  assign p1_prod__504_comb = {{8{p1_concat_135228_comb[23]}}, p1_concat_135228_comb};
  assign p1_prod__507_comb = {{7{p1_concat_135229_comb[24]}}, p1_concat_135229_comb};
  assign p1_prod__509_comb = {{8{p1_concat_135230_comb[23]}}, p1_concat_135230_comb};
  assign p1_concat_135807_comb = {p1_smul_58094_NarrowedMult__comb, p1_smul_57330_TrailingBits___160_comb};
  assign p1_prod__57_comb = {{7{p1_concat_135233_comb[24]}}, p1_concat_135233_comb};
  assign p1_prod__62_comb = {{7{p1_concat_135234_comb[24]}}, p1_concat_135234_comb};
  assign p1_concat_135812_comb = {p1_smul_58108_NarrowedMult__comb, p1_smul_57330_TrailingBits___163_comb};
  assign p1_concat_135813_comb = {p1_smul_58110_NarrowedMult__comb, p1_smul_57330_TrailingBits___164_comb};
  assign p1_prod__106_comb = {{7{p1_concat_135239_comb[24]}}, p1_concat_135239_comb};
  assign p1_prod__126_comb = {{7{p1_concat_135240_comb[24]}}, p1_concat_135240_comb};
  assign p1_concat_135818_comb = {p1_smul_58124_NarrowedMult__comb, p1_smul_57330_TrailingBits___167_comb};
  assign p1_concat_135819_comb = {p1_smul_58142_NarrowedMult__comb, p1_smul_57330_TrailingBits___172_comb};
  assign p1_prod__234_comb = {{7{p1_concat_135245_comb[24]}}, p1_concat_135245_comb};
  assign p1_prod__254_comb = {{7{p1_concat_135246_comb[24]}}, p1_concat_135246_comb};
  assign p1_concat_135824_comb = {p1_smul_58156_NarrowedMult__comb, p1_smul_57330_TrailingBits___175_comb};
  assign p1_concat_135825_comb = {p1_smul_58158_NarrowedMult__comb, p1_smul_57330_TrailingBits___176_comb};
  assign p1_prod__298_comb = {{7{p1_concat_135251_comb[24]}}, p1_concat_135251_comb};
  assign p1_prod__318_comb = {{7{p1_concat_135252_comb[24]}}, p1_concat_135252_comb};
  assign p1_concat_135830_comb = {p1_smul_58172_NarrowedMult__comb, p1_smul_57330_TrailingBits___179_comb};
  assign p1_concat_135831_comb = {p1_smul_58190_NarrowedMult__comb, p1_smul_57330_TrailingBits___184_comb};
  assign p1_prod__426_comb = {{7{p1_concat_135257_comb[24]}}, p1_concat_135257_comb};
  assign p1_prod__446_comb = {{7{p1_concat_135258_comb[24]}}, p1_concat_135258_comb};
  assign p1_concat_135836_comb = {p1_smul_58204_NarrowedMult__comb, p1_smul_57330_TrailingBits___187_comb};
  assign p1_concat_135837_comb = {p1_smul_58206_NarrowedMult__comb, p1_smul_57330_TrailingBits___188_comb};
  assign p1_prod__490_comb = {{7{p1_concat_135263_comb[24]}}, p1_concat_135263_comb};
  assign p1_prod__510_comb = {{7{p1_concat_135264_comb[24]}}, p1_concat_135264_comb};
  assign p1_concat_135842_comb = {p1_smul_58220_NarrowedMult__comb, p1_smul_57330_TrailingBits___191_comb};
  assign p1_shifted__16_comb = {~p1_array_index_133927_comb[7], p1_array_index_133927_comb[6:0], p1_smul_57326_TrailingBits___144_comb};
  assign p1_smul_57326_TrailingBits___16_comb = 8'h00;
  assign p1_shifted__17_comb = {~p1_array_index_133928_comb[7], p1_array_index_133928_comb[6:0], p1_smul_57326_TrailingBits___145_comb};
  assign p1_smul_57326_TrailingBits___17_comb = 8'h00;
  assign p1_shifted__18_comb = {~p1_array_index_133923_comb[7], p1_array_index_133923_comb[6:0], p1_smul_57326_TrailingBits___146_comb};
  assign p1_smul_57326_TrailingBits___18_comb = 8'h00;
  assign p1_shifted__19_comb = {~p1_array_index_133929_comb[7], p1_array_index_133929_comb[6:0], p1_smul_57326_TrailingBits___147_comb};
  assign p1_smul_57326_TrailingBits___19_comb = 8'h00;
  assign p1_shifted__20_comb = {~p1_array_index_133930_comb[7], p1_array_index_133930_comb[6:0], p1_smul_57326_TrailingBits___148_comb};
  assign p1_smul_57326_TrailingBits___20_comb = 8'h00;
  assign p1_shifted__21_comb = {~p1_array_index_133924_comb[7], p1_array_index_133924_comb[6:0], p1_smul_57326_TrailingBits___149_comb};
  assign p1_smul_57326_TrailingBits___21_comb = 8'h00;
  assign p1_shifted__22_comb = {~p1_array_index_133931_comb[7], p1_array_index_133931_comb[6:0], p1_smul_57326_TrailingBits___150_comb};
  assign p1_smul_57326_TrailingBits___22_comb = 8'h00;
  assign p1_shifted__23_comb = {~p1_array_index_133932_comb[7], p1_array_index_133932_comb[6:0], p1_smul_57326_TrailingBits___151_comb};
  assign p1_smul_57326_TrailingBits___23_comb = 8'h00;
  assign p1_shifted__40_comb = {~p1_array_index_133933_comb[7], p1_array_index_133933_comb[6:0], p1_smul_57326_TrailingBits___168_comb};
  assign p1_smul_57326_TrailingBits___40_comb = 8'h00;
  assign p1_shifted__41_comb = {~p1_array_index_133934_comb[7], p1_array_index_133934_comb[6:0], p1_smul_57326_TrailingBits___169_comb};
  assign p1_smul_57326_TrailingBits___41_comb = 8'h00;
  assign p1_shifted__42_comb = {~p1_array_index_133925_comb[7], p1_array_index_133925_comb[6:0], p1_smul_57326_TrailingBits___170_comb};
  assign p1_smul_57326_TrailingBits___42_comb = 8'h00;
  assign p1_shifted__43_comb = {~p1_array_index_133935_comb[7], p1_array_index_133935_comb[6:0], p1_smul_57326_TrailingBits___171_comb};
  assign p1_smul_57326_TrailingBits___43_comb = 8'h00;
  assign p1_shifted__44_comb = {~p1_array_index_133936_comb[7], p1_array_index_133936_comb[6:0], p1_smul_57326_TrailingBits___172_comb};
  assign p1_smul_57326_TrailingBits___44_comb = 8'h00;
  assign p1_shifted__45_comb = {~p1_array_index_133926_comb[7], p1_array_index_133926_comb[6:0], p1_smul_57326_TrailingBits___173_comb};
  assign p1_smul_57326_TrailingBits___45_comb = 8'h00;
  assign p1_shifted__46_comb = {~p1_array_index_133937_comb[7], p1_array_index_133937_comb[6:0], p1_smul_57326_TrailingBits___174_comb};
  assign p1_smul_57326_TrailingBits___46_comb = 8'h00;
  assign p1_shifted__47_comb = {~p1_array_index_133938_comb[7], p1_array_index_133938_comb[6:0], p1_smul_57326_TrailingBits___175_comb};
  assign p1_smul_57326_TrailingBits___47_comb = 8'h00;
  assign p1_or_135911_comb = p1_prod__135_comb | 32'h0000_0080;
  assign p1_prod__139_comb = {{9{p1_concat_135317_comb[22]}}, p1_concat_135317_comb};
  assign p1_prod__144_comb = {{9{p1_concat_135318_comb[22]}}, p1_concat_135318_comb};
  assign p1_or_135918_comb = p1_prod__150_comb | 32'h0000_0080;
  assign p1_or_135925_comb = p1_prod__327_comb | 32'h0000_0080;
  assign p1_prod__331_comb = {{9{p1_concat_135323_comb[22]}}, p1_concat_135323_comb};
  assign p1_prod__336_comb = {{9{p1_concat_135324_comb[22]}}, p1_concat_135324_comb};
  assign p1_or_135932_comb = p1_prod__342_comb | 32'h0000_0080;
  assign p1_or_135937_comb = p1_prod__133_comb | 32'h0000_0080;
  assign p1_or_135944_comb = p1_prod__145_comb | 32'h0000_0080;
  assign p1_or_135947_comb = p1_prod__151_comb | 32'h0000_0080;
  assign p1_or_135954_comb = p1_prod__171_comb | 32'h0000_0080;
  assign p1_or_135957_comb = p1_prod__325_comb | 32'h0000_0080;
  assign p1_or_135964_comb = p1_prod__337_comb | 32'h0000_0080;
  assign p1_or_135967_comb = p1_prod__343_comb | 32'h0000_0080;
  assign p1_or_135974_comb = p1_prod__363_comb | 32'h0000_0080;
  assign p1_prod__141_comb = {{9{p1_concat_135351_comb[22]}}, p1_concat_135351_comb};
  assign p1_or_135981_comb = p1_prod__152_comb | 32'h0000_0080;
  assign p1_or_135984_comb = p1_prod__159_comb | 32'h0000_0080;
  assign p1_prod__172_comb = {{9{p1_concat_135356_comb[22]}}, p1_concat_135356_comb};
  assign p1_prod__333_comb = {{9{p1_concat_135357_comb[22]}}, p1_concat_135357_comb};
  assign p1_or_135995_comb = p1_prod__344_comb | 32'h0000_0080;
  assign p1_or_135998_comb = p1_prod__351_comb | 32'h0000_0080;
  assign p1_prod__364_comb = {{9{p1_concat_135362_comb[22]}}, p1_concat_135362_comb};
  assign p1_or_136021_comb = p1_prod__148_comb | 32'h0000_0080;
  assign p1_prod__161_comb = {{9{p1_concat_135365_comb[22]}}, p1_concat_135365_comb};
  assign p1_prod__179_comb = {{9{p1_concat_135366_comb[22]}}, p1_concat_135366_comb};
  assign p1_or_136032_comb = p1_prod__186_comb | 32'h0000_0080;
  assign p1_or_136035_comb = p1_prod__340_comb | 32'h0000_0080;
  assign p1_prod__353_comb = {{9{p1_concat_135371_comb[22]}}, p1_concat_135371_comb};
  assign p1_prod__371_comb = {{9{p1_concat_135372_comb[22]}}, p1_concat_135372_comb};
  assign p1_or_136046_comb = p1_prod__378_comb | 32'h0000_0080;
  assign p1_or_136051_comb = p1_prod__162_comb | 32'h0000_0080;
  assign p1_or_136056_comb = p1_prod__175_comb | 32'h0000_0080;
  assign p1_or_136059_comb = p1_prod__180_comb | 32'h0000_0080;
  assign p1_or_136064_comb = p1_prod__187_comb | 32'h0000_0080;
  assign p1_or_136071_comb = p1_prod__354_comb | 32'h0000_0080;
  assign p1_or_136076_comb = p1_prod__367_comb | 32'h0000_0080;
  assign p1_or_136079_comb = p1_prod__372_comb | 32'h0000_0080;
  assign p1_or_136084_comb = p1_prod__379_comb | 32'h0000_0080;
  assign p1_prod__163_comb = {{9{p1_concat_135399_comb[22]}}, p1_concat_135399_comb};
  assign p1_or_136091_comb = p1_prod__170_comb | 32'h0000_0080;
  assign p1_or_136098_comb = p1_prod__190_comb | 32'h0000_0080;
  assign p1_prod__191_comb = {{9{p1_concat_135404_comb[22]}}, p1_concat_135404_comb};
  assign p1_prod__355_comb = {{9{p1_concat_135405_comb[22]}}, p1_concat_135405_comb};
  assign p1_or_136105_comb = p1_prod__362_comb | 32'h0000_0080;
  assign p1_or_136112_comb = p1_prod__382_comb | 32'h0000_0080;
  assign p1_prod__383_comb = {{9{p1_concat_135410_comb[22]}}, p1_concat_135410_comb};
  assign p1_shifted_comb = {~p1_array_index_133951_comb[7], p1_array_index_133951_comb[6:0], p1_smul_57326_TrailingBits___128_comb};
  assign p1_smul_57326_TrailingBits__comb = 8'h00;
  assign p1_shifted__1_comb = {~p1_array_index_133952_comb[7], p1_array_index_133952_comb[6:0], p1_smul_57326_TrailingBits___129_comb};
  assign p1_smul_57326_TrailingBits___1_comb = 8'h00;
  assign p1_shifted__2_comb = {~p1_array_index_133939_comb[7], p1_array_index_133939_comb[6:0], p1_smul_57326_TrailingBits___130_comb};
  assign p1_smul_57326_TrailingBits___2_comb = 8'h00;
  assign p1_shifted__3_comb = {~p1_array_index_133953_comb[7], p1_array_index_133953_comb[6:0], p1_smul_57326_TrailingBits___131_comb};
  assign p1_smul_57326_TrailingBits___3_comb = 8'h00;
  assign p1_shifted__4_comb = {~p1_array_index_133954_comb[7], p1_array_index_133954_comb[6:0], p1_smul_57326_TrailingBits___132_comb};
  assign p1_smul_57326_TrailingBits___4_comb = 8'h00;
  assign p1_shifted__5_comb = {~p1_array_index_133940_comb[7], p1_array_index_133940_comb[6:0], p1_smul_57326_TrailingBits___133_comb};
  assign p1_smul_57326_TrailingBits___5_comb = 8'h00;
  assign p1_shifted__6_comb = {~p1_array_index_133955_comb[7], p1_array_index_133955_comb[6:0], p1_smul_57326_TrailingBits___134_comb};
  assign p1_smul_57326_TrailingBits___6_comb = 8'h00;
  assign p1_shifted__7_comb = {~p1_array_index_133956_comb[7], p1_array_index_133956_comb[6:0], p1_smul_57326_TrailingBits___135_comb};
  assign p1_smul_57326_TrailingBits___7_comb = 8'h00;
  assign p1_shifted__8_comb = {~p1_array_index_133957_comb[7], p1_array_index_133957_comb[6:0], p1_smul_57326_TrailingBits___136_comb};
  assign p1_smul_57326_TrailingBits___8_comb = 8'h00;
  assign p1_shifted__9_comb = {~p1_array_index_133958_comb[7], p1_array_index_133958_comb[6:0], p1_smul_57326_TrailingBits___137_comb};
  assign p1_smul_57326_TrailingBits___9_comb = 8'h00;
  assign p1_shifted__10_comb = {~p1_array_index_133941_comb[7], p1_array_index_133941_comb[6:0], p1_smul_57326_TrailingBits___138_comb};
  assign p1_smul_57326_TrailingBits___10_comb = 8'h00;
  assign p1_shifted__11_comb = {~p1_array_index_133959_comb[7], p1_array_index_133959_comb[6:0], p1_smul_57326_TrailingBits___139_comb};
  assign p1_smul_57326_TrailingBits___11_comb = 8'h00;
  assign p1_shifted__12_comb = {~p1_array_index_133960_comb[7], p1_array_index_133960_comb[6:0], p1_smul_57326_TrailingBits___140_comb};
  assign p1_smul_57326_TrailingBits___12_comb = 8'h00;
  assign p1_shifted__13_comb = {~p1_array_index_133942_comb[7], p1_array_index_133942_comb[6:0], p1_smul_57326_TrailingBits___141_comb};
  assign p1_smul_57326_TrailingBits___13_comb = 8'h00;
  assign p1_shifted__14_comb = {~p1_array_index_133961_comb[7], p1_array_index_133961_comb[6:0], p1_smul_57326_TrailingBits___142_comb};
  assign p1_smul_57326_TrailingBits___14_comb = 8'h00;
  assign p1_shifted__15_comb = {~p1_array_index_133962_comb[7], p1_array_index_133962_comb[6:0], p1_smul_57326_TrailingBits___143_comb};
  assign p1_smul_57326_TrailingBits___15_comb = 8'h00;
  assign p1_shifted__24_comb = {~p1_array_index_133963_comb[7], p1_array_index_133963_comb[6:0], p1_smul_57326_TrailingBits___152_comb};
  assign p1_smul_57326_TrailingBits___24_comb = 8'h00;
  assign p1_shifted__25_comb = {~p1_array_index_133964_comb[7], p1_array_index_133964_comb[6:0], p1_smul_57326_TrailingBits___153_comb};
  assign p1_smul_57326_TrailingBits___25_comb = 8'h00;
  assign p1_shifted__26_comb = {~p1_array_index_133943_comb[7], p1_array_index_133943_comb[6:0], p1_smul_57326_TrailingBits___154_comb};
  assign p1_smul_57326_TrailingBits___26_comb = 8'h00;
  assign p1_shifted__27_comb = {~p1_array_index_133965_comb[7], p1_array_index_133965_comb[6:0], p1_smul_57326_TrailingBits___155_comb};
  assign p1_smul_57326_TrailingBits___27_comb = 8'h00;
  assign p1_shifted__28_comb = {~p1_array_index_133966_comb[7], p1_array_index_133966_comb[6:0], p1_smul_57326_TrailingBits___156_comb};
  assign p1_smul_57326_TrailingBits___28_comb = 8'h00;
  assign p1_shifted__29_comb = {~p1_array_index_133944_comb[7], p1_array_index_133944_comb[6:0], p1_smul_57326_TrailingBits___157_comb};
  assign p1_smul_57326_TrailingBits___29_comb = 8'h00;
  assign p1_shifted__30_comb = {~p1_array_index_133967_comb[7], p1_array_index_133967_comb[6:0], p1_smul_57326_TrailingBits___158_comb};
  assign p1_smul_57326_TrailingBits___30_comb = 8'h00;
  assign p1_shifted__31_comb = {~p1_array_index_133968_comb[7], p1_array_index_133968_comb[6:0], p1_smul_57326_TrailingBits___159_comb};
  assign p1_smul_57326_TrailingBits___31_comb = 8'h00;
  assign p1_shifted__32_comb = {~p1_array_index_133969_comb[7], p1_array_index_133969_comb[6:0], p1_smul_57326_TrailingBits___160_comb};
  assign p1_smul_57326_TrailingBits___32_comb = 8'h00;
  assign p1_shifted__33_comb = {~p1_array_index_133970_comb[7], p1_array_index_133970_comb[6:0], p1_smul_57326_TrailingBits___161_comb};
  assign p1_smul_57326_TrailingBits___33_comb = 8'h00;
  assign p1_shifted__34_comb = {~p1_array_index_133945_comb[7], p1_array_index_133945_comb[6:0], p1_smul_57326_TrailingBits___162_comb};
  assign p1_smul_57326_TrailingBits___34_comb = 8'h00;
  assign p1_shifted__35_comb = {~p1_array_index_133971_comb[7], p1_array_index_133971_comb[6:0], p1_smul_57326_TrailingBits___163_comb};
  assign p1_smul_57326_TrailingBits___35_comb = 8'h00;
  assign p1_shifted__36_comb = {~p1_array_index_133972_comb[7], p1_array_index_133972_comb[6:0], p1_smul_57326_TrailingBits___164_comb};
  assign p1_smul_57326_TrailingBits___36_comb = 8'h00;
  assign p1_shifted__37_comb = {~p1_array_index_133946_comb[7], p1_array_index_133946_comb[6:0], p1_smul_57326_TrailingBits___165_comb};
  assign p1_smul_57326_TrailingBits___37_comb = 8'h00;
  assign p1_shifted__38_comb = {~p1_array_index_133973_comb[7], p1_array_index_133973_comb[6:0], p1_smul_57326_TrailingBits___166_comb};
  assign p1_smul_57326_TrailingBits___38_comb = 8'h00;
  assign p1_shifted__39_comb = {~p1_array_index_133974_comb[7], p1_array_index_133974_comb[6:0], p1_smul_57326_TrailingBits___167_comb};
  assign p1_smul_57326_TrailingBits___39_comb = 8'h00;
  assign p1_shifted__48_comb = {~p1_array_index_133975_comb[7], p1_array_index_133975_comb[6:0], p1_smul_57326_TrailingBits___176_comb};
  assign p1_smul_57326_TrailingBits___48_comb = 8'h00;
  assign p1_shifted__49_comb = {~p1_array_index_133976_comb[7], p1_array_index_133976_comb[6:0], p1_smul_57326_TrailingBits___177_comb};
  assign p1_smul_57326_TrailingBits___49_comb = 8'h00;
  assign p1_shifted__50_comb = {~p1_array_index_133947_comb[7], p1_array_index_133947_comb[6:0], p1_smul_57326_TrailingBits___178_comb};
  assign p1_smul_57326_TrailingBits___50_comb = 8'h00;
  assign p1_shifted__51_comb = {~p1_array_index_133977_comb[7], p1_array_index_133977_comb[6:0], p1_smul_57326_TrailingBits___179_comb};
  assign p1_smul_57326_TrailingBits___51_comb = 8'h00;
  assign p1_shifted__52_comb = {~p1_array_index_133978_comb[7], p1_array_index_133978_comb[6:0], p1_smul_57326_TrailingBits___180_comb};
  assign p1_smul_57326_TrailingBits___52_comb = 8'h00;
  assign p1_shifted__53_comb = {~p1_array_index_133948_comb[7], p1_array_index_133948_comb[6:0], p1_smul_57326_TrailingBits___181_comb};
  assign p1_smul_57326_TrailingBits___53_comb = 8'h00;
  assign p1_shifted__54_comb = {~p1_array_index_133979_comb[7], p1_array_index_133979_comb[6:0], p1_smul_57326_TrailingBits___182_comb};
  assign p1_smul_57326_TrailingBits___54_comb = 8'h00;
  assign p1_shifted__55_comb = {~p1_array_index_133980_comb[7], p1_array_index_133980_comb[6:0], p1_smul_57326_TrailingBits___183_comb};
  assign p1_smul_57326_TrailingBits___55_comb = 8'h00;
  assign p1_shifted__56_comb = {~p1_array_index_133981_comb[7], p1_array_index_133981_comb[6:0], p1_smul_57326_TrailingBits___184_comb};
  assign p1_smul_57326_TrailingBits___56_comb = 8'h00;
  assign p1_shifted__57_comb = {~p1_array_index_133982_comb[7], p1_array_index_133982_comb[6:0], p1_smul_57326_TrailingBits___185_comb};
  assign p1_smul_57326_TrailingBits___57_comb = 8'h00;
  assign p1_shifted__58_comb = {~p1_array_index_133949_comb[7], p1_array_index_133949_comb[6:0], p1_smul_57326_TrailingBits___186_comb};
  assign p1_smul_57326_TrailingBits___58_comb = 8'h00;
  assign p1_shifted__59_comb = {~p1_array_index_133983_comb[7], p1_array_index_133983_comb[6:0], p1_smul_57326_TrailingBits___187_comb};
  assign p1_smul_57326_TrailingBits___59_comb = 8'h00;
  assign p1_shifted__60_comb = {~p1_array_index_133984_comb[7], p1_array_index_133984_comb[6:0], p1_smul_57326_TrailingBits___188_comb};
  assign p1_smul_57326_TrailingBits___60_comb = 8'h00;
  assign p1_shifted__61_comb = {~p1_array_index_133950_comb[7], p1_array_index_133950_comb[6:0], p1_smul_57326_TrailingBits___189_comb};
  assign p1_smul_57326_TrailingBits___61_comb = 8'h00;
  assign p1_shifted__62_comb = {~p1_array_index_133985_comb[7], p1_array_index_133985_comb[6:0], p1_smul_57326_TrailingBits___190_comb};
  assign p1_smul_57326_TrailingBits___62_comb = 8'h00;
  assign p1_shifted__63_comb = {~p1_array_index_133986_comb[7], p1_array_index_133986_comb[6:0], p1_smul_57326_TrailingBits___191_comb};
  assign p1_smul_57326_TrailingBits___63_comb = 8'h00;
  assign p1_or_136311_comb = p1_prod__10_comb | 32'h0000_0080;
  assign p1_prod__11_comb = {{9{p1_concat_135557_comb[22]}}, p1_concat_135557_comb};
  assign p1_prod__12_comb = {{9{p1_concat_135558_comb[22]}}, p1_concat_135558_comb};
  assign p1_or_136318_comb = p1_prod__13_comb | 32'h0000_0080;
  assign p1_or_136325_comb = p1_prod__71_comb | 32'h0000_0080;
  assign p1_prod__75_comb = {{9{p1_concat_135563_comb[22]}}, p1_concat_135563_comb};
  assign p1_prod__80_comb = {{9{p1_concat_135564_comb[22]}}, p1_concat_135564_comb};
  assign p1_or_136332_comb = p1_prod__86_comb | 32'h0000_0080;
  assign p1_or_136339_comb = p1_prod__199_comb | 32'h0000_0080;
  assign p1_prod__203_comb = {{9{p1_concat_135569_comb[22]}}, p1_concat_135569_comb};
  assign p1_prod__208_comb = {{9{p1_concat_135570_comb[22]}}, p1_concat_135570_comb};
  assign p1_or_136346_comb = p1_prod__214_comb | 32'h0000_0080;
  assign p1_or_136353_comb = p1_prod__263_comb | 32'h0000_0080;
  assign p1_prod__267_comb = {{9{p1_concat_135575_comb[22]}}, p1_concat_135575_comb};
  assign p1_prod__272_comb = {{9{p1_concat_135576_comb[22]}}, p1_concat_135576_comb};
  assign p1_or_136360_comb = p1_prod__278_comb | 32'h0000_0080;
  assign p1_or_136367_comb = p1_prod__391_comb | 32'h0000_0080;
  assign p1_prod__395_comb = {{9{p1_concat_135581_comb[22]}}, p1_concat_135581_comb};
  assign p1_prod__400_comb = {{9{p1_concat_135582_comb[22]}}, p1_concat_135582_comb};
  assign p1_or_136374_comb = p1_prod__406_comb | 32'h0000_0080;
  assign p1_or_136381_comb = p1_prod__455_comb | 32'h0000_0080;
  assign p1_prod__459_comb = {{9{p1_concat_135587_comb[22]}}, p1_concat_135587_comb};
  assign p1_prod__464_comb = {{9{p1_concat_135588_comb[22]}}, p1_concat_135588_comb};
  assign p1_or_136388_comb = p1_prod__470_comb | 32'h0000_0080;
  assign p1_or_136393_comb = p1_prod__16_comb | 32'h0000_0080;
  assign p1_or_136400_comb = p1_prod__19_comb | 32'h0000_0080;
  assign p1_or_136403_comb = p1_prod__20_comb | 32'h0000_0080;
  assign p1_or_136410_comb = p1_prod__23_comb | 32'h0000_0080;
  assign p1_or_136413_comb = p1_prod__69_comb | 32'h0000_0080;
  assign p1_or_136420_comb = p1_prod__81_comb | 32'h0000_0080;
  assign p1_or_136423_comb = p1_prod__87_comb | 32'h0000_0080;
  assign p1_or_136430_comb = p1_prod__107_comb | 32'h0000_0080;
  assign p1_or_136433_comb = p1_prod__197_comb | 32'h0000_0080;
  assign p1_or_136440_comb = p1_prod__209_comb | 32'h0000_0080;
  assign p1_or_136443_comb = p1_prod__215_comb | 32'h0000_0080;
  assign p1_or_136450_comb = p1_prod__235_comb | 32'h0000_0080;
  assign p1_or_136453_comb = p1_prod__261_comb | 32'h0000_0080;
  assign p1_or_136460_comb = p1_prod__273_comb | 32'h0000_0080;
  assign p1_or_136463_comb = p1_prod__279_comb | 32'h0000_0080;
  assign p1_or_136470_comb = p1_prod__299_comb | 32'h0000_0080;
  assign p1_or_136473_comb = p1_prod__389_comb | 32'h0000_0080;
  assign p1_or_136480_comb = p1_prod__401_comb | 32'h0000_0080;
  assign p1_or_136483_comb = p1_prod__407_comb | 32'h0000_0080;
  assign p1_or_136490_comb = p1_prod__427_comb | 32'h0000_0080;
  assign p1_or_136493_comb = p1_prod__453_comb | 32'h0000_0080;
  assign p1_or_136500_comb = p1_prod__465_comb | 32'h0000_0080;
  assign p1_or_136503_comb = p1_prod__471_comb | 32'h0000_0080;
  assign p1_or_136510_comb = p1_prod__491_comb | 32'h0000_0080;
  assign p1_prod__25_comb = {{9{p1_concat_135663_comb[22]}}, p1_concat_135663_comb};
  assign p1_or_136517_comb = p1_prod__27_comb | 32'h0000_0080;
  assign p1_or_136520_comb = p1_prod__28_comb | 32'h0000_0080;
  assign p1_prod__30_comb = {{9{p1_concat_135668_comb[22]}}, p1_concat_135668_comb};
  assign p1_prod__77_comb = {{9{p1_concat_135669_comb[22]}}, p1_concat_135669_comb};
  assign p1_or_136531_comb = p1_prod__88_comb | 32'h0000_0080;
  assign p1_or_136534_comb = p1_prod__95_comb | 32'h0000_0080;
  assign p1_prod__108_comb = {{9{p1_concat_135674_comb[22]}}, p1_concat_135674_comb};
  assign p1_prod__205_comb = {{9{p1_concat_135675_comb[22]}}, p1_concat_135675_comb};
  assign p1_or_136545_comb = p1_prod__216_comb | 32'h0000_0080;
  assign p1_or_136548_comb = p1_prod__223_comb | 32'h0000_0080;
  assign p1_prod__236_comb = {{9{p1_concat_135680_comb[22]}}, p1_concat_135680_comb};
  assign p1_prod__269_comb = {{9{p1_concat_135681_comb[22]}}, p1_concat_135681_comb};
  assign p1_or_136559_comb = p1_prod__280_comb | 32'h0000_0080;
  assign p1_or_136562_comb = p1_prod__287_comb | 32'h0000_0080;
  assign p1_prod__300_comb = {{9{p1_concat_135686_comb[22]}}, p1_concat_135686_comb};
  assign p1_prod__397_comb = {{9{p1_concat_135687_comb[22]}}, p1_concat_135687_comb};
  assign p1_or_136573_comb = p1_prod__408_comb | 32'h0000_0080;
  assign p1_or_136576_comb = p1_prod__415_comb | 32'h0000_0080;
  assign p1_prod__428_comb = {{9{p1_concat_135692_comb[22]}}, p1_concat_135692_comb};
  assign p1_prod__461_comb = {{9{p1_concat_135693_comb[22]}}, p1_concat_135693_comb};
  assign p1_or_136587_comb = p1_prod__472_comb | 32'h0000_0080;
  assign p1_or_136590_comb = p1_prod__479_comb | 32'h0000_0080;
  assign p1_prod__492_comb = {{9{p1_concat_135698_comb[22]}}, p1_concat_135698_comb};
  assign p1_or_136645_comb = p1_prod__40_comb | 32'h0000_0080;
  assign p1_prod__42_comb = {{9{p1_concat_135701_comb[22]}}, p1_concat_135701_comb};
  assign p1_prod__45_comb = {{9{p1_concat_135702_comb[22]}}, p1_concat_135702_comb};
  assign p1_or_136656_comb = p1_prod__47_comb | 32'h0000_0080;
  assign p1_or_136659_comb = p1_prod__84_comb | 32'h0000_0080;
  assign p1_prod__97_comb = {{9{p1_concat_135707_comb[22]}}, p1_concat_135707_comb};
  assign p1_prod__115_comb = {{9{p1_concat_135708_comb[22]}}, p1_concat_135708_comb};
  assign p1_or_136670_comb = p1_prod__122_comb | 32'h0000_0080;
  assign p1_or_136673_comb = p1_prod__212_comb | 32'h0000_0080;
  assign p1_prod__225_comb = {{9{p1_concat_135713_comb[22]}}, p1_concat_135713_comb};
  assign p1_prod__243_comb = {{9{p1_concat_135714_comb[22]}}, p1_concat_135714_comb};
  assign p1_or_136684_comb = p1_prod__250_comb | 32'h0000_0080;
  assign p1_or_136687_comb = p1_prod__276_comb | 32'h0000_0080;
  assign p1_prod__289_comb = {{9{p1_concat_135719_comb[22]}}, p1_concat_135719_comb};
  assign p1_prod__307_comb = {{9{p1_concat_135720_comb[22]}}, p1_concat_135720_comb};
  assign p1_or_136698_comb = p1_prod__314_comb | 32'h0000_0080;
  assign p1_or_136701_comb = p1_prod__404_comb | 32'h0000_0080;
  assign p1_prod__417_comb = {{9{p1_concat_135725_comb[22]}}, p1_concat_135725_comb};
  assign p1_prod__435_comb = {{9{p1_concat_135726_comb[22]}}, p1_concat_135726_comb};
  assign p1_or_136712_comb = p1_prod__442_comb | 32'h0000_0080;
  assign p1_or_136715_comb = p1_prod__468_comb | 32'h0000_0080;
  assign p1_prod__481_comb = {{9{p1_concat_135731_comb[22]}}, p1_concat_135731_comb};
  assign p1_prod__499_comb = {{9{p1_concat_135732_comb[22]}}, p1_concat_135732_comb};
  assign p1_or_136726_comb = p1_prod__506_comb | 32'h0000_0080;
  assign p1_or_136731_comb = p1_prod__49_comb | 32'h0000_0080;
  assign p1_or_136736_comb = p1_prod__51_comb | 32'h0000_0080;
  assign p1_or_136739_comb = p1_prod__52_comb | 32'h0000_0080;
  assign p1_or_136744_comb = p1_prod__54_comb | 32'h0000_0080;
  assign p1_or_136751_comb = p1_prod__98_comb | 32'h0000_0080;
  assign p1_or_136756_comb = p1_prod__111_comb | 32'h0000_0080;
  assign p1_or_136759_comb = p1_prod__116_comb | 32'h0000_0080;
  assign p1_or_136764_comb = p1_prod__123_comb | 32'h0000_0080;
  assign p1_or_136771_comb = p1_prod__226_comb | 32'h0000_0080;
  assign p1_or_136776_comb = p1_prod__239_comb | 32'h0000_0080;
  assign p1_or_136779_comb = p1_prod__244_comb | 32'h0000_0080;
  assign p1_or_136784_comb = p1_prod__251_comb | 32'h0000_0080;
  assign p1_or_136791_comb = p1_prod__290_comb | 32'h0000_0080;
  assign p1_or_136796_comb = p1_prod__303_comb | 32'h0000_0080;
  assign p1_or_136799_comb = p1_prod__308_comb | 32'h0000_0080;
  assign p1_or_136804_comb = p1_prod__315_comb | 32'h0000_0080;
  assign p1_or_136811_comb = p1_prod__418_comb | 32'h0000_0080;
  assign p1_or_136816_comb = p1_prod__431_comb | 32'h0000_0080;
  assign p1_or_136819_comb = p1_prod__436_comb | 32'h0000_0080;
  assign p1_or_136824_comb = p1_prod__443_comb | 32'h0000_0080;
  assign p1_or_136831_comb = p1_prod__482_comb | 32'h0000_0080;
  assign p1_or_136836_comb = p1_prod__495_comb | 32'h0000_0080;
  assign p1_or_136839_comb = p1_prod__500_comb | 32'h0000_0080;
  assign p1_or_136844_comb = p1_prod__507_comb | 32'h0000_0080;
  assign p1_prod__56_comb = {{9{p1_concat_135807_comb[22]}}, p1_concat_135807_comb};
  assign p1_or_136851_comb = p1_prod__57_comb | 32'h0000_0080;
  assign p1_or_136858_comb = p1_prod__62_comb | 32'h0000_0080;
  assign p1_prod__63_comb = {{9{p1_concat_135812_comb[22]}}, p1_concat_135812_comb};
  assign p1_prod__99_comb = {{9{p1_concat_135813_comb[22]}}, p1_concat_135813_comb};
  assign p1_or_136865_comb = p1_prod__106_comb | 32'h0000_0080;
  assign p1_or_136872_comb = p1_prod__126_comb | 32'h0000_0080;
  assign p1_prod__127_comb = {{9{p1_concat_135818_comb[22]}}, p1_concat_135818_comb};
  assign p1_prod__227_comb = {{9{p1_concat_135819_comb[22]}}, p1_concat_135819_comb};
  assign p1_or_136879_comb = p1_prod__234_comb | 32'h0000_0080;
  assign p1_or_136886_comb = p1_prod__254_comb | 32'h0000_0080;
  assign p1_prod__255_comb = {{9{p1_concat_135824_comb[22]}}, p1_concat_135824_comb};
  assign p1_prod__291_comb = {{9{p1_concat_135825_comb[22]}}, p1_concat_135825_comb};
  assign p1_or_136893_comb = p1_prod__298_comb | 32'h0000_0080;
  assign p1_or_136900_comb = p1_prod__318_comb | 32'h0000_0080;
  assign p1_prod__319_comb = {{9{p1_concat_135830_comb[22]}}, p1_concat_135830_comb};
  assign p1_prod__419_comb = {{9{p1_concat_135831_comb[22]}}, p1_concat_135831_comb};
  assign p1_or_136907_comb = p1_prod__426_comb | 32'h0000_0080;
  assign p1_or_136914_comb = p1_prod__446_comb | 32'h0000_0080;
  assign p1_prod__447_comb = {{9{p1_concat_135836_comb[22]}}, p1_concat_135836_comb};
  assign p1_prod__483_comb = {{9{p1_concat_135837_comb[22]}}, p1_concat_135837_comb};
  assign p1_or_136921_comb = p1_prod__490_comb | 32'h0000_0080;
  assign p1_or_136928_comb = p1_prod__510_comb | 32'h0000_0080;
  assign p1_prod__511_comb = {{9{p1_concat_135842_comb[22]}}, p1_concat_135842_comb};
  assign p1_smul_57358_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__16_squeezed_comb, 9'h0fb);
  assign p1_smul_57360_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__17_squeezed_comb, 9'h0d5);
  assign p1_or_136986_comb = p1_prod__139_comb | 32'h0000_0080;
  assign p1_or_136987_comb = p1_prod__144_comb | 32'h0000_0080;
  assign p1_smul_57370_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__22_squeezed_comb, 9'h12b);
  assign p1_smul_57372_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__23_squeezed_comb, 9'h105);
  assign p1_smul_57406_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__40_squeezed_comb, 9'h0fb);
  assign p1_smul_57408_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__41_squeezed_comb, 9'h0d5);
  assign p1_or_137002_comb = p1_prod__331_comb | 32'h0000_0080;
  assign p1_or_137003_comb = p1_prod__336_comb | 32'h0000_0080;
  assign p1_smul_57418_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__46_squeezed_comb, 9'h12b);
  assign p1_smul_57420_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__47_squeezed_comb, 9'h105);
  assign p1_smul_57614_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__16_squeezed_comb, 9'h0d5);
  assign p1_or_137053_comb = p1_prod__141_comb | 32'h0000_0080;
  assign p1_smul_57618_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__18_squeezed_comb, 9'h105);
  assign p1_smul_57624_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__21_squeezed_comb, 9'h0fb);
  assign p1_or_137064_comb = p1_prod__172_comb | 32'h0000_0080;
  assign p1_smul_57628_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__23_squeezed_comb, 9'h12b);
  assign p1_smul_57662_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__40_squeezed_comb, 9'h0d5);
  assign p1_or_137069_comb = p1_prod__333_comb | 32'h0000_0080;
  assign p1_smul_57666_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__42_squeezed_comb, 9'h105);
  assign p1_smul_57672_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__45_squeezed_comb, 9'h0fb);
  assign p1_or_137080_comb = p1_prod__364_comb | 32'h0000_0080;
  assign p1_smul_57676_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__47_squeezed_comb, 9'h12b);
  assign p1_smul_57742_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__16_squeezed_comb, 9'h0b5);
  assign p1_smul_57744_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__17_squeezed_comb, 9'h14b);
  assign p1_smul_57746_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__18_squeezed_comb, 9'h14b);
  assign p1_smul_57748_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__19_squeezed_comb, 9'h0b5);
  assign p1_smul_57750_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__20_squeezed_comb, 9'h0b5);
  assign p1_smul_57752_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__21_squeezed_comb, 9'h14b);
  assign p1_smul_57754_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__22_squeezed_comb, 9'h14b);
  assign p1_smul_57756_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__23_squeezed_comb, 9'h0b5);
  assign p1_smul_57790_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__40_squeezed_comb, 9'h0b5);
  assign p1_smul_57792_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__41_squeezed_comb, 9'h14b);
  assign p1_smul_57794_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__42_squeezed_comb, 9'h14b);
  assign p1_smul_57796_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__43_squeezed_comb, 9'h0b5);
  assign p1_smul_57798_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__44_squeezed_comb, 9'h0b5);
  assign p1_smul_57800_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__45_squeezed_comb, 9'h14b);
  assign p1_smul_57802_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__46_squeezed_comb, 9'h14b);
  assign p1_smul_57804_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__47_squeezed_comb, 9'h0b5);
  assign p1_smul_57872_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__17_squeezed_comb, 9'h105);
  assign p1_or_137120_comb = p1_prod__161_comb | 32'h0000_0080;
  assign p1_smul_57876_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__19_squeezed_comb, 9'h0d5);
  assign p1_smul_57878_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__20_squeezed_comb, 9'h0d5);
  assign p1_or_137125_comb = p1_prod__179_comb | 32'h0000_0080;
  assign p1_smul_57882_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__22_squeezed_comb, 9'h105);
  assign p1_smul_57920_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__41_squeezed_comb, 9'h105);
  assign p1_or_137136_comb = p1_prod__353_comb | 32'h0000_0080;
  assign p1_smul_57924_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__43_squeezed_comb, 9'h0d5);
  assign p1_smul_57926_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__44_squeezed_comb, 9'h0d5);
  assign p1_or_137141_comb = p1_prod__371_comb | 32'h0000_0080;
  assign p1_smul_57930_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__46_squeezed_comb, 9'h105);
  assign p1_or_137187_comb = p1_prod__163_comb | 32'h0000_0080;
  assign p1_smul_58130_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__18_squeezed_comb, 9'h0d5);
  assign p1_smul_58132_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__19_squeezed_comb, 9'h105);
  assign p1_smul_58134_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__20_squeezed_comb, 9'h105);
  assign p1_smul_58136_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__21_squeezed_comb, 9'h0d5);
  assign p1_or_137202_comb = p1_prod__191_comb | 32'h0000_0080;
  assign p1_or_137203_comb = p1_prod__355_comb | 32'h0000_0080;
  assign p1_smul_58178_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__42_squeezed_comb, 9'h0d5);
  assign p1_smul_58180_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__43_squeezed_comb, 9'h105);
  assign p1_smul_58182_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__44_squeezed_comb, 9'h105);
  assign p1_smul_58184_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__45_squeezed_comb, 9'h0d5);
  assign p1_or_137218_comb = p1_prod__383_comb | 32'h0000_0080;
  assign p1_smul_57326_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted_squeezed_comb, 9'h0fb);
  assign p1_smul_57328_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__1_squeezed_comb, 9'h0d5);
  assign p1_or_137370_comb = p1_prod__11_comb | 32'h0000_0080;
  assign p1_or_137371_comb = p1_prod__12_comb | 32'h0000_0080;
  assign p1_smul_57338_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__6_squeezed_comb, 9'h12b);
  assign p1_smul_57340_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__7_squeezed_comb, 9'h105);
  assign p1_smul_57342_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__8_squeezed_comb, 9'h0fb);
  assign p1_smul_57344_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__9_squeezed_comb, 9'h0d5);
  assign p1_or_137386_comb = p1_prod__75_comb | 32'h0000_0080;
  assign p1_or_137387_comb = p1_prod__80_comb | 32'h0000_0080;
  assign p1_smul_57354_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__14_squeezed_comb, 9'h12b);
  assign p1_smul_57356_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__15_squeezed_comb, 9'h105);
  assign p1_smul_57374_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__24_squeezed_comb, 9'h0fb);
  assign p1_smul_57376_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__25_squeezed_comb, 9'h0d5);
  assign p1_or_137402_comb = p1_prod__203_comb | 32'h0000_0080;
  assign p1_or_137403_comb = p1_prod__208_comb | 32'h0000_0080;
  assign p1_smul_57386_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__30_squeezed_comb, 9'h12b);
  assign p1_smul_57388_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__31_squeezed_comb, 9'h105);
  assign p1_smul_57390_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__32_squeezed_comb, 9'h0fb);
  assign p1_smul_57392_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__33_squeezed_comb, 9'h0d5);
  assign p1_or_137418_comb = p1_prod__267_comb | 32'h0000_0080;
  assign p1_or_137419_comb = p1_prod__272_comb | 32'h0000_0080;
  assign p1_smul_57402_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__38_squeezed_comb, 9'h12b);
  assign p1_smul_57404_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__39_squeezed_comb, 9'h105);
  assign p1_smul_57422_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__48_squeezed_comb, 9'h0fb);
  assign p1_smul_57424_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__49_squeezed_comb, 9'h0d5);
  assign p1_or_137434_comb = p1_prod__395_comb | 32'h0000_0080;
  assign p1_or_137435_comb = p1_prod__400_comb | 32'h0000_0080;
  assign p1_smul_57434_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__54_squeezed_comb, 9'h12b);
  assign p1_smul_57436_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__55_squeezed_comb, 9'h105);
  assign p1_smul_57438_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__56_squeezed_comb, 9'h0fb);
  assign p1_smul_57440_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__57_squeezed_comb, 9'h0d5);
  assign p1_or_137450_comb = p1_prod__459_comb | 32'h0000_0080;
  assign p1_or_137451_comb = p1_prod__464_comb | 32'h0000_0080;
  assign p1_smul_57450_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__62_squeezed_comb, 9'h12b);
  assign p1_smul_57452_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__63_squeezed_comb, 9'h105);
  assign p1_smul_57582_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted_squeezed_comb, 9'h0d5);
  assign p1_or_137581_comb = p1_prod__25_comb | 32'h0000_0080;
  assign p1_smul_57586_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__2_squeezed_comb, 9'h105);
  assign p1_smul_57592_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__5_squeezed_comb, 9'h0fb);
  assign p1_or_137592_comb = p1_prod__30_comb | 32'h0000_0080;
  assign p1_smul_57596_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__7_squeezed_comb, 9'h12b);
  assign p1_smul_57598_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__8_squeezed_comb, 9'h0d5);
  assign p1_or_137597_comb = p1_prod__77_comb | 32'h0000_0080;
  assign p1_smul_57602_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__10_squeezed_comb, 9'h105);
  assign p1_smul_57608_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__13_squeezed_comb, 9'h0fb);
  assign p1_or_137608_comb = p1_prod__108_comb | 32'h0000_0080;
  assign p1_smul_57612_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__15_squeezed_comb, 9'h12b);
  assign p1_smul_57630_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__24_squeezed_comb, 9'h0d5);
  assign p1_or_137613_comb = p1_prod__205_comb | 32'h0000_0080;
  assign p1_smul_57634_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__26_squeezed_comb, 9'h105);
  assign p1_smul_57640_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__29_squeezed_comb, 9'h0fb);
  assign p1_or_137624_comb = p1_prod__236_comb | 32'h0000_0080;
  assign p1_smul_57644_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__31_squeezed_comb, 9'h12b);
  assign p1_smul_57646_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__32_squeezed_comb, 9'h0d5);
  assign p1_or_137629_comb = p1_prod__269_comb | 32'h0000_0080;
  assign p1_smul_57650_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__34_squeezed_comb, 9'h105);
  assign p1_smul_57656_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__37_squeezed_comb, 9'h0fb);
  assign p1_or_137640_comb = p1_prod__300_comb | 32'h0000_0080;
  assign p1_smul_57660_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__39_squeezed_comb, 9'h12b);
  assign p1_smul_57678_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__48_squeezed_comb, 9'h0d5);
  assign p1_or_137645_comb = p1_prod__397_comb | 32'h0000_0080;
  assign p1_smul_57682_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__50_squeezed_comb, 9'h105);
  assign p1_smul_57688_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__53_squeezed_comb, 9'h0fb);
  assign p1_or_137656_comb = p1_prod__428_comb | 32'h0000_0080;
  assign p1_smul_57692_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__55_squeezed_comb, 9'h12b);
  assign p1_smul_57694_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__56_squeezed_comb, 9'h0d5);
  assign p1_or_137661_comb = p1_prod__461_comb | 32'h0000_0080;
  assign p1_smul_57698_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__58_squeezed_comb, 9'h105);
  assign p1_smul_57704_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__61_squeezed_comb, 9'h0fb);
  assign p1_or_137672_comb = p1_prod__492_comb | 32'h0000_0080;
  assign p1_smul_57708_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__63_squeezed_comb, 9'h12b);
  assign p1_smul_57710_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted_squeezed_comb, 9'h0b5);
  assign p1_smul_57712_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__1_squeezed_comb, 9'h14b);
  assign p1_smul_57714_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__2_squeezed_comb, 9'h14b);
  assign p1_smul_57716_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__3_squeezed_comb, 9'h0b5);
  assign p1_smul_57718_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__4_squeezed_comb, 9'h0b5);
  assign p1_smul_57720_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__5_squeezed_comb, 9'h14b);
  assign p1_smul_57722_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__6_squeezed_comb, 9'h14b);
  assign p1_smul_57724_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__7_squeezed_comb, 9'h0b5);
  assign p1_smul_57726_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__8_squeezed_comb, 9'h0b5);
  assign p1_smul_57728_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__9_squeezed_comb, 9'h14b);
  assign p1_smul_57730_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__10_squeezed_comb, 9'h14b);
  assign p1_smul_57732_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__11_squeezed_comb, 9'h0b5);
  assign p1_smul_57734_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__12_squeezed_comb, 9'h0b5);
  assign p1_smul_57736_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__13_squeezed_comb, 9'h14b);
  assign p1_smul_57738_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__14_squeezed_comb, 9'h14b);
  assign p1_smul_57740_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__15_squeezed_comb, 9'h0b5);
  assign p1_smul_57758_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__24_squeezed_comb, 9'h0b5);
  assign p1_smul_57760_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__25_squeezed_comb, 9'h14b);
  assign p1_smul_57762_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__26_squeezed_comb, 9'h14b);
  assign p1_smul_57764_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__27_squeezed_comb, 9'h0b5);
  assign p1_smul_57766_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__28_squeezed_comb, 9'h0b5);
  assign p1_smul_57768_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__29_squeezed_comb, 9'h14b);
  assign p1_smul_57770_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__30_squeezed_comb, 9'h14b);
  assign p1_smul_57772_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__31_squeezed_comb, 9'h0b5);
  assign p1_smul_57774_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__32_squeezed_comb, 9'h0b5);
  assign p1_smul_57776_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__33_squeezed_comb, 9'h14b);
  assign p1_smul_57778_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__34_squeezed_comb, 9'h14b);
  assign p1_smul_57780_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__35_squeezed_comb, 9'h0b5);
  assign p1_smul_57782_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__36_squeezed_comb, 9'h0b5);
  assign p1_smul_57784_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__37_squeezed_comb, 9'h14b);
  assign p1_smul_57786_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__38_squeezed_comb, 9'h14b);
  assign p1_smul_57788_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__39_squeezed_comb, 9'h0b5);
  assign p1_smul_57806_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__48_squeezed_comb, 9'h0b5);
  assign p1_smul_57808_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__49_squeezed_comb, 9'h14b);
  assign p1_smul_57810_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__50_squeezed_comb, 9'h14b);
  assign p1_smul_57812_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__51_squeezed_comb, 9'h0b5);
  assign p1_smul_57814_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__52_squeezed_comb, 9'h0b5);
  assign p1_smul_57816_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__53_squeezed_comb, 9'h14b);
  assign p1_smul_57818_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__54_squeezed_comb, 9'h14b);
  assign p1_smul_57820_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__55_squeezed_comb, 9'h0b5);
  assign p1_smul_57822_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__56_squeezed_comb, 9'h0b5);
  assign p1_smul_57824_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__57_squeezed_comb, 9'h14b);
  assign p1_smul_57826_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__58_squeezed_comb, 9'h14b);
  assign p1_smul_57828_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__59_squeezed_comb, 9'h0b5);
  assign p1_smul_57830_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__60_squeezed_comb, 9'h0b5);
  assign p1_smul_57832_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__61_squeezed_comb, 9'h14b);
  assign p1_smul_57834_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__62_squeezed_comb, 9'h14b);
  assign p1_smul_57836_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__63_squeezed_comb, 9'h0b5);
  assign p1_smul_57840_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__1_squeezed_comb, 9'h105);
  assign p1_or_137776_comb = p1_prod__42_comb | 32'h0000_0080;
  assign p1_smul_57844_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__3_squeezed_comb, 9'h0d5);
  assign p1_smul_57846_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__4_squeezed_comb, 9'h0d5);
  assign p1_or_137781_comb = p1_prod__45_comb | 32'h0000_0080;
  assign p1_smul_57850_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__6_squeezed_comb, 9'h105);
  assign p1_smul_57856_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__9_squeezed_comb, 9'h105);
  assign p1_or_137792_comb = p1_prod__97_comb | 32'h0000_0080;
  assign p1_smul_57860_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__11_squeezed_comb, 9'h0d5);
  assign p1_smul_57862_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__12_squeezed_comb, 9'h0d5);
  assign p1_or_137797_comb = p1_prod__115_comb | 32'h0000_0080;
  assign p1_smul_57866_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__14_squeezed_comb, 9'h105);
  assign p1_smul_57888_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__25_squeezed_comb, 9'h105);
  assign p1_or_137808_comb = p1_prod__225_comb | 32'h0000_0080;
  assign p1_smul_57892_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__27_squeezed_comb, 9'h0d5);
  assign p1_smul_57894_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__28_squeezed_comb, 9'h0d5);
  assign p1_or_137813_comb = p1_prod__243_comb | 32'h0000_0080;
  assign p1_smul_57898_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__30_squeezed_comb, 9'h105);
  assign p1_smul_57904_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__33_squeezed_comb, 9'h105);
  assign p1_or_137824_comb = p1_prod__289_comb | 32'h0000_0080;
  assign p1_smul_57908_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__35_squeezed_comb, 9'h0d5);
  assign p1_smul_57910_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__36_squeezed_comb, 9'h0d5);
  assign p1_or_137829_comb = p1_prod__307_comb | 32'h0000_0080;
  assign p1_smul_57914_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__38_squeezed_comb, 9'h105);
  assign p1_smul_57936_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__49_squeezed_comb, 9'h105);
  assign p1_or_137840_comb = p1_prod__417_comb | 32'h0000_0080;
  assign p1_smul_57940_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__51_squeezed_comb, 9'h0d5);
  assign p1_smul_57942_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__52_squeezed_comb, 9'h0d5);
  assign p1_or_137845_comb = p1_prod__435_comb | 32'h0000_0080;
  assign p1_smul_57946_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__54_squeezed_comb, 9'h105);
  assign p1_smul_57952_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__57_squeezed_comb, 9'h105);
  assign p1_or_137856_comb = p1_prod__481_comb | 32'h0000_0080;
  assign p1_smul_57956_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__59_squeezed_comb, 9'h0d5);
  assign p1_smul_57958_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__60_squeezed_comb, 9'h0d5);
  assign p1_or_137861_comb = p1_prod__499_comb | 32'h0000_0080;
  assign p1_smul_57962_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__62_squeezed_comb, 9'h105);
  assign p1_or_137987_comb = p1_prod__56_comb | 32'h0000_0080;
  assign p1_smul_58098_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__2_squeezed_comb, 9'h0d5);
  assign p1_smul_58100_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__3_squeezed_comb, 9'h105);
  assign p1_smul_58102_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__4_squeezed_comb, 9'h105);
  assign p1_smul_58104_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__5_squeezed_comb, 9'h0d5);
  assign p1_or_138002_comb = p1_prod__63_comb | 32'h0000_0080;
  assign p1_or_138003_comb = p1_prod__99_comb | 32'h0000_0080;
  assign p1_smul_58114_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__10_squeezed_comb, 9'h0d5);
  assign p1_smul_58116_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__11_squeezed_comb, 9'h105);
  assign p1_smul_58118_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__12_squeezed_comb, 9'h105);
  assign p1_smul_58120_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__13_squeezed_comb, 9'h0d5);
  assign p1_or_138018_comb = p1_prod__127_comb | 32'h0000_0080;
  assign p1_or_138019_comb = p1_prod__227_comb | 32'h0000_0080;
  assign p1_smul_58146_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__26_squeezed_comb, 9'h0d5);
  assign p1_smul_58148_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__27_squeezed_comb, 9'h105);
  assign p1_smul_58150_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__28_squeezed_comb, 9'h105);
  assign p1_smul_58152_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__29_squeezed_comb, 9'h0d5);
  assign p1_or_138034_comb = p1_prod__255_comb | 32'h0000_0080;
  assign p1_or_138035_comb = p1_prod__291_comb | 32'h0000_0080;
  assign p1_smul_58162_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__34_squeezed_comb, 9'h0d5);
  assign p1_smul_58164_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__35_squeezed_comb, 9'h105);
  assign p1_smul_58166_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__36_squeezed_comb, 9'h105);
  assign p1_smul_58168_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__37_squeezed_comb, 9'h0d5);
  assign p1_or_138050_comb = p1_prod__319_comb | 32'h0000_0080;
  assign p1_or_138051_comb = p1_prod__419_comb | 32'h0000_0080;
  assign p1_smul_58194_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__50_squeezed_comb, 9'h0d5);
  assign p1_smul_58196_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__51_squeezed_comb, 9'h105);
  assign p1_smul_58198_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__52_squeezed_comb, 9'h105);
  assign p1_smul_58200_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__53_squeezed_comb, 9'h0d5);
  assign p1_or_138066_comb = p1_prod__447_comb | 32'h0000_0080;
  assign p1_or_138067_comb = p1_prod__483_comb | 32'h0000_0080;
  assign p1_smul_58210_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__58_squeezed_comb, 9'h0d5);
  assign p1_smul_58212_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__59_squeezed_comb, 9'h105);
  assign p1_smul_58214_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__60_squeezed_comb, 9'h105);
  assign p1_smul_58216_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__61_squeezed_comb, 9'h0d5);
  assign p1_or_138082_comb = p1_prod__511_comb | 32'h0000_0080;
  assign p1_sel_138083_comb = $signed(p1_shifted__16_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__16_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__16_squeezed_comb, p1_smul_57326_TrailingBits___16_comb};
  assign p1_sel_138084_comb = $signed(p1_shifted__17_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__17_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__17_squeezed_comb, p1_smul_57326_TrailingBits___17_comb};
  assign p1_sel_138085_comb = $signed(p1_shifted__18_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__18_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__18_squeezed_comb, p1_smul_57326_TrailingBits___18_comb};
  assign p1_sel_138086_comb = $signed(p1_shifted__19_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__19_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__19_squeezed_comb, p1_smul_57326_TrailingBits___19_comb};
  assign p1_sel_138087_comb = $signed(p1_shifted__20_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__20_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__20_squeezed_comb, p1_smul_57326_TrailingBits___20_comb};
  assign p1_sel_138088_comb = $signed(p1_shifted__21_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__21_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__21_squeezed_comb, p1_smul_57326_TrailingBits___21_comb};
  assign p1_sel_138089_comb = $signed(p1_shifted__22_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__22_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__22_squeezed_comb, p1_smul_57326_TrailingBits___22_comb};
  assign p1_sel_138090_comb = $signed(p1_shifted__23_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__23_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__23_squeezed_comb, p1_smul_57326_TrailingBits___23_comb};
  assign p1_sel_138091_comb = $signed(p1_shifted__40_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__40_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__40_squeezed_comb, p1_smul_57326_TrailingBits___40_comb};
  assign p1_sel_138092_comb = $signed(p1_shifted__41_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__41_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__41_squeezed_comb, p1_smul_57326_TrailingBits___41_comb};
  assign p1_sel_138093_comb = $signed(p1_shifted__42_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__42_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__42_squeezed_comb, p1_smul_57326_TrailingBits___42_comb};
  assign p1_sel_138094_comb = $signed(p1_shifted__43_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__43_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__43_squeezed_comb, p1_smul_57326_TrailingBits___43_comb};
  assign p1_sel_138095_comb = $signed(p1_shifted__44_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__44_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__44_squeezed_comb, p1_smul_57326_TrailingBits___44_comb};
  assign p1_sel_138096_comb = $signed(p1_shifted__45_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__45_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__45_squeezed_comb, p1_smul_57326_TrailingBits___45_comb};
  assign p1_sel_138097_comb = $signed(p1_shifted__46_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__46_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__46_squeezed_comb, p1_smul_57326_TrailingBits___46_comb};
  assign p1_sel_138098_comb = $signed(p1_shifted__47_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__47_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__47_squeezed_comb, p1_smul_57326_TrailingBits___47_comb};
  assign p1_sel_138547_comb = $signed(p1_shifted_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted_squeezed_comb, p1_smul_57326_TrailingBits__comb};
  assign p1_sel_138548_comb = $signed(p1_shifted__1_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__1_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__1_squeezed_comb, p1_smul_57326_TrailingBits___1_comb};
  assign p1_sel_138549_comb = $signed(p1_shifted__2_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__2_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__2_squeezed_comb, p1_smul_57326_TrailingBits___2_comb};
  assign p1_sel_138550_comb = $signed(p1_shifted__3_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__3_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__3_squeezed_comb, p1_smul_57326_TrailingBits___3_comb};
  assign p1_sel_138551_comb = $signed(p1_shifted__4_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__4_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__4_squeezed_comb, p1_smul_57326_TrailingBits___4_comb};
  assign p1_sel_138552_comb = $signed(p1_shifted__5_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__5_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__5_squeezed_comb, p1_smul_57326_TrailingBits___5_comb};
  assign p1_sel_138553_comb = $signed(p1_shifted__6_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__6_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__6_squeezed_comb, p1_smul_57326_TrailingBits___6_comb};
  assign p1_sel_138554_comb = $signed(p1_shifted__7_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__7_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__7_squeezed_comb, p1_smul_57326_TrailingBits___7_comb};
  assign p1_sel_138555_comb = $signed(p1_shifted__8_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__8_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__8_squeezed_comb, p1_smul_57326_TrailingBits___8_comb};
  assign p1_sel_138556_comb = $signed(p1_shifted__9_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__9_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__9_squeezed_comb, p1_smul_57326_TrailingBits___9_comb};
  assign p1_sel_138557_comb = $signed(p1_shifted__10_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__10_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__10_squeezed_comb, p1_smul_57326_TrailingBits___10_comb};
  assign p1_sel_138558_comb = $signed(p1_shifted__11_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__11_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__11_squeezed_comb, p1_smul_57326_TrailingBits___11_comb};
  assign p1_sel_138559_comb = $signed(p1_shifted__12_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__12_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__12_squeezed_comb, p1_smul_57326_TrailingBits___12_comb};
  assign p1_sel_138560_comb = $signed(p1_shifted__13_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__13_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__13_squeezed_comb, p1_smul_57326_TrailingBits___13_comb};
  assign p1_sel_138561_comb = $signed(p1_shifted__14_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__14_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__14_squeezed_comb, p1_smul_57326_TrailingBits___14_comb};
  assign p1_sel_138562_comb = $signed(p1_shifted__15_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__15_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__15_squeezed_comb, p1_smul_57326_TrailingBits___15_comb};
  assign p1_sel_138563_comb = $signed(p1_shifted__24_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__24_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__24_squeezed_comb, p1_smul_57326_TrailingBits___24_comb};
  assign p1_sel_138564_comb = $signed(p1_shifted__25_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__25_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__25_squeezed_comb, p1_smul_57326_TrailingBits___25_comb};
  assign p1_sel_138565_comb = $signed(p1_shifted__26_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__26_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__26_squeezed_comb, p1_smul_57326_TrailingBits___26_comb};
  assign p1_sel_138566_comb = $signed(p1_shifted__27_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__27_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__27_squeezed_comb, p1_smul_57326_TrailingBits___27_comb};
  assign p1_sel_138567_comb = $signed(p1_shifted__28_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__28_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__28_squeezed_comb, p1_smul_57326_TrailingBits___28_comb};
  assign p1_sel_138568_comb = $signed(p1_shifted__29_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__29_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__29_squeezed_comb, p1_smul_57326_TrailingBits___29_comb};
  assign p1_sel_138569_comb = $signed(p1_shifted__30_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__30_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__30_squeezed_comb, p1_smul_57326_TrailingBits___30_comb};
  assign p1_sel_138570_comb = $signed(p1_shifted__31_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__31_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__31_squeezed_comb, p1_smul_57326_TrailingBits___31_comb};
  assign p1_sel_138571_comb = $signed(p1_shifted__32_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__32_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__32_squeezed_comb, p1_smul_57326_TrailingBits___32_comb};
  assign p1_sel_138572_comb = $signed(p1_shifted__33_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__33_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__33_squeezed_comb, p1_smul_57326_TrailingBits___33_comb};
  assign p1_sel_138573_comb = $signed(p1_shifted__34_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__34_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__34_squeezed_comb, p1_smul_57326_TrailingBits___34_comb};
  assign p1_sel_138574_comb = $signed(p1_shifted__35_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__35_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__35_squeezed_comb, p1_smul_57326_TrailingBits___35_comb};
  assign p1_sel_138575_comb = $signed(p1_shifted__36_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__36_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__36_squeezed_comb, p1_smul_57326_TrailingBits___36_comb};
  assign p1_sel_138576_comb = $signed(p1_shifted__37_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__37_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__37_squeezed_comb, p1_smul_57326_TrailingBits___37_comb};
  assign p1_sel_138577_comb = $signed(p1_shifted__38_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__38_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__38_squeezed_comb, p1_smul_57326_TrailingBits___38_comb};
  assign p1_sel_138578_comb = $signed(p1_shifted__39_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__39_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__39_squeezed_comb, p1_smul_57326_TrailingBits___39_comb};
  assign p1_sel_138579_comb = $signed(p1_shifted__48_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__48_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__48_squeezed_comb, p1_smul_57326_TrailingBits___48_comb};
  assign p1_sel_138580_comb = $signed(p1_shifted__49_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__49_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__49_squeezed_comb, p1_smul_57326_TrailingBits___49_comb};
  assign p1_sel_138581_comb = $signed(p1_shifted__50_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__50_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__50_squeezed_comb, p1_smul_57326_TrailingBits___50_comb};
  assign p1_sel_138582_comb = $signed(p1_shifted__51_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__51_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__51_squeezed_comb, p1_smul_57326_TrailingBits___51_comb};
  assign p1_sel_138583_comb = $signed(p1_shifted__52_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__52_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__52_squeezed_comb, p1_smul_57326_TrailingBits___52_comb};
  assign p1_sel_138584_comb = $signed(p1_shifted__53_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__53_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__53_squeezed_comb, p1_smul_57326_TrailingBits___53_comb};
  assign p1_sel_138585_comb = $signed(p1_shifted__54_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__54_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__54_squeezed_comb, p1_smul_57326_TrailingBits___54_comb};
  assign p1_sel_138586_comb = $signed(p1_shifted__55_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__55_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__55_squeezed_comb, p1_smul_57326_TrailingBits___55_comb};
  assign p1_sel_138587_comb = $signed(p1_shifted__56_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__56_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__56_squeezed_comb, p1_smul_57326_TrailingBits___56_comb};
  assign p1_sel_138588_comb = $signed(p1_shifted__57_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__57_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__57_squeezed_comb, p1_smul_57326_TrailingBits___57_comb};
  assign p1_sel_138589_comb = $signed(p1_shifted__58_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__58_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__58_squeezed_comb, p1_smul_57326_TrailingBits___58_comb};
  assign p1_sel_138590_comb = $signed(p1_shifted__59_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__59_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__59_squeezed_comb, p1_smul_57326_TrailingBits___59_comb};
  assign p1_sel_138591_comb = $signed(p1_shifted__60_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__60_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__60_squeezed_comb, p1_smul_57326_TrailingBits___60_comb};
  assign p1_sel_138592_comb = $signed(p1_shifted__61_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__61_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__61_squeezed_comb, p1_smul_57326_TrailingBits___61_comb};
  assign p1_sel_138593_comb = $signed(p1_shifted__62_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__62_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__62_squeezed_comb, p1_smul_57326_TrailingBits___62_comb};
  assign p1_sel_138594_comb = $signed(p1_shifted__63_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__63_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__63_squeezed_comb, p1_smul_57326_TrailingBits___63_comb};
  assign p1_add_141347_comb = {{1{p1_sel_138083_comb[15]}}, p1_sel_138083_comb} + {{1{p1_sel_138084_comb[15]}}, p1_sel_138084_comb};
  assign p1_add_141348_comb = {{1{p1_sel_138085_comb[15]}}, p1_sel_138085_comb} + {{1{p1_sel_138086_comb[15]}}, p1_sel_138086_comb};
  assign p1_add_141349_comb = {{1{p1_sel_138087_comb[15]}}, p1_sel_138087_comb} + {{1{p1_sel_138088_comb[15]}}, p1_sel_138088_comb};
  assign p1_add_141350_comb = {{1{p1_sel_138089_comb[15]}}, p1_sel_138089_comb} + {{1{p1_sel_138090_comb[15]}}, p1_sel_138090_comb};
  assign p1_add_141351_comb = {{1{p1_sel_138091_comb[15]}}, p1_sel_138091_comb} + {{1{p1_sel_138092_comb[15]}}, p1_sel_138092_comb};
  assign p1_add_141352_comb = {{1{p1_sel_138093_comb[15]}}, p1_sel_138093_comb} + {{1{p1_sel_138094_comb[15]}}, p1_sel_138094_comb};
  assign p1_add_141353_comb = {{1{p1_sel_138095_comb[15]}}, p1_sel_138095_comb} + {{1{p1_sel_138096_comb[15]}}, p1_sel_138096_comb};
  assign p1_add_141354_comb = {{1{p1_sel_138097_comb[15]}}, p1_sel_138097_comb} + {{1{p1_sel_138098_comb[15]}}, p1_sel_138098_comb};
  assign p1_sel_141355_comb = $signed(p1_smul_57358_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57358_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57358_NarrowedMult__comb[15:0]);
  assign p1_sel_141356_comb = $signed(p1_smul_57360_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57360_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57360_NarrowedMult__comb[15:0]);
  assign p1_sel_141357_comb = $signed(p1_or_135911_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__135_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_135911_comb[23:9], 1'h0};
  assign p1_sel_141358_comb = $signed(p1_or_136986_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_136986_comb[23:9], 1'h0};
  assign p1_sel_141359_comb = $signed(p1_or_136987_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_136987_comb[23:9], 1'h0};
  assign p1_sel_141360_comb = $signed(p1_or_135918_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__150_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_135918_comb[23:9], 1'h0};
  assign p1_sel_141361_comb = $signed(p1_smul_57370_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57370_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57370_NarrowedMult__comb[15:0]);
  assign p1_sel_141362_comb = $signed(p1_smul_57372_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57372_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57372_NarrowedMult__comb[15:0]);
  assign p1_sel_141363_comb = $signed(p1_smul_57406_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57406_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57406_NarrowedMult__comb[15:0]);
  assign p1_sel_141364_comb = $signed(p1_smul_57408_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57408_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57408_NarrowedMult__comb[15:0]);
  assign p1_sel_141365_comb = $signed(p1_or_135925_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__327_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_135925_comb[23:9], 1'h0};
  assign p1_sel_141366_comb = $signed(p1_or_137002_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137002_comb[23:9], 1'h0};
  assign p1_sel_141367_comb = $signed(p1_or_137003_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137003_comb[23:9], 1'h0};
  assign p1_sel_141368_comb = $signed(p1_or_135932_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__342_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_135932_comb[23:9], 1'h0};
  assign p1_sel_141369_comb = $signed(p1_smul_57418_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57418_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57418_NarrowedMult__comb[15:0]);
  assign p1_sel_141370_comb = $signed(p1_smul_57420_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57420_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57420_NarrowedMult__comb[15:0]);
  assign p1_sel_141371_comb = $signed(p1_or_135937_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__133_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_135937_comb[23:10], 2'h0};
  assign p1_sel_141372_comb = $signed(p1_prod__136_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__136_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57488_NarrowedMult__comb, 1'h0};
  assign p1_sel_141373_comb = $signed(p1_prod__140_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__140_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57490_NarrowedMult__comb, 1'h0};
  assign p1_sel_141374_comb = $signed(p1_or_135944_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__145_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_135944_comb[23:10], 2'h0};
  assign p1_sel_141375_comb = $signed(p1_or_135947_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__151_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_135947_comb[23:10], 2'h0};
  assign p1_sel_141376_comb = $signed(p1_prod__158_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__158_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57496_NarrowedMult__comb, 1'h0};
  assign p1_sel_141377_comb = $signed(p1_prod__165_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__165_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57498_NarrowedMult__comb, 1'h0};
  assign p1_sel_141378_comb = $signed(p1_or_135954_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__171_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_135954_comb[23:10], 2'h0};
  assign p1_sel_141379_comb = $signed(p1_or_135957_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__325_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_135957_comb[23:10], 2'h0};
  assign p1_sel_141380_comb = $signed(p1_prod__328_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__328_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57536_NarrowedMult__comb, 1'h0};
  assign p1_sel_141381_comb = $signed(p1_prod__332_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__332_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57538_NarrowedMult__comb, 1'h0};
  assign p1_sel_141382_comb = $signed(p1_or_135964_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__337_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_135964_comb[23:10], 2'h0};
  assign p1_sel_141383_comb = $signed(p1_or_135967_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__343_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_135967_comb[23:10], 2'h0};
  assign p1_sel_141384_comb = $signed(p1_prod__350_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__350_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57544_NarrowedMult__comb, 1'h0};
  assign p1_sel_141385_comb = $signed(p1_prod__357_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__357_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57546_NarrowedMult__comb, 1'h0};
  assign p1_sel_141386_comb = $signed(p1_or_135974_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__363_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_135974_comb[23:10], 2'h0};
  assign p1_sel_141387_comb = $signed(p1_smul_57614_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57614_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57614_NarrowedMult__comb[15:0]);
  assign p1_sel_141388_comb = $signed(p1_or_137053_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137053_comb[23:9], 1'h0};
  assign p1_sel_141389_comb = $signed(p1_smul_57618_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57618_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57618_NarrowedMult__comb[15:0]);
  assign p1_sel_141390_comb = $signed(p1_or_135981_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__152_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_135981_comb[23:9], 1'h0};
  assign p1_sel_141391_comb = $signed(p1_or_135984_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__159_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_135984_comb[23:9], 1'h0};
  assign p1_sel_141392_comb = $signed(p1_smul_57624_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57624_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57624_NarrowedMult__comb[15:0]);
  assign p1_sel_141393_comb = $signed(p1_or_137064_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137064_comb[23:9], 1'h0};
  assign p1_sel_141394_comb = $signed(p1_smul_57628_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57628_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57628_NarrowedMult__comb[15:0]);
  assign p1_sel_141395_comb = $signed(p1_smul_57662_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57662_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57662_NarrowedMult__comb[15:0]);
  assign p1_sel_141396_comb = $signed(p1_or_137069_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137069_comb[23:9], 1'h0};
  assign p1_sel_141397_comb = $signed(p1_smul_57666_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57666_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57666_NarrowedMult__comb[15:0]);
  assign p1_sel_141398_comb = $signed(p1_or_135995_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__344_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_135995_comb[23:9], 1'h0};
  assign p1_sel_141399_comb = $signed(p1_or_135998_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__351_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_135998_comb[23:9], 1'h0};
  assign p1_sel_141400_comb = $signed(p1_smul_57672_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57672_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57672_NarrowedMult__comb[15:0]);
  assign p1_sel_141401_comb = $signed(p1_or_137080_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137080_comb[23:9], 1'h0};
  assign p1_sel_141402_comb = $signed(p1_smul_57676_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57676_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57676_NarrowedMult__comb[15:0]);
  assign p1_sel_141403_comb = $signed(p1_smul_57742_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57742_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57742_NarrowedMult__comb[15:0]);
  assign p1_sel_141404_comb = $signed(p1_smul_57744_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57744_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57744_NarrowedMult__comb[15:0]);
  assign p1_sel_141405_comb = $signed(p1_smul_57746_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57746_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57746_NarrowedMult__comb[15:0]);
  assign p1_sel_141406_comb = $signed(p1_smul_57748_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57748_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57748_NarrowedMult__comb[15:0]);
  assign p1_sel_141407_comb = $signed(p1_smul_57750_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57750_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57750_NarrowedMult__comb[15:0]);
  assign p1_sel_141408_comb = $signed(p1_smul_57752_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57752_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57752_NarrowedMult__comb[15:0]);
  assign p1_sel_141409_comb = $signed(p1_smul_57754_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57754_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57754_NarrowedMult__comb[15:0]);
  assign p1_sel_141410_comb = $signed(p1_smul_57756_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57756_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57756_NarrowedMult__comb[15:0]);
  assign p1_sel_141411_comb = $signed(p1_smul_57790_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57790_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57790_NarrowedMult__comb[15:0]);
  assign p1_sel_141412_comb = $signed(p1_smul_57792_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57792_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57792_NarrowedMult__comb[15:0]);
  assign p1_sel_141413_comb = $signed(p1_smul_57794_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57794_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57794_NarrowedMult__comb[15:0]);
  assign p1_sel_141414_comb = $signed(p1_smul_57796_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57796_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57796_NarrowedMult__comb[15:0]);
  assign p1_sel_141415_comb = $signed(p1_smul_57798_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57798_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57798_NarrowedMult__comb[15:0]);
  assign p1_sel_141416_comb = $signed(p1_smul_57800_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57800_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57800_NarrowedMult__comb[15:0]);
  assign p1_sel_141417_comb = $signed(p1_smul_57802_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57802_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57802_NarrowedMult__comb[15:0]);
  assign p1_sel_141418_comb = $signed(p1_smul_57804_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57804_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57804_NarrowedMult__comb[15:0]);
  assign p1_sel_141419_comb = $signed(p1_or_136021_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__148_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136021_comb[23:9], 1'h0};
  assign p1_sel_141420_comb = $signed(p1_smul_57872_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57872_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57872_NarrowedMult__comb[15:0]);
  assign p1_sel_141421_comb = $signed(p1_or_137120_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137120_comb[23:9], 1'h0};
  assign p1_sel_141422_comb = $signed(p1_smul_57876_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57876_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57876_NarrowedMult__comb[15:0]);
  assign p1_sel_141423_comb = $signed(p1_smul_57878_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57878_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57878_NarrowedMult__comb[15:0]);
  assign p1_sel_141424_comb = $signed(p1_or_137125_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137125_comb[23:9], 1'h0};
  assign p1_sel_141425_comb = $signed(p1_smul_57882_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57882_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57882_NarrowedMult__comb[15:0]);
  assign p1_sel_141426_comb = $signed(p1_or_136032_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__186_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136032_comb[23:9], 1'h0};
  assign p1_sel_141427_comb = $signed(p1_or_136035_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__340_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136035_comb[23:9], 1'h0};
  assign p1_sel_141428_comb = $signed(p1_smul_57920_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57920_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57920_NarrowedMult__comb[15:0]);
  assign p1_sel_141429_comb = $signed(p1_or_137136_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137136_comb[23:9], 1'h0};
  assign p1_sel_141430_comb = $signed(p1_smul_57924_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57924_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57924_NarrowedMult__comb[15:0]);
  assign p1_sel_141431_comb = $signed(p1_smul_57926_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57926_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57926_NarrowedMult__comb[15:0]);
  assign p1_sel_141432_comb = $signed(p1_or_137141_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137141_comb[23:9], 1'h0};
  assign p1_sel_141433_comb = $signed(p1_smul_57930_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57930_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57930_NarrowedMult__comb[15:0]);
  assign p1_sel_141434_comb = $signed(p1_or_136046_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__378_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136046_comb[23:9], 1'h0};
  assign p1_sel_141435_comb = $signed(p1_prod__155_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__155_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57998_NarrowedMult__comb, 1'h0};
  assign p1_sel_141436_comb = $signed(p1_or_136051_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__162_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136051_comb[23:10], 2'h0};
  assign p1_sel_141437_comb = $signed(p1_prod__169_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__169_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58002_NarrowedMult__comb, 1'h0};
  assign p1_sel_141438_comb = $signed(p1_or_136056_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__175_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136056_comb[23:10], 2'h0};
  assign p1_sel_141439_comb = $signed(p1_or_136059_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__180_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136059_comb[23:10], 2'h0};
  assign p1_sel_141440_comb = $signed(p1_prod__184_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__184_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58008_NarrowedMult__comb, 1'h0};
  assign p1_sel_141441_comb = $signed(p1_or_136064_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__187_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136064_comb[23:10], 2'h0};
  assign p1_sel_141442_comb = $signed(p1_prod__189_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__189_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58012_NarrowedMult__comb, 1'h0};
  assign p1_sel_141443_comb = $signed(p1_prod__347_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__347_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58046_NarrowedMult__comb, 1'h0};
  assign p1_sel_141444_comb = $signed(p1_or_136071_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__354_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136071_comb[23:10], 2'h0};
  assign p1_sel_141445_comb = $signed(p1_prod__361_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__361_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58050_NarrowedMult__comb, 1'h0};
  assign p1_sel_141446_comb = $signed(p1_or_136076_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__367_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136076_comb[23:10], 2'h0};
  assign p1_sel_141447_comb = $signed(p1_or_136079_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__372_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136079_comb[23:10], 2'h0};
  assign p1_sel_141448_comb = $signed(p1_prod__376_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__376_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58056_NarrowedMult__comb, 1'h0};
  assign p1_sel_141449_comb = $signed(p1_or_136084_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__379_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136084_comb[23:10], 2'h0};
  assign p1_sel_141450_comb = $signed(p1_prod__381_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__381_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58060_NarrowedMult__comb, 1'h0};
  assign p1_sel_141451_comb = $signed(p1_or_137187_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137187_comb[23:9], 1'h0};
  assign p1_sel_141452_comb = $signed(p1_or_136091_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__170_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136091_comb[23:9], 1'h0};
  assign p1_sel_141453_comb = $signed(p1_smul_58130_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58130_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58130_NarrowedMult__comb[15:0]);
  assign p1_sel_141454_comb = $signed(p1_smul_58132_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58132_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58132_NarrowedMult__comb[15:0]);
  assign p1_sel_141455_comb = $signed(p1_smul_58134_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58134_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58134_NarrowedMult__comb[15:0]);
  assign p1_sel_141456_comb = $signed(p1_smul_58136_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58136_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58136_NarrowedMult__comb[15:0]);
  assign p1_sel_141457_comb = $signed(p1_or_136098_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__190_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136098_comb[23:9], 1'h0};
  assign p1_sel_141458_comb = $signed(p1_or_137202_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137202_comb[23:9], 1'h0};
  assign p1_sel_141459_comb = $signed(p1_or_137203_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137203_comb[23:9], 1'h0};
  assign p1_sel_141460_comb = $signed(p1_or_136105_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__362_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136105_comb[23:9], 1'h0};
  assign p1_sel_141461_comb = $signed(p1_smul_58178_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58178_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58178_NarrowedMult__comb[15:0]);
  assign p1_sel_141462_comb = $signed(p1_smul_58180_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58180_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58180_NarrowedMult__comb[15:0]);
  assign p1_sel_141463_comb = $signed(p1_smul_58182_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58182_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58182_NarrowedMult__comb[15:0]);
  assign p1_sel_141464_comb = $signed(p1_smul_58184_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58184_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58184_NarrowedMult__comb[15:0]);
  assign p1_sel_141465_comb = $signed(p1_or_136112_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__382_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136112_comb[23:9], 1'h0};
  assign p1_sel_141466_comb = $signed(p1_or_137218_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137218_comb[23:9], 1'h0};
  assign p1_add_141467_comb = {{1{p1_sel_138547_comb[15]}}, p1_sel_138547_comb} + {{1{p1_sel_138548_comb[15]}}, p1_sel_138548_comb};
  assign p1_add_141468_comb = {{1{p1_sel_138549_comb[15]}}, p1_sel_138549_comb} + {{1{p1_sel_138550_comb[15]}}, p1_sel_138550_comb};
  assign p1_add_141469_comb = {{1{p1_sel_138551_comb[15]}}, p1_sel_138551_comb} + {{1{p1_sel_138552_comb[15]}}, p1_sel_138552_comb};
  assign p1_add_141470_comb = {{1{p1_sel_138553_comb[15]}}, p1_sel_138553_comb} + {{1{p1_sel_138554_comb[15]}}, p1_sel_138554_comb};
  assign p1_add_141471_comb = {{1{p1_sel_138555_comb[15]}}, p1_sel_138555_comb} + {{1{p1_sel_138556_comb[15]}}, p1_sel_138556_comb};
  assign p1_add_141472_comb = {{1{p1_sel_138557_comb[15]}}, p1_sel_138557_comb} + {{1{p1_sel_138558_comb[15]}}, p1_sel_138558_comb};
  assign p1_add_141473_comb = {{1{p1_sel_138559_comb[15]}}, p1_sel_138559_comb} + {{1{p1_sel_138560_comb[15]}}, p1_sel_138560_comb};
  assign p1_add_141474_comb = {{1{p1_sel_138561_comb[15]}}, p1_sel_138561_comb} + {{1{p1_sel_138562_comb[15]}}, p1_sel_138562_comb};
  assign p1_add_141475_comb = {{1{p1_sel_138563_comb[15]}}, p1_sel_138563_comb} + {{1{p1_sel_138564_comb[15]}}, p1_sel_138564_comb};
  assign p1_add_141476_comb = {{1{p1_sel_138565_comb[15]}}, p1_sel_138565_comb} + {{1{p1_sel_138566_comb[15]}}, p1_sel_138566_comb};
  assign p1_add_141477_comb = {{1{p1_sel_138567_comb[15]}}, p1_sel_138567_comb} + {{1{p1_sel_138568_comb[15]}}, p1_sel_138568_comb};
  assign p1_add_141478_comb = {{1{p1_sel_138569_comb[15]}}, p1_sel_138569_comb} + {{1{p1_sel_138570_comb[15]}}, p1_sel_138570_comb};
  assign p1_add_141479_comb = {{1{p1_sel_138571_comb[15]}}, p1_sel_138571_comb} + {{1{p1_sel_138572_comb[15]}}, p1_sel_138572_comb};
  assign p1_add_141480_comb = {{1{p1_sel_138573_comb[15]}}, p1_sel_138573_comb} + {{1{p1_sel_138574_comb[15]}}, p1_sel_138574_comb};
  assign p1_add_141481_comb = {{1{p1_sel_138575_comb[15]}}, p1_sel_138575_comb} + {{1{p1_sel_138576_comb[15]}}, p1_sel_138576_comb};
  assign p1_add_141482_comb = {{1{p1_sel_138577_comb[15]}}, p1_sel_138577_comb} + {{1{p1_sel_138578_comb[15]}}, p1_sel_138578_comb};
  assign p1_add_141483_comb = {{1{p1_sel_138579_comb[15]}}, p1_sel_138579_comb} + {{1{p1_sel_138580_comb[15]}}, p1_sel_138580_comb};
  assign p1_add_141484_comb = {{1{p1_sel_138581_comb[15]}}, p1_sel_138581_comb} + {{1{p1_sel_138582_comb[15]}}, p1_sel_138582_comb};
  assign p1_add_141485_comb = {{1{p1_sel_138583_comb[15]}}, p1_sel_138583_comb} + {{1{p1_sel_138584_comb[15]}}, p1_sel_138584_comb};
  assign p1_add_141486_comb = {{1{p1_sel_138585_comb[15]}}, p1_sel_138585_comb} + {{1{p1_sel_138586_comb[15]}}, p1_sel_138586_comb};
  assign p1_add_141487_comb = {{1{p1_sel_138587_comb[15]}}, p1_sel_138587_comb} + {{1{p1_sel_138588_comb[15]}}, p1_sel_138588_comb};
  assign p1_add_141488_comb = {{1{p1_sel_138589_comb[15]}}, p1_sel_138589_comb} + {{1{p1_sel_138590_comb[15]}}, p1_sel_138590_comb};
  assign p1_add_141489_comb = {{1{p1_sel_138591_comb[15]}}, p1_sel_138591_comb} + {{1{p1_sel_138592_comb[15]}}, p1_sel_138592_comb};
  assign p1_add_141490_comb = {{1{p1_sel_138593_comb[15]}}, p1_sel_138593_comb} + {{1{p1_sel_138594_comb[15]}}, p1_sel_138594_comb};
  assign p1_sel_141491_comb = $signed(p1_smul_57326_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57326_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57326_NarrowedMult__comb[15:0]);
  assign p1_sel_141492_comb = $signed(p1_smul_57328_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57328_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57328_NarrowedMult__comb[15:0]);
  assign p1_sel_141493_comb = $signed(p1_or_136311_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__10_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136311_comb[23:9], 1'h0};
  assign p1_sel_141494_comb = $signed(p1_or_137370_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137370_comb[23:9], 1'h0};
  assign p1_sel_141495_comb = $signed(p1_or_137371_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137371_comb[23:9], 1'h0};
  assign p1_sel_141496_comb = $signed(p1_or_136318_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__13_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136318_comb[23:9], 1'h0};
  assign p1_sel_141497_comb = $signed(p1_smul_57338_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57338_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57338_NarrowedMult__comb[15:0]);
  assign p1_sel_141498_comb = $signed(p1_smul_57340_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57340_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57340_NarrowedMult__comb[15:0]);
  assign p1_sel_141499_comb = $signed(p1_smul_57342_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57342_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57342_NarrowedMult__comb[15:0]);
  assign p1_sel_141500_comb = $signed(p1_smul_57344_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57344_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57344_NarrowedMult__comb[15:0]);
  assign p1_sel_141501_comb = $signed(p1_or_136325_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__71_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136325_comb[23:9], 1'h0};
  assign p1_sel_141502_comb = $signed(p1_or_137386_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137386_comb[23:9], 1'h0};
  assign p1_sel_141503_comb = $signed(p1_or_137387_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137387_comb[23:9], 1'h0};
  assign p1_sel_141504_comb = $signed(p1_or_136332_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__86_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136332_comb[23:9], 1'h0};
  assign p1_sel_141505_comb = $signed(p1_smul_57354_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57354_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57354_NarrowedMult__comb[15:0]);
  assign p1_sel_141506_comb = $signed(p1_smul_57356_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57356_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57356_NarrowedMult__comb[15:0]);
  assign p1_sel_141507_comb = $signed(p1_smul_57374_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57374_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57374_NarrowedMult__comb[15:0]);
  assign p1_sel_141508_comb = $signed(p1_smul_57376_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57376_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57376_NarrowedMult__comb[15:0]);
  assign p1_sel_141509_comb = $signed(p1_or_136339_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__199_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136339_comb[23:9], 1'h0};
  assign p1_sel_141510_comb = $signed(p1_or_137402_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137402_comb[23:9], 1'h0};
  assign p1_sel_141511_comb = $signed(p1_or_137403_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137403_comb[23:9], 1'h0};
  assign p1_sel_141512_comb = $signed(p1_or_136346_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__214_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136346_comb[23:9], 1'h0};
  assign p1_sel_141513_comb = $signed(p1_smul_57386_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57386_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57386_NarrowedMult__comb[15:0]);
  assign p1_sel_141514_comb = $signed(p1_smul_57388_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57388_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57388_NarrowedMult__comb[15:0]);
  assign p1_sel_141515_comb = $signed(p1_smul_57390_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57390_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57390_NarrowedMult__comb[15:0]);
  assign p1_sel_141516_comb = $signed(p1_smul_57392_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57392_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57392_NarrowedMult__comb[15:0]);
  assign p1_sel_141517_comb = $signed(p1_or_136353_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__263_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136353_comb[23:9], 1'h0};
  assign p1_sel_141518_comb = $signed(p1_or_137418_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137418_comb[23:9], 1'h0};
  assign p1_sel_141519_comb = $signed(p1_or_137419_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137419_comb[23:9], 1'h0};
  assign p1_sel_141520_comb = $signed(p1_or_136360_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__278_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136360_comb[23:9], 1'h0};
  assign p1_sel_141521_comb = $signed(p1_smul_57402_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57402_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57402_NarrowedMult__comb[15:0]);
  assign p1_sel_141522_comb = $signed(p1_smul_57404_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57404_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57404_NarrowedMult__comb[15:0]);
  assign p1_sel_141523_comb = $signed(p1_smul_57422_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57422_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57422_NarrowedMult__comb[15:0]);
  assign p1_sel_141524_comb = $signed(p1_smul_57424_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57424_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57424_NarrowedMult__comb[15:0]);
  assign p1_sel_141525_comb = $signed(p1_or_136367_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__391_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136367_comb[23:9], 1'h0};
  assign p1_sel_141526_comb = $signed(p1_or_137434_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137434_comb[23:9], 1'h0};
  assign p1_sel_141527_comb = $signed(p1_or_137435_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137435_comb[23:9], 1'h0};
  assign p1_sel_141528_comb = $signed(p1_or_136374_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__406_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136374_comb[23:9], 1'h0};
  assign p1_sel_141529_comb = $signed(p1_smul_57434_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57434_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57434_NarrowedMult__comb[15:0]);
  assign p1_sel_141530_comb = $signed(p1_smul_57436_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57436_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57436_NarrowedMult__comb[15:0]);
  assign p1_sel_141531_comb = $signed(p1_smul_57438_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57438_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57438_NarrowedMult__comb[15:0]);
  assign p1_sel_141532_comb = $signed(p1_smul_57440_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57440_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57440_NarrowedMult__comb[15:0]);
  assign p1_sel_141533_comb = $signed(p1_or_136381_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__455_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136381_comb[23:9], 1'h0};
  assign p1_sel_141534_comb = $signed(p1_or_137450_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137450_comb[23:9], 1'h0};
  assign p1_sel_141535_comb = $signed(p1_or_137451_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137451_comb[23:9], 1'h0};
  assign p1_sel_141536_comb = $signed(p1_or_136388_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__470_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136388_comb[23:9], 1'h0};
  assign p1_sel_141537_comb = $signed(p1_smul_57450_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57450_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57450_NarrowedMult__comb[15:0]);
  assign p1_sel_141538_comb = $signed(p1_smul_57452_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57452_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57452_NarrowedMult__comb[15:0]);
  assign p1_sel_141539_comb = $signed(p1_or_136393_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__16_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136393_comb[23:10], 2'h0};
  assign p1_sel_141540_comb = $signed(p1_prod__17_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__17_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57456_NarrowedMult__comb, 1'h0};
  assign p1_sel_141541_comb = $signed(p1_prod__18_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__18_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57458_NarrowedMult__comb, 1'h0};
  assign p1_sel_141542_comb = $signed(p1_or_136400_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__19_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136400_comb[23:10], 2'h0};
  assign p1_sel_141543_comb = $signed(p1_or_136403_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__20_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136403_comb[23:10], 2'h0};
  assign p1_sel_141544_comb = $signed(p1_prod__21_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__21_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57464_NarrowedMult__comb, 1'h0};
  assign p1_sel_141545_comb = $signed(p1_prod__22_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__22_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57466_NarrowedMult__comb, 1'h0};
  assign p1_sel_141546_comb = $signed(p1_or_136410_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__23_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136410_comb[23:10], 2'h0};
  assign p1_sel_141547_comb = $signed(p1_or_136413_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__69_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136413_comb[23:10], 2'h0};
  assign p1_sel_141548_comb = $signed(p1_prod__72_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__72_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57472_NarrowedMult__comb, 1'h0};
  assign p1_sel_141549_comb = $signed(p1_prod__76_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__76_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57474_NarrowedMult__comb, 1'h0};
  assign p1_sel_141550_comb = $signed(p1_or_136420_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__81_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136420_comb[23:10], 2'h0};
  assign p1_sel_141551_comb = $signed(p1_or_136423_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__87_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136423_comb[23:10], 2'h0};
  assign p1_sel_141552_comb = $signed(p1_prod__94_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__94_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57480_NarrowedMult__comb, 1'h0};
  assign p1_sel_141553_comb = $signed(p1_prod__101_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__101_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57482_NarrowedMult__comb, 1'h0};
  assign p1_sel_141554_comb = $signed(p1_or_136430_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__107_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136430_comb[23:10], 2'h0};
  assign p1_sel_141555_comb = $signed(p1_or_136433_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__197_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136433_comb[23:10], 2'h0};
  assign p1_sel_141556_comb = $signed(p1_prod__200_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__200_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57504_NarrowedMult__comb, 1'h0};
  assign p1_sel_141557_comb = $signed(p1_prod__204_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__204_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57506_NarrowedMult__comb, 1'h0};
  assign p1_sel_141558_comb = $signed(p1_or_136440_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__209_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136440_comb[23:10], 2'h0};
  assign p1_sel_141559_comb = $signed(p1_or_136443_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__215_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136443_comb[23:10], 2'h0};
  assign p1_sel_141560_comb = $signed(p1_prod__222_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__222_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57512_NarrowedMult__comb, 1'h0};
  assign p1_sel_141561_comb = $signed(p1_prod__229_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__229_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57514_NarrowedMult__comb, 1'h0};
  assign p1_sel_141562_comb = $signed(p1_or_136450_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__235_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136450_comb[23:10], 2'h0};
  assign p1_sel_141563_comb = $signed(p1_or_136453_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__261_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136453_comb[23:10], 2'h0};
  assign p1_sel_141564_comb = $signed(p1_prod__264_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__264_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57520_NarrowedMult__comb, 1'h0};
  assign p1_sel_141565_comb = $signed(p1_prod__268_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__268_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57522_NarrowedMult__comb, 1'h0};
  assign p1_sel_141566_comb = $signed(p1_or_136460_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__273_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136460_comb[23:10], 2'h0};
  assign p1_sel_141567_comb = $signed(p1_or_136463_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__279_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136463_comb[23:10], 2'h0};
  assign p1_sel_141568_comb = $signed(p1_prod__286_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__286_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57528_NarrowedMult__comb, 1'h0};
  assign p1_sel_141569_comb = $signed(p1_prod__293_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__293_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57530_NarrowedMult__comb, 1'h0};
  assign p1_sel_141570_comb = $signed(p1_or_136470_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__299_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136470_comb[23:10], 2'h0};
  assign p1_sel_141571_comb = $signed(p1_or_136473_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__389_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136473_comb[23:10], 2'h0};
  assign p1_sel_141572_comb = $signed(p1_prod__392_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__392_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57552_NarrowedMult__comb, 1'h0};
  assign p1_sel_141573_comb = $signed(p1_prod__396_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__396_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57554_NarrowedMult__comb, 1'h0};
  assign p1_sel_141574_comb = $signed(p1_or_136480_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__401_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136480_comb[23:10], 2'h0};
  assign p1_sel_141575_comb = $signed(p1_or_136483_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__407_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136483_comb[23:10], 2'h0};
  assign p1_sel_141576_comb = $signed(p1_prod__414_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__414_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57560_NarrowedMult__comb, 1'h0};
  assign p1_sel_141577_comb = $signed(p1_prod__421_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__421_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57562_NarrowedMult__comb, 1'h0};
  assign p1_sel_141578_comb = $signed(p1_or_136490_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__427_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136490_comb[23:10], 2'h0};
  assign p1_sel_141579_comb = $signed(p1_or_136493_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__453_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136493_comb[23:10], 2'h0};
  assign p1_sel_141580_comb = $signed(p1_prod__456_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__456_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57568_NarrowedMult__comb, 1'h0};
  assign p1_sel_141581_comb = $signed(p1_prod__460_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__460_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57570_NarrowedMult__comb, 1'h0};
  assign p1_sel_141582_comb = $signed(p1_or_136500_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__465_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136500_comb[23:10], 2'h0};
  assign p1_sel_141583_comb = $signed(p1_or_136503_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__471_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136503_comb[23:10], 2'h0};
  assign p1_sel_141584_comb = $signed(p1_prod__478_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__478_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57576_NarrowedMult__comb, 1'h0};
  assign p1_sel_141585_comb = $signed(p1_prod__485_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__485_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57578_NarrowedMult__comb, 1'h0};
  assign p1_sel_141586_comb = $signed(p1_or_136510_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__491_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136510_comb[23:10], 2'h0};
  assign p1_sel_141587_comb = $signed(p1_smul_57582_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57582_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57582_NarrowedMult__comb[15:0]);
  assign p1_sel_141588_comb = $signed(p1_or_137581_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137581_comb[23:9], 1'h0};
  assign p1_sel_141589_comb = $signed(p1_smul_57586_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57586_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57586_NarrowedMult__comb[15:0]);
  assign p1_sel_141590_comb = $signed(p1_or_136517_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__27_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136517_comb[23:9], 1'h0};
  assign p1_sel_141591_comb = $signed(p1_or_136520_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__28_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136520_comb[23:9], 1'h0};
  assign p1_sel_141592_comb = $signed(p1_smul_57592_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57592_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57592_NarrowedMult__comb[15:0]);
  assign p1_sel_141593_comb = $signed(p1_or_137592_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137592_comb[23:9], 1'h0};
  assign p1_sel_141594_comb = $signed(p1_smul_57596_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57596_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57596_NarrowedMult__comb[15:0]);
  assign p1_sel_141595_comb = $signed(p1_smul_57598_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57598_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57598_NarrowedMult__comb[15:0]);
  assign p1_sel_141596_comb = $signed(p1_or_137597_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137597_comb[23:9], 1'h0};
  assign p1_sel_141597_comb = $signed(p1_smul_57602_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57602_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57602_NarrowedMult__comb[15:0]);
  assign p1_sel_141598_comb = $signed(p1_or_136531_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__88_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136531_comb[23:9], 1'h0};
  assign p1_sel_141599_comb = $signed(p1_or_136534_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__95_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136534_comb[23:9], 1'h0};
  assign p1_sel_141600_comb = $signed(p1_smul_57608_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57608_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57608_NarrowedMult__comb[15:0]);
  assign p1_sel_141601_comb = $signed(p1_or_137608_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137608_comb[23:9], 1'h0};
  assign p1_sel_141602_comb = $signed(p1_smul_57612_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57612_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57612_NarrowedMult__comb[15:0]);
  assign p1_sel_141603_comb = $signed(p1_smul_57630_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57630_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57630_NarrowedMult__comb[15:0]);
  assign p1_sel_141604_comb = $signed(p1_or_137613_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137613_comb[23:9], 1'h0};
  assign p1_sel_141605_comb = $signed(p1_smul_57634_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57634_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57634_NarrowedMult__comb[15:0]);
  assign p1_sel_141606_comb = $signed(p1_or_136545_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__216_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136545_comb[23:9], 1'h0};
  assign p1_sel_141607_comb = $signed(p1_or_136548_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__223_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136548_comb[23:9], 1'h0};
  assign p1_sel_141608_comb = $signed(p1_smul_57640_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57640_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57640_NarrowedMult__comb[15:0]);
  assign p1_sel_141609_comb = $signed(p1_or_137624_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137624_comb[23:9], 1'h0};
  assign p1_sel_141610_comb = $signed(p1_smul_57644_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57644_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57644_NarrowedMult__comb[15:0]);
  assign p1_sel_141611_comb = $signed(p1_smul_57646_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57646_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57646_NarrowedMult__comb[15:0]);
  assign p1_sel_141612_comb = $signed(p1_or_137629_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137629_comb[23:9], 1'h0};
  assign p1_sel_141613_comb = $signed(p1_smul_57650_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57650_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57650_NarrowedMult__comb[15:0]);
  assign p1_sel_141614_comb = $signed(p1_or_136559_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__280_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136559_comb[23:9], 1'h0};
  assign p1_sel_141615_comb = $signed(p1_or_136562_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__287_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136562_comb[23:9], 1'h0};
  assign p1_sel_141616_comb = $signed(p1_smul_57656_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57656_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57656_NarrowedMult__comb[15:0]);
  assign p1_sel_141617_comb = $signed(p1_or_137640_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137640_comb[23:9], 1'h0};
  assign p1_sel_141618_comb = $signed(p1_smul_57660_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57660_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57660_NarrowedMult__comb[15:0]);
  assign p1_sel_141619_comb = $signed(p1_smul_57678_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57678_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57678_NarrowedMult__comb[15:0]);
  assign p1_sel_141620_comb = $signed(p1_or_137645_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137645_comb[23:9], 1'h0};
  assign p1_sel_141621_comb = $signed(p1_smul_57682_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57682_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57682_NarrowedMult__comb[15:0]);
  assign p1_sel_141622_comb = $signed(p1_or_136573_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__408_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136573_comb[23:9], 1'h0};
  assign p1_sel_141623_comb = $signed(p1_or_136576_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__415_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136576_comb[23:9], 1'h0};
  assign p1_sel_141624_comb = $signed(p1_smul_57688_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57688_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57688_NarrowedMult__comb[15:0]);
  assign p1_sel_141625_comb = $signed(p1_or_137656_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137656_comb[23:9], 1'h0};
  assign p1_sel_141626_comb = $signed(p1_smul_57692_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57692_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57692_NarrowedMult__comb[15:0]);
  assign p1_sel_141627_comb = $signed(p1_smul_57694_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57694_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57694_NarrowedMult__comb[15:0]);
  assign p1_sel_141628_comb = $signed(p1_or_137661_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137661_comb[23:9], 1'h0};
  assign p1_sel_141629_comb = $signed(p1_smul_57698_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57698_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57698_NarrowedMult__comb[15:0]);
  assign p1_sel_141630_comb = $signed(p1_or_136587_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__472_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136587_comb[23:9], 1'h0};
  assign p1_sel_141631_comb = $signed(p1_or_136590_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__479_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136590_comb[23:9], 1'h0};
  assign p1_sel_141632_comb = $signed(p1_smul_57704_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57704_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57704_NarrowedMult__comb[15:0]);
  assign p1_sel_141633_comb = $signed(p1_or_137672_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137672_comb[23:9], 1'h0};
  assign p1_sel_141634_comb = $signed(p1_smul_57708_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57708_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57708_NarrowedMult__comb[15:0]);
  assign p1_sel_141635_comb = $signed(p1_smul_57710_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57710_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57710_NarrowedMult__comb[15:0]);
  assign p1_sel_141636_comb = $signed(p1_smul_57712_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57712_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57712_NarrowedMult__comb[15:0]);
  assign p1_sel_141637_comb = $signed(p1_smul_57714_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57714_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57714_NarrowedMult__comb[15:0]);
  assign p1_sel_141638_comb = $signed(p1_smul_57716_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57716_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57716_NarrowedMult__comb[15:0]);
  assign p1_sel_141639_comb = $signed(p1_smul_57718_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57718_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57718_NarrowedMult__comb[15:0]);
  assign p1_sel_141640_comb = $signed(p1_smul_57720_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57720_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57720_NarrowedMult__comb[15:0]);
  assign p1_sel_141641_comb = $signed(p1_smul_57722_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57722_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57722_NarrowedMult__comb[15:0]);
  assign p1_sel_141642_comb = $signed(p1_smul_57724_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57724_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57724_NarrowedMult__comb[15:0]);
  assign p1_sel_141643_comb = $signed(p1_smul_57726_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57726_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57726_NarrowedMult__comb[15:0]);
  assign p1_sel_141644_comb = $signed(p1_smul_57728_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57728_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57728_NarrowedMult__comb[15:0]);
  assign p1_sel_141645_comb = $signed(p1_smul_57730_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57730_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57730_NarrowedMult__comb[15:0]);
  assign p1_sel_141646_comb = $signed(p1_smul_57732_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57732_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57732_NarrowedMult__comb[15:0]);
  assign p1_sel_141647_comb = $signed(p1_smul_57734_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57734_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57734_NarrowedMult__comb[15:0]);
  assign p1_sel_141648_comb = $signed(p1_smul_57736_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57736_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57736_NarrowedMult__comb[15:0]);
  assign p1_sel_141649_comb = $signed(p1_smul_57738_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57738_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57738_NarrowedMult__comb[15:0]);
  assign p1_sel_141650_comb = $signed(p1_smul_57740_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57740_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57740_NarrowedMult__comb[15:0]);
  assign p1_sel_141651_comb = $signed(p1_smul_57758_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57758_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57758_NarrowedMult__comb[15:0]);
  assign p1_sel_141652_comb = $signed(p1_smul_57760_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57760_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57760_NarrowedMult__comb[15:0]);
  assign p1_sel_141653_comb = $signed(p1_smul_57762_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57762_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57762_NarrowedMult__comb[15:0]);
  assign p1_sel_141654_comb = $signed(p1_smul_57764_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57764_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57764_NarrowedMult__comb[15:0]);
  assign p1_sel_141655_comb = $signed(p1_smul_57766_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57766_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57766_NarrowedMult__comb[15:0]);
  assign p1_sel_141656_comb = $signed(p1_smul_57768_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57768_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57768_NarrowedMult__comb[15:0]);
  assign p1_sel_141657_comb = $signed(p1_smul_57770_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57770_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57770_NarrowedMult__comb[15:0]);
  assign p1_sel_141658_comb = $signed(p1_smul_57772_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57772_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57772_NarrowedMult__comb[15:0]);
  assign p1_sel_141659_comb = $signed(p1_smul_57774_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57774_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57774_NarrowedMult__comb[15:0]);
  assign p1_sel_141660_comb = $signed(p1_smul_57776_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57776_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57776_NarrowedMult__comb[15:0]);
  assign p1_sel_141661_comb = $signed(p1_smul_57778_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57778_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57778_NarrowedMult__comb[15:0]);
  assign p1_sel_141662_comb = $signed(p1_smul_57780_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57780_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57780_NarrowedMult__comb[15:0]);
  assign p1_sel_141663_comb = $signed(p1_smul_57782_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57782_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57782_NarrowedMult__comb[15:0]);
  assign p1_sel_141664_comb = $signed(p1_smul_57784_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57784_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57784_NarrowedMult__comb[15:0]);
  assign p1_sel_141665_comb = $signed(p1_smul_57786_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57786_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57786_NarrowedMult__comb[15:0]);
  assign p1_sel_141666_comb = $signed(p1_smul_57788_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57788_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57788_NarrowedMult__comb[15:0]);
  assign p1_sel_141667_comb = $signed(p1_smul_57806_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57806_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57806_NarrowedMult__comb[15:0]);
  assign p1_sel_141668_comb = $signed(p1_smul_57808_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57808_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57808_NarrowedMult__comb[15:0]);
  assign p1_sel_141669_comb = $signed(p1_smul_57810_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57810_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57810_NarrowedMult__comb[15:0]);
  assign p1_sel_141670_comb = $signed(p1_smul_57812_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57812_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57812_NarrowedMult__comb[15:0]);
  assign p1_sel_141671_comb = $signed(p1_smul_57814_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57814_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57814_NarrowedMult__comb[15:0]);
  assign p1_sel_141672_comb = $signed(p1_smul_57816_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57816_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57816_NarrowedMult__comb[15:0]);
  assign p1_sel_141673_comb = $signed(p1_smul_57818_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57818_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57818_NarrowedMult__comb[15:0]);
  assign p1_sel_141674_comb = $signed(p1_smul_57820_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57820_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57820_NarrowedMult__comb[15:0]);
  assign p1_sel_141675_comb = $signed(p1_smul_57822_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57822_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57822_NarrowedMult__comb[15:0]);
  assign p1_sel_141676_comb = $signed(p1_smul_57824_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57824_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57824_NarrowedMult__comb[15:0]);
  assign p1_sel_141677_comb = $signed(p1_smul_57826_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57826_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57826_NarrowedMult__comb[15:0]);
  assign p1_sel_141678_comb = $signed(p1_smul_57828_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57828_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57828_NarrowedMult__comb[15:0]);
  assign p1_sel_141679_comb = $signed(p1_smul_57830_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57830_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57830_NarrowedMult__comb[15:0]);
  assign p1_sel_141680_comb = $signed(p1_smul_57832_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57832_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57832_NarrowedMult__comb[15:0]);
  assign p1_sel_141681_comb = $signed(p1_smul_57834_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57834_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57834_NarrowedMult__comb[15:0]);
  assign p1_sel_141682_comb = $signed(p1_smul_57836_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57836_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57836_NarrowedMult__comb[15:0]);
  assign p1_sel_141683_comb = $signed(p1_or_136645_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__40_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136645_comb[23:9], 1'h0};
  assign p1_sel_141684_comb = $signed(p1_smul_57840_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57840_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57840_NarrowedMult__comb[15:0]);
  assign p1_sel_141685_comb = $signed(p1_or_137776_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137776_comb[23:9], 1'h0};
  assign p1_sel_141686_comb = $signed(p1_smul_57844_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57844_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57844_NarrowedMult__comb[15:0]);
  assign p1_sel_141687_comb = $signed(p1_smul_57846_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57846_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57846_NarrowedMult__comb[15:0]);
  assign p1_sel_141688_comb = $signed(p1_or_137781_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137781_comb[23:9], 1'h0};
  assign p1_sel_141689_comb = $signed(p1_smul_57850_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57850_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57850_NarrowedMult__comb[15:0]);
  assign p1_sel_141690_comb = $signed(p1_or_136656_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__47_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136656_comb[23:9], 1'h0};
  assign p1_sel_141691_comb = $signed(p1_or_136659_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__84_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136659_comb[23:9], 1'h0};
  assign p1_sel_141692_comb = $signed(p1_smul_57856_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57856_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57856_NarrowedMult__comb[15:0]);
  assign p1_sel_141693_comb = $signed(p1_or_137792_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137792_comb[23:9], 1'h0};
  assign p1_sel_141694_comb = $signed(p1_smul_57860_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57860_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57860_NarrowedMult__comb[15:0]);
  assign p1_sel_141695_comb = $signed(p1_smul_57862_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57862_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57862_NarrowedMult__comb[15:0]);
  assign p1_sel_141696_comb = $signed(p1_or_137797_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137797_comb[23:9], 1'h0};
  assign p1_sel_141697_comb = $signed(p1_smul_57866_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57866_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57866_NarrowedMult__comb[15:0]);
  assign p1_sel_141698_comb = $signed(p1_or_136670_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__122_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136670_comb[23:9], 1'h0};
  assign p1_sel_141699_comb = $signed(p1_or_136673_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__212_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136673_comb[23:9], 1'h0};
  assign p1_sel_141700_comb = $signed(p1_smul_57888_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57888_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57888_NarrowedMult__comb[15:0]);
  assign p1_sel_141701_comb = $signed(p1_or_137808_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137808_comb[23:9], 1'h0};
  assign p1_sel_141702_comb = $signed(p1_smul_57892_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57892_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57892_NarrowedMult__comb[15:0]);
  assign p1_sel_141703_comb = $signed(p1_smul_57894_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57894_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57894_NarrowedMult__comb[15:0]);
  assign p1_sel_141704_comb = $signed(p1_or_137813_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137813_comb[23:9], 1'h0};
  assign p1_sel_141705_comb = $signed(p1_smul_57898_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57898_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57898_NarrowedMult__comb[15:0]);
  assign p1_sel_141706_comb = $signed(p1_or_136684_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__250_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136684_comb[23:9], 1'h0};
  assign p1_sel_141707_comb = $signed(p1_or_136687_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__276_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136687_comb[23:9], 1'h0};
  assign p1_sel_141708_comb = $signed(p1_smul_57904_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57904_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57904_NarrowedMult__comb[15:0]);
  assign p1_sel_141709_comb = $signed(p1_or_137824_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137824_comb[23:9], 1'h0};
  assign p1_sel_141710_comb = $signed(p1_smul_57908_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57908_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57908_NarrowedMult__comb[15:0]);
  assign p1_sel_141711_comb = $signed(p1_smul_57910_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57910_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57910_NarrowedMult__comb[15:0]);
  assign p1_sel_141712_comb = $signed(p1_or_137829_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137829_comb[23:9], 1'h0};
  assign p1_sel_141713_comb = $signed(p1_smul_57914_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57914_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57914_NarrowedMult__comb[15:0]);
  assign p1_sel_141714_comb = $signed(p1_or_136698_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__314_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136698_comb[23:9], 1'h0};
  assign p1_sel_141715_comb = $signed(p1_or_136701_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__404_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136701_comb[23:9], 1'h0};
  assign p1_sel_141716_comb = $signed(p1_smul_57936_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57936_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57936_NarrowedMult__comb[15:0]);
  assign p1_sel_141717_comb = $signed(p1_or_137840_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137840_comb[23:9], 1'h0};
  assign p1_sel_141718_comb = $signed(p1_smul_57940_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57940_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57940_NarrowedMult__comb[15:0]);
  assign p1_sel_141719_comb = $signed(p1_smul_57942_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57942_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57942_NarrowedMult__comb[15:0]);
  assign p1_sel_141720_comb = $signed(p1_or_137845_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137845_comb[23:9], 1'h0};
  assign p1_sel_141721_comb = $signed(p1_smul_57946_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57946_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57946_NarrowedMult__comb[15:0]);
  assign p1_sel_141722_comb = $signed(p1_or_136712_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__442_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136712_comb[23:9], 1'h0};
  assign p1_sel_141723_comb = $signed(p1_or_136715_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__468_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136715_comb[23:9], 1'h0};
  assign p1_sel_141724_comb = $signed(p1_smul_57952_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57952_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57952_NarrowedMult__comb[15:0]);
  assign p1_sel_141725_comb = $signed(p1_or_137856_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137856_comb[23:9], 1'h0};
  assign p1_sel_141726_comb = $signed(p1_smul_57956_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57956_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57956_NarrowedMult__comb[15:0]);
  assign p1_sel_141727_comb = $signed(p1_smul_57958_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57958_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57958_NarrowedMult__comb[15:0]);
  assign p1_sel_141728_comb = $signed(p1_or_137861_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137861_comb[23:9], 1'h0};
  assign p1_sel_141729_comb = $signed(p1_smul_57962_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_57962_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_57962_NarrowedMult__comb[15:0]);
  assign p1_sel_141730_comb = $signed(p1_or_136726_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__506_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136726_comb[23:9], 1'h0};
  assign p1_sel_141731_comb = $signed(p1_prod__48_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__48_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57966_NarrowedMult__comb, 1'h0};
  assign p1_sel_141732_comb = $signed(p1_or_136731_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__49_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136731_comb[23:10], 2'h0};
  assign p1_sel_141733_comb = $signed(p1_prod__50_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__50_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57970_NarrowedMult__comb, 1'h0};
  assign p1_sel_141734_comb = $signed(p1_or_136736_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__51_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136736_comb[23:10], 2'h0};
  assign p1_sel_141735_comb = $signed(p1_or_136739_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__52_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136739_comb[23:10], 2'h0};
  assign p1_sel_141736_comb = $signed(p1_prod__53_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__53_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57976_NarrowedMult__comb, 1'h0};
  assign p1_sel_141737_comb = $signed(p1_or_136744_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__54_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136744_comb[23:10], 2'h0};
  assign p1_sel_141738_comb = $signed(p1_prod__55_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__55_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57980_NarrowedMult__comb, 1'h0};
  assign p1_sel_141739_comb = $signed(p1_prod__91_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__91_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57982_NarrowedMult__comb, 1'h0};
  assign p1_sel_141740_comb = $signed(p1_or_136751_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__98_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136751_comb[23:10], 2'h0};
  assign p1_sel_141741_comb = $signed(p1_prod__105_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__105_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57986_NarrowedMult__comb, 1'h0};
  assign p1_sel_141742_comb = $signed(p1_or_136756_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__111_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136756_comb[23:10], 2'h0};
  assign p1_sel_141743_comb = $signed(p1_or_136759_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__116_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136759_comb[23:10], 2'h0};
  assign p1_sel_141744_comb = $signed(p1_prod__120_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__120_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57992_NarrowedMult__comb, 1'h0};
  assign p1_sel_141745_comb = $signed(p1_or_136764_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__123_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136764_comb[23:10], 2'h0};
  assign p1_sel_141746_comb = $signed(p1_prod__125_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__125_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_57996_NarrowedMult__comb, 1'h0};
  assign p1_sel_141747_comb = $signed(p1_prod__219_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__219_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58014_NarrowedMult__comb, 1'h0};
  assign p1_sel_141748_comb = $signed(p1_or_136771_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__226_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136771_comb[23:10], 2'h0};
  assign p1_sel_141749_comb = $signed(p1_prod__233_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__233_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58018_NarrowedMult__comb, 1'h0};
  assign p1_sel_141750_comb = $signed(p1_or_136776_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__239_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136776_comb[23:10], 2'h0};
  assign p1_sel_141751_comb = $signed(p1_or_136779_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__244_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136779_comb[23:10], 2'h0};
  assign p1_sel_141752_comb = $signed(p1_prod__248_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__248_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58024_NarrowedMult__comb, 1'h0};
  assign p1_sel_141753_comb = $signed(p1_or_136784_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__251_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136784_comb[23:10], 2'h0};
  assign p1_sel_141754_comb = $signed(p1_prod__253_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__253_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58028_NarrowedMult__comb, 1'h0};
  assign p1_sel_141755_comb = $signed(p1_prod__283_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__283_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58030_NarrowedMult__comb, 1'h0};
  assign p1_sel_141756_comb = $signed(p1_or_136791_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__290_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136791_comb[23:10], 2'h0};
  assign p1_sel_141757_comb = $signed(p1_prod__297_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__297_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58034_NarrowedMult__comb, 1'h0};
  assign p1_sel_141758_comb = $signed(p1_or_136796_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__303_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136796_comb[23:10], 2'h0};
  assign p1_sel_141759_comb = $signed(p1_or_136799_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__308_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136799_comb[23:10], 2'h0};
  assign p1_sel_141760_comb = $signed(p1_prod__312_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__312_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58040_NarrowedMult__comb, 1'h0};
  assign p1_sel_141761_comb = $signed(p1_or_136804_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__315_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136804_comb[23:10], 2'h0};
  assign p1_sel_141762_comb = $signed(p1_prod__317_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__317_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58044_NarrowedMult__comb, 1'h0};
  assign p1_sel_141763_comb = $signed(p1_prod__411_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__411_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58062_NarrowedMult__comb, 1'h0};
  assign p1_sel_141764_comb = $signed(p1_or_136811_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__418_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136811_comb[23:10], 2'h0};
  assign p1_sel_141765_comb = $signed(p1_prod__425_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__425_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58066_NarrowedMult__comb, 1'h0};
  assign p1_sel_141766_comb = $signed(p1_or_136816_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__431_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136816_comb[23:10], 2'h0};
  assign p1_sel_141767_comb = $signed(p1_or_136819_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__436_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136819_comb[23:10], 2'h0};
  assign p1_sel_141768_comb = $signed(p1_prod__440_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__440_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58072_NarrowedMult__comb, 1'h0};
  assign p1_sel_141769_comb = $signed(p1_or_136824_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__443_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136824_comb[23:10], 2'h0};
  assign p1_sel_141770_comb = $signed(p1_prod__445_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__445_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58076_NarrowedMult__comb, 1'h0};
  assign p1_sel_141771_comb = $signed(p1_prod__475_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__475_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58078_NarrowedMult__comb, 1'h0};
  assign p1_sel_141772_comb = $signed(p1_or_136831_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__482_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136831_comb[23:10], 2'h0};
  assign p1_sel_141773_comb = $signed(p1_prod__489_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__489_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58082_NarrowedMult__comb, 1'h0};
  assign p1_sel_141774_comb = $signed(p1_or_136836_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__495_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136836_comb[23:10], 2'h0};
  assign p1_sel_141775_comb = $signed(p1_or_136839_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__500_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136839_comb[23:10], 2'h0};
  assign p1_sel_141776_comb = $signed(p1_prod__504_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__504_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58088_NarrowedMult__comb, 1'h0};
  assign p1_sel_141777_comb = $signed(p1_or_136844_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__507_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_136844_comb[23:10], 2'h0};
  assign p1_sel_141778_comb = $signed(p1_prod__509_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__509_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58092_NarrowedMult__comb, 1'h0};
  assign p1_sel_141779_comb = $signed(p1_or_137987_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_137987_comb[23:9], 1'h0};
  assign p1_sel_141780_comb = $signed(p1_or_136851_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__57_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136851_comb[23:9], 1'h0};
  assign p1_sel_141781_comb = $signed(p1_smul_58098_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58098_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58098_NarrowedMult__comb[15:0]);
  assign p1_sel_141782_comb = $signed(p1_smul_58100_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58100_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58100_NarrowedMult__comb[15:0]);
  assign p1_sel_141783_comb = $signed(p1_smul_58102_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58102_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58102_NarrowedMult__comb[15:0]);
  assign p1_sel_141784_comb = $signed(p1_smul_58104_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58104_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58104_NarrowedMult__comb[15:0]);
  assign p1_sel_141785_comb = $signed(p1_or_136858_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__62_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136858_comb[23:9], 1'h0};
  assign p1_sel_141786_comb = $signed(p1_or_138002_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138002_comb[23:9], 1'h0};
  assign p1_sel_141787_comb = $signed(p1_or_138003_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138003_comb[23:9], 1'h0};
  assign p1_sel_141788_comb = $signed(p1_or_136865_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__106_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136865_comb[23:9], 1'h0};
  assign p1_sel_141789_comb = $signed(p1_smul_58114_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58114_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58114_NarrowedMult__comb[15:0]);
  assign p1_sel_141790_comb = $signed(p1_smul_58116_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58116_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58116_NarrowedMult__comb[15:0]);
  assign p1_sel_141791_comb = $signed(p1_smul_58118_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58118_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58118_NarrowedMult__comb[15:0]);
  assign p1_sel_141792_comb = $signed(p1_smul_58120_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58120_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58120_NarrowedMult__comb[15:0]);
  assign p1_sel_141793_comb = $signed(p1_or_136872_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__126_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136872_comb[23:9], 1'h0};
  assign p1_sel_141794_comb = $signed(p1_or_138018_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138018_comb[23:9], 1'h0};
  assign p1_sel_141795_comb = $signed(p1_or_138019_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138019_comb[23:9], 1'h0};
  assign p1_sel_141796_comb = $signed(p1_or_136879_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__234_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136879_comb[23:9], 1'h0};
  assign p1_sel_141797_comb = $signed(p1_smul_58146_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58146_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58146_NarrowedMult__comb[15:0]);
  assign p1_sel_141798_comb = $signed(p1_smul_58148_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58148_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58148_NarrowedMult__comb[15:0]);
  assign p1_sel_141799_comb = $signed(p1_smul_58150_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58150_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58150_NarrowedMult__comb[15:0]);
  assign p1_sel_141800_comb = $signed(p1_smul_58152_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58152_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58152_NarrowedMult__comb[15:0]);
  assign p1_sel_141801_comb = $signed(p1_or_136886_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__254_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136886_comb[23:9], 1'h0};
  assign p1_sel_141802_comb = $signed(p1_or_138034_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138034_comb[23:9], 1'h0};
  assign p1_sel_141803_comb = $signed(p1_or_138035_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138035_comb[23:9], 1'h0};
  assign p1_sel_141804_comb = $signed(p1_or_136893_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__298_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136893_comb[23:9], 1'h0};
  assign p1_sel_141805_comb = $signed(p1_smul_58162_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58162_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58162_NarrowedMult__comb[15:0]);
  assign p1_sel_141806_comb = $signed(p1_smul_58164_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58164_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58164_NarrowedMult__comb[15:0]);
  assign p1_sel_141807_comb = $signed(p1_smul_58166_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58166_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58166_NarrowedMult__comb[15:0]);
  assign p1_sel_141808_comb = $signed(p1_smul_58168_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58168_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58168_NarrowedMult__comb[15:0]);
  assign p1_sel_141809_comb = $signed(p1_or_136900_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__318_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136900_comb[23:9], 1'h0};
  assign p1_sel_141810_comb = $signed(p1_or_138050_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138050_comb[23:9], 1'h0};
  assign p1_sel_141811_comb = $signed(p1_or_138051_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138051_comb[23:9], 1'h0};
  assign p1_sel_141812_comb = $signed(p1_or_136907_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__426_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136907_comb[23:9], 1'h0};
  assign p1_sel_141813_comb = $signed(p1_smul_58194_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58194_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58194_NarrowedMult__comb[15:0]);
  assign p1_sel_141814_comb = $signed(p1_smul_58196_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58196_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58196_NarrowedMult__comb[15:0]);
  assign p1_sel_141815_comb = $signed(p1_smul_58198_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58198_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58198_NarrowedMult__comb[15:0]);
  assign p1_sel_141816_comb = $signed(p1_smul_58200_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58200_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58200_NarrowedMult__comb[15:0]);
  assign p1_sel_141817_comb = $signed(p1_or_136914_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__446_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136914_comb[23:9], 1'h0};
  assign p1_sel_141818_comb = $signed(p1_or_138066_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138066_comb[23:9], 1'h0};
  assign p1_sel_141819_comb = $signed(p1_or_138067_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138067_comb[23:9], 1'h0};
  assign p1_sel_141820_comb = $signed(p1_or_136921_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__490_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136921_comb[23:9], 1'h0};
  assign p1_sel_141821_comb = $signed(p1_smul_58210_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58210_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58210_NarrowedMult__comb[15:0]);
  assign p1_sel_141822_comb = $signed(p1_smul_58212_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58212_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58212_NarrowedMult__comb[15:0]);
  assign p1_sel_141823_comb = $signed(p1_smul_58214_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58214_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58214_NarrowedMult__comb[15:0]);
  assign p1_sel_141824_comb = $signed(p1_smul_58216_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58216_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58216_NarrowedMult__comb[15:0]);
  assign p1_sel_141825_comb = $signed(p1_or_136928_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__510_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_136928_comb[23:9], 1'h0};
  assign p1_sel_141826_comb = $signed(p1_or_138082_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_138082_comb[23:9], 1'h0};
  assign p1_sum__989_comb = {{15{p1_add_141347_comb[16]}}, p1_add_141347_comb};
  assign p1_sum__990_comb = {{15{p1_add_141348_comb[16]}}, p1_add_141348_comb};
  assign p1_sum__991_comb = {{15{p1_add_141349_comb[16]}}, p1_add_141349_comb};
  assign p1_sum__992_comb = {{15{p1_add_141350_comb[16]}}, p1_add_141350_comb};
  assign p1_sum__884_comb = {{15{p1_add_141351_comb[16]}}, p1_add_141351_comb};
  assign p1_sum__885_comb = {{15{p1_add_141352_comb[16]}}, p1_add_141352_comb};
  assign p1_sum__886_comb = {{15{p1_add_141353_comb[16]}}, p1_add_141353_comb};
  assign p1_sum__887_comb = {{15{p1_add_141354_comb[16]}}, p1_add_141354_comb};
  assign p1_sum__1017_comb = {{15{p1_add_141467_comb[16]}}, p1_add_141467_comb};
  assign p1_sum__1018_comb = {{15{p1_add_141468_comb[16]}}, p1_add_141468_comb};
  assign p1_sum__1019_comb = {{15{p1_add_141469_comb[16]}}, p1_add_141469_comb};
  assign p1_sum__1020_comb = {{15{p1_add_141470_comb[16]}}, p1_add_141470_comb};
  assign p1_sum__1010_comb = {{15{p1_add_141471_comb[16]}}, p1_add_141471_comb};
  assign p1_sum__1011_comb = {{15{p1_add_141472_comb[16]}}, p1_add_141472_comb};
  assign p1_sum__1012_comb = {{15{p1_add_141473_comb[16]}}, p1_add_141473_comb};
  assign p1_sum__1013_comb = {{15{p1_add_141474_comb[16]}}, p1_add_141474_comb};
  assign p1_sum__961_comb = {{15{p1_add_141475_comb[16]}}, p1_add_141475_comb};
  assign p1_sum__962_comb = {{15{p1_add_141476_comb[16]}}, p1_add_141476_comb};
  assign p1_sum__963_comb = {{15{p1_add_141477_comb[16]}}, p1_add_141477_comb};
  assign p1_sum__964_comb = {{15{p1_add_141478_comb[16]}}, p1_add_141478_comb};
  assign p1_sum__926_comb = {{15{p1_add_141479_comb[16]}}, p1_add_141479_comb};
  assign p1_sum__927_comb = {{15{p1_add_141480_comb[16]}}, p1_add_141480_comb};
  assign p1_sum__928_comb = {{15{p1_add_141481_comb[16]}}, p1_add_141481_comb};
  assign p1_sum__929_comb = {{15{p1_add_141482_comb[16]}}, p1_add_141482_comb};
  assign p1_sum__835_comb = {{15{p1_add_141483_comb[16]}}, p1_add_141483_comb};
  assign p1_sum__836_comb = {{15{p1_add_141484_comb[16]}}, p1_add_141484_comb};
  assign p1_sum__837_comb = {{15{p1_add_141485_comb[16]}}, p1_add_141485_comb};
  assign p1_sum__838_comb = {{15{p1_add_141486_comb[16]}}, p1_add_141486_comb};
  assign p1_sum__779_comb = {{15{p1_add_141487_comb[16]}}, p1_add_141487_comb};
  assign p1_sum__780_comb = {{15{p1_add_141488_comb[16]}}, p1_add_141488_comb};
  assign p1_sum__781_comb = {{15{p1_add_141489_comb[16]}}, p1_add_141489_comb};
  assign p1_sum__782_comb = {{15{p1_add_141490_comb[16]}}, p1_add_141490_comb};
  assign p1_sum__993_comb = p1_sum__989_comb + p1_sum__990_comb;
  assign p1_sum__994_comb = p1_sum__991_comb + p1_sum__992_comb;
  assign p1_sum__888_comb = p1_sum__884_comb + p1_sum__885_comb;
  assign p1_sum__889_comb = p1_sum__886_comb + p1_sum__887_comb;
  assign p1_add_142311_comb = {{1{p1_sel_141355_comb[15]}}, p1_sel_141355_comb} + {{1{p1_sel_141356_comb[15]}}, p1_sel_141356_comb};
  assign p1_add_142312_comb = {{1{p1_sel_141357_comb[15]}}, p1_sel_141357_comb} + {{1{p1_sel_141358_comb[15]}}, p1_sel_141358_comb};
  assign p1_add_142313_comb = {{1{p1_sel_141359_comb[15]}}, p1_sel_141359_comb} + {{1{p1_sel_141360_comb[15]}}, p1_sel_141360_comb};
  assign p1_add_142314_comb = {{1{p1_sel_141361_comb[15]}}, p1_sel_141361_comb} + {{1{p1_sel_141362_comb[15]}}, p1_sel_141362_comb};
  assign p1_add_142315_comb = {{1{p1_sel_141363_comb[15]}}, p1_sel_141363_comb} + {{1{p1_sel_141364_comb[15]}}, p1_sel_141364_comb};
  assign p1_add_142316_comb = {{1{p1_sel_141365_comb[15]}}, p1_sel_141365_comb} + {{1{p1_sel_141366_comb[15]}}, p1_sel_141366_comb};
  assign p1_add_142317_comb = {{1{p1_sel_141367_comb[15]}}, p1_sel_141367_comb} + {{1{p1_sel_141368_comb[15]}}, p1_sel_141368_comb};
  assign p1_add_142318_comb = {{1{p1_sel_141369_comb[15]}}, p1_sel_141369_comb} + {{1{p1_sel_141370_comb[15]}}, p1_sel_141370_comb};
  assign p1_add_142319_comb = {{1{p1_sel_141371_comb[15]}}, p1_sel_141371_comb} + {{1{p1_sel_141372_comb[15]}}, p1_sel_141372_comb};
  assign p1_add_142320_comb = {{1{p1_sel_141373_comb[15]}}, p1_sel_141373_comb} + {{1{p1_sel_141374_comb[15]}}, p1_sel_141374_comb};
  assign p1_add_142321_comb = {{1{p1_sel_141375_comb[15]}}, p1_sel_141375_comb} + {{1{p1_sel_141376_comb[15]}}, p1_sel_141376_comb};
  assign p1_add_142322_comb = {{1{p1_sel_141377_comb[15]}}, p1_sel_141377_comb} + {{1{p1_sel_141378_comb[15]}}, p1_sel_141378_comb};
  assign p1_add_142323_comb = {{1{p1_sel_141379_comb[15]}}, p1_sel_141379_comb} + {{1{p1_sel_141380_comb[15]}}, p1_sel_141380_comb};
  assign p1_add_142324_comb = {{1{p1_sel_141381_comb[15]}}, p1_sel_141381_comb} + {{1{p1_sel_141382_comb[15]}}, p1_sel_141382_comb};
  assign p1_add_142325_comb = {{1{p1_sel_141383_comb[15]}}, p1_sel_141383_comb} + {{1{p1_sel_141384_comb[15]}}, p1_sel_141384_comb};
  assign p1_add_142326_comb = {{1{p1_sel_141385_comb[15]}}, p1_sel_141385_comb} + {{1{p1_sel_141386_comb[15]}}, p1_sel_141386_comb};
  assign p1_add_142327_comb = {{1{p1_sel_141387_comb[15]}}, p1_sel_141387_comb} + {{1{p1_sel_141388_comb[15]}}, p1_sel_141388_comb};
  assign p1_add_142328_comb = {{1{p1_sel_141389_comb[15]}}, p1_sel_141389_comb} + {{1{p1_sel_141390_comb[15]}}, p1_sel_141390_comb};
  assign p1_add_142329_comb = {{1{p1_sel_141391_comb[15]}}, p1_sel_141391_comb} + {{1{p1_sel_141392_comb[15]}}, p1_sel_141392_comb};
  assign p1_add_142330_comb = {{1{p1_sel_141393_comb[15]}}, p1_sel_141393_comb} + {{1{p1_sel_141394_comb[15]}}, p1_sel_141394_comb};
  assign p1_add_142331_comb = {{1{p1_sel_141395_comb[15]}}, p1_sel_141395_comb} + {{1{p1_sel_141396_comb[15]}}, p1_sel_141396_comb};
  assign p1_add_142332_comb = {{1{p1_sel_141397_comb[15]}}, p1_sel_141397_comb} + {{1{p1_sel_141398_comb[15]}}, p1_sel_141398_comb};
  assign p1_add_142333_comb = {{1{p1_sel_141399_comb[15]}}, p1_sel_141399_comb} + {{1{p1_sel_141400_comb[15]}}, p1_sel_141400_comb};
  assign p1_add_142334_comb = {{1{p1_sel_141401_comb[15]}}, p1_sel_141401_comb} + {{1{p1_sel_141402_comb[15]}}, p1_sel_141402_comb};
  assign p1_add_142335_comb = {{1{p1_sel_141403_comb[15]}}, p1_sel_141403_comb} + {{1{p1_sel_141404_comb[15]}}, p1_sel_141404_comb};
  assign p1_add_142336_comb = {{1{p1_sel_141405_comb[15]}}, p1_sel_141405_comb} + {{1{p1_sel_141406_comb[15]}}, p1_sel_141406_comb};
  assign p1_add_142337_comb = {{1{p1_sel_141407_comb[15]}}, p1_sel_141407_comb} + {{1{p1_sel_141408_comb[15]}}, p1_sel_141408_comb};
  assign p1_add_142338_comb = {{1{p1_sel_141409_comb[15]}}, p1_sel_141409_comb} + {{1{p1_sel_141410_comb[15]}}, p1_sel_141410_comb};
  assign p1_add_142339_comb = {{1{p1_sel_141411_comb[15]}}, p1_sel_141411_comb} + {{1{p1_sel_141412_comb[15]}}, p1_sel_141412_comb};
  assign p1_add_142340_comb = {{1{p1_sel_141413_comb[15]}}, p1_sel_141413_comb} + {{1{p1_sel_141414_comb[15]}}, p1_sel_141414_comb};
  assign p1_add_142341_comb = {{1{p1_sel_141415_comb[15]}}, p1_sel_141415_comb} + {{1{p1_sel_141416_comb[15]}}, p1_sel_141416_comb};
  assign p1_add_142342_comb = {{1{p1_sel_141417_comb[15]}}, p1_sel_141417_comb} + {{1{p1_sel_141418_comb[15]}}, p1_sel_141418_comb};
  assign p1_add_142343_comb = {{1{p1_sel_141419_comb[15]}}, p1_sel_141419_comb} + {{1{p1_sel_141420_comb[15]}}, p1_sel_141420_comb};
  assign p1_add_142344_comb = {{1{p1_sel_141421_comb[15]}}, p1_sel_141421_comb} + {{1{p1_sel_141422_comb[15]}}, p1_sel_141422_comb};
  assign p1_add_142345_comb = {{1{p1_sel_141423_comb[15]}}, p1_sel_141423_comb} + {{1{p1_sel_141424_comb[15]}}, p1_sel_141424_comb};
  assign p1_add_142346_comb = {{1{p1_sel_141425_comb[15]}}, p1_sel_141425_comb} + {{1{p1_sel_141426_comb[15]}}, p1_sel_141426_comb};
  assign p1_add_142347_comb = {{1{p1_sel_141427_comb[15]}}, p1_sel_141427_comb} + {{1{p1_sel_141428_comb[15]}}, p1_sel_141428_comb};
  assign p1_add_142348_comb = {{1{p1_sel_141429_comb[15]}}, p1_sel_141429_comb} + {{1{p1_sel_141430_comb[15]}}, p1_sel_141430_comb};
  assign p1_add_142349_comb = {{1{p1_sel_141431_comb[15]}}, p1_sel_141431_comb} + {{1{p1_sel_141432_comb[15]}}, p1_sel_141432_comb};
  assign p1_add_142350_comb = {{1{p1_sel_141433_comb[15]}}, p1_sel_141433_comb} + {{1{p1_sel_141434_comb[15]}}, p1_sel_141434_comb};
  assign p1_add_142351_comb = {{1{p1_sel_141435_comb[15]}}, p1_sel_141435_comb} + {{1{p1_sel_141436_comb[15]}}, p1_sel_141436_comb};
  assign p1_add_142352_comb = {{1{p1_sel_141437_comb[15]}}, p1_sel_141437_comb} + {{1{p1_sel_141438_comb[15]}}, p1_sel_141438_comb};
  assign p1_add_142353_comb = {{1{p1_sel_141439_comb[15]}}, p1_sel_141439_comb} + {{1{p1_sel_141440_comb[15]}}, p1_sel_141440_comb};
  assign p1_add_142354_comb = {{1{p1_sel_141441_comb[15]}}, p1_sel_141441_comb} + {{1{p1_sel_141442_comb[15]}}, p1_sel_141442_comb};
  assign p1_add_142355_comb = {{1{p1_sel_141443_comb[15]}}, p1_sel_141443_comb} + {{1{p1_sel_141444_comb[15]}}, p1_sel_141444_comb};
  assign p1_add_142356_comb = {{1{p1_sel_141445_comb[15]}}, p1_sel_141445_comb} + {{1{p1_sel_141446_comb[15]}}, p1_sel_141446_comb};
  assign p1_add_142357_comb = {{1{p1_sel_141447_comb[15]}}, p1_sel_141447_comb} + {{1{p1_sel_141448_comb[15]}}, p1_sel_141448_comb};
  assign p1_add_142358_comb = {{1{p1_sel_141449_comb[15]}}, p1_sel_141449_comb} + {{1{p1_sel_141450_comb[15]}}, p1_sel_141450_comb};
  assign p1_add_142359_comb = {{1{p1_sel_141451_comb[15]}}, p1_sel_141451_comb} + {{1{p1_sel_141452_comb[15]}}, p1_sel_141452_comb};
  assign p1_add_142360_comb = {{1{p1_sel_141453_comb[15]}}, p1_sel_141453_comb} + {{1{p1_sel_141454_comb[15]}}, p1_sel_141454_comb};
  assign p1_add_142361_comb = {{1{p1_sel_141455_comb[15]}}, p1_sel_141455_comb} + {{1{p1_sel_141456_comb[15]}}, p1_sel_141456_comb};
  assign p1_add_142362_comb = {{1{p1_sel_141457_comb[15]}}, p1_sel_141457_comb} + {{1{p1_sel_141458_comb[15]}}, p1_sel_141458_comb};
  assign p1_add_142363_comb = {{1{p1_sel_141459_comb[15]}}, p1_sel_141459_comb} + {{1{p1_sel_141460_comb[15]}}, p1_sel_141460_comb};
  assign p1_add_142364_comb = {{1{p1_sel_141461_comb[15]}}, p1_sel_141461_comb} + {{1{p1_sel_141462_comb[15]}}, p1_sel_141462_comb};
  assign p1_add_142365_comb = {{1{p1_sel_141463_comb[15]}}, p1_sel_141463_comb} + {{1{p1_sel_141464_comb[15]}}, p1_sel_141464_comb};
  assign p1_add_142366_comb = {{1{p1_sel_141465_comb[15]}}, p1_sel_141465_comb} + {{1{p1_sel_141466_comb[15]}}, p1_sel_141466_comb};
  assign p1_sum__1021_comb = p1_sum__1017_comb + p1_sum__1018_comb;
  assign p1_sum__1022_comb = p1_sum__1019_comb + p1_sum__1020_comb;
  assign p1_sum__1014_comb = p1_sum__1010_comb + p1_sum__1011_comb;
  assign p1_sum__1015_comb = p1_sum__1012_comb + p1_sum__1013_comb;
  assign p1_sum__965_comb = p1_sum__961_comb + p1_sum__962_comb;
  assign p1_sum__966_comb = p1_sum__963_comb + p1_sum__964_comb;
  assign p1_sum__930_comb = p1_sum__926_comb + p1_sum__927_comb;
  assign p1_sum__931_comb = p1_sum__928_comb + p1_sum__929_comb;
  assign p1_sum__839_comb = p1_sum__835_comb + p1_sum__836_comb;
  assign p1_sum__840_comb = p1_sum__837_comb + p1_sum__838_comb;
  assign p1_sum__783_comb = p1_sum__779_comb + p1_sum__780_comb;
  assign p1_sum__784_comb = p1_sum__781_comb + p1_sum__782_comb;
  assign p1_add_142379_comb = {{1{p1_sel_141491_comb[15]}}, p1_sel_141491_comb} + {{1{p1_sel_141492_comb[15]}}, p1_sel_141492_comb};
  assign p1_add_142380_comb = {{1{p1_sel_141493_comb[15]}}, p1_sel_141493_comb} + {{1{p1_sel_141494_comb[15]}}, p1_sel_141494_comb};
  assign p1_add_142381_comb = {{1{p1_sel_141495_comb[15]}}, p1_sel_141495_comb} + {{1{p1_sel_141496_comb[15]}}, p1_sel_141496_comb};
  assign p1_add_142382_comb = {{1{p1_sel_141497_comb[15]}}, p1_sel_141497_comb} + {{1{p1_sel_141498_comb[15]}}, p1_sel_141498_comb};
  assign p1_add_142383_comb = {{1{p1_sel_141499_comb[15]}}, p1_sel_141499_comb} + {{1{p1_sel_141500_comb[15]}}, p1_sel_141500_comb};
  assign p1_add_142384_comb = {{1{p1_sel_141501_comb[15]}}, p1_sel_141501_comb} + {{1{p1_sel_141502_comb[15]}}, p1_sel_141502_comb};
  assign p1_add_142385_comb = {{1{p1_sel_141503_comb[15]}}, p1_sel_141503_comb} + {{1{p1_sel_141504_comb[15]}}, p1_sel_141504_comb};
  assign p1_add_142386_comb = {{1{p1_sel_141505_comb[15]}}, p1_sel_141505_comb} + {{1{p1_sel_141506_comb[15]}}, p1_sel_141506_comb};
  assign p1_add_142387_comb = {{1{p1_sel_141507_comb[15]}}, p1_sel_141507_comb} + {{1{p1_sel_141508_comb[15]}}, p1_sel_141508_comb};
  assign p1_add_142388_comb = {{1{p1_sel_141509_comb[15]}}, p1_sel_141509_comb} + {{1{p1_sel_141510_comb[15]}}, p1_sel_141510_comb};
  assign p1_add_142389_comb = {{1{p1_sel_141511_comb[15]}}, p1_sel_141511_comb} + {{1{p1_sel_141512_comb[15]}}, p1_sel_141512_comb};
  assign p1_add_142390_comb = {{1{p1_sel_141513_comb[15]}}, p1_sel_141513_comb} + {{1{p1_sel_141514_comb[15]}}, p1_sel_141514_comb};
  assign p1_add_142391_comb = {{1{p1_sel_141515_comb[15]}}, p1_sel_141515_comb} + {{1{p1_sel_141516_comb[15]}}, p1_sel_141516_comb};
  assign p1_add_142392_comb = {{1{p1_sel_141517_comb[15]}}, p1_sel_141517_comb} + {{1{p1_sel_141518_comb[15]}}, p1_sel_141518_comb};
  assign p1_add_142393_comb = {{1{p1_sel_141519_comb[15]}}, p1_sel_141519_comb} + {{1{p1_sel_141520_comb[15]}}, p1_sel_141520_comb};
  assign p1_add_142394_comb = {{1{p1_sel_141521_comb[15]}}, p1_sel_141521_comb} + {{1{p1_sel_141522_comb[15]}}, p1_sel_141522_comb};
  assign p1_add_142395_comb = {{1{p1_sel_141523_comb[15]}}, p1_sel_141523_comb} + {{1{p1_sel_141524_comb[15]}}, p1_sel_141524_comb};
  assign p1_add_142396_comb = {{1{p1_sel_141525_comb[15]}}, p1_sel_141525_comb} + {{1{p1_sel_141526_comb[15]}}, p1_sel_141526_comb};
  assign p1_add_142397_comb = {{1{p1_sel_141527_comb[15]}}, p1_sel_141527_comb} + {{1{p1_sel_141528_comb[15]}}, p1_sel_141528_comb};
  assign p1_add_142398_comb = {{1{p1_sel_141529_comb[15]}}, p1_sel_141529_comb} + {{1{p1_sel_141530_comb[15]}}, p1_sel_141530_comb};
  assign p1_add_142399_comb = {{1{p1_sel_141531_comb[15]}}, p1_sel_141531_comb} + {{1{p1_sel_141532_comb[15]}}, p1_sel_141532_comb};
  assign p1_add_142400_comb = {{1{p1_sel_141533_comb[15]}}, p1_sel_141533_comb} + {{1{p1_sel_141534_comb[15]}}, p1_sel_141534_comb};
  assign p1_add_142401_comb = {{1{p1_sel_141535_comb[15]}}, p1_sel_141535_comb} + {{1{p1_sel_141536_comb[15]}}, p1_sel_141536_comb};
  assign p1_add_142402_comb = {{1{p1_sel_141537_comb[15]}}, p1_sel_141537_comb} + {{1{p1_sel_141538_comb[15]}}, p1_sel_141538_comb};
  assign p1_add_142403_comb = {{1{p1_sel_141539_comb[15]}}, p1_sel_141539_comb} + {{1{p1_sel_141540_comb[15]}}, p1_sel_141540_comb};
  assign p1_add_142404_comb = {{1{p1_sel_141541_comb[15]}}, p1_sel_141541_comb} + {{1{p1_sel_141542_comb[15]}}, p1_sel_141542_comb};
  assign p1_add_142405_comb = {{1{p1_sel_141543_comb[15]}}, p1_sel_141543_comb} + {{1{p1_sel_141544_comb[15]}}, p1_sel_141544_comb};
  assign p1_add_142406_comb = {{1{p1_sel_141545_comb[15]}}, p1_sel_141545_comb} + {{1{p1_sel_141546_comb[15]}}, p1_sel_141546_comb};
  assign p1_add_142407_comb = {{1{p1_sel_141547_comb[15]}}, p1_sel_141547_comb} + {{1{p1_sel_141548_comb[15]}}, p1_sel_141548_comb};
  assign p1_add_142408_comb = {{1{p1_sel_141549_comb[15]}}, p1_sel_141549_comb} + {{1{p1_sel_141550_comb[15]}}, p1_sel_141550_comb};
  assign p1_add_142409_comb = {{1{p1_sel_141551_comb[15]}}, p1_sel_141551_comb} + {{1{p1_sel_141552_comb[15]}}, p1_sel_141552_comb};
  assign p1_add_142410_comb = {{1{p1_sel_141553_comb[15]}}, p1_sel_141553_comb} + {{1{p1_sel_141554_comb[15]}}, p1_sel_141554_comb};
  assign p1_add_142411_comb = {{1{p1_sel_141555_comb[15]}}, p1_sel_141555_comb} + {{1{p1_sel_141556_comb[15]}}, p1_sel_141556_comb};
  assign p1_add_142412_comb = {{1{p1_sel_141557_comb[15]}}, p1_sel_141557_comb} + {{1{p1_sel_141558_comb[15]}}, p1_sel_141558_comb};
  assign p1_add_142413_comb = {{1{p1_sel_141559_comb[15]}}, p1_sel_141559_comb} + {{1{p1_sel_141560_comb[15]}}, p1_sel_141560_comb};
  assign p1_add_142414_comb = {{1{p1_sel_141561_comb[15]}}, p1_sel_141561_comb} + {{1{p1_sel_141562_comb[15]}}, p1_sel_141562_comb};
  assign p1_add_142415_comb = {{1{p1_sel_141563_comb[15]}}, p1_sel_141563_comb} + {{1{p1_sel_141564_comb[15]}}, p1_sel_141564_comb};
  assign p1_add_142416_comb = {{1{p1_sel_141565_comb[15]}}, p1_sel_141565_comb} + {{1{p1_sel_141566_comb[15]}}, p1_sel_141566_comb};
  assign p1_add_142417_comb = {{1{p1_sel_141567_comb[15]}}, p1_sel_141567_comb} + {{1{p1_sel_141568_comb[15]}}, p1_sel_141568_comb};
  assign p1_add_142418_comb = {{1{p1_sel_141569_comb[15]}}, p1_sel_141569_comb} + {{1{p1_sel_141570_comb[15]}}, p1_sel_141570_comb};
  assign p1_add_142419_comb = {{1{p1_sel_141571_comb[15]}}, p1_sel_141571_comb} + {{1{p1_sel_141572_comb[15]}}, p1_sel_141572_comb};
  assign p1_add_142420_comb = {{1{p1_sel_141573_comb[15]}}, p1_sel_141573_comb} + {{1{p1_sel_141574_comb[15]}}, p1_sel_141574_comb};
  assign p1_add_142421_comb = {{1{p1_sel_141575_comb[15]}}, p1_sel_141575_comb} + {{1{p1_sel_141576_comb[15]}}, p1_sel_141576_comb};
  assign p1_add_142422_comb = {{1{p1_sel_141577_comb[15]}}, p1_sel_141577_comb} + {{1{p1_sel_141578_comb[15]}}, p1_sel_141578_comb};
  assign p1_add_142423_comb = {{1{p1_sel_141579_comb[15]}}, p1_sel_141579_comb} + {{1{p1_sel_141580_comb[15]}}, p1_sel_141580_comb};
  assign p1_add_142424_comb = {{1{p1_sel_141581_comb[15]}}, p1_sel_141581_comb} + {{1{p1_sel_141582_comb[15]}}, p1_sel_141582_comb};
  assign p1_add_142425_comb = {{1{p1_sel_141583_comb[15]}}, p1_sel_141583_comb} + {{1{p1_sel_141584_comb[15]}}, p1_sel_141584_comb};
  assign p1_add_142426_comb = {{1{p1_sel_141585_comb[15]}}, p1_sel_141585_comb} + {{1{p1_sel_141586_comb[15]}}, p1_sel_141586_comb};
  assign p1_add_142427_comb = {{1{p1_sel_141587_comb[15]}}, p1_sel_141587_comb} + {{1{p1_sel_141588_comb[15]}}, p1_sel_141588_comb};
  assign p1_add_142428_comb = {{1{p1_sel_141589_comb[15]}}, p1_sel_141589_comb} + {{1{p1_sel_141590_comb[15]}}, p1_sel_141590_comb};
  assign p1_add_142429_comb = {{1{p1_sel_141591_comb[15]}}, p1_sel_141591_comb} + {{1{p1_sel_141592_comb[15]}}, p1_sel_141592_comb};
  assign p1_add_142430_comb = {{1{p1_sel_141593_comb[15]}}, p1_sel_141593_comb} + {{1{p1_sel_141594_comb[15]}}, p1_sel_141594_comb};
  assign p1_add_142431_comb = {{1{p1_sel_141595_comb[15]}}, p1_sel_141595_comb} + {{1{p1_sel_141596_comb[15]}}, p1_sel_141596_comb};
  assign p1_add_142432_comb = {{1{p1_sel_141597_comb[15]}}, p1_sel_141597_comb} + {{1{p1_sel_141598_comb[15]}}, p1_sel_141598_comb};
  assign p1_add_142433_comb = {{1{p1_sel_141599_comb[15]}}, p1_sel_141599_comb} + {{1{p1_sel_141600_comb[15]}}, p1_sel_141600_comb};
  assign p1_add_142434_comb = {{1{p1_sel_141601_comb[15]}}, p1_sel_141601_comb} + {{1{p1_sel_141602_comb[15]}}, p1_sel_141602_comb};
  assign p1_add_142435_comb = {{1{p1_sel_141603_comb[15]}}, p1_sel_141603_comb} + {{1{p1_sel_141604_comb[15]}}, p1_sel_141604_comb};
  assign p1_add_142436_comb = {{1{p1_sel_141605_comb[15]}}, p1_sel_141605_comb} + {{1{p1_sel_141606_comb[15]}}, p1_sel_141606_comb};
  assign p1_add_142437_comb = {{1{p1_sel_141607_comb[15]}}, p1_sel_141607_comb} + {{1{p1_sel_141608_comb[15]}}, p1_sel_141608_comb};
  assign p1_add_142438_comb = {{1{p1_sel_141609_comb[15]}}, p1_sel_141609_comb} + {{1{p1_sel_141610_comb[15]}}, p1_sel_141610_comb};
  assign p1_add_142439_comb = {{1{p1_sel_141611_comb[15]}}, p1_sel_141611_comb} + {{1{p1_sel_141612_comb[15]}}, p1_sel_141612_comb};
  assign p1_add_142440_comb = {{1{p1_sel_141613_comb[15]}}, p1_sel_141613_comb} + {{1{p1_sel_141614_comb[15]}}, p1_sel_141614_comb};
  assign p1_add_142441_comb = {{1{p1_sel_141615_comb[15]}}, p1_sel_141615_comb} + {{1{p1_sel_141616_comb[15]}}, p1_sel_141616_comb};
  assign p1_add_142442_comb = {{1{p1_sel_141617_comb[15]}}, p1_sel_141617_comb} + {{1{p1_sel_141618_comb[15]}}, p1_sel_141618_comb};
  assign p1_add_142443_comb = {{1{p1_sel_141619_comb[15]}}, p1_sel_141619_comb} + {{1{p1_sel_141620_comb[15]}}, p1_sel_141620_comb};
  assign p1_add_142444_comb = {{1{p1_sel_141621_comb[15]}}, p1_sel_141621_comb} + {{1{p1_sel_141622_comb[15]}}, p1_sel_141622_comb};
  assign p1_add_142445_comb = {{1{p1_sel_141623_comb[15]}}, p1_sel_141623_comb} + {{1{p1_sel_141624_comb[15]}}, p1_sel_141624_comb};
  assign p1_add_142446_comb = {{1{p1_sel_141625_comb[15]}}, p1_sel_141625_comb} + {{1{p1_sel_141626_comb[15]}}, p1_sel_141626_comb};
  assign p1_add_142447_comb = {{1{p1_sel_141627_comb[15]}}, p1_sel_141627_comb} + {{1{p1_sel_141628_comb[15]}}, p1_sel_141628_comb};
  assign p1_add_142448_comb = {{1{p1_sel_141629_comb[15]}}, p1_sel_141629_comb} + {{1{p1_sel_141630_comb[15]}}, p1_sel_141630_comb};
  assign p1_add_142449_comb = {{1{p1_sel_141631_comb[15]}}, p1_sel_141631_comb} + {{1{p1_sel_141632_comb[15]}}, p1_sel_141632_comb};
  assign p1_add_142450_comb = {{1{p1_sel_141633_comb[15]}}, p1_sel_141633_comb} + {{1{p1_sel_141634_comb[15]}}, p1_sel_141634_comb};
  assign p1_add_142451_comb = {{1{p1_sel_141635_comb[15]}}, p1_sel_141635_comb} + {{1{p1_sel_141636_comb[15]}}, p1_sel_141636_comb};
  assign p1_add_142452_comb = {{1{p1_sel_141637_comb[15]}}, p1_sel_141637_comb} + {{1{p1_sel_141638_comb[15]}}, p1_sel_141638_comb};
  assign p1_add_142453_comb = {{1{p1_sel_141639_comb[15]}}, p1_sel_141639_comb} + {{1{p1_sel_141640_comb[15]}}, p1_sel_141640_comb};
  assign p1_add_142454_comb = {{1{p1_sel_141641_comb[15]}}, p1_sel_141641_comb} + {{1{p1_sel_141642_comb[15]}}, p1_sel_141642_comb};
  assign p1_add_142455_comb = {{1{p1_sel_141643_comb[15]}}, p1_sel_141643_comb} + {{1{p1_sel_141644_comb[15]}}, p1_sel_141644_comb};
  assign p1_add_142456_comb = {{1{p1_sel_141645_comb[15]}}, p1_sel_141645_comb} + {{1{p1_sel_141646_comb[15]}}, p1_sel_141646_comb};
  assign p1_add_142457_comb = {{1{p1_sel_141647_comb[15]}}, p1_sel_141647_comb} + {{1{p1_sel_141648_comb[15]}}, p1_sel_141648_comb};
  assign p1_add_142458_comb = {{1{p1_sel_141649_comb[15]}}, p1_sel_141649_comb} + {{1{p1_sel_141650_comb[15]}}, p1_sel_141650_comb};
  assign p1_add_142459_comb = {{1{p1_sel_141651_comb[15]}}, p1_sel_141651_comb} + {{1{p1_sel_141652_comb[15]}}, p1_sel_141652_comb};
  assign p1_add_142460_comb = {{1{p1_sel_141653_comb[15]}}, p1_sel_141653_comb} + {{1{p1_sel_141654_comb[15]}}, p1_sel_141654_comb};
  assign p1_add_142461_comb = {{1{p1_sel_141655_comb[15]}}, p1_sel_141655_comb} + {{1{p1_sel_141656_comb[15]}}, p1_sel_141656_comb};
  assign p1_add_142462_comb = {{1{p1_sel_141657_comb[15]}}, p1_sel_141657_comb} + {{1{p1_sel_141658_comb[15]}}, p1_sel_141658_comb};
  assign p1_add_142463_comb = {{1{p1_sel_141659_comb[15]}}, p1_sel_141659_comb} + {{1{p1_sel_141660_comb[15]}}, p1_sel_141660_comb};
  assign p1_add_142464_comb = {{1{p1_sel_141661_comb[15]}}, p1_sel_141661_comb} + {{1{p1_sel_141662_comb[15]}}, p1_sel_141662_comb};
  assign p1_add_142465_comb = {{1{p1_sel_141663_comb[15]}}, p1_sel_141663_comb} + {{1{p1_sel_141664_comb[15]}}, p1_sel_141664_comb};
  assign p1_add_142466_comb = {{1{p1_sel_141665_comb[15]}}, p1_sel_141665_comb} + {{1{p1_sel_141666_comb[15]}}, p1_sel_141666_comb};
  assign p1_add_142467_comb = {{1{p1_sel_141667_comb[15]}}, p1_sel_141667_comb} + {{1{p1_sel_141668_comb[15]}}, p1_sel_141668_comb};
  assign p1_add_142468_comb = {{1{p1_sel_141669_comb[15]}}, p1_sel_141669_comb} + {{1{p1_sel_141670_comb[15]}}, p1_sel_141670_comb};
  assign p1_add_142469_comb = {{1{p1_sel_141671_comb[15]}}, p1_sel_141671_comb} + {{1{p1_sel_141672_comb[15]}}, p1_sel_141672_comb};
  assign p1_add_142470_comb = {{1{p1_sel_141673_comb[15]}}, p1_sel_141673_comb} + {{1{p1_sel_141674_comb[15]}}, p1_sel_141674_comb};
  assign p1_add_142471_comb = {{1{p1_sel_141675_comb[15]}}, p1_sel_141675_comb} + {{1{p1_sel_141676_comb[15]}}, p1_sel_141676_comb};
  assign p1_add_142472_comb = {{1{p1_sel_141677_comb[15]}}, p1_sel_141677_comb} + {{1{p1_sel_141678_comb[15]}}, p1_sel_141678_comb};
  assign p1_add_142473_comb = {{1{p1_sel_141679_comb[15]}}, p1_sel_141679_comb} + {{1{p1_sel_141680_comb[15]}}, p1_sel_141680_comb};
  assign p1_add_142474_comb = {{1{p1_sel_141681_comb[15]}}, p1_sel_141681_comb} + {{1{p1_sel_141682_comb[15]}}, p1_sel_141682_comb};
  assign p1_add_142475_comb = {{1{p1_sel_141683_comb[15]}}, p1_sel_141683_comb} + {{1{p1_sel_141684_comb[15]}}, p1_sel_141684_comb};
  assign p1_add_142476_comb = {{1{p1_sel_141685_comb[15]}}, p1_sel_141685_comb} + {{1{p1_sel_141686_comb[15]}}, p1_sel_141686_comb};
  assign p1_add_142477_comb = {{1{p1_sel_141687_comb[15]}}, p1_sel_141687_comb} + {{1{p1_sel_141688_comb[15]}}, p1_sel_141688_comb};
  assign p1_add_142478_comb = {{1{p1_sel_141689_comb[15]}}, p1_sel_141689_comb} + {{1{p1_sel_141690_comb[15]}}, p1_sel_141690_comb};
  assign p1_add_142479_comb = {{1{p1_sel_141691_comb[15]}}, p1_sel_141691_comb} + {{1{p1_sel_141692_comb[15]}}, p1_sel_141692_comb};
  assign p1_add_142480_comb = {{1{p1_sel_141693_comb[15]}}, p1_sel_141693_comb} + {{1{p1_sel_141694_comb[15]}}, p1_sel_141694_comb};
  assign p1_add_142481_comb = {{1{p1_sel_141695_comb[15]}}, p1_sel_141695_comb} + {{1{p1_sel_141696_comb[15]}}, p1_sel_141696_comb};
  assign p1_add_142482_comb = {{1{p1_sel_141697_comb[15]}}, p1_sel_141697_comb} + {{1{p1_sel_141698_comb[15]}}, p1_sel_141698_comb};
  assign p1_add_142483_comb = {{1{p1_sel_141699_comb[15]}}, p1_sel_141699_comb} + {{1{p1_sel_141700_comb[15]}}, p1_sel_141700_comb};
  assign p1_add_142484_comb = {{1{p1_sel_141701_comb[15]}}, p1_sel_141701_comb} + {{1{p1_sel_141702_comb[15]}}, p1_sel_141702_comb};
  assign p1_add_142485_comb = {{1{p1_sel_141703_comb[15]}}, p1_sel_141703_comb} + {{1{p1_sel_141704_comb[15]}}, p1_sel_141704_comb};
  assign p1_add_142486_comb = {{1{p1_sel_141705_comb[15]}}, p1_sel_141705_comb} + {{1{p1_sel_141706_comb[15]}}, p1_sel_141706_comb};
  assign p1_add_142487_comb = {{1{p1_sel_141707_comb[15]}}, p1_sel_141707_comb} + {{1{p1_sel_141708_comb[15]}}, p1_sel_141708_comb};
  assign p1_add_142488_comb = {{1{p1_sel_141709_comb[15]}}, p1_sel_141709_comb} + {{1{p1_sel_141710_comb[15]}}, p1_sel_141710_comb};
  assign p1_add_142489_comb = {{1{p1_sel_141711_comb[15]}}, p1_sel_141711_comb} + {{1{p1_sel_141712_comb[15]}}, p1_sel_141712_comb};
  assign p1_add_142490_comb = {{1{p1_sel_141713_comb[15]}}, p1_sel_141713_comb} + {{1{p1_sel_141714_comb[15]}}, p1_sel_141714_comb};
  assign p1_add_142491_comb = {{1{p1_sel_141715_comb[15]}}, p1_sel_141715_comb} + {{1{p1_sel_141716_comb[15]}}, p1_sel_141716_comb};
  assign p1_add_142492_comb = {{1{p1_sel_141717_comb[15]}}, p1_sel_141717_comb} + {{1{p1_sel_141718_comb[15]}}, p1_sel_141718_comb};
  assign p1_add_142493_comb = {{1{p1_sel_141719_comb[15]}}, p1_sel_141719_comb} + {{1{p1_sel_141720_comb[15]}}, p1_sel_141720_comb};
  assign p1_add_142494_comb = {{1{p1_sel_141721_comb[15]}}, p1_sel_141721_comb} + {{1{p1_sel_141722_comb[15]}}, p1_sel_141722_comb};
  assign p1_add_142495_comb = {{1{p1_sel_141723_comb[15]}}, p1_sel_141723_comb} + {{1{p1_sel_141724_comb[15]}}, p1_sel_141724_comb};
  assign p1_add_142496_comb = {{1{p1_sel_141725_comb[15]}}, p1_sel_141725_comb} + {{1{p1_sel_141726_comb[15]}}, p1_sel_141726_comb};
  assign p1_add_142497_comb = {{1{p1_sel_141727_comb[15]}}, p1_sel_141727_comb} + {{1{p1_sel_141728_comb[15]}}, p1_sel_141728_comb};
  assign p1_add_142498_comb = {{1{p1_sel_141729_comb[15]}}, p1_sel_141729_comb} + {{1{p1_sel_141730_comb[15]}}, p1_sel_141730_comb};
  assign p1_add_142499_comb = {{1{p1_sel_141731_comb[15]}}, p1_sel_141731_comb} + {{1{p1_sel_141732_comb[15]}}, p1_sel_141732_comb};
  assign p1_add_142500_comb = {{1{p1_sel_141733_comb[15]}}, p1_sel_141733_comb} + {{1{p1_sel_141734_comb[15]}}, p1_sel_141734_comb};
  assign p1_add_142501_comb = {{1{p1_sel_141735_comb[15]}}, p1_sel_141735_comb} + {{1{p1_sel_141736_comb[15]}}, p1_sel_141736_comb};
  assign p1_add_142502_comb = {{1{p1_sel_141737_comb[15]}}, p1_sel_141737_comb} + {{1{p1_sel_141738_comb[15]}}, p1_sel_141738_comb};
  assign p1_add_142503_comb = {{1{p1_sel_141739_comb[15]}}, p1_sel_141739_comb} + {{1{p1_sel_141740_comb[15]}}, p1_sel_141740_comb};
  assign p1_add_142504_comb = {{1{p1_sel_141741_comb[15]}}, p1_sel_141741_comb} + {{1{p1_sel_141742_comb[15]}}, p1_sel_141742_comb};
  assign p1_add_142505_comb = {{1{p1_sel_141743_comb[15]}}, p1_sel_141743_comb} + {{1{p1_sel_141744_comb[15]}}, p1_sel_141744_comb};
  assign p1_add_142506_comb = {{1{p1_sel_141745_comb[15]}}, p1_sel_141745_comb} + {{1{p1_sel_141746_comb[15]}}, p1_sel_141746_comb};
  assign p1_add_142507_comb = {{1{p1_sel_141747_comb[15]}}, p1_sel_141747_comb} + {{1{p1_sel_141748_comb[15]}}, p1_sel_141748_comb};
  assign p1_add_142508_comb = {{1{p1_sel_141749_comb[15]}}, p1_sel_141749_comb} + {{1{p1_sel_141750_comb[15]}}, p1_sel_141750_comb};
  assign p1_add_142509_comb = {{1{p1_sel_141751_comb[15]}}, p1_sel_141751_comb} + {{1{p1_sel_141752_comb[15]}}, p1_sel_141752_comb};
  assign p1_add_142510_comb = {{1{p1_sel_141753_comb[15]}}, p1_sel_141753_comb} + {{1{p1_sel_141754_comb[15]}}, p1_sel_141754_comb};
  assign p1_add_142511_comb = {{1{p1_sel_141755_comb[15]}}, p1_sel_141755_comb} + {{1{p1_sel_141756_comb[15]}}, p1_sel_141756_comb};
  assign p1_add_142512_comb = {{1{p1_sel_141757_comb[15]}}, p1_sel_141757_comb} + {{1{p1_sel_141758_comb[15]}}, p1_sel_141758_comb};
  assign p1_add_142513_comb = {{1{p1_sel_141759_comb[15]}}, p1_sel_141759_comb} + {{1{p1_sel_141760_comb[15]}}, p1_sel_141760_comb};
  assign p1_add_142514_comb = {{1{p1_sel_141761_comb[15]}}, p1_sel_141761_comb} + {{1{p1_sel_141762_comb[15]}}, p1_sel_141762_comb};
  assign p1_add_142515_comb = {{1{p1_sel_141763_comb[15]}}, p1_sel_141763_comb} + {{1{p1_sel_141764_comb[15]}}, p1_sel_141764_comb};
  assign p1_add_142516_comb = {{1{p1_sel_141765_comb[15]}}, p1_sel_141765_comb} + {{1{p1_sel_141766_comb[15]}}, p1_sel_141766_comb};
  assign p1_add_142517_comb = {{1{p1_sel_141767_comb[15]}}, p1_sel_141767_comb} + {{1{p1_sel_141768_comb[15]}}, p1_sel_141768_comb};
  assign p1_add_142518_comb = {{1{p1_sel_141769_comb[15]}}, p1_sel_141769_comb} + {{1{p1_sel_141770_comb[15]}}, p1_sel_141770_comb};
  assign p1_add_142519_comb = {{1{p1_sel_141771_comb[15]}}, p1_sel_141771_comb} + {{1{p1_sel_141772_comb[15]}}, p1_sel_141772_comb};
  assign p1_add_142520_comb = {{1{p1_sel_141773_comb[15]}}, p1_sel_141773_comb} + {{1{p1_sel_141774_comb[15]}}, p1_sel_141774_comb};
  assign p1_add_142521_comb = {{1{p1_sel_141775_comb[15]}}, p1_sel_141775_comb} + {{1{p1_sel_141776_comb[15]}}, p1_sel_141776_comb};
  assign p1_add_142522_comb = {{1{p1_sel_141777_comb[15]}}, p1_sel_141777_comb} + {{1{p1_sel_141778_comb[15]}}, p1_sel_141778_comb};
  assign p1_add_142523_comb = {{1{p1_sel_141779_comb[15]}}, p1_sel_141779_comb} + {{1{p1_sel_141780_comb[15]}}, p1_sel_141780_comb};
  assign p1_add_142524_comb = {{1{p1_sel_141781_comb[15]}}, p1_sel_141781_comb} + {{1{p1_sel_141782_comb[15]}}, p1_sel_141782_comb};
  assign p1_add_142525_comb = {{1{p1_sel_141783_comb[15]}}, p1_sel_141783_comb} + {{1{p1_sel_141784_comb[15]}}, p1_sel_141784_comb};
  assign p1_add_142526_comb = {{1{p1_sel_141785_comb[15]}}, p1_sel_141785_comb} + {{1{p1_sel_141786_comb[15]}}, p1_sel_141786_comb};
  assign p1_add_142527_comb = {{1{p1_sel_141787_comb[15]}}, p1_sel_141787_comb} + {{1{p1_sel_141788_comb[15]}}, p1_sel_141788_comb};
  assign p1_add_142528_comb = {{1{p1_sel_141789_comb[15]}}, p1_sel_141789_comb} + {{1{p1_sel_141790_comb[15]}}, p1_sel_141790_comb};
  assign p1_add_142529_comb = {{1{p1_sel_141791_comb[15]}}, p1_sel_141791_comb} + {{1{p1_sel_141792_comb[15]}}, p1_sel_141792_comb};
  assign p1_add_142530_comb = {{1{p1_sel_141793_comb[15]}}, p1_sel_141793_comb} + {{1{p1_sel_141794_comb[15]}}, p1_sel_141794_comb};
  assign p1_add_142531_comb = {{1{p1_sel_141795_comb[15]}}, p1_sel_141795_comb} + {{1{p1_sel_141796_comb[15]}}, p1_sel_141796_comb};
  assign p1_add_142532_comb = {{1{p1_sel_141797_comb[15]}}, p1_sel_141797_comb} + {{1{p1_sel_141798_comb[15]}}, p1_sel_141798_comb};
  assign p1_add_142533_comb = {{1{p1_sel_141799_comb[15]}}, p1_sel_141799_comb} + {{1{p1_sel_141800_comb[15]}}, p1_sel_141800_comb};
  assign p1_add_142534_comb = {{1{p1_sel_141801_comb[15]}}, p1_sel_141801_comb} + {{1{p1_sel_141802_comb[15]}}, p1_sel_141802_comb};
  assign p1_add_142535_comb = {{1{p1_sel_141803_comb[15]}}, p1_sel_141803_comb} + {{1{p1_sel_141804_comb[15]}}, p1_sel_141804_comb};
  assign p1_add_142536_comb = {{1{p1_sel_141805_comb[15]}}, p1_sel_141805_comb} + {{1{p1_sel_141806_comb[15]}}, p1_sel_141806_comb};
  assign p1_add_142537_comb = {{1{p1_sel_141807_comb[15]}}, p1_sel_141807_comb} + {{1{p1_sel_141808_comb[15]}}, p1_sel_141808_comb};
  assign p1_add_142538_comb = {{1{p1_sel_141809_comb[15]}}, p1_sel_141809_comb} + {{1{p1_sel_141810_comb[15]}}, p1_sel_141810_comb};
  assign p1_add_142539_comb = {{1{p1_sel_141811_comb[15]}}, p1_sel_141811_comb} + {{1{p1_sel_141812_comb[15]}}, p1_sel_141812_comb};
  assign p1_add_142540_comb = {{1{p1_sel_141813_comb[15]}}, p1_sel_141813_comb} + {{1{p1_sel_141814_comb[15]}}, p1_sel_141814_comb};
  assign p1_add_142541_comb = {{1{p1_sel_141815_comb[15]}}, p1_sel_141815_comb} + {{1{p1_sel_141816_comb[15]}}, p1_sel_141816_comb};
  assign p1_add_142542_comb = {{1{p1_sel_141817_comb[15]}}, p1_sel_141817_comb} + {{1{p1_sel_141818_comb[15]}}, p1_sel_141818_comb};
  assign p1_add_142543_comb = {{1{p1_sel_141819_comb[15]}}, p1_sel_141819_comb} + {{1{p1_sel_141820_comb[15]}}, p1_sel_141820_comb};
  assign p1_add_142544_comb = {{1{p1_sel_141821_comb[15]}}, p1_sel_141821_comb} + {{1{p1_sel_141822_comb[15]}}, p1_sel_141822_comb};
  assign p1_add_142545_comb = {{1{p1_sel_141823_comb[15]}}, p1_sel_141823_comb} + {{1{p1_sel_141824_comb[15]}}, p1_sel_141824_comb};
  assign p1_add_142546_comb = {{1{p1_sel_141825_comb[15]}}, p1_sel_141825_comb} + {{1{p1_sel_141826_comb[15]}}, p1_sel_141826_comb};
  assign p1_sum__995_comb = p1_sum__993_comb + p1_sum__994_comb;
  assign p1_sum__890_comb = p1_sum__888_comb + p1_sum__889_comb;
  assign p1_sum__1784_comb = {{8{p1_add_142311_comb[16]}}, p1_add_142311_comb};
  assign p1_sum__1785_comb = {{8{p1_add_142312_comb[16]}}, p1_add_142312_comb};
  assign p1_sum__1786_comb = {{8{p1_add_142313_comb[16]}}, p1_add_142313_comb};
  assign p1_sum__1787_comb = {{8{p1_add_142314_comb[16]}}, p1_add_142314_comb};
  assign p1_sum__1724_comb = {{8{p1_add_142315_comb[16]}}, p1_add_142315_comb};
  assign p1_sum__1725_comb = {{8{p1_add_142316_comb[16]}}, p1_add_142316_comb};
  assign p1_sum__1726_comb = {{8{p1_add_142317_comb[16]}}, p1_add_142317_comb};
  assign p1_sum__1727_comb = {{8{p1_add_142318_comb[16]}}, p1_add_142318_comb};
  assign p1_sum__1772_comb = {{8{p1_add_142319_comb[16]}}, p1_add_142319_comb};
  assign p1_sum__1773_comb = {{8{p1_add_142320_comb[16]}}, p1_add_142320_comb};
  assign p1_sum__1774_comb = {{8{p1_add_142321_comb[16]}}, p1_add_142321_comb};
  assign p1_sum__1775_comb = {{8{p1_add_142322_comb[16]}}, p1_add_142322_comb};
  assign p1_sum__1700_comb = {{8{p1_add_142323_comb[16]}}, p1_add_142323_comb};
  assign p1_sum__1701_comb = {{8{p1_add_142324_comb[16]}}, p1_add_142324_comb};
  assign p1_sum__1702_comb = {{8{p1_add_142325_comb[16]}}, p1_add_142325_comb};
  assign p1_sum__1703_comb = {{8{p1_add_142326_comb[16]}}, p1_add_142326_comb};
  assign p1_sum__1756_comb = {{8{p1_add_142327_comb[16]}}, p1_add_142327_comb};
  assign p1_sum__1757_comb = {{8{p1_add_142328_comb[16]}}, p1_add_142328_comb};
  assign p1_sum__1758_comb = {{8{p1_add_142329_comb[16]}}, p1_add_142329_comb};
  assign p1_sum__1759_comb = {{8{p1_add_142330_comb[16]}}, p1_add_142330_comb};
  assign p1_sum__1676_comb = {{8{p1_add_142331_comb[16]}}, p1_add_142331_comb};
  assign p1_sum__1677_comb = {{8{p1_add_142332_comb[16]}}, p1_add_142332_comb};
  assign p1_sum__1678_comb = {{8{p1_add_142333_comb[16]}}, p1_add_142333_comb};
  assign p1_sum__1679_comb = {{8{p1_add_142334_comb[16]}}, p1_add_142334_comb};
  assign p1_sum__1736_comb = {{8{p1_add_142335_comb[16]}}, p1_add_142335_comb};
  assign p1_sum__1737_comb = {{8{p1_add_142336_comb[16]}}, p1_add_142336_comb};
  assign p1_sum__1738_comb = {{8{p1_add_142337_comb[16]}}, p1_add_142337_comb};
  assign p1_sum__1739_comb = {{8{p1_add_142338_comb[16]}}, p1_add_142338_comb};
  assign p1_sum__1652_comb = {{8{p1_add_142339_comb[16]}}, p1_add_142339_comb};
  assign p1_sum__1653_comb = {{8{p1_add_142340_comb[16]}}, p1_add_142340_comb};
  assign p1_sum__1654_comb = {{8{p1_add_142341_comb[16]}}, p1_add_142341_comb};
  assign p1_sum__1655_comb = {{8{p1_add_142342_comb[16]}}, p1_add_142342_comb};
  assign p1_sum__1712_comb = {{8{p1_add_142343_comb[16]}}, p1_add_142343_comb};
  assign p1_sum__1713_comb = {{8{p1_add_142344_comb[16]}}, p1_add_142344_comb};
  assign p1_sum__1714_comb = {{8{p1_add_142345_comb[16]}}, p1_add_142345_comb};
  assign p1_sum__1715_comb = {{8{p1_add_142346_comb[16]}}, p1_add_142346_comb};
  assign p1_sum__1632_comb = {{8{p1_add_142347_comb[16]}}, p1_add_142347_comb};
  assign p1_sum__1633_comb = {{8{p1_add_142348_comb[16]}}, p1_add_142348_comb};
  assign p1_sum__1634_comb = {{8{p1_add_142349_comb[16]}}, p1_add_142349_comb};
  assign p1_sum__1635_comb = {{8{p1_add_142350_comb[16]}}, p1_add_142350_comb};
  assign p1_sum__1688_comb = {{8{p1_add_142351_comb[16]}}, p1_add_142351_comb};
  assign p1_sum__1689_comb = {{8{p1_add_142352_comb[16]}}, p1_add_142352_comb};
  assign p1_sum__1690_comb = {{8{p1_add_142353_comb[16]}}, p1_add_142353_comb};
  assign p1_sum__1691_comb = {{8{p1_add_142354_comb[16]}}, p1_add_142354_comb};
  assign p1_sum__1616_comb = {{8{p1_add_142355_comb[16]}}, p1_add_142355_comb};
  assign p1_sum__1617_comb = {{8{p1_add_142356_comb[16]}}, p1_add_142356_comb};
  assign p1_sum__1618_comb = {{8{p1_add_142357_comb[16]}}, p1_add_142357_comb};
  assign p1_sum__1619_comb = {{8{p1_add_142358_comb[16]}}, p1_add_142358_comb};
  assign p1_sum__1664_comb = {{8{p1_add_142359_comb[16]}}, p1_add_142359_comb};
  assign p1_sum__1665_comb = {{8{p1_add_142360_comb[16]}}, p1_add_142360_comb};
  assign p1_sum__1666_comb = {{8{p1_add_142361_comb[16]}}, p1_add_142361_comb};
  assign p1_sum__1667_comb = {{8{p1_add_142362_comb[16]}}, p1_add_142362_comb};
  assign p1_sum__1604_comb = {{8{p1_add_142363_comb[16]}}, p1_add_142363_comb};
  assign p1_sum__1605_comb = {{8{p1_add_142364_comb[16]}}, p1_add_142364_comb};
  assign p1_sum__1606_comb = {{8{p1_add_142365_comb[16]}}, p1_add_142365_comb};
  assign p1_sum__1607_comb = {{8{p1_add_142366_comb[16]}}, p1_add_142366_comb};
  assign p1_sum__1023_comb = p1_sum__1021_comb + p1_sum__1022_comb;
  assign p1_sum__1016_comb = p1_sum__1014_comb + p1_sum__1015_comb;
  assign p1_sum__967_comb = p1_sum__965_comb + p1_sum__966_comb;
  assign p1_sum__932_comb = p1_sum__930_comb + p1_sum__931_comb;
  assign p1_sum__841_comb = p1_sum__839_comb + p1_sum__840_comb;
  assign p1_sum__785_comb = p1_sum__783_comb + p1_sum__784_comb;
  assign p1_sum__1804_comb = {{8{p1_add_142379_comb[16]}}, p1_add_142379_comb};
  assign p1_sum__1805_comb = {{8{p1_add_142380_comb[16]}}, p1_add_142380_comb};
  assign p1_sum__1806_comb = {{8{p1_add_142381_comb[16]}}, p1_add_142381_comb};
  assign p1_sum__1807_comb = {{8{p1_add_142382_comb[16]}}, p1_add_142382_comb};
  assign p1_sum__1796_comb = {{8{p1_add_142383_comb[16]}}, p1_add_142383_comb};
  assign p1_sum__1797_comb = {{8{p1_add_142384_comb[16]}}, p1_add_142384_comb};
  assign p1_sum__1798_comb = {{8{p1_add_142385_comb[16]}}, p1_add_142385_comb};
  assign p1_sum__1799_comb = {{8{p1_add_142386_comb[16]}}, p1_add_142386_comb};
  assign p1_sum__1768_comb = {{8{p1_add_142387_comb[16]}}, p1_add_142387_comb};
  assign p1_sum__1769_comb = {{8{p1_add_142388_comb[16]}}, p1_add_142388_comb};
  assign p1_sum__1770_comb = {{8{p1_add_142389_comb[16]}}, p1_add_142389_comb};
  assign p1_sum__1771_comb = {{8{p1_add_142390_comb[16]}}, p1_add_142390_comb};
  assign p1_sum__1748_comb = {{8{p1_add_142391_comb[16]}}, p1_add_142391_comb};
  assign p1_sum__1749_comb = {{8{p1_add_142392_comb[16]}}, p1_add_142392_comb};
  assign p1_sum__1750_comb = {{8{p1_add_142393_comb[16]}}, p1_add_142393_comb};
  assign p1_sum__1751_comb = {{8{p1_add_142394_comb[16]}}, p1_add_142394_comb};
  assign p1_sum__1696_comb = {{8{p1_add_142395_comb[16]}}, p1_add_142395_comb};
  assign p1_sum__1697_comb = {{8{p1_add_142396_comb[16]}}, p1_add_142396_comb};
  assign p1_sum__1698_comb = {{8{p1_add_142397_comb[16]}}, p1_add_142397_comb};
  assign p1_sum__1699_comb = {{8{p1_add_142398_comb[16]}}, p1_add_142398_comb};
  assign p1_sum__1668_comb = {{8{p1_add_142399_comb[16]}}, p1_add_142399_comb};
  assign p1_sum__1669_comb = {{8{p1_add_142400_comb[16]}}, p1_add_142400_comb};
  assign p1_sum__1670_comb = {{8{p1_add_142401_comb[16]}}, p1_add_142401_comb};
  assign p1_sum__1671_comb = {{8{p1_add_142402_comb[16]}}, p1_add_142402_comb};
  assign p1_sum__1800_comb = {{8{p1_add_142403_comb[16]}}, p1_add_142403_comb};
  assign p1_sum__1801_comb = {{8{p1_add_142404_comb[16]}}, p1_add_142404_comb};
  assign p1_sum__1802_comb = {{8{p1_add_142405_comb[16]}}, p1_add_142405_comb};
  assign p1_sum__1803_comb = {{8{p1_add_142406_comb[16]}}, p1_add_142406_comb};
  assign p1_sum__1788_comb = {{8{p1_add_142407_comb[16]}}, p1_add_142407_comb};
  assign p1_sum__1789_comb = {{8{p1_add_142408_comb[16]}}, p1_add_142408_comb};
  assign p1_sum__1790_comb = {{8{p1_add_142409_comb[16]}}, p1_add_142409_comb};
  assign p1_sum__1791_comb = {{8{p1_add_142410_comb[16]}}, p1_add_142410_comb};
  assign p1_sum__1752_comb = {{8{p1_add_142411_comb[16]}}, p1_add_142411_comb};
  assign p1_sum__1753_comb = {{8{p1_add_142412_comb[16]}}, p1_add_142412_comb};
  assign p1_sum__1754_comb = {{8{p1_add_142413_comb[16]}}, p1_add_142413_comb};
  assign p1_sum__1755_comb = {{8{p1_add_142414_comb[16]}}, p1_add_142414_comb};
  assign p1_sum__1728_comb = {{8{p1_add_142415_comb[16]}}, p1_add_142415_comb};
  assign p1_sum__1729_comb = {{8{p1_add_142416_comb[16]}}, p1_add_142416_comb};
  assign p1_sum__1730_comb = {{8{p1_add_142417_comb[16]}}, p1_add_142417_comb};
  assign p1_sum__1731_comb = {{8{p1_add_142418_comb[16]}}, p1_add_142418_comb};
  assign p1_sum__1672_comb = {{8{p1_add_142419_comb[16]}}, p1_add_142419_comb};
  assign p1_sum__1673_comb = {{8{p1_add_142420_comb[16]}}, p1_add_142420_comb};
  assign p1_sum__1674_comb = {{8{p1_add_142421_comb[16]}}, p1_add_142421_comb};
  assign p1_sum__1675_comb = {{8{p1_add_142422_comb[16]}}, p1_add_142422_comb};
  assign p1_sum__1644_comb = {{8{p1_add_142423_comb[16]}}, p1_add_142423_comb};
  assign p1_sum__1645_comb = {{8{p1_add_142424_comb[16]}}, p1_add_142424_comb};
  assign p1_sum__1646_comb = {{8{p1_add_142425_comb[16]}}, p1_add_142425_comb};
  assign p1_sum__1647_comb = {{8{p1_add_142426_comb[16]}}, p1_add_142426_comb};
  assign p1_sum__1792_comb = {{8{p1_add_142427_comb[16]}}, p1_add_142427_comb};
  assign p1_sum__1793_comb = {{8{p1_add_142428_comb[16]}}, p1_add_142428_comb};
  assign p1_sum__1794_comb = {{8{p1_add_142429_comb[16]}}, p1_add_142429_comb};
  assign p1_sum__1795_comb = {{8{p1_add_142430_comb[16]}}, p1_add_142430_comb};
  assign p1_sum__1776_comb = {{8{p1_add_142431_comb[16]}}, p1_add_142431_comb};
  assign p1_sum__1777_comb = {{8{p1_add_142432_comb[16]}}, p1_add_142432_comb};
  assign p1_sum__1778_comb = {{8{p1_add_142433_comb[16]}}, p1_add_142433_comb};
  assign p1_sum__1779_comb = {{8{p1_add_142434_comb[16]}}, p1_add_142434_comb};
  assign p1_sum__1732_comb = {{8{p1_add_142435_comb[16]}}, p1_add_142435_comb};
  assign p1_sum__1733_comb = {{8{p1_add_142436_comb[16]}}, p1_add_142436_comb};
  assign p1_sum__1734_comb = {{8{p1_add_142437_comb[16]}}, p1_add_142437_comb};
  assign p1_sum__1735_comb = {{8{p1_add_142438_comb[16]}}, p1_add_142438_comb};
  assign p1_sum__1704_comb = {{8{p1_add_142439_comb[16]}}, p1_add_142439_comb};
  assign p1_sum__1705_comb = {{8{p1_add_142440_comb[16]}}, p1_add_142440_comb};
  assign p1_sum__1706_comb = {{8{p1_add_142441_comb[16]}}, p1_add_142441_comb};
  assign p1_sum__1707_comb = {{8{p1_add_142442_comb[16]}}, p1_add_142442_comb};
  assign p1_sum__1648_comb = {{8{p1_add_142443_comb[16]}}, p1_add_142443_comb};
  assign p1_sum__1649_comb = {{8{p1_add_142444_comb[16]}}, p1_add_142444_comb};
  assign p1_sum__1650_comb = {{8{p1_add_142445_comb[16]}}, p1_add_142445_comb};
  assign p1_sum__1651_comb = {{8{p1_add_142446_comb[16]}}, p1_add_142446_comb};
  assign p1_sum__1624_comb = {{8{p1_add_142447_comb[16]}}, p1_add_142447_comb};
  assign p1_sum__1625_comb = {{8{p1_add_142448_comb[16]}}, p1_add_142448_comb};
  assign p1_sum__1626_comb = {{8{p1_add_142449_comb[16]}}, p1_add_142449_comb};
  assign p1_sum__1627_comb = {{8{p1_add_142450_comb[16]}}, p1_add_142450_comb};
  assign p1_sum__1780_comb = {{8{p1_add_142451_comb[16]}}, p1_add_142451_comb};
  assign p1_sum__1781_comb = {{8{p1_add_142452_comb[16]}}, p1_add_142452_comb};
  assign p1_sum__1782_comb = {{8{p1_add_142453_comb[16]}}, p1_add_142453_comb};
  assign p1_sum__1783_comb = {{8{p1_add_142454_comb[16]}}, p1_add_142454_comb};
  assign p1_sum__1760_comb = {{8{p1_add_142455_comb[16]}}, p1_add_142455_comb};
  assign p1_sum__1761_comb = {{8{p1_add_142456_comb[16]}}, p1_add_142456_comb};
  assign p1_sum__1762_comb = {{8{p1_add_142457_comb[16]}}, p1_add_142457_comb};
  assign p1_sum__1763_comb = {{8{p1_add_142458_comb[16]}}, p1_add_142458_comb};
  assign p1_sum__1708_comb = {{8{p1_add_142459_comb[16]}}, p1_add_142459_comb};
  assign p1_sum__1709_comb = {{8{p1_add_142460_comb[16]}}, p1_add_142460_comb};
  assign p1_sum__1710_comb = {{8{p1_add_142461_comb[16]}}, p1_add_142461_comb};
  assign p1_sum__1711_comb = {{8{p1_add_142462_comb[16]}}, p1_add_142462_comb};
  assign p1_sum__1680_comb = {{8{p1_add_142463_comb[16]}}, p1_add_142463_comb};
  assign p1_sum__1681_comb = {{8{p1_add_142464_comb[16]}}, p1_add_142464_comb};
  assign p1_sum__1682_comb = {{8{p1_add_142465_comb[16]}}, p1_add_142465_comb};
  assign p1_sum__1683_comb = {{8{p1_add_142466_comb[16]}}, p1_add_142466_comb};
  assign p1_sum__1628_comb = {{8{p1_add_142467_comb[16]}}, p1_add_142467_comb};
  assign p1_sum__1629_comb = {{8{p1_add_142468_comb[16]}}, p1_add_142468_comb};
  assign p1_sum__1630_comb = {{8{p1_add_142469_comb[16]}}, p1_add_142469_comb};
  assign p1_sum__1631_comb = {{8{p1_add_142470_comb[16]}}, p1_add_142470_comb};
  assign p1_sum__1608_comb = {{8{p1_add_142471_comb[16]}}, p1_add_142471_comb};
  assign p1_sum__1609_comb = {{8{p1_add_142472_comb[16]}}, p1_add_142472_comb};
  assign p1_sum__1610_comb = {{8{p1_add_142473_comb[16]}}, p1_add_142473_comb};
  assign p1_sum__1611_comb = {{8{p1_add_142474_comb[16]}}, p1_add_142474_comb};
  assign p1_sum__1764_comb = {{8{p1_add_142475_comb[16]}}, p1_add_142475_comb};
  assign p1_sum__1765_comb = {{8{p1_add_142476_comb[16]}}, p1_add_142476_comb};
  assign p1_sum__1766_comb = {{8{p1_add_142477_comb[16]}}, p1_add_142477_comb};
  assign p1_sum__1767_comb = {{8{p1_add_142478_comb[16]}}, p1_add_142478_comb};
  assign p1_sum__1740_comb = {{8{p1_add_142479_comb[16]}}, p1_add_142479_comb};
  assign p1_sum__1741_comb = {{8{p1_add_142480_comb[16]}}, p1_add_142480_comb};
  assign p1_sum__1742_comb = {{8{p1_add_142481_comb[16]}}, p1_add_142481_comb};
  assign p1_sum__1743_comb = {{8{p1_add_142482_comb[16]}}, p1_add_142482_comb};
  assign p1_sum__1684_comb = {{8{p1_add_142483_comb[16]}}, p1_add_142483_comb};
  assign p1_sum__1685_comb = {{8{p1_add_142484_comb[16]}}, p1_add_142484_comb};
  assign p1_sum__1686_comb = {{8{p1_add_142485_comb[16]}}, p1_add_142485_comb};
  assign p1_sum__1687_comb = {{8{p1_add_142486_comb[16]}}, p1_add_142486_comb};
  assign p1_sum__1656_comb = {{8{p1_add_142487_comb[16]}}, p1_add_142487_comb};
  assign p1_sum__1657_comb = {{8{p1_add_142488_comb[16]}}, p1_add_142488_comb};
  assign p1_sum__1658_comb = {{8{p1_add_142489_comb[16]}}, p1_add_142489_comb};
  assign p1_sum__1659_comb = {{8{p1_add_142490_comb[16]}}, p1_add_142490_comb};
  assign p1_sum__1612_comb = {{8{p1_add_142491_comb[16]}}, p1_add_142491_comb};
  assign p1_sum__1613_comb = {{8{p1_add_142492_comb[16]}}, p1_add_142492_comb};
  assign p1_sum__1614_comb = {{8{p1_add_142493_comb[16]}}, p1_add_142493_comb};
  assign p1_sum__1615_comb = {{8{p1_add_142494_comb[16]}}, p1_add_142494_comb};
  assign p1_sum__1596_comb = {{8{p1_add_142495_comb[16]}}, p1_add_142495_comb};
  assign p1_sum__1597_comb = {{8{p1_add_142496_comb[16]}}, p1_add_142496_comb};
  assign p1_sum__1598_comb = {{8{p1_add_142497_comb[16]}}, p1_add_142497_comb};
  assign p1_sum__1599_comb = {{8{p1_add_142498_comb[16]}}, p1_add_142498_comb};
  assign p1_sum__1744_comb = {{8{p1_add_142499_comb[16]}}, p1_add_142499_comb};
  assign p1_sum__1745_comb = {{8{p1_add_142500_comb[16]}}, p1_add_142500_comb};
  assign p1_sum__1746_comb = {{8{p1_add_142501_comb[16]}}, p1_add_142501_comb};
  assign p1_sum__1747_comb = {{8{p1_add_142502_comb[16]}}, p1_add_142502_comb};
  assign p1_sum__1716_comb = {{8{p1_add_142503_comb[16]}}, p1_add_142503_comb};
  assign p1_sum__1717_comb = {{8{p1_add_142504_comb[16]}}, p1_add_142504_comb};
  assign p1_sum__1718_comb = {{8{p1_add_142505_comb[16]}}, p1_add_142505_comb};
  assign p1_sum__1719_comb = {{8{p1_add_142506_comb[16]}}, p1_add_142506_comb};
  assign p1_sum__1660_comb = {{8{p1_add_142507_comb[16]}}, p1_add_142507_comb};
  assign p1_sum__1661_comb = {{8{p1_add_142508_comb[16]}}, p1_add_142508_comb};
  assign p1_sum__1662_comb = {{8{p1_add_142509_comb[16]}}, p1_add_142509_comb};
  assign p1_sum__1663_comb = {{8{p1_add_142510_comb[16]}}, p1_add_142510_comb};
  assign p1_sum__1636_comb = {{8{p1_add_142511_comb[16]}}, p1_add_142511_comb};
  assign p1_sum__1637_comb = {{8{p1_add_142512_comb[16]}}, p1_add_142512_comb};
  assign p1_sum__1638_comb = {{8{p1_add_142513_comb[16]}}, p1_add_142513_comb};
  assign p1_sum__1639_comb = {{8{p1_add_142514_comb[16]}}, p1_add_142514_comb};
  assign p1_sum__1600_comb = {{8{p1_add_142515_comb[16]}}, p1_add_142515_comb};
  assign p1_sum__1601_comb = {{8{p1_add_142516_comb[16]}}, p1_add_142516_comb};
  assign p1_sum__1602_comb = {{8{p1_add_142517_comb[16]}}, p1_add_142517_comb};
  assign p1_sum__1603_comb = {{8{p1_add_142518_comb[16]}}, p1_add_142518_comb};
  assign p1_sum__1588_comb = {{8{p1_add_142519_comb[16]}}, p1_add_142519_comb};
  assign p1_sum__1589_comb = {{8{p1_add_142520_comb[16]}}, p1_add_142520_comb};
  assign p1_sum__1590_comb = {{8{p1_add_142521_comb[16]}}, p1_add_142521_comb};
  assign p1_sum__1591_comb = {{8{p1_add_142522_comb[16]}}, p1_add_142522_comb};
  assign p1_sum__1720_comb = {{8{p1_add_142523_comb[16]}}, p1_add_142523_comb};
  assign p1_sum__1721_comb = {{8{p1_add_142524_comb[16]}}, p1_add_142524_comb};
  assign p1_sum__1722_comb = {{8{p1_add_142525_comb[16]}}, p1_add_142525_comb};
  assign p1_sum__1723_comb = {{8{p1_add_142526_comb[16]}}, p1_add_142526_comb};
  assign p1_sum__1692_comb = {{8{p1_add_142527_comb[16]}}, p1_add_142527_comb};
  assign p1_sum__1693_comb = {{8{p1_add_142528_comb[16]}}, p1_add_142528_comb};
  assign p1_sum__1694_comb = {{8{p1_add_142529_comb[16]}}, p1_add_142529_comb};
  assign p1_sum__1695_comb = {{8{p1_add_142530_comb[16]}}, p1_add_142530_comb};
  assign p1_sum__1640_comb = {{8{p1_add_142531_comb[16]}}, p1_add_142531_comb};
  assign p1_sum__1641_comb = {{8{p1_add_142532_comb[16]}}, p1_add_142532_comb};
  assign p1_sum__1642_comb = {{8{p1_add_142533_comb[16]}}, p1_add_142533_comb};
  assign p1_sum__1643_comb = {{8{p1_add_142534_comb[16]}}, p1_add_142534_comb};
  assign p1_sum__1620_comb = {{8{p1_add_142535_comb[16]}}, p1_add_142535_comb};
  assign p1_sum__1621_comb = {{8{p1_add_142536_comb[16]}}, p1_add_142536_comb};
  assign p1_sum__1622_comb = {{8{p1_add_142537_comb[16]}}, p1_add_142537_comb};
  assign p1_sum__1623_comb = {{8{p1_add_142538_comb[16]}}, p1_add_142538_comb};
  assign p1_sum__1592_comb = {{8{p1_add_142539_comb[16]}}, p1_add_142539_comb};
  assign p1_sum__1593_comb = {{8{p1_add_142540_comb[16]}}, p1_add_142540_comb};
  assign p1_sum__1594_comb = {{8{p1_add_142541_comb[16]}}, p1_add_142541_comb};
  assign p1_sum__1595_comb = {{8{p1_add_142542_comb[16]}}, p1_add_142542_comb};
  assign p1_sum__1584_comb = {{8{p1_add_142543_comb[16]}}, p1_add_142543_comb};
  assign p1_sum__1585_comb = {{8{p1_add_142544_comb[16]}}, p1_add_142544_comb};
  assign p1_sum__1586_comb = {{8{p1_add_142545_comb[16]}}, p1_add_142545_comb};
  assign p1_sum__1587_comb = {{8{p1_add_142546_comb[16]}}, p1_add_142546_comb};
  assign p1_umul_142787_comb = umul32b_32b_x_7b(p1_sum__995_comb, 7'h5b);
  assign p1_umul_142788_comb = umul32b_32b_x_7b(p1_sum__890_comb, 7'h5b);
  assign p1_sum__1348_comb = p1_sum__1784_comb + p1_sum__1785_comb;
  assign p1_sum__1349_comb = p1_sum__1786_comb + p1_sum__1787_comb;
  assign p1_sum__1318_comb = p1_sum__1724_comb + p1_sum__1725_comb;
  assign p1_sum__1319_comb = p1_sum__1726_comb + p1_sum__1727_comb;
  assign p1_sum__1342_comb = p1_sum__1772_comb + p1_sum__1773_comb;
  assign p1_sum__1343_comb = p1_sum__1774_comb + p1_sum__1775_comb;
  assign p1_sum__1306_comb = p1_sum__1700_comb + p1_sum__1701_comb;
  assign p1_sum__1307_comb = p1_sum__1702_comb + p1_sum__1703_comb;
  assign p1_sum__1334_comb = p1_sum__1756_comb + p1_sum__1757_comb;
  assign p1_sum__1335_comb = p1_sum__1758_comb + p1_sum__1759_comb;
  assign p1_sum__1294_comb = p1_sum__1676_comb + p1_sum__1677_comb;
  assign p1_sum__1295_comb = p1_sum__1678_comb + p1_sum__1679_comb;
  assign p1_sum__1324_comb = p1_sum__1736_comb + p1_sum__1737_comb;
  assign p1_sum__1325_comb = p1_sum__1738_comb + p1_sum__1739_comb;
  assign p1_sum__1282_comb = p1_sum__1652_comb + p1_sum__1653_comb;
  assign p1_sum__1283_comb = p1_sum__1654_comb + p1_sum__1655_comb;
  assign p1_sum__1312_comb = p1_sum__1712_comb + p1_sum__1713_comb;
  assign p1_sum__1313_comb = p1_sum__1714_comb + p1_sum__1715_comb;
  assign p1_sum__1272_comb = p1_sum__1632_comb + p1_sum__1633_comb;
  assign p1_sum__1273_comb = p1_sum__1634_comb + p1_sum__1635_comb;
  assign p1_sum__1300_comb = p1_sum__1688_comb + p1_sum__1689_comb;
  assign p1_sum__1301_comb = p1_sum__1690_comb + p1_sum__1691_comb;
  assign p1_sum__1264_comb = p1_sum__1616_comb + p1_sum__1617_comb;
  assign p1_sum__1265_comb = p1_sum__1618_comb + p1_sum__1619_comb;
  assign p1_sum__1288_comb = p1_sum__1664_comb + p1_sum__1665_comb;
  assign p1_sum__1289_comb = p1_sum__1666_comb + p1_sum__1667_comb;
  assign p1_sum__1258_comb = p1_sum__1604_comb + p1_sum__1605_comb;
  assign p1_sum__1259_comb = p1_sum__1606_comb + p1_sum__1607_comb;
  assign p1_umul_142817_comb = umul32b_32b_x_7b(p1_sum__1023_comb, 7'h5b);
  assign p1_umul_142818_comb = umul32b_32b_x_7b(p1_sum__1016_comb, 7'h5b);
  assign p1_umul_142819_comb = umul32b_32b_x_7b(p1_sum__967_comb, 7'h5b);
  assign p1_umul_142820_comb = umul32b_32b_x_7b(p1_sum__932_comb, 7'h5b);
  assign p1_umul_142821_comb = umul32b_32b_x_7b(p1_sum__841_comb, 7'h5b);
  assign p1_umul_142822_comb = umul32b_32b_x_7b(p1_sum__785_comb, 7'h5b);
  assign p1_sum__1358_comb = p1_sum__1804_comb + p1_sum__1805_comb;
  assign p1_sum__1359_comb = p1_sum__1806_comb + p1_sum__1807_comb;
  assign p1_sum__1354_comb = p1_sum__1796_comb + p1_sum__1797_comb;
  assign p1_sum__1355_comb = p1_sum__1798_comb + p1_sum__1799_comb;
  assign p1_sum__1340_comb = p1_sum__1768_comb + p1_sum__1769_comb;
  assign p1_sum__1341_comb = p1_sum__1770_comb + p1_sum__1771_comb;
  assign p1_sum__1330_comb = p1_sum__1748_comb + p1_sum__1749_comb;
  assign p1_sum__1331_comb = p1_sum__1750_comb + p1_sum__1751_comb;
  assign p1_sum__1304_comb = p1_sum__1696_comb + p1_sum__1697_comb;
  assign p1_sum__1305_comb = p1_sum__1698_comb + p1_sum__1699_comb;
  assign p1_sum__1290_comb = p1_sum__1668_comb + p1_sum__1669_comb;
  assign p1_sum__1291_comb = p1_sum__1670_comb + p1_sum__1671_comb;
  assign p1_sum__1356_comb = p1_sum__1800_comb + p1_sum__1801_comb;
  assign p1_sum__1357_comb = p1_sum__1802_comb + p1_sum__1803_comb;
  assign p1_sum__1350_comb = p1_sum__1788_comb + p1_sum__1789_comb;
  assign p1_sum__1351_comb = p1_sum__1790_comb + p1_sum__1791_comb;
  assign p1_sum__1332_comb = p1_sum__1752_comb + p1_sum__1753_comb;
  assign p1_sum__1333_comb = p1_sum__1754_comb + p1_sum__1755_comb;
  assign p1_sum__1320_comb = p1_sum__1728_comb + p1_sum__1729_comb;
  assign p1_sum__1321_comb = p1_sum__1730_comb + p1_sum__1731_comb;
  assign p1_sum__1292_comb = p1_sum__1672_comb + p1_sum__1673_comb;
  assign p1_sum__1293_comb = p1_sum__1674_comb + p1_sum__1675_comb;
  assign p1_sum__1278_comb = p1_sum__1644_comb + p1_sum__1645_comb;
  assign p1_sum__1279_comb = p1_sum__1646_comb + p1_sum__1647_comb;
  assign p1_sum__1352_comb = p1_sum__1792_comb + p1_sum__1793_comb;
  assign p1_sum__1353_comb = p1_sum__1794_comb + p1_sum__1795_comb;
  assign p1_sum__1344_comb = p1_sum__1776_comb + p1_sum__1777_comb;
  assign p1_sum__1345_comb = p1_sum__1778_comb + p1_sum__1779_comb;
  assign p1_sum__1322_comb = p1_sum__1732_comb + p1_sum__1733_comb;
  assign p1_sum__1323_comb = p1_sum__1734_comb + p1_sum__1735_comb;
  assign p1_sum__1308_comb = p1_sum__1704_comb + p1_sum__1705_comb;
  assign p1_sum__1309_comb = p1_sum__1706_comb + p1_sum__1707_comb;
  assign p1_sum__1280_comb = p1_sum__1648_comb + p1_sum__1649_comb;
  assign p1_sum__1281_comb = p1_sum__1650_comb + p1_sum__1651_comb;
  assign p1_sum__1268_comb = p1_sum__1624_comb + p1_sum__1625_comb;
  assign p1_sum__1269_comb = p1_sum__1626_comb + p1_sum__1627_comb;
  assign p1_sum__1346_comb = p1_sum__1780_comb + p1_sum__1781_comb;
  assign p1_sum__1347_comb = p1_sum__1782_comb + p1_sum__1783_comb;
  assign p1_sum__1336_comb = p1_sum__1760_comb + p1_sum__1761_comb;
  assign p1_sum__1337_comb = p1_sum__1762_comb + p1_sum__1763_comb;
  assign p1_sum__1310_comb = p1_sum__1708_comb + p1_sum__1709_comb;
  assign p1_sum__1311_comb = p1_sum__1710_comb + p1_sum__1711_comb;
  assign p1_sum__1296_comb = p1_sum__1680_comb + p1_sum__1681_comb;
  assign p1_sum__1297_comb = p1_sum__1682_comb + p1_sum__1683_comb;
  assign p1_sum__1270_comb = p1_sum__1628_comb + p1_sum__1629_comb;
  assign p1_sum__1271_comb = p1_sum__1630_comb + p1_sum__1631_comb;
  assign p1_sum__1260_comb = p1_sum__1608_comb + p1_sum__1609_comb;
  assign p1_sum__1261_comb = p1_sum__1610_comb + p1_sum__1611_comb;
  assign p1_sum__1338_comb = p1_sum__1764_comb + p1_sum__1765_comb;
  assign p1_sum__1339_comb = p1_sum__1766_comb + p1_sum__1767_comb;
  assign p1_sum__1326_comb = p1_sum__1740_comb + p1_sum__1741_comb;
  assign p1_sum__1327_comb = p1_sum__1742_comb + p1_sum__1743_comb;
  assign p1_sum__1298_comb = p1_sum__1684_comb + p1_sum__1685_comb;
  assign p1_sum__1299_comb = p1_sum__1686_comb + p1_sum__1687_comb;
  assign p1_sum__1284_comb = p1_sum__1656_comb + p1_sum__1657_comb;
  assign p1_sum__1285_comb = p1_sum__1658_comb + p1_sum__1659_comb;
  assign p1_sum__1262_comb = p1_sum__1612_comb + p1_sum__1613_comb;
  assign p1_sum__1263_comb = p1_sum__1614_comb + p1_sum__1615_comb;
  assign p1_sum__1254_comb = p1_sum__1596_comb + p1_sum__1597_comb;
  assign p1_sum__1255_comb = p1_sum__1598_comb + p1_sum__1599_comb;
  assign p1_sum__1328_comb = p1_sum__1744_comb + p1_sum__1745_comb;
  assign p1_sum__1329_comb = p1_sum__1746_comb + p1_sum__1747_comb;
  assign p1_sum__1314_comb = p1_sum__1716_comb + p1_sum__1717_comb;
  assign p1_sum__1315_comb = p1_sum__1718_comb + p1_sum__1719_comb;
  assign p1_sum__1286_comb = p1_sum__1660_comb + p1_sum__1661_comb;
  assign p1_sum__1287_comb = p1_sum__1662_comb + p1_sum__1663_comb;
  assign p1_sum__1274_comb = p1_sum__1636_comb + p1_sum__1637_comb;
  assign p1_sum__1275_comb = p1_sum__1638_comb + p1_sum__1639_comb;
  assign p1_sum__1256_comb = p1_sum__1600_comb + p1_sum__1601_comb;
  assign p1_sum__1257_comb = p1_sum__1602_comb + p1_sum__1603_comb;
  assign p1_sum__1250_comb = p1_sum__1588_comb + p1_sum__1589_comb;
  assign p1_sum__1251_comb = p1_sum__1590_comb + p1_sum__1591_comb;
  assign p1_sum__1316_comb = p1_sum__1720_comb + p1_sum__1721_comb;
  assign p1_sum__1317_comb = p1_sum__1722_comb + p1_sum__1723_comb;
  assign p1_sum__1302_comb = p1_sum__1692_comb + p1_sum__1693_comb;
  assign p1_sum__1303_comb = p1_sum__1694_comb + p1_sum__1695_comb;
  assign p1_sum__1276_comb = p1_sum__1640_comb + p1_sum__1641_comb;
  assign p1_sum__1277_comb = p1_sum__1642_comb + p1_sum__1643_comb;
  assign p1_sum__1266_comb = p1_sum__1620_comb + p1_sum__1621_comb;
  assign p1_sum__1267_comb = p1_sum__1622_comb + p1_sum__1623_comb;
  assign p1_sum__1252_comb = p1_sum__1592_comb + p1_sum__1593_comb;
  assign p1_sum__1253_comb = p1_sum__1594_comb + p1_sum__1595_comb;
  assign p1_sum__1248_comb = p1_sum__1584_comb + p1_sum__1585_comb;
  assign p1_sum__1249_comb = p1_sum__1586_comb + p1_sum__1587_comb;
  assign p1_sum__1130_comb = p1_sum__1348_comb + p1_sum__1349_comb;
  assign p1_sum__1115_comb = p1_sum__1318_comb + p1_sum__1319_comb;
  assign p1_sum__1127_comb = p1_sum__1342_comb + p1_sum__1343_comb;
  assign p1_sum__1109_comb = p1_sum__1306_comb + p1_sum__1307_comb;
  assign p1_sum__1123_comb = p1_sum__1334_comb + p1_sum__1335_comb;
  assign p1_sum__1103_comb = p1_sum__1294_comb + p1_sum__1295_comb;
  assign p1_sum__1118_comb = p1_sum__1324_comb + p1_sum__1325_comb;
  assign p1_sum__1097_comb = p1_sum__1282_comb + p1_sum__1283_comb;
  assign p1_sum__1112_comb = p1_sum__1312_comb + p1_sum__1313_comb;
  assign p1_sum__1092_comb = p1_sum__1272_comb + p1_sum__1273_comb;
  assign p1_sum__1106_comb = p1_sum__1300_comb + p1_sum__1301_comb;
  assign p1_sum__1088_comb = p1_sum__1264_comb + p1_sum__1265_comb;
  assign p1_sum__1100_comb = p1_sum__1288_comb + p1_sum__1289_comb;
  assign p1_sum__1085_comb = p1_sum__1258_comb + p1_sum__1259_comb;
  assign p1_sum__1135_comb = p1_sum__1358_comb + p1_sum__1359_comb;
  assign p1_sum__1133_comb = p1_sum__1354_comb + p1_sum__1355_comb;
  assign p1_sum__1126_comb = p1_sum__1340_comb + p1_sum__1341_comb;
  assign p1_sum__1121_comb = p1_sum__1330_comb + p1_sum__1331_comb;
  assign p1_sum__1108_comb = p1_sum__1304_comb + p1_sum__1305_comb;
  assign p1_sum__1101_comb = p1_sum__1290_comb + p1_sum__1291_comb;
  assign p1_sum__1134_comb = p1_sum__1356_comb + p1_sum__1357_comb;
  assign p1_sum__1131_comb = p1_sum__1350_comb + p1_sum__1351_comb;
  assign p1_sum__1122_comb = p1_sum__1332_comb + p1_sum__1333_comb;
  assign p1_sum__1116_comb = p1_sum__1320_comb + p1_sum__1321_comb;
  assign p1_sum__1102_comb = p1_sum__1292_comb + p1_sum__1293_comb;
  assign p1_sum__1095_comb = p1_sum__1278_comb + p1_sum__1279_comb;
  assign p1_sum__1132_comb = p1_sum__1352_comb + p1_sum__1353_comb;
  assign p1_sum__1128_comb = p1_sum__1344_comb + p1_sum__1345_comb;
  assign p1_sum__1117_comb = p1_sum__1322_comb + p1_sum__1323_comb;
  assign p1_sum__1110_comb = p1_sum__1308_comb + p1_sum__1309_comb;
  assign p1_sum__1096_comb = p1_sum__1280_comb + p1_sum__1281_comb;
  assign p1_sum__1090_comb = p1_sum__1268_comb + p1_sum__1269_comb;
  assign p1_sum__1129_comb = p1_sum__1346_comb + p1_sum__1347_comb;
  assign p1_sum__1124_comb = p1_sum__1336_comb + p1_sum__1337_comb;
  assign p1_sum__1111_comb = p1_sum__1310_comb + p1_sum__1311_comb;
  assign p1_sum__1104_comb = p1_sum__1296_comb + p1_sum__1297_comb;
  assign p1_sum__1091_comb = p1_sum__1270_comb + p1_sum__1271_comb;
  assign p1_sum__1086_comb = p1_sum__1260_comb + p1_sum__1261_comb;
  assign p1_sum__1125_comb = p1_sum__1338_comb + p1_sum__1339_comb;
  assign p1_sum__1119_comb = p1_sum__1326_comb + p1_sum__1327_comb;
  assign p1_sum__1105_comb = p1_sum__1298_comb + p1_sum__1299_comb;
  assign p1_sum__1098_comb = p1_sum__1284_comb + p1_sum__1285_comb;
  assign p1_sum__1087_comb = p1_sum__1262_comb + p1_sum__1263_comb;
  assign p1_sum__1083_comb = p1_sum__1254_comb + p1_sum__1255_comb;
  assign p1_sum__1120_comb = p1_sum__1328_comb + p1_sum__1329_comb;
  assign p1_sum__1113_comb = p1_sum__1314_comb + p1_sum__1315_comb;
  assign p1_sum__1099_comb = p1_sum__1286_comb + p1_sum__1287_comb;
  assign p1_sum__1093_comb = p1_sum__1274_comb + p1_sum__1275_comb;
  assign p1_sum__1084_comb = p1_sum__1256_comb + p1_sum__1257_comb;
  assign p1_sum__1081_comb = p1_sum__1250_comb + p1_sum__1251_comb;
  assign p1_sum__1114_comb = p1_sum__1316_comb + p1_sum__1317_comb;
  assign p1_sum__1107_comb = p1_sum__1302_comb + p1_sum__1303_comb;
  assign p1_sum__1094_comb = p1_sum__1276_comb + p1_sum__1277_comb;
  assign p1_sum__1089_comb = p1_sum__1266_comb + p1_sum__1267_comb;
  assign p1_sum__1082_comb = p1_sum__1252_comb + p1_sum__1253_comb;
  assign p1_sum__1080_comb = p1_sum__1248_comb + p1_sum__1249_comb;
  assign p1_add_143035_comb = p1_umul_142787_comb[31:7] + 25'h000_0001;
  assign p1_add_143036_comb = p1_umul_142788_comb[31:7] + 25'h000_0001;
  assign p1_add_143037_comb = p1_sum__1130_comb + 25'h000_0001;
  assign p1_add_143038_comb = p1_sum__1115_comb + 25'h000_0001;
  assign p1_add_143039_comb = p1_sum__1127_comb + 25'h000_0001;
  assign p1_add_143040_comb = p1_sum__1109_comb + 25'h000_0001;
  assign p1_add_143041_comb = p1_sum__1123_comb + 25'h000_0001;
  assign p1_add_143042_comb = p1_sum__1103_comb + 25'h000_0001;
  assign p1_add_143043_comb = p1_sum__1118_comb + 25'h000_0001;
  assign p1_add_143044_comb = p1_sum__1097_comb + 25'h000_0001;
  assign p1_add_143045_comb = p1_sum__1112_comb + 25'h000_0001;
  assign p1_add_143046_comb = p1_sum__1092_comb + 25'h000_0001;
  assign p1_add_143047_comb = p1_sum__1106_comb + 25'h000_0001;
  assign p1_add_143048_comb = p1_sum__1088_comb + 25'h000_0001;
  assign p1_add_143049_comb = p1_sum__1100_comb + 25'h000_0001;
  assign p1_add_143050_comb = p1_sum__1085_comb + 25'h000_0001;
  assign p1_add_143051_comb = p1_umul_142817_comb[31:7] + 25'h000_0001;
  assign p1_add_143052_comb = p1_umul_142818_comb[31:7] + 25'h000_0001;
  assign p1_add_143053_comb = p1_umul_142819_comb[31:7] + 25'h000_0001;
  assign p1_add_143054_comb = p1_umul_142820_comb[31:7] + 25'h000_0001;
  assign p1_add_143055_comb = p1_umul_142821_comb[31:7] + 25'h000_0001;
  assign p1_add_143056_comb = p1_umul_142822_comb[31:7] + 25'h000_0001;
  assign p1_add_143057_comb = p1_sum__1135_comb + 25'h000_0001;
  assign p1_add_143058_comb = p1_sum__1133_comb + 25'h000_0001;
  assign p1_add_143059_comb = p1_sum__1126_comb + 25'h000_0001;
  assign p1_add_143060_comb = p1_sum__1121_comb + 25'h000_0001;
  assign p1_add_143061_comb = p1_sum__1108_comb + 25'h000_0001;
  assign p1_add_143062_comb = p1_sum__1101_comb + 25'h000_0001;
  assign p1_add_143063_comb = p1_sum__1134_comb + 25'h000_0001;
  assign p1_add_143064_comb = p1_sum__1131_comb + 25'h000_0001;
  assign p1_add_143065_comb = p1_sum__1122_comb + 25'h000_0001;
  assign p1_add_143066_comb = p1_sum__1116_comb + 25'h000_0001;
  assign p1_add_143067_comb = p1_sum__1102_comb + 25'h000_0001;
  assign p1_add_143068_comb = p1_sum__1095_comb + 25'h000_0001;
  assign p1_add_143069_comb = p1_sum__1132_comb + 25'h000_0001;
  assign p1_add_143070_comb = p1_sum__1128_comb + 25'h000_0001;
  assign p1_add_143071_comb = p1_sum__1117_comb + 25'h000_0001;
  assign p1_add_143072_comb = p1_sum__1110_comb + 25'h000_0001;
  assign p1_add_143073_comb = p1_sum__1096_comb + 25'h000_0001;
  assign p1_add_143074_comb = p1_sum__1090_comb + 25'h000_0001;
  assign p1_add_143075_comb = p1_sum__1129_comb + 25'h000_0001;
  assign p1_add_143076_comb = p1_sum__1124_comb + 25'h000_0001;
  assign p1_add_143077_comb = p1_sum__1111_comb + 25'h000_0001;
  assign p1_add_143078_comb = p1_sum__1104_comb + 25'h000_0001;
  assign p1_add_143079_comb = p1_sum__1091_comb + 25'h000_0001;
  assign p1_add_143080_comb = p1_sum__1086_comb + 25'h000_0001;
  assign p1_add_143081_comb = p1_sum__1125_comb + 25'h000_0001;
  assign p1_add_143082_comb = p1_sum__1119_comb + 25'h000_0001;
  assign p1_add_143083_comb = p1_sum__1105_comb + 25'h000_0001;
  assign p1_add_143084_comb = p1_sum__1098_comb + 25'h000_0001;
  assign p1_add_143085_comb = p1_sum__1087_comb + 25'h000_0001;
  assign p1_add_143086_comb = p1_sum__1083_comb + 25'h000_0001;
  assign p1_add_143087_comb = p1_sum__1120_comb + 25'h000_0001;
  assign p1_add_143088_comb = p1_sum__1113_comb + 25'h000_0001;
  assign p1_add_143089_comb = p1_sum__1099_comb + 25'h000_0001;
  assign p1_add_143090_comb = p1_sum__1093_comb + 25'h000_0001;
  assign p1_add_143091_comb = p1_sum__1084_comb + 25'h000_0001;
  assign p1_add_143092_comb = p1_sum__1081_comb + 25'h000_0001;
  assign p1_add_143093_comb = p1_sum__1114_comb + 25'h000_0001;
  assign p1_add_143094_comb = p1_sum__1107_comb + 25'h000_0001;
  assign p1_add_143095_comb = p1_sum__1094_comb + 25'h000_0001;
  assign p1_add_143096_comb = p1_sum__1089_comb + 25'h000_0001;
  assign p1_add_143097_comb = p1_sum__1082_comb + 25'h000_0001;
  assign p1_add_143098_comb = p1_sum__1080_comb + 25'h000_0001;
  assign p1_clipped__256_comb = $signed(p1_add_143035_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143035_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143035_comb[16:8]);
  assign p1_clipped__259_comb = $signed(p1_add_143036_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143036_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143036_comb[16:8]);
  assign p1_clipped__260_comb = $signed(p1_add_143037_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143037_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143037_comb[16:8]);
  assign p1_clipped__263_comb = $signed(p1_add_143038_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143038_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143038_comb[16:8]);
  assign p1_clipped__264_comb = $signed(p1_add_143039_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143039_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143039_comb[16:8]);
  assign p1_clipped__267_comb = $signed(p1_add_143040_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143040_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143040_comb[16:8]);
  assign p1_clipped__268_comb = $signed(p1_add_143041_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143041_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143041_comb[16:8]);
  assign p1_clipped__271_comb = $signed(p1_add_143042_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143042_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143042_comb[16:8]);
  assign p1_clipped__272_comb = $signed(p1_add_143043_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143043_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143043_comb[16:8]);
  assign p1_clipped__275_comb = $signed(p1_add_143044_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143044_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143044_comb[16:8]);
  assign p1_clipped__276_comb = $signed(p1_add_143045_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143045_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143045_comb[16:8]);
  assign p1_clipped__279_comb = $signed(p1_add_143046_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143046_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143046_comb[16:8]);
  assign p1_clipped__280_comb = $signed(p1_add_143047_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143047_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143047_comb[16:8]);
  assign p1_clipped__283_comb = $signed(p1_add_143048_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143048_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143048_comb[16:8]);
  assign p1_clipped__284_comb = $signed(p1_add_143049_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143049_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143049_comb[16:8]);
  assign p1_clipped__287_comb = $signed(p1_add_143050_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143050_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143050_comb[16:8]);
  assign p1_clipped__288_comb = $signed(p1_add_143051_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143051_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143051_comb[16:8]);
  assign p1_clipped__289_comb = $signed(p1_add_143052_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143052_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143052_comb[16:8]);
  assign p1_clipped__257_comb = $signed(p1_add_143053_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143053_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143053_comb[16:8]);
  assign p1_clipped__258_comb = $signed(p1_add_143054_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143054_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143054_comb[16:8]);
  assign p1_clipped__290_comb = $signed(p1_add_143055_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143055_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143055_comb[16:8]);
  assign p1_clipped__291_comb = $signed(p1_add_143056_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143056_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143056_comb[16:8]);
  assign p1_clipped__292_comb = $signed(p1_add_143057_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143057_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143057_comb[16:8]);
  assign p1_clipped__293_comb = $signed(p1_add_143058_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143058_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143058_comb[16:8]);
  assign p1_clipped__261_comb = $signed(p1_add_143059_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143059_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143059_comb[16:8]);
  assign p1_clipped__262_comb = $signed(p1_add_143060_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143060_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143060_comb[16:8]);
  assign p1_clipped__294_comb = $signed(p1_add_143061_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143061_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143061_comb[16:8]);
  assign p1_clipped__295_comb = $signed(p1_add_143062_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143062_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143062_comb[16:8]);
  assign p1_clipped__296_comb = $signed(p1_add_143063_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143063_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143063_comb[16:8]);
  assign p1_clipped__297_comb = $signed(p1_add_143064_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143064_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143064_comb[16:8]);
  assign p1_clipped__265_comb = $signed(p1_add_143065_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143065_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143065_comb[16:8]);
  assign p1_clipped__266_comb = $signed(p1_add_143066_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143066_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143066_comb[16:8]);
  assign p1_clipped__298_comb = $signed(p1_add_143067_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143067_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143067_comb[16:8]);
  assign p1_clipped__299_comb = $signed(p1_add_143068_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143068_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143068_comb[16:8]);
  assign p1_clipped__300_comb = $signed(p1_add_143069_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143069_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143069_comb[16:8]);
  assign p1_clipped__301_comb = $signed(p1_add_143070_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143070_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143070_comb[16:8]);
  assign p1_clipped__269_comb = $signed(p1_add_143071_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143071_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143071_comb[16:8]);
  assign p1_clipped__270_comb = $signed(p1_add_143072_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143072_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143072_comb[16:8]);
  assign p1_clipped__302_comb = $signed(p1_add_143073_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143073_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143073_comb[16:8]);
  assign p1_clipped__303_comb = $signed(p1_add_143074_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143074_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143074_comb[16:8]);
  assign p1_clipped__304_comb = $signed(p1_add_143075_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143075_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143075_comb[16:8]);
  assign p1_clipped__305_comb = $signed(p1_add_143076_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143076_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143076_comb[16:8]);
  assign p1_clipped__273_comb = $signed(p1_add_143077_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143077_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143077_comb[16:8]);
  assign p1_clipped__274_comb = $signed(p1_add_143078_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143078_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143078_comb[16:8]);
  assign p1_clipped__306_comb = $signed(p1_add_143079_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143079_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143079_comb[16:8]);
  assign p1_clipped__307_comb = $signed(p1_add_143080_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143080_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143080_comb[16:8]);
  assign p1_clipped__308_comb = $signed(p1_add_143081_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143081_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143081_comb[16:8]);
  assign p1_clipped__309_comb = $signed(p1_add_143082_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143082_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143082_comb[16:8]);
  assign p1_clipped__277_comb = $signed(p1_add_143083_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143083_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143083_comb[16:8]);
  assign p1_clipped__278_comb = $signed(p1_add_143084_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143084_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143084_comb[16:8]);
  assign p1_clipped__310_comb = $signed(p1_add_143085_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143085_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143085_comb[16:8]);
  assign p1_clipped__311_comb = $signed(p1_add_143086_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143086_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143086_comb[16:8]);
  assign p1_clipped__312_comb = $signed(p1_add_143087_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143087_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143087_comb[16:8]);
  assign p1_clipped__313_comb = $signed(p1_add_143088_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143088_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143088_comb[16:8]);
  assign p1_clipped__281_comb = $signed(p1_add_143089_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143089_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143089_comb[16:8]);
  assign p1_clipped__282_comb = $signed(p1_add_143090_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143090_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143090_comb[16:8]);
  assign p1_clipped__314_comb = $signed(p1_add_143091_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143091_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143091_comb[16:8]);
  assign p1_clipped__315_comb = $signed(p1_add_143092_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143092_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143092_comb[16:8]);
  assign p1_clipped__316_comb = $signed(p1_add_143093_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143093_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143093_comb[16:8]);
  assign p1_clipped__317_comb = $signed(p1_add_143094_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143094_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143094_comb[16:8]);
  assign p1_clipped__285_comb = $signed(p1_add_143095_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143095_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143095_comb[16:8]);
  assign p1_clipped__286_comb = $signed(p1_add_143096_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143096_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143096_comb[16:8]);
  assign p1_clipped__318_comb = $signed(p1_add_143097_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143097_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143097_comb[16:8]);
  assign p1_clipped__319_comb = $signed(p1_add_143098_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_143098_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_143098_comb[16:8]);
  assign p1_add_143867_comb = {{1{p1_clipped__256_comb[8]}}, p1_clipped__256_comb} + 10'h001;
  assign p1_add_143868_comb = {{1{p1_clipped__259_comb[8]}}, p1_clipped__259_comb} + 10'h001;
  assign p1_add_143869_comb = {{1{p1_clipped__260_comb[8]}}, p1_clipped__260_comb} + 10'h001;
  assign p1_add_143870_comb = {{1{p1_clipped__263_comb[8]}}, p1_clipped__263_comb} + 10'h001;
  assign p1_add_143871_comb = {{1{p1_clipped__264_comb[8]}}, p1_clipped__264_comb} + 10'h001;
  assign p1_add_143872_comb = {{1{p1_clipped__267_comb[8]}}, p1_clipped__267_comb} + 10'h001;
  assign p1_add_143873_comb = {{1{p1_clipped__268_comb[8]}}, p1_clipped__268_comb} + 10'h001;
  assign p1_add_143874_comb = {{1{p1_clipped__271_comb[8]}}, p1_clipped__271_comb} + 10'h001;
  assign p1_add_143875_comb = {{1{p1_clipped__272_comb[8]}}, p1_clipped__272_comb} + 10'h001;
  assign p1_add_143876_comb = {{1{p1_clipped__275_comb[8]}}, p1_clipped__275_comb} + 10'h001;
  assign p1_add_143877_comb = {{1{p1_clipped__276_comb[8]}}, p1_clipped__276_comb} + 10'h001;
  assign p1_add_143878_comb = {{1{p1_clipped__279_comb[8]}}, p1_clipped__279_comb} + 10'h001;
  assign p1_add_143879_comb = {{1{p1_clipped__280_comb[8]}}, p1_clipped__280_comb} + 10'h001;
  assign p1_add_143880_comb = {{1{p1_clipped__283_comb[8]}}, p1_clipped__283_comb} + 10'h001;
  assign p1_add_143881_comb = {{1{p1_clipped__284_comb[8]}}, p1_clipped__284_comb} + 10'h001;
  assign p1_add_143882_comb = {{1{p1_clipped__287_comb[8]}}, p1_clipped__287_comb} + 10'h001;
  assign p1_add_143883_comb = {{1{p1_clipped__288_comb[8]}}, p1_clipped__288_comb} + 10'h001;
  assign p1_add_143884_comb = {{1{p1_clipped__289_comb[8]}}, p1_clipped__289_comb} + 10'h001;
  assign p1_add_143885_comb = {{1{p1_clipped__257_comb[8]}}, p1_clipped__257_comb} + 10'h001;
  assign p1_add_143886_comb = {{1{p1_clipped__258_comb[8]}}, p1_clipped__258_comb} + 10'h001;
  assign p1_add_143887_comb = {{1{p1_clipped__290_comb[8]}}, p1_clipped__290_comb} + 10'h001;
  assign p1_add_143888_comb = {{1{p1_clipped__291_comb[8]}}, p1_clipped__291_comb} + 10'h001;
  assign p1_add_143889_comb = {{1{p1_clipped__292_comb[8]}}, p1_clipped__292_comb} + 10'h001;
  assign p1_add_143890_comb = {{1{p1_clipped__293_comb[8]}}, p1_clipped__293_comb} + 10'h001;
  assign p1_add_143891_comb = {{1{p1_clipped__261_comb[8]}}, p1_clipped__261_comb} + 10'h001;
  assign p1_add_143892_comb = {{1{p1_clipped__262_comb[8]}}, p1_clipped__262_comb} + 10'h001;
  assign p1_add_143893_comb = {{1{p1_clipped__294_comb[8]}}, p1_clipped__294_comb} + 10'h001;
  assign p1_add_143894_comb = {{1{p1_clipped__295_comb[8]}}, p1_clipped__295_comb} + 10'h001;
  assign p1_add_143895_comb = {{1{p1_clipped__296_comb[8]}}, p1_clipped__296_comb} + 10'h001;
  assign p1_add_143896_comb = {{1{p1_clipped__297_comb[8]}}, p1_clipped__297_comb} + 10'h001;
  assign p1_add_143897_comb = {{1{p1_clipped__265_comb[8]}}, p1_clipped__265_comb} + 10'h001;
  assign p1_add_143898_comb = {{1{p1_clipped__266_comb[8]}}, p1_clipped__266_comb} + 10'h001;
  assign p1_add_143899_comb = {{1{p1_clipped__298_comb[8]}}, p1_clipped__298_comb} + 10'h001;
  assign p1_add_143900_comb = {{1{p1_clipped__299_comb[8]}}, p1_clipped__299_comb} + 10'h001;
  assign p1_add_143901_comb = {{1{p1_clipped__300_comb[8]}}, p1_clipped__300_comb} + 10'h001;
  assign p1_add_143902_comb = {{1{p1_clipped__301_comb[8]}}, p1_clipped__301_comb} + 10'h001;
  assign p1_add_143903_comb = {{1{p1_clipped__269_comb[8]}}, p1_clipped__269_comb} + 10'h001;
  assign p1_add_143904_comb = {{1{p1_clipped__270_comb[8]}}, p1_clipped__270_comb} + 10'h001;
  assign p1_add_143905_comb = {{1{p1_clipped__302_comb[8]}}, p1_clipped__302_comb} + 10'h001;
  assign p1_add_143906_comb = {{1{p1_clipped__303_comb[8]}}, p1_clipped__303_comb} + 10'h001;
  assign p1_add_143907_comb = {{1{p1_clipped__304_comb[8]}}, p1_clipped__304_comb} + 10'h001;
  assign p1_add_143908_comb = {{1{p1_clipped__305_comb[8]}}, p1_clipped__305_comb} + 10'h001;
  assign p1_add_143909_comb = {{1{p1_clipped__273_comb[8]}}, p1_clipped__273_comb} + 10'h001;
  assign p1_add_143910_comb = {{1{p1_clipped__274_comb[8]}}, p1_clipped__274_comb} + 10'h001;
  assign p1_add_143911_comb = {{1{p1_clipped__306_comb[8]}}, p1_clipped__306_comb} + 10'h001;
  assign p1_add_143912_comb = {{1{p1_clipped__307_comb[8]}}, p1_clipped__307_comb} + 10'h001;
  assign p1_add_143913_comb = {{1{p1_clipped__308_comb[8]}}, p1_clipped__308_comb} + 10'h001;
  assign p1_add_143914_comb = {{1{p1_clipped__309_comb[8]}}, p1_clipped__309_comb} + 10'h001;
  assign p1_add_143915_comb = {{1{p1_clipped__277_comb[8]}}, p1_clipped__277_comb} + 10'h001;
  assign p1_add_143916_comb = {{1{p1_clipped__278_comb[8]}}, p1_clipped__278_comb} + 10'h001;
  assign p1_add_143917_comb = {{1{p1_clipped__310_comb[8]}}, p1_clipped__310_comb} + 10'h001;
  assign p1_add_143918_comb = {{1{p1_clipped__311_comb[8]}}, p1_clipped__311_comb} + 10'h001;
  assign p1_add_143919_comb = {{1{p1_clipped__312_comb[8]}}, p1_clipped__312_comb} + 10'h001;
  assign p1_add_143920_comb = {{1{p1_clipped__313_comb[8]}}, p1_clipped__313_comb} + 10'h001;
  assign p1_add_143921_comb = {{1{p1_clipped__281_comb[8]}}, p1_clipped__281_comb} + 10'h001;
  assign p1_add_143922_comb = {{1{p1_clipped__282_comb[8]}}, p1_clipped__282_comb} + 10'h001;
  assign p1_add_143923_comb = {{1{p1_clipped__314_comb[8]}}, p1_clipped__314_comb} + 10'h001;
  assign p1_add_143924_comb = {{1{p1_clipped__315_comb[8]}}, p1_clipped__315_comb} + 10'h001;
  assign p1_add_143925_comb = {{1{p1_clipped__316_comb[8]}}, p1_clipped__316_comb} + 10'h001;
  assign p1_add_143926_comb = {{1{p1_clipped__317_comb[8]}}, p1_clipped__317_comb} + 10'h001;
  assign p1_add_143927_comb = {{1{p1_clipped__285_comb[8]}}, p1_clipped__285_comb} + 10'h001;
  assign p1_add_143928_comb = {{1{p1_clipped__286_comb[8]}}, p1_clipped__286_comb} + 10'h001;
  assign p1_add_143929_comb = {{1{p1_clipped__318_comb[8]}}, p1_clipped__318_comb} + 10'h001;
  assign p1_add_143930_comb = {{1{p1_clipped__319_comb[8]}}, p1_clipped__319_comb} + 10'h001;
  assign p1_bit_slice_143931_comb = p1_add_143867_comb[9:8];
  assign p1_bit_slice_143932_comb = p1_add_143868_comb[9:8];
  assign p1_bit_slice_143933_comb = p1_add_143869_comb[9:8];
  assign p1_bit_slice_143934_comb = p1_add_143870_comb[9:8];
  assign p1_bit_slice_143935_comb = p1_add_143871_comb[9:8];
  assign p1_bit_slice_143936_comb = p1_add_143872_comb[9:8];
  assign p1_bit_slice_143937_comb = p1_add_143873_comb[9:8];
  assign p1_bit_slice_143938_comb = p1_add_143874_comb[9:8];
  assign p1_bit_slice_143939_comb = p1_add_143875_comb[9:8];
  assign p1_bit_slice_143940_comb = p1_add_143876_comb[9:8];
  assign p1_bit_slice_143941_comb = p1_add_143877_comb[9:8];
  assign p1_bit_slice_143942_comb = p1_add_143878_comb[9:8];
  assign p1_bit_slice_143943_comb = p1_add_143879_comb[9:8];
  assign p1_bit_slice_143944_comb = p1_add_143880_comb[9:8];
  assign p1_bit_slice_143945_comb = p1_add_143881_comb[9:8];
  assign p1_bit_slice_143946_comb = p1_add_143882_comb[9:8];
  assign p1_bit_slice_143947_comb = p1_add_143883_comb[9:8];
  assign p1_bit_slice_143948_comb = p1_add_143884_comb[9:8];
  assign p1_bit_slice_143949_comb = p1_add_143885_comb[9:8];
  assign p1_bit_slice_143950_comb = p1_add_143886_comb[9:8];
  assign p1_bit_slice_143951_comb = p1_add_143887_comb[9:8];
  assign p1_bit_slice_143952_comb = p1_add_143888_comb[9:8];
  assign p1_bit_slice_143953_comb = p1_add_143889_comb[9:8];
  assign p1_bit_slice_143954_comb = p1_add_143890_comb[9:8];
  assign p1_bit_slice_143955_comb = p1_add_143891_comb[9:8];
  assign p1_bit_slice_143956_comb = p1_add_143892_comb[9:8];
  assign p1_bit_slice_143957_comb = p1_add_143893_comb[9:8];
  assign p1_bit_slice_143958_comb = p1_add_143894_comb[9:8];
  assign p1_bit_slice_143959_comb = p1_add_143895_comb[9:8];
  assign p1_bit_slice_143960_comb = p1_add_143896_comb[9:8];
  assign p1_bit_slice_143961_comb = p1_add_143897_comb[9:8];
  assign p1_bit_slice_143962_comb = p1_add_143898_comb[9:8];
  assign p1_bit_slice_143963_comb = p1_add_143899_comb[9:8];
  assign p1_bit_slice_143964_comb = p1_add_143900_comb[9:8];
  assign p1_bit_slice_143965_comb = p1_add_143901_comb[9:8];
  assign p1_bit_slice_143966_comb = p1_add_143902_comb[9:8];
  assign p1_bit_slice_143967_comb = p1_add_143903_comb[9:8];
  assign p1_bit_slice_143968_comb = p1_add_143904_comb[9:8];
  assign p1_bit_slice_143969_comb = p1_add_143905_comb[9:8];
  assign p1_bit_slice_143970_comb = p1_add_143906_comb[9:8];
  assign p1_bit_slice_143971_comb = p1_add_143907_comb[9:8];
  assign p1_bit_slice_143972_comb = p1_add_143908_comb[9:8];
  assign p1_bit_slice_143973_comb = p1_add_143909_comb[9:8];
  assign p1_bit_slice_143974_comb = p1_add_143910_comb[9:8];
  assign p1_bit_slice_143975_comb = p1_add_143911_comb[9:8];
  assign p1_bit_slice_143976_comb = p1_add_143912_comb[9:8];
  assign p1_bit_slice_143977_comb = p1_add_143913_comb[9:8];
  assign p1_bit_slice_143978_comb = p1_add_143914_comb[9:8];
  assign p1_bit_slice_143979_comb = p1_add_143915_comb[9:8];
  assign p1_bit_slice_143980_comb = p1_add_143916_comb[9:8];
  assign p1_bit_slice_143981_comb = p1_add_143917_comb[9:8];
  assign p1_bit_slice_143982_comb = p1_add_143918_comb[9:8];
  assign p1_bit_slice_143983_comb = p1_add_143919_comb[9:8];
  assign p1_bit_slice_143984_comb = p1_add_143920_comb[9:8];
  assign p1_bit_slice_143985_comb = p1_add_143921_comb[9:8];
  assign p1_bit_slice_143986_comb = p1_add_143922_comb[9:8];
  assign p1_bit_slice_143987_comb = p1_add_143923_comb[9:8];
  assign p1_bit_slice_143988_comb = p1_add_143924_comb[9:8];
  assign p1_bit_slice_143989_comb = p1_add_143925_comb[9:8];
  assign p1_bit_slice_143990_comb = p1_add_143926_comb[9:8];
  assign p1_bit_slice_143991_comb = p1_add_143927_comb[9:8];
  assign p1_bit_slice_143992_comb = p1_add_143928_comb[9:8];
  assign p1_bit_slice_143993_comb = p1_add_143929_comb[9:8];
  assign p1_bit_slice_143994_comb = p1_add_143930_comb[9:8];
  assign p1_add_144123_comb = {{1{p1_bit_slice_143931_comb[1]}}, p1_bit_slice_143931_comb} + 3'h1;
  assign p1_add_144124_comb = {{1{p1_bit_slice_143932_comb[1]}}, p1_bit_slice_143932_comb} + 3'h1;
  assign p1_add_144125_comb = {{1{p1_bit_slice_143933_comb[1]}}, p1_bit_slice_143933_comb} + 3'h1;
  assign p1_add_144126_comb = {{1{p1_bit_slice_143934_comb[1]}}, p1_bit_slice_143934_comb} + 3'h1;
  assign p1_add_144127_comb = {{1{p1_bit_slice_143935_comb[1]}}, p1_bit_slice_143935_comb} + 3'h1;
  assign p1_add_144128_comb = {{1{p1_bit_slice_143936_comb[1]}}, p1_bit_slice_143936_comb} + 3'h1;
  assign p1_add_144129_comb = {{1{p1_bit_slice_143937_comb[1]}}, p1_bit_slice_143937_comb} + 3'h1;
  assign p1_add_144130_comb = {{1{p1_bit_slice_143938_comb[1]}}, p1_bit_slice_143938_comb} + 3'h1;
  assign p1_add_144131_comb = {{1{p1_bit_slice_143939_comb[1]}}, p1_bit_slice_143939_comb} + 3'h1;
  assign p1_add_144132_comb = {{1{p1_bit_slice_143940_comb[1]}}, p1_bit_slice_143940_comb} + 3'h1;
  assign p1_add_144133_comb = {{1{p1_bit_slice_143941_comb[1]}}, p1_bit_slice_143941_comb} + 3'h1;
  assign p1_add_144134_comb = {{1{p1_bit_slice_143942_comb[1]}}, p1_bit_slice_143942_comb} + 3'h1;
  assign p1_add_144135_comb = {{1{p1_bit_slice_143943_comb[1]}}, p1_bit_slice_143943_comb} + 3'h1;
  assign p1_add_144136_comb = {{1{p1_bit_slice_143944_comb[1]}}, p1_bit_slice_143944_comb} + 3'h1;
  assign p1_add_144137_comb = {{1{p1_bit_slice_143945_comb[1]}}, p1_bit_slice_143945_comb} + 3'h1;
  assign p1_add_144138_comb = {{1{p1_bit_slice_143946_comb[1]}}, p1_bit_slice_143946_comb} + 3'h1;
  assign p1_add_144139_comb = {{1{p1_bit_slice_143947_comb[1]}}, p1_bit_slice_143947_comb} + 3'h1;
  assign p1_add_144140_comb = {{1{p1_bit_slice_143948_comb[1]}}, p1_bit_slice_143948_comb} + 3'h1;
  assign p1_add_144141_comb = {{1{p1_bit_slice_143949_comb[1]}}, p1_bit_slice_143949_comb} + 3'h1;
  assign p1_add_144142_comb = {{1{p1_bit_slice_143950_comb[1]}}, p1_bit_slice_143950_comb} + 3'h1;
  assign p1_add_144143_comb = {{1{p1_bit_slice_143951_comb[1]}}, p1_bit_slice_143951_comb} + 3'h1;
  assign p1_add_144144_comb = {{1{p1_bit_slice_143952_comb[1]}}, p1_bit_slice_143952_comb} + 3'h1;
  assign p1_add_144145_comb = {{1{p1_bit_slice_143953_comb[1]}}, p1_bit_slice_143953_comb} + 3'h1;
  assign p1_add_144146_comb = {{1{p1_bit_slice_143954_comb[1]}}, p1_bit_slice_143954_comb} + 3'h1;
  assign p1_add_144147_comb = {{1{p1_bit_slice_143955_comb[1]}}, p1_bit_slice_143955_comb} + 3'h1;
  assign p1_add_144148_comb = {{1{p1_bit_slice_143956_comb[1]}}, p1_bit_slice_143956_comb} + 3'h1;
  assign p1_add_144149_comb = {{1{p1_bit_slice_143957_comb[1]}}, p1_bit_slice_143957_comb} + 3'h1;
  assign p1_add_144150_comb = {{1{p1_bit_slice_143958_comb[1]}}, p1_bit_slice_143958_comb} + 3'h1;
  assign p1_add_144151_comb = {{1{p1_bit_slice_143959_comb[1]}}, p1_bit_slice_143959_comb} + 3'h1;
  assign p1_add_144152_comb = {{1{p1_bit_slice_143960_comb[1]}}, p1_bit_slice_143960_comb} + 3'h1;
  assign p1_add_144153_comb = {{1{p1_bit_slice_143961_comb[1]}}, p1_bit_slice_143961_comb} + 3'h1;
  assign p1_add_144154_comb = {{1{p1_bit_slice_143962_comb[1]}}, p1_bit_slice_143962_comb} + 3'h1;
  assign p1_add_144155_comb = {{1{p1_bit_slice_143963_comb[1]}}, p1_bit_slice_143963_comb} + 3'h1;
  assign p1_add_144156_comb = {{1{p1_bit_slice_143964_comb[1]}}, p1_bit_slice_143964_comb} + 3'h1;
  assign p1_add_144157_comb = {{1{p1_bit_slice_143965_comb[1]}}, p1_bit_slice_143965_comb} + 3'h1;
  assign p1_add_144158_comb = {{1{p1_bit_slice_143966_comb[1]}}, p1_bit_slice_143966_comb} + 3'h1;
  assign p1_add_144159_comb = {{1{p1_bit_slice_143967_comb[1]}}, p1_bit_slice_143967_comb} + 3'h1;
  assign p1_add_144160_comb = {{1{p1_bit_slice_143968_comb[1]}}, p1_bit_slice_143968_comb} + 3'h1;
  assign p1_add_144161_comb = {{1{p1_bit_slice_143969_comb[1]}}, p1_bit_slice_143969_comb} + 3'h1;
  assign p1_add_144162_comb = {{1{p1_bit_slice_143970_comb[1]}}, p1_bit_slice_143970_comb} + 3'h1;
  assign p1_add_144163_comb = {{1{p1_bit_slice_143971_comb[1]}}, p1_bit_slice_143971_comb} + 3'h1;
  assign p1_add_144164_comb = {{1{p1_bit_slice_143972_comb[1]}}, p1_bit_slice_143972_comb} + 3'h1;
  assign p1_add_144165_comb = {{1{p1_bit_slice_143973_comb[1]}}, p1_bit_slice_143973_comb} + 3'h1;
  assign p1_add_144166_comb = {{1{p1_bit_slice_143974_comb[1]}}, p1_bit_slice_143974_comb} + 3'h1;
  assign p1_add_144167_comb = {{1{p1_bit_slice_143975_comb[1]}}, p1_bit_slice_143975_comb} + 3'h1;
  assign p1_add_144168_comb = {{1{p1_bit_slice_143976_comb[1]}}, p1_bit_slice_143976_comb} + 3'h1;
  assign p1_add_144169_comb = {{1{p1_bit_slice_143977_comb[1]}}, p1_bit_slice_143977_comb} + 3'h1;
  assign p1_add_144170_comb = {{1{p1_bit_slice_143978_comb[1]}}, p1_bit_slice_143978_comb} + 3'h1;
  assign p1_add_144171_comb = {{1{p1_bit_slice_143979_comb[1]}}, p1_bit_slice_143979_comb} + 3'h1;
  assign p1_add_144172_comb = {{1{p1_bit_slice_143980_comb[1]}}, p1_bit_slice_143980_comb} + 3'h1;
  assign p1_add_144173_comb = {{1{p1_bit_slice_143981_comb[1]}}, p1_bit_slice_143981_comb} + 3'h1;
  assign p1_add_144174_comb = {{1{p1_bit_slice_143982_comb[1]}}, p1_bit_slice_143982_comb} + 3'h1;
  assign p1_add_144175_comb = {{1{p1_bit_slice_143983_comb[1]}}, p1_bit_slice_143983_comb} + 3'h1;
  assign p1_add_144176_comb = {{1{p1_bit_slice_143984_comb[1]}}, p1_bit_slice_143984_comb} + 3'h1;
  assign p1_add_144177_comb = {{1{p1_bit_slice_143985_comb[1]}}, p1_bit_slice_143985_comb} + 3'h1;
  assign p1_add_144178_comb = {{1{p1_bit_slice_143986_comb[1]}}, p1_bit_slice_143986_comb} + 3'h1;
  assign p1_add_144179_comb = {{1{p1_bit_slice_143987_comb[1]}}, p1_bit_slice_143987_comb} + 3'h1;
  assign p1_add_144180_comb = {{1{p1_bit_slice_143988_comb[1]}}, p1_bit_slice_143988_comb} + 3'h1;
  assign p1_add_144181_comb = {{1{p1_bit_slice_143989_comb[1]}}, p1_bit_slice_143989_comb} + 3'h1;
  assign p1_add_144182_comb = {{1{p1_bit_slice_143990_comb[1]}}, p1_bit_slice_143990_comb} + 3'h1;
  assign p1_add_144183_comb = {{1{p1_bit_slice_143991_comb[1]}}, p1_bit_slice_143991_comb} + 3'h1;
  assign p1_add_144184_comb = {{1{p1_bit_slice_143992_comb[1]}}, p1_bit_slice_143992_comb} + 3'h1;
  assign p1_add_144185_comb = {{1{p1_bit_slice_143993_comb[1]}}, p1_bit_slice_143993_comb} + 3'h1;
  assign p1_add_144186_comb = {{1{p1_bit_slice_143994_comb[1]}}, p1_bit_slice_143994_comb} + 3'h1;
  assign p1_clipped__40_comb = p1_add_144123_comb[1] ? 8'hff : {p1_add_144123_comb[0], p1_add_143867_comb[7:1]};
  assign p1_clipped__88_comb = p1_add_144124_comb[1] ? 8'hff : {p1_add_144124_comb[0], p1_add_143868_comb[7:1]};
  assign p1_clipped__41_comb = p1_add_144125_comb[1] ? 8'hff : {p1_add_144125_comb[0], p1_add_143869_comb[7:1]};
  assign p1_clipped__89_comb = p1_add_144126_comb[1] ? 8'hff : {p1_add_144126_comb[0], p1_add_143870_comb[7:1]};
  assign p1_clipped__42_comb = p1_add_144127_comb[1] ? 8'hff : {p1_add_144127_comb[0], p1_add_143871_comb[7:1]};
  assign p1_clipped__90_comb = p1_add_144128_comb[1] ? 8'hff : {p1_add_144128_comb[0], p1_add_143872_comb[7:1]};
  assign p1_clipped__43_comb = p1_add_144129_comb[1] ? 8'hff : {p1_add_144129_comb[0], p1_add_143873_comb[7:1]};
  assign p1_clipped__91_comb = p1_add_144130_comb[1] ? 8'hff : {p1_add_144130_comb[0], p1_add_143874_comb[7:1]};
  assign p1_clipped__44_comb = p1_add_144131_comb[1] ? 8'hff : {p1_add_144131_comb[0], p1_add_143875_comb[7:1]};
  assign p1_clipped__92_comb = p1_add_144132_comb[1] ? 8'hff : {p1_add_144132_comb[0], p1_add_143876_comb[7:1]};
  assign p1_clipped__45_comb = p1_add_144133_comb[1] ? 8'hff : {p1_add_144133_comb[0], p1_add_143877_comb[7:1]};
  assign p1_clipped__93_comb = p1_add_144134_comb[1] ? 8'hff : {p1_add_144134_comb[0], p1_add_143878_comb[7:1]};
  assign p1_clipped__46_comb = p1_add_144135_comb[1] ? 8'hff : {p1_add_144135_comb[0], p1_add_143879_comb[7:1]};
  assign p1_clipped__94_comb = p1_add_144136_comb[1] ? 8'hff : {p1_add_144136_comb[0], p1_add_143880_comb[7:1]};
  assign p1_clipped__47_comb = p1_add_144137_comb[1] ? 8'hff : {p1_add_144137_comb[0], p1_add_143881_comb[7:1]};
  assign p1_clipped__95_comb = p1_add_144138_comb[1] ? 8'hff : {p1_add_144138_comb[0], p1_add_143882_comb[7:1]};
  assign p1_clipped__8_comb = p1_add_144139_comb[1] ? 8'hff : {p1_add_144139_comb[0], p1_add_143883_comb[7:1]};
  assign p1_clipped__24_comb = p1_add_144140_comb[1] ? 8'hff : {p1_add_144140_comb[0], p1_add_143884_comb[7:1]};
  assign p1_clipped__56_comb = p1_add_144141_comb[1] ? 8'hff : {p1_add_144141_comb[0], p1_add_143885_comb[7:1]};
  assign p1_clipped__72_comb = p1_add_144142_comb[1] ? 8'hff : {p1_add_144142_comb[0], p1_add_143886_comb[7:1]};
  assign p1_clipped__104_comb = p1_add_144143_comb[1] ? 8'hff : {p1_add_144143_comb[0], p1_add_143887_comb[7:1]};
  assign p1_clipped__120_comb = p1_add_144144_comb[1] ? 8'hff : {p1_add_144144_comb[0], p1_add_143888_comb[7:1]};
  assign p1_clipped__9_comb = p1_add_144145_comb[1] ? 8'hff : {p1_add_144145_comb[0], p1_add_143889_comb[7:1]};
  assign p1_clipped__25_comb = p1_add_144146_comb[1] ? 8'hff : {p1_add_144146_comb[0], p1_add_143890_comb[7:1]};
  assign p1_clipped__57_comb = p1_add_144147_comb[1] ? 8'hff : {p1_add_144147_comb[0], p1_add_143891_comb[7:1]};
  assign p1_clipped__73_comb = p1_add_144148_comb[1] ? 8'hff : {p1_add_144148_comb[0], p1_add_143892_comb[7:1]};
  assign p1_clipped__105_comb = p1_add_144149_comb[1] ? 8'hff : {p1_add_144149_comb[0], p1_add_143893_comb[7:1]};
  assign p1_clipped__121_comb = p1_add_144150_comb[1] ? 8'hff : {p1_add_144150_comb[0], p1_add_143894_comb[7:1]};
  assign p1_clipped__10_comb = p1_add_144151_comb[1] ? 8'hff : {p1_add_144151_comb[0], p1_add_143895_comb[7:1]};
  assign p1_clipped__26_comb = p1_add_144152_comb[1] ? 8'hff : {p1_add_144152_comb[0], p1_add_143896_comb[7:1]};
  assign p1_clipped__58_comb = p1_add_144153_comb[1] ? 8'hff : {p1_add_144153_comb[0], p1_add_143897_comb[7:1]};
  assign p1_clipped__74_comb = p1_add_144154_comb[1] ? 8'hff : {p1_add_144154_comb[0], p1_add_143898_comb[7:1]};
  assign p1_clipped__106_comb = p1_add_144155_comb[1] ? 8'hff : {p1_add_144155_comb[0], p1_add_143899_comb[7:1]};
  assign p1_clipped__122_comb = p1_add_144156_comb[1] ? 8'hff : {p1_add_144156_comb[0], p1_add_143900_comb[7:1]};
  assign p1_clipped__11_comb = p1_add_144157_comb[1] ? 8'hff : {p1_add_144157_comb[0], p1_add_143901_comb[7:1]};
  assign p1_clipped__27_comb = p1_add_144158_comb[1] ? 8'hff : {p1_add_144158_comb[0], p1_add_143902_comb[7:1]};
  assign p1_clipped__59_comb = p1_add_144159_comb[1] ? 8'hff : {p1_add_144159_comb[0], p1_add_143903_comb[7:1]};
  assign p1_clipped__75_comb = p1_add_144160_comb[1] ? 8'hff : {p1_add_144160_comb[0], p1_add_143904_comb[7:1]};
  assign p1_clipped__107_comb = p1_add_144161_comb[1] ? 8'hff : {p1_add_144161_comb[0], p1_add_143905_comb[7:1]};
  assign p1_clipped__123_comb = p1_add_144162_comb[1] ? 8'hff : {p1_add_144162_comb[0], p1_add_143906_comb[7:1]};
  assign p1_clipped__12_comb = p1_add_144163_comb[1] ? 8'hff : {p1_add_144163_comb[0], p1_add_143907_comb[7:1]};
  assign p1_clipped__28_comb = p1_add_144164_comb[1] ? 8'hff : {p1_add_144164_comb[0], p1_add_143908_comb[7:1]};
  assign p1_clipped__60_comb = p1_add_144165_comb[1] ? 8'hff : {p1_add_144165_comb[0], p1_add_143909_comb[7:1]};
  assign p1_clipped__76_comb = p1_add_144166_comb[1] ? 8'hff : {p1_add_144166_comb[0], p1_add_143910_comb[7:1]};
  assign p1_clipped__108_comb = p1_add_144167_comb[1] ? 8'hff : {p1_add_144167_comb[0], p1_add_143911_comb[7:1]};
  assign p1_clipped__124_comb = p1_add_144168_comb[1] ? 8'hff : {p1_add_144168_comb[0], p1_add_143912_comb[7:1]};
  assign p1_clipped__13_comb = p1_add_144169_comb[1] ? 8'hff : {p1_add_144169_comb[0], p1_add_143913_comb[7:1]};
  assign p1_clipped__29_comb = p1_add_144170_comb[1] ? 8'hff : {p1_add_144170_comb[0], p1_add_143914_comb[7:1]};
  assign p1_clipped__61_comb = p1_add_144171_comb[1] ? 8'hff : {p1_add_144171_comb[0], p1_add_143915_comb[7:1]};
  assign p1_clipped__77_comb = p1_add_144172_comb[1] ? 8'hff : {p1_add_144172_comb[0], p1_add_143916_comb[7:1]};
  assign p1_clipped__109_comb = p1_add_144173_comb[1] ? 8'hff : {p1_add_144173_comb[0], p1_add_143917_comb[7:1]};
  assign p1_clipped__125_comb = p1_add_144174_comb[1] ? 8'hff : {p1_add_144174_comb[0], p1_add_143918_comb[7:1]};
  assign p1_clipped__14_comb = p1_add_144175_comb[1] ? 8'hff : {p1_add_144175_comb[0], p1_add_143919_comb[7:1]};
  assign p1_clipped__30_comb = p1_add_144176_comb[1] ? 8'hff : {p1_add_144176_comb[0], p1_add_143920_comb[7:1]};
  assign p1_clipped__62_comb = p1_add_144177_comb[1] ? 8'hff : {p1_add_144177_comb[0], p1_add_143921_comb[7:1]};
  assign p1_clipped__78_comb = p1_add_144178_comb[1] ? 8'hff : {p1_add_144178_comb[0], p1_add_143922_comb[7:1]};
  assign p1_clipped__110_comb = p1_add_144179_comb[1] ? 8'hff : {p1_add_144179_comb[0], p1_add_143923_comb[7:1]};
  assign p1_clipped__126_comb = p1_add_144180_comb[1] ? 8'hff : {p1_add_144180_comb[0], p1_add_143924_comb[7:1]};
  assign p1_clipped__15_comb = p1_add_144181_comb[1] ? 8'hff : {p1_add_144181_comb[0], p1_add_143925_comb[7:1]};
  assign p1_clipped__31_comb = p1_add_144182_comb[1] ? 8'hff : {p1_add_144182_comb[0], p1_add_143926_comb[7:1]};
  assign p1_clipped__63_comb = p1_add_144183_comb[1] ? 8'hff : {p1_add_144183_comb[0], p1_add_143927_comb[7:1]};
  assign p1_clipped__79_comb = p1_add_144184_comb[1] ? 8'hff : {p1_add_144184_comb[0], p1_add_143928_comb[7:1]};
  assign p1_clipped__111_comb = p1_add_144185_comb[1] ? 8'hff : {p1_add_144185_comb[0], p1_add_143929_comb[7:1]};
  assign p1_clipped__127_comb = p1_add_144186_comb[1] ? 8'hff : {p1_add_144186_comb[0], p1_add_143930_comb[7:1]};
  assign p1_shifted__66_squeezed_comb = {~p1_clipped__40_comb[7], p1_clipped__40_comb[6:0]};
  assign p1_shifted__69_squeezed_comb = {~p1_clipped__88_comb[7], p1_clipped__88_comb[6:0]};
  assign p1_shifted__74_squeezed_comb = {~p1_clipped__41_comb[7], p1_clipped__41_comb[6:0]};
  assign p1_shifted__77_squeezed_comb = {~p1_clipped__89_comb[7], p1_clipped__89_comb[6:0]};
  assign p1_shifted__82_squeezed_comb = {~p1_clipped__42_comb[7], p1_clipped__42_comb[6:0]};
  assign p1_shifted__85_squeezed_comb = {~p1_clipped__90_comb[7], p1_clipped__90_comb[6:0]};
  assign p1_shifted__90_squeezed_comb = {~p1_clipped__43_comb[7], p1_clipped__43_comb[6:0]};
  assign p1_shifted__93_squeezed_comb = {~p1_clipped__91_comb[7], p1_clipped__91_comb[6:0]};
  assign p1_shifted__98_squeezed_comb = {~p1_clipped__44_comb[7], p1_clipped__44_comb[6:0]};
  assign p1_shifted__101_squeezed_comb = {~p1_clipped__92_comb[7], p1_clipped__92_comb[6:0]};
  assign p1_shifted__106_squeezed_comb = {~p1_clipped__45_comb[7], p1_clipped__45_comb[6:0]};
  assign p1_shifted__109_squeezed_comb = {~p1_clipped__93_comb[7], p1_clipped__93_comb[6:0]};
  assign p1_shifted__114_squeezed_comb = {~p1_clipped__46_comb[7], p1_clipped__46_comb[6:0]};
  assign p1_shifted__117_squeezed_comb = {~p1_clipped__94_comb[7], p1_clipped__94_comb[6:0]};
  assign p1_shifted__122_squeezed_comb = {~p1_clipped__47_comb[7], p1_clipped__47_comb[6:0]};
  assign p1_shifted__125_squeezed_comb = {~p1_clipped__95_comb[7], p1_clipped__95_comb[6:0]};
  assign p1_shifted__64_squeezed_comb = {~p1_clipped__8_comb[7], p1_clipped__8_comb[6:0]};
  assign p1_shifted__65_squeezed_comb = {~p1_clipped__24_comb[7], p1_clipped__24_comb[6:0]};
  assign p1_shifted__67_squeezed_comb = {~p1_clipped__56_comb[7], p1_clipped__56_comb[6:0]};
  assign p1_shifted__68_squeezed_comb = {~p1_clipped__72_comb[7], p1_clipped__72_comb[6:0]};
  assign p1_shifted__70_squeezed_comb = {~p1_clipped__104_comb[7], p1_clipped__104_comb[6:0]};
  assign p1_shifted__71_squeezed_comb = {~p1_clipped__120_comb[7], p1_clipped__120_comb[6:0]};
  assign p1_shifted__72_squeezed_comb = {~p1_clipped__9_comb[7], p1_clipped__9_comb[6:0]};
  assign p1_shifted__73_squeezed_comb = {~p1_clipped__25_comb[7], p1_clipped__25_comb[6:0]};
  assign p1_shifted__75_squeezed_comb = {~p1_clipped__57_comb[7], p1_clipped__57_comb[6:0]};
  assign p1_shifted__76_squeezed_comb = {~p1_clipped__73_comb[7], p1_clipped__73_comb[6:0]};
  assign p1_shifted__78_squeezed_comb = {~p1_clipped__105_comb[7], p1_clipped__105_comb[6:0]};
  assign p1_shifted__79_squeezed_comb = {~p1_clipped__121_comb[7], p1_clipped__121_comb[6:0]};
  assign p1_shifted__80_squeezed_comb = {~p1_clipped__10_comb[7], p1_clipped__10_comb[6:0]};
  assign p1_shifted__81_squeezed_comb = {~p1_clipped__26_comb[7], p1_clipped__26_comb[6:0]};
  assign p1_shifted__83_squeezed_comb = {~p1_clipped__58_comb[7], p1_clipped__58_comb[6:0]};
  assign p1_shifted__84_squeezed_comb = {~p1_clipped__74_comb[7], p1_clipped__74_comb[6:0]};
  assign p1_shifted__86_squeezed_comb = {~p1_clipped__106_comb[7], p1_clipped__106_comb[6:0]};
  assign p1_shifted__87_squeezed_comb = {~p1_clipped__122_comb[7], p1_clipped__122_comb[6:0]};
  assign p1_shifted__88_squeezed_comb = {~p1_clipped__11_comb[7], p1_clipped__11_comb[6:0]};
  assign p1_shifted__89_squeezed_comb = {~p1_clipped__27_comb[7], p1_clipped__27_comb[6:0]};
  assign p1_shifted__91_squeezed_comb = {~p1_clipped__59_comb[7], p1_clipped__59_comb[6:0]};
  assign p1_shifted__92_squeezed_comb = {~p1_clipped__75_comb[7], p1_clipped__75_comb[6:0]};
  assign p1_shifted__94_squeezed_comb = {~p1_clipped__107_comb[7], p1_clipped__107_comb[6:0]};
  assign p1_shifted__95_squeezed_comb = {~p1_clipped__123_comb[7], p1_clipped__123_comb[6:0]};
  assign p1_shifted__96_squeezed_comb = {~p1_clipped__12_comb[7], p1_clipped__12_comb[6:0]};
  assign p1_shifted__97_squeezed_comb = {~p1_clipped__28_comb[7], p1_clipped__28_comb[6:0]};
  assign p1_shifted__99_squeezed_comb = {~p1_clipped__60_comb[7], p1_clipped__60_comb[6:0]};
  assign p1_shifted__100_squeezed_comb = {~p1_clipped__76_comb[7], p1_clipped__76_comb[6:0]};
  assign p1_shifted__102_squeezed_comb = {~p1_clipped__108_comb[7], p1_clipped__108_comb[6:0]};
  assign p1_shifted__103_squeezed_comb = {~p1_clipped__124_comb[7], p1_clipped__124_comb[6:0]};
  assign p1_shifted__104_squeezed_comb = {~p1_clipped__13_comb[7], p1_clipped__13_comb[6:0]};
  assign p1_shifted__105_squeezed_comb = {~p1_clipped__29_comb[7], p1_clipped__29_comb[6:0]};
  assign p1_shifted__107_squeezed_comb = {~p1_clipped__61_comb[7], p1_clipped__61_comb[6:0]};
  assign p1_shifted__108_squeezed_comb = {~p1_clipped__77_comb[7], p1_clipped__77_comb[6:0]};
  assign p1_shifted__110_squeezed_comb = {~p1_clipped__109_comb[7], p1_clipped__109_comb[6:0]};
  assign p1_shifted__111_squeezed_comb = {~p1_clipped__125_comb[7], p1_clipped__125_comb[6:0]};
  assign p1_shifted__112_squeezed_comb = {~p1_clipped__14_comb[7], p1_clipped__14_comb[6:0]};
  assign p1_shifted__113_squeezed_comb = {~p1_clipped__30_comb[7], p1_clipped__30_comb[6:0]};
  assign p1_shifted__115_squeezed_comb = {~p1_clipped__62_comb[7], p1_clipped__62_comb[6:0]};
  assign p1_shifted__116_squeezed_comb = {~p1_clipped__78_comb[7], p1_clipped__78_comb[6:0]};
  assign p1_shifted__118_squeezed_comb = {~p1_clipped__110_comb[7], p1_clipped__110_comb[6:0]};
  assign p1_shifted__119_squeezed_comb = {~p1_clipped__126_comb[7], p1_clipped__126_comb[6:0]};
  assign p1_shifted__120_squeezed_comb = {~p1_clipped__15_comb[7], p1_clipped__15_comb[6:0]};
  assign p1_shifted__121_squeezed_comb = {~p1_clipped__31_comb[7], p1_clipped__31_comb[6:0]};
  assign p1_shifted__123_squeezed_comb = {~p1_clipped__63_comb[7], p1_clipped__63_comb[6:0]};
  assign p1_shifted__124_squeezed_comb = {~p1_clipped__79_comb[7], p1_clipped__79_comb[6:0]};
  assign p1_shifted__126_squeezed_comb = {~p1_clipped__111_comb[7], p1_clipped__111_comb[6:0]};
  assign p1_shifted__127_squeezed_comb = {~p1_clipped__127_comb[7], p1_clipped__127_comb[6:0]};
  assign p1_smul_58226_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__66_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___192_comb = 9'h000;
  assign p1_smul_58232_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__69_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___195_comb = 9'h000;
  assign p1_smul_58242_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__74_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___196_comb = 9'h000;
  assign p1_smul_58248_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__77_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___199_comb = 9'h000;
  assign p1_smul_58258_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__82_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___200_comb = 9'h000;
  assign p1_smul_58264_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__85_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___203_comb = 9'h000;
  assign p1_smul_58274_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__90_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___204_comb = 9'h000;
  assign p1_smul_58280_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__93_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___207_comb = 9'h000;
  assign p1_smul_58290_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__98_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___208_comb = 9'h000;
  assign p1_smul_58296_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__101_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___211_comb = 9'h000;
  assign p1_smul_58306_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__106_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___212_comb = 9'h000;
  assign p1_smul_58312_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__109_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___215_comb = 9'h000;
  assign p1_smul_58322_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__114_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___216_comb = 9'h000;
  assign p1_smul_58328_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__117_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___219_comb = 9'h000;
  assign p1_smul_58338_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__122_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___220_comb = 9'h000;
  assign p1_smul_58344_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__125_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___223_comb = 9'h000;
  assign p1_smul_58350_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__64_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___64_comb = 10'h000;
  assign p1_smul_58352_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__65_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___224_comb = 9'h000;
  assign p1_smul_58354_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__66_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___225_comb = 9'h000;
  assign p1_smul_58356_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__67_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___65_comb = 10'h000;
  assign p1_smul_58358_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__68_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___66_comb = 10'h000;
  assign p1_smul_58360_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__69_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___226_comb = 9'h000;
  assign p1_smul_58362_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__70_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___227_comb = 9'h000;
  assign p1_smul_58364_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__71_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___67_comb = 10'h000;
  assign p1_smul_58366_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__72_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___68_comb = 10'h000;
  assign p1_smul_58368_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__73_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___228_comb = 9'h000;
  assign p1_smul_58370_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__74_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___229_comb = 9'h000;
  assign p1_smul_58372_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__75_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___69_comb = 10'h000;
  assign p1_smul_58374_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__76_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___70_comb = 10'h000;
  assign p1_smul_58376_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__77_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___230_comb = 9'h000;
  assign p1_smul_58378_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__78_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___231_comb = 9'h000;
  assign p1_smul_58380_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__79_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___71_comb = 10'h000;
  assign p1_smul_58382_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__80_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___72_comb = 10'h000;
  assign p1_smul_58384_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__81_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___232_comb = 9'h000;
  assign p1_smul_58386_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__82_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___233_comb = 9'h000;
  assign p1_smul_58388_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__83_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___73_comb = 10'h000;
  assign p1_smul_58390_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__84_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___74_comb = 10'h000;
  assign p1_smul_58392_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__85_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___234_comb = 9'h000;
  assign p1_smul_58394_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__86_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___235_comb = 9'h000;
  assign p1_smul_58396_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__87_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___75_comb = 10'h000;
  assign p1_smul_58398_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__88_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___76_comb = 10'h000;
  assign p1_smul_58400_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__89_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___236_comb = 9'h000;
  assign p1_smul_58402_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__90_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___237_comb = 9'h000;
  assign p1_smul_58404_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__91_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___77_comb = 10'h000;
  assign p1_smul_58406_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__92_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___78_comb = 10'h000;
  assign p1_smul_58408_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__93_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___238_comb = 9'h000;
  assign p1_smul_58410_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__94_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___239_comb = 9'h000;
  assign p1_smul_58412_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__95_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___79_comb = 10'h000;
  assign p1_smul_58414_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__96_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___80_comb = 10'h000;
  assign p1_smul_58416_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__97_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___240_comb = 9'h000;
  assign p1_smul_58418_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__98_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___241_comb = 9'h000;
  assign p1_smul_58420_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__99_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___81_comb = 10'h000;
  assign p1_smul_58422_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__100_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___82_comb = 10'h000;
  assign p1_smul_58424_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__101_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___242_comb = 9'h000;
  assign p1_smul_58426_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__102_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___243_comb = 9'h000;
  assign p1_smul_58428_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__103_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___83_comb = 10'h000;
  assign p1_smul_58430_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__104_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___84_comb = 10'h000;
  assign p1_smul_58432_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__105_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___244_comb = 9'h000;
  assign p1_smul_58434_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__106_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___245_comb = 9'h000;
  assign p1_smul_58436_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__107_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___85_comb = 10'h000;
  assign p1_smul_58438_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__108_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___86_comb = 10'h000;
  assign p1_smul_58440_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__109_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___246_comb = 9'h000;
  assign p1_smul_58442_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__110_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___247_comb = 9'h000;
  assign p1_smul_58444_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__111_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___87_comb = 10'h000;
  assign p1_smul_58446_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__112_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___88_comb = 10'h000;
  assign p1_smul_58448_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__113_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___248_comb = 9'h000;
  assign p1_smul_58450_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__114_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___249_comb = 9'h000;
  assign p1_smul_58452_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__115_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___89_comb = 10'h000;
  assign p1_smul_58454_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__116_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___90_comb = 10'h000;
  assign p1_smul_58456_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__117_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___250_comb = 9'h000;
  assign p1_smul_58458_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__118_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___251_comb = 9'h000;
  assign p1_smul_58460_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__119_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___91_comb = 10'h000;
  assign p1_smul_58462_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__120_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___92_comb = 10'h000;
  assign p1_smul_58464_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__121_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___252_comb = 9'h000;
  assign p1_smul_58466_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__122_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___253_comb = 9'h000;
  assign p1_smul_58468_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__123_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___93_comb = 10'h000;
  assign p1_smul_58470_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__124_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___94_comb = 10'h000;
  assign p1_smul_58472_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__125_squeezed_comb, 7'h4f);
  assign p1_smul_57330_TrailingBits___254_comb = 9'h000;
  assign p1_smul_58474_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__126_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___255_comb = 9'h000;
  assign p1_smul_58476_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__127_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___95_comb = 10'h000;
  assign p1_smul_58484_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__67_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___257_comb = 9'h000;
  assign p1_smul_58486_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__68_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___258_comb = 9'h000;
  assign p1_smul_58500_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__75_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___261_comb = 9'h000;
  assign p1_smul_58502_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__76_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___262_comb = 9'h000;
  assign p1_smul_58516_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__83_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___265_comb = 9'h000;
  assign p1_smul_58518_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__84_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___266_comb = 9'h000;
  assign p1_smul_58532_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__91_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___269_comb = 9'h000;
  assign p1_smul_58534_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__92_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___270_comb = 9'h000;
  assign p1_smul_58548_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__99_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___273_comb = 9'h000;
  assign p1_smul_58550_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__100_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___274_comb = 9'h000;
  assign p1_smul_58564_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__107_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___277_comb = 9'h000;
  assign p1_smul_58566_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__108_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___278_comb = 9'h000;
  assign p1_smul_58580_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__115_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___281_comb = 9'h000;
  assign p1_smul_58582_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__116_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___282_comb = 9'h000;
  assign p1_smul_58596_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__123_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___285_comb = 9'h000;
  assign p1_smul_58598_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__124_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___286_comb = 9'h000;
  assign p1_smul_58734_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__64_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___288_comb = 9'h000;
  assign p1_smul_58748_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__71_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___291_comb = 9'h000;
  assign p1_smul_58750_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__72_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___292_comb = 9'h000;
  assign p1_smul_58764_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__79_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___295_comb = 9'h000;
  assign p1_smul_58766_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__80_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___296_comb = 9'h000;
  assign p1_smul_58780_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__87_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___299_comb = 9'h000;
  assign p1_smul_58782_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__88_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___300_comb = 9'h000;
  assign p1_smul_58796_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__95_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___303_comb = 9'h000;
  assign p1_smul_58798_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__96_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___304_comb = 9'h000;
  assign p1_smul_58812_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__103_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___307_comb = 9'h000;
  assign p1_smul_58814_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__104_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___308_comb = 9'h000;
  assign p1_smul_58828_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__111_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___311_comb = 9'h000;
  assign p1_smul_58830_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__112_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___312_comb = 9'h000;
  assign p1_smul_58844_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__119_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___315_comb = 9'h000;
  assign p1_smul_58846_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__120_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___316_comb = 9'h000;
  assign p1_smul_58860_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__127_squeezed_comb, 8'h47);
  assign p1_smul_57330_TrailingBits___319_comb = 9'h000;
  assign p1_smul_58862_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__64_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___320_comb = 9'h000;
  assign p1_smul_58864_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__65_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___96_comb = 10'h000;
  assign p1_smul_58866_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__66_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___321_comb = 9'h000;
  assign p1_smul_58868_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__67_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___97_comb = 10'h000;
  assign p1_smul_58870_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__68_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___98_comb = 10'h000;
  assign p1_smul_58872_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__69_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___322_comb = 9'h000;
  assign p1_smul_58874_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__70_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___99_comb = 10'h000;
  assign p1_smul_58876_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__71_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___323_comb = 9'h000;
  assign p1_smul_58878_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__72_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___324_comb = 9'h000;
  assign p1_smul_58880_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__73_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___100_comb = 10'h000;
  assign p1_smul_58882_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__74_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___325_comb = 9'h000;
  assign p1_smul_58884_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__75_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___101_comb = 10'h000;
  assign p1_smul_58886_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__76_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___102_comb = 10'h000;
  assign p1_smul_58888_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__77_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___326_comb = 9'h000;
  assign p1_smul_58890_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__78_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___103_comb = 10'h000;
  assign p1_smul_58892_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__79_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___327_comb = 9'h000;
  assign p1_smul_58894_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__80_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___328_comb = 9'h000;
  assign p1_smul_58896_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__81_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___104_comb = 10'h000;
  assign p1_smul_58898_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__82_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___329_comb = 9'h000;
  assign p1_smul_58900_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__83_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___105_comb = 10'h000;
  assign p1_smul_58902_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__84_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___106_comb = 10'h000;
  assign p1_smul_58904_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__85_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___330_comb = 9'h000;
  assign p1_smul_58906_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__86_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___107_comb = 10'h000;
  assign p1_smul_58908_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__87_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___331_comb = 9'h000;
  assign p1_smul_58910_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__88_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___332_comb = 9'h000;
  assign p1_smul_58912_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__89_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___108_comb = 10'h000;
  assign p1_smul_58914_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__90_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___333_comb = 9'h000;
  assign p1_smul_58916_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__91_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___109_comb = 10'h000;
  assign p1_smul_58918_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__92_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___110_comb = 10'h000;
  assign p1_smul_58920_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__93_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___334_comb = 9'h000;
  assign p1_smul_58922_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__94_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___111_comb = 10'h000;
  assign p1_smul_58924_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__95_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___335_comb = 9'h000;
  assign p1_smul_58926_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__96_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___336_comb = 9'h000;
  assign p1_smul_58928_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__97_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___112_comb = 10'h000;
  assign p1_smul_58930_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__98_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___337_comb = 9'h000;
  assign p1_smul_58932_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__99_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___113_comb = 10'h000;
  assign p1_smul_58934_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__100_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___114_comb = 10'h000;
  assign p1_smul_58936_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__101_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___338_comb = 9'h000;
  assign p1_smul_58938_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__102_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___115_comb = 10'h000;
  assign p1_smul_58940_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__103_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___339_comb = 9'h000;
  assign p1_smul_58942_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__104_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___340_comb = 9'h000;
  assign p1_smul_58944_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__105_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___116_comb = 10'h000;
  assign p1_smul_58946_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__106_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___341_comb = 9'h000;
  assign p1_smul_58948_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__107_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___117_comb = 10'h000;
  assign p1_smul_58950_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__108_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___118_comb = 10'h000;
  assign p1_smul_58952_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__109_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___342_comb = 9'h000;
  assign p1_smul_58954_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__110_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___119_comb = 10'h000;
  assign p1_smul_58956_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__111_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___343_comb = 9'h000;
  assign p1_smul_58958_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__112_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___344_comb = 9'h000;
  assign p1_smul_58960_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__113_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___120_comb = 10'h000;
  assign p1_smul_58962_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__114_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___345_comb = 9'h000;
  assign p1_smul_58964_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__115_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___121_comb = 10'h000;
  assign p1_smul_58966_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__116_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___122_comb = 10'h000;
  assign p1_smul_58968_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__117_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___346_comb = 9'h000;
  assign p1_smul_58970_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__118_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___123_comb = 10'h000;
  assign p1_smul_58972_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__119_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___347_comb = 9'h000;
  assign p1_smul_58974_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__120_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___348_comb = 9'h000;
  assign p1_smul_58976_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__121_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___124_comb = 10'h000;
  assign p1_smul_58978_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__122_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___349_comb = 9'h000;
  assign p1_smul_58980_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__123_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___125_comb = 10'h000;
  assign p1_smul_58982_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__124_squeezed_comb, 7'h3b);
  assign p1_smul_57454_TrailingBits___126_comb = 10'h000;
  assign p1_smul_58984_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__125_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___350_comb = 9'h000;
  assign p1_smul_58986_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__126_squeezed_comb, 7'h45);
  assign p1_smul_57454_TrailingBits___127_comb = 10'h000;
  assign p1_smul_58988_NarrowedMult__comb = smul15b_8b_x_7b(p1_shifted__127_squeezed_comb, 7'h31);
  assign p1_smul_57330_TrailingBits___351_comb = 9'h000;
  assign p1_smul_58992_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__65_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___353_comb = 9'h000;
  assign p1_smul_59002_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__70_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___354_comb = 9'h000;
  assign p1_smul_59008_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__73_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___357_comb = 9'h000;
  assign p1_smul_59018_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__78_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___358_comb = 9'h000;
  assign p1_smul_59024_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__81_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___361_comb = 9'h000;
  assign p1_smul_59034_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__86_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___362_comb = 9'h000;
  assign p1_smul_59040_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__89_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___365_comb = 9'h000;
  assign p1_smul_59050_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__94_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___366_comb = 9'h000;
  assign p1_smul_59056_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__97_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___369_comb = 9'h000;
  assign p1_smul_59066_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__102_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___370_comb = 9'h000;
  assign p1_smul_59072_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__105_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___373_comb = 9'h000;
  assign p1_smul_59082_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__110_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___374_comb = 9'h000;
  assign p1_smul_59088_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__113_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___377_comb = 9'h000;
  assign p1_smul_59098_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__118_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___378_comb = 9'h000;
  assign p1_smul_59104_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__121_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___381_comb = 9'h000;
  assign p1_smul_59114_NarrowedMult__comb = smul16b_8b_x_8b(p1_shifted__126_squeezed_comb, 8'hb9);
  assign p1_smul_57330_TrailingBits___382_comb = 9'h000;
  assign p1_concat_145531_comb = {p1_smul_58226_NarrowedMult__comb, p1_smul_57330_TrailingBits___192_comb};
  assign p1_smul_58228_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__67_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___193_comb = 9'h000;
  assign p1_smul_58230_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__68_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___194_comb = 9'h000;
  assign p1_concat_145536_comb = {p1_smul_58232_NarrowedMult__comb, p1_smul_57330_TrailingBits___195_comb};
  assign p1_concat_145537_comb = {p1_smul_58242_NarrowedMult__comb, p1_smul_57330_TrailingBits___196_comb};
  assign p1_smul_58244_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__75_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___197_comb = 9'h000;
  assign p1_smul_58246_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__76_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___198_comb = 9'h000;
  assign p1_concat_145542_comb = {p1_smul_58248_NarrowedMult__comb, p1_smul_57330_TrailingBits___199_comb};
  assign p1_concat_145543_comb = {p1_smul_58258_NarrowedMult__comb, p1_smul_57330_TrailingBits___200_comb};
  assign p1_smul_58260_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__83_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___201_comb = 9'h000;
  assign p1_smul_58262_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__84_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___202_comb = 9'h000;
  assign p1_concat_145548_comb = {p1_smul_58264_NarrowedMult__comb, p1_smul_57330_TrailingBits___203_comb};
  assign p1_concat_145549_comb = {p1_smul_58274_NarrowedMult__comb, p1_smul_57330_TrailingBits___204_comb};
  assign p1_smul_58276_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__91_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___205_comb = 9'h000;
  assign p1_smul_58278_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__92_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___206_comb = 9'h000;
  assign p1_concat_145554_comb = {p1_smul_58280_NarrowedMult__comb, p1_smul_57330_TrailingBits___207_comb};
  assign p1_concat_145555_comb = {p1_smul_58290_NarrowedMult__comb, p1_smul_57330_TrailingBits___208_comb};
  assign p1_smul_58292_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__99_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___209_comb = 9'h000;
  assign p1_smul_58294_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__100_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___210_comb = 9'h000;
  assign p1_concat_145560_comb = {p1_smul_58296_NarrowedMult__comb, p1_smul_57330_TrailingBits___211_comb};
  assign p1_concat_145561_comb = {p1_smul_58306_NarrowedMult__comb, p1_smul_57330_TrailingBits___212_comb};
  assign p1_smul_58308_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__107_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___213_comb = 9'h000;
  assign p1_smul_58310_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__108_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___214_comb = 9'h000;
  assign p1_concat_145566_comb = {p1_smul_58312_NarrowedMult__comb, p1_smul_57330_TrailingBits___215_comb};
  assign p1_concat_145567_comb = {p1_smul_58322_NarrowedMult__comb, p1_smul_57330_TrailingBits___216_comb};
  assign p1_smul_58324_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__115_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___217_comb = 9'h000;
  assign p1_smul_58326_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__116_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___218_comb = 9'h000;
  assign p1_concat_145572_comb = {p1_smul_58328_NarrowedMult__comb, p1_smul_57330_TrailingBits___219_comb};
  assign p1_concat_145573_comb = {p1_smul_58338_NarrowedMult__comb, p1_smul_57330_TrailingBits___220_comb};
  assign p1_smul_58340_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__123_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___221_comb = 9'h000;
  assign p1_smul_58342_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__124_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___222_comb = 9'h000;
  assign p1_concat_145578_comb = {p1_smul_58344_NarrowedMult__comb, p1_smul_57330_TrailingBits___223_comb};
  assign p1_concat_145579_comb = {p1_smul_58350_NarrowedMult__comb, p1_smul_57454_TrailingBits___64_comb};
  assign p1_concat_145580_comb = {p1_smul_58352_NarrowedMult__comb, p1_smul_57330_TrailingBits___224_comb};
  assign p1_concat_145581_comb = {p1_smul_58354_NarrowedMult__comb, p1_smul_57330_TrailingBits___225_comb};
  assign p1_concat_145582_comb = {p1_smul_58356_NarrowedMult__comb, p1_smul_57454_TrailingBits___65_comb};
  assign p1_concat_145583_comb = {p1_smul_58358_NarrowedMult__comb, p1_smul_57454_TrailingBits___66_comb};
  assign p1_concat_145584_comb = {p1_smul_58360_NarrowedMult__comb, p1_smul_57330_TrailingBits___226_comb};
  assign p1_concat_145585_comb = {p1_smul_58362_NarrowedMult__comb, p1_smul_57330_TrailingBits___227_comb};
  assign p1_concat_145586_comb = {p1_smul_58364_NarrowedMult__comb, p1_smul_57454_TrailingBits___67_comb};
  assign p1_concat_145587_comb = {p1_smul_58366_NarrowedMult__comb, p1_smul_57454_TrailingBits___68_comb};
  assign p1_concat_145588_comb = {p1_smul_58368_NarrowedMult__comb, p1_smul_57330_TrailingBits___228_comb};
  assign p1_concat_145589_comb = {p1_smul_58370_NarrowedMult__comb, p1_smul_57330_TrailingBits___229_comb};
  assign p1_concat_145590_comb = {p1_smul_58372_NarrowedMult__comb, p1_smul_57454_TrailingBits___69_comb};
  assign p1_concat_145591_comb = {p1_smul_58374_NarrowedMult__comb, p1_smul_57454_TrailingBits___70_comb};
  assign p1_concat_145592_comb = {p1_smul_58376_NarrowedMult__comb, p1_smul_57330_TrailingBits___230_comb};
  assign p1_concat_145593_comb = {p1_smul_58378_NarrowedMult__comb, p1_smul_57330_TrailingBits___231_comb};
  assign p1_concat_145594_comb = {p1_smul_58380_NarrowedMult__comb, p1_smul_57454_TrailingBits___71_comb};
  assign p1_concat_145595_comb = {p1_smul_58382_NarrowedMult__comb, p1_smul_57454_TrailingBits___72_comb};
  assign p1_concat_145596_comb = {p1_smul_58384_NarrowedMult__comb, p1_smul_57330_TrailingBits___232_comb};
  assign p1_concat_145597_comb = {p1_smul_58386_NarrowedMult__comb, p1_smul_57330_TrailingBits___233_comb};
  assign p1_concat_145598_comb = {p1_smul_58388_NarrowedMult__comb, p1_smul_57454_TrailingBits___73_comb};
  assign p1_concat_145599_comb = {p1_smul_58390_NarrowedMult__comb, p1_smul_57454_TrailingBits___74_comb};
  assign p1_concat_145600_comb = {p1_smul_58392_NarrowedMult__comb, p1_smul_57330_TrailingBits___234_comb};
  assign p1_concat_145601_comb = {p1_smul_58394_NarrowedMult__comb, p1_smul_57330_TrailingBits___235_comb};
  assign p1_concat_145602_comb = {p1_smul_58396_NarrowedMult__comb, p1_smul_57454_TrailingBits___75_comb};
  assign p1_concat_145603_comb = {p1_smul_58398_NarrowedMult__comb, p1_smul_57454_TrailingBits___76_comb};
  assign p1_concat_145604_comb = {p1_smul_58400_NarrowedMult__comb, p1_smul_57330_TrailingBits___236_comb};
  assign p1_concat_145605_comb = {p1_smul_58402_NarrowedMult__comb, p1_smul_57330_TrailingBits___237_comb};
  assign p1_concat_145606_comb = {p1_smul_58404_NarrowedMult__comb, p1_smul_57454_TrailingBits___77_comb};
  assign p1_concat_145607_comb = {p1_smul_58406_NarrowedMult__comb, p1_smul_57454_TrailingBits___78_comb};
  assign p1_concat_145608_comb = {p1_smul_58408_NarrowedMult__comb, p1_smul_57330_TrailingBits___238_comb};
  assign p1_concat_145609_comb = {p1_smul_58410_NarrowedMult__comb, p1_smul_57330_TrailingBits___239_comb};
  assign p1_concat_145610_comb = {p1_smul_58412_NarrowedMult__comb, p1_smul_57454_TrailingBits___79_comb};
  assign p1_concat_145611_comb = {p1_smul_58414_NarrowedMult__comb, p1_smul_57454_TrailingBits___80_comb};
  assign p1_concat_145612_comb = {p1_smul_58416_NarrowedMult__comb, p1_smul_57330_TrailingBits___240_comb};
  assign p1_concat_145613_comb = {p1_smul_58418_NarrowedMult__comb, p1_smul_57330_TrailingBits___241_comb};
  assign p1_concat_145614_comb = {p1_smul_58420_NarrowedMult__comb, p1_smul_57454_TrailingBits___81_comb};
  assign p1_concat_145615_comb = {p1_smul_58422_NarrowedMult__comb, p1_smul_57454_TrailingBits___82_comb};
  assign p1_concat_145616_comb = {p1_smul_58424_NarrowedMult__comb, p1_smul_57330_TrailingBits___242_comb};
  assign p1_concat_145617_comb = {p1_smul_58426_NarrowedMult__comb, p1_smul_57330_TrailingBits___243_comb};
  assign p1_concat_145618_comb = {p1_smul_58428_NarrowedMult__comb, p1_smul_57454_TrailingBits___83_comb};
  assign p1_concat_145619_comb = {p1_smul_58430_NarrowedMult__comb, p1_smul_57454_TrailingBits___84_comb};
  assign p1_concat_145620_comb = {p1_smul_58432_NarrowedMult__comb, p1_smul_57330_TrailingBits___244_comb};
  assign p1_concat_145621_comb = {p1_smul_58434_NarrowedMult__comb, p1_smul_57330_TrailingBits___245_comb};
  assign p1_concat_145622_comb = {p1_smul_58436_NarrowedMult__comb, p1_smul_57454_TrailingBits___85_comb};
  assign p1_concat_145623_comb = {p1_smul_58438_NarrowedMult__comb, p1_smul_57454_TrailingBits___86_comb};
  assign p1_concat_145624_comb = {p1_smul_58440_NarrowedMult__comb, p1_smul_57330_TrailingBits___246_comb};
  assign p1_concat_145625_comb = {p1_smul_58442_NarrowedMult__comb, p1_smul_57330_TrailingBits___247_comb};
  assign p1_concat_145626_comb = {p1_smul_58444_NarrowedMult__comb, p1_smul_57454_TrailingBits___87_comb};
  assign p1_concat_145627_comb = {p1_smul_58446_NarrowedMult__comb, p1_smul_57454_TrailingBits___88_comb};
  assign p1_concat_145628_comb = {p1_smul_58448_NarrowedMult__comb, p1_smul_57330_TrailingBits___248_comb};
  assign p1_concat_145629_comb = {p1_smul_58450_NarrowedMult__comb, p1_smul_57330_TrailingBits___249_comb};
  assign p1_concat_145630_comb = {p1_smul_58452_NarrowedMult__comb, p1_smul_57454_TrailingBits___89_comb};
  assign p1_concat_145631_comb = {p1_smul_58454_NarrowedMult__comb, p1_smul_57454_TrailingBits___90_comb};
  assign p1_concat_145632_comb = {p1_smul_58456_NarrowedMult__comb, p1_smul_57330_TrailingBits___250_comb};
  assign p1_concat_145633_comb = {p1_smul_58458_NarrowedMult__comb, p1_smul_57330_TrailingBits___251_comb};
  assign p1_concat_145634_comb = {p1_smul_58460_NarrowedMult__comb, p1_smul_57454_TrailingBits___91_comb};
  assign p1_concat_145635_comb = {p1_smul_58462_NarrowedMult__comb, p1_smul_57454_TrailingBits___92_comb};
  assign p1_concat_145636_comb = {p1_smul_58464_NarrowedMult__comb, p1_smul_57330_TrailingBits___252_comb};
  assign p1_concat_145637_comb = {p1_smul_58466_NarrowedMult__comb, p1_smul_57330_TrailingBits___253_comb};
  assign p1_concat_145638_comb = {p1_smul_58468_NarrowedMult__comb, p1_smul_57454_TrailingBits___93_comb};
  assign p1_concat_145639_comb = {p1_smul_58470_NarrowedMult__comb, p1_smul_57454_TrailingBits___94_comb};
  assign p1_concat_145640_comb = {p1_smul_58472_NarrowedMult__comb, p1_smul_57330_TrailingBits___254_comb};
  assign p1_concat_145641_comb = {p1_smul_58474_NarrowedMult__comb, p1_smul_57330_TrailingBits___255_comb};
  assign p1_concat_145642_comb = {p1_smul_58476_NarrowedMult__comb, p1_smul_57454_TrailingBits___95_comb};
  assign p1_smul_58480_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__65_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___256_comb = 9'h000;
  assign p1_concat_145645_comb = {p1_smul_58484_NarrowedMult__comb, p1_smul_57330_TrailingBits___257_comb};
  assign p1_concat_145646_comb = {p1_smul_58486_NarrowedMult__comb, p1_smul_57330_TrailingBits___258_comb};
  assign p1_smul_58490_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__70_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___259_comb = 9'h000;
  assign p1_smul_58496_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__73_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___260_comb = 9'h000;
  assign p1_concat_145651_comb = {p1_smul_58500_NarrowedMult__comb, p1_smul_57330_TrailingBits___261_comb};
  assign p1_concat_145652_comb = {p1_smul_58502_NarrowedMult__comb, p1_smul_57330_TrailingBits___262_comb};
  assign p1_smul_58506_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__78_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___263_comb = 9'h000;
  assign p1_smul_58512_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__81_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___264_comb = 9'h000;
  assign p1_concat_145657_comb = {p1_smul_58516_NarrowedMult__comb, p1_smul_57330_TrailingBits___265_comb};
  assign p1_concat_145658_comb = {p1_smul_58518_NarrowedMult__comb, p1_smul_57330_TrailingBits___266_comb};
  assign p1_smul_58522_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__86_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___267_comb = 9'h000;
  assign p1_smul_58528_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__89_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___268_comb = 9'h000;
  assign p1_concat_145663_comb = {p1_smul_58532_NarrowedMult__comb, p1_smul_57330_TrailingBits___269_comb};
  assign p1_concat_145664_comb = {p1_smul_58534_NarrowedMult__comb, p1_smul_57330_TrailingBits___270_comb};
  assign p1_smul_58538_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__94_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___271_comb = 9'h000;
  assign p1_smul_58544_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__97_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___272_comb = 9'h000;
  assign p1_concat_145669_comb = {p1_smul_58548_NarrowedMult__comb, p1_smul_57330_TrailingBits___273_comb};
  assign p1_concat_145670_comb = {p1_smul_58550_NarrowedMult__comb, p1_smul_57330_TrailingBits___274_comb};
  assign p1_smul_58554_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__102_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___275_comb = 9'h000;
  assign p1_smul_58560_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__105_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___276_comb = 9'h000;
  assign p1_concat_145675_comb = {p1_smul_58564_NarrowedMult__comb, p1_smul_57330_TrailingBits___277_comb};
  assign p1_concat_145676_comb = {p1_smul_58566_NarrowedMult__comb, p1_smul_57330_TrailingBits___278_comb};
  assign p1_smul_58570_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__110_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___279_comb = 9'h000;
  assign p1_smul_58576_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__113_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___280_comb = 9'h000;
  assign p1_concat_145681_comb = {p1_smul_58580_NarrowedMult__comb, p1_smul_57330_TrailingBits___281_comb};
  assign p1_concat_145682_comb = {p1_smul_58582_NarrowedMult__comb, p1_smul_57330_TrailingBits___282_comb};
  assign p1_smul_58586_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__118_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___283_comb = 9'h000;
  assign p1_smul_58592_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__121_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___284_comb = 9'h000;
  assign p1_concat_145687_comb = {p1_smul_58596_NarrowedMult__comb, p1_smul_57330_TrailingBits___285_comb};
  assign p1_concat_145688_comb = {p1_smul_58598_NarrowedMult__comb, p1_smul_57330_TrailingBits___286_comb};
  assign p1_smul_58602_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__126_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___287_comb = 9'h000;
  assign p1_concat_145691_comb = {p1_smul_58734_NarrowedMult__comb, p1_smul_57330_TrailingBits___288_comb};
  assign p1_smul_58738_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__66_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___289_comb = 9'h000;
  assign p1_smul_58744_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__69_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___290_comb = 9'h000;
  assign p1_concat_145696_comb = {p1_smul_58748_NarrowedMult__comb, p1_smul_57330_TrailingBits___291_comb};
  assign p1_concat_145697_comb = {p1_smul_58750_NarrowedMult__comb, p1_smul_57330_TrailingBits___292_comb};
  assign p1_smul_58754_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__74_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___293_comb = 9'h000;
  assign p1_smul_58760_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__77_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___294_comb = 9'h000;
  assign p1_concat_145702_comb = {p1_smul_58764_NarrowedMult__comb, p1_smul_57330_TrailingBits___295_comb};
  assign p1_concat_145703_comb = {p1_smul_58766_NarrowedMult__comb, p1_smul_57330_TrailingBits___296_comb};
  assign p1_smul_58770_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__82_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___297_comb = 9'h000;
  assign p1_smul_58776_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__85_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___298_comb = 9'h000;
  assign p1_concat_145708_comb = {p1_smul_58780_NarrowedMult__comb, p1_smul_57330_TrailingBits___299_comb};
  assign p1_concat_145709_comb = {p1_smul_58782_NarrowedMult__comb, p1_smul_57330_TrailingBits___300_comb};
  assign p1_smul_58786_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__90_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___301_comb = 9'h000;
  assign p1_smul_58792_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__93_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___302_comb = 9'h000;
  assign p1_concat_145714_comb = {p1_smul_58796_NarrowedMult__comb, p1_smul_57330_TrailingBits___303_comb};
  assign p1_concat_145715_comb = {p1_smul_58798_NarrowedMult__comb, p1_smul_57330_TrailingBits___304_comb};
  assign p1_smul_58802_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__98_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___305_comb = 9'h000;
  assign p1_smul_58808_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__101_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___306_comb = 9'h000;
  assign p1_concat_145720_comb = {p1_smul_58812_NarrowedMult__comb, p1_smul_57330_TrailingBits___307_comb};
  assign p1_concat_145721_comb = {p1_smul_58814_NarrowedMult__comb, p1_smul_57330_TrailingBits___308_comb};
  assign p1_smul_58818_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__106_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___309_comb = 9'h000;
  assign p1_smul_58824_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__109_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___310_comb = 9'h000;
  assign p1_concat_145726_comb = {p1_smul_58828_NarrowedMult__comb, p1_smul_57330_TrailingBits___311_comb};
  assign p1_concat_145727_comb = {p1_smul_58830_NarrowedMult__comb, p1_smul_57330_TrailingBits___312_comb};
  assign p1_smul_58834_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__114_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___313_comb = 9'h000;
  assign p1_smul_58840_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__117_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___314_comb = 9'h000;
  assign p1_concat_145732_comb = {p1_smul_58844_NarrowedMult__comb, p1_smul_57330_TrailingBits___315_comb};
  assign p1_concat_145733_comb = {p1_smul_58846_NarrowedMult__comb, p1_smul_57330_TrailingBits___316_comb};
  assign p1_smul_58850_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__122_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___317_comb = 9'h000;
  assign p1_smul_58856_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__125_squeezed_comb, 6'h27);
  assign p1_smul_57330_TrailingBits___318_comb = 9'h000;
  assign p1_concat_145738_comb = {p1_smul_58860_NarrowedMult__comb, p1_smul_57330_TrailingBits___319_comb};
  assign p1_concat_145739_comb = {p1_smul_58862_NarrowedMult__comb, p1_smul_57330_TrailingBits___320_comb};
  assign p1_concat_145740_comb = {p1_smul_58864_NarrowedMult__comb, p1_smul_57454_TrailingBits___96_comb};
  assign p1_concat_145741_comb = {p1_smul_58866_NarrowedMult__comb, p1_smul_57330_TrailingBits___321_comb};
  assign p1_concat_145742_comb = {p1_smul_58868_NarrowedMult__comb, p1_smul_57454_TrailingBits___97_comb};
  assign p1_concat_145743_comb = {p1_smul_58870_NarrowedMult__comb, p1_smul_57454_TrailingBits___98_comb};
  assign p1_concat_145744_comb = {p1_smul_58872_NarrowedMult__comb, p1_smul_57330_TrailingBits___322_comb};
  assign p1_concat_145745_comb = {p1_smul_58874_NarrowedMult__comb, p1_smul_57454_TrailingBits___99_comb};
  assign p1_concat_145746_comb = {p1_smul_58876_NarrowedMult__comb, p1_smul_57330_TrailingBits___323_comb};
  assign p1_concat_145747_comb = {p1_smul_58878_NarrowedMult__comb, p1_smul_57330_TrailingBits___324_comb};
  assign p1_concat_145748_comb = {p1_smul_58880_NarrowedMult__comb, p1_smul_57454_TrailingBits___100_comb};
  assign p1_concat_145749_comb = {p1_smul_58882_NarrowedMult__comb, p1_smul_57330_TrailingBits___325_comb};
  assign p1_concat_145750_comb = {p1_smul_58884_NarrowedMult__comb, p1_smul_57454_TrailingBits___101_comb};
  assign p1_concat_145751_comb = {p1_smul_58886_NarrowedMult__comb, p1_smul_57454_TrailingBits___102_comb};
  assign p1_concat_145752_comb = {p1_smul_58888_NarrowedMult__comb, p1_smul_57330_TrailingBits___326_comb};
  assign p1_concat_145753_comb = {p1_smul_58890_NarrowedMult__comb, p1_smul_57454_TrailingBits___103_comb};
  assign p1_concat_145754_comb = {p1_smul_58892_NarrowedMult__comb, p1_smul_57330_TrailingBits___327_comb};
  assign p1_concat_145755_comb = {p1_smul_58894_NarrowedMult__comb, p1_smul_57330_TrailingBits___328_comb};
  assign p1_concat_145756_comb = {p1_smul_58896_NarrowedMult__comb, p1_smul_57454_TrailingBits___104_comb};
  assign p1_concat_145757_comb = {p1_smul_58898_NarrowedMult__comb, p1_smul_57330_TrailingBits___329_comb};
  assign p1_concat_145758_comb = {p1_smul_58900_NarrowedMult__comb, p1_smul_57454_TrailingBits___105_comb};
  assign p1_concat_145759_comb = {p1_smul_58902_NarrowedMult__comb, p1_smul_57454_TrailingBits___106_comb};
  assign p1_concat_145760_comb = {p1_smul_58904_NarrowedMult__comb, p1_smul_57330_TrailingBits___330_comb};
  assign p1_concat_145761_comb = {p1_smul_58906_NarrowedMult__comb, p1_smul_57454_TrailingBits___107_comb};
  assign p1_concat_145762_comb = {p1_smul_58908_NarrowedMult__comb, p1_smul_57330_TrailingBits___331_comb};
  assign p1_concat_145763_comb = {p1_smul_58910_NarrowedMult__comb, p1_smul_57330_TrailingBits___332_comb};
  assign p1_concat_145764_comb = {p1_smul_58912_NarrowedMult__comb, p1_smul_57454_TrailingBits___108_comb};
  assign p1_concat_145765_comb = {p1_smul_58914_NarrowedMult__comb, p1_smul_57330_TrailingBits___333_comb};
  assign p1_concat_145766_comb = {p1_smul_58916_NarrowedMult__comb, p1_smul_57454_TrailingBits___109_comb};
  assign p1_concat_145767_comb = {p1_smul_58918_NarrowedMult__comb, p1_smul_57454_TrailingBits___110_comb};
  assign p1_concat_145768_comb = {p1_smul_58920_NarrowedMult__comb, p1_smul_57330_TrailingBits___334_comb};
  assign p1_concat_145769_comb = {p1_smul_58922_NarrowedMult__comb, p1_smul_57454_TrailingBits___111_comb};
  assign p1_concat_145770_comb = {p1_smul_58924_NarrowedMult__comb, p1_smul_57330_TrailingBits___335_comb};
  assign p1_concat_145771_comb = {p1_smul_58926_NarrowedMult__comb, p1_smul_57330_TrailingBits___336_comb};
  assign p1_concat_145772_comb = {p1_smul_58928_NarrowedMult__comb, p1_smul_57454_TrailingBits___112_comb};
  assign p1_concat_145773_comb = {p1_smul_58930_NarrowedMult__comb, p1_smul_57330_TrailingBits___337_comb};
  assign p1_concat_145774_comb = {p1_smul_58932_NarrowedMult__comb, p1_smul_57454_TrailingBits___113_comb};
  assign p1_concat_145775_comb = {p1_smul_58934_NarrowedMult__comb, p1_smul_57454_TrailingBits___114_comb};
  assign p1_concat_145776_comb = {p1_smul_58936_NarrowedMult__comb, p1_smul_57330_TrailingBits___338_comb};
  assign p1_concat_145777_comb = {p1_smul_58938_NarrowedMult__comb, p1_smul_57454_TrailingBits___115_comb};
  assign p1_concat_145778_comb = {p1_smul_58940_NarrowedMult__comb, p1_smul_57330_TrailingBits___339_comb};
  assign p1_concat_145779_comb = {p1_smul_58942_NarrowedMult__comb, p1_smul_57330_TrailingBits___340_comb};
  assign p1_concat_145780_comb = {p1_smul_58944_NarrowedMult__comb, p1_smul_57454_TrailingBits___116_comb};
  assign p1_concat_145781_comb = {p1_smul_58946_NarrowedMult__comb, p1_smul_57330_TrailingBits___341_comb};
  assign p1_concat_145782_comb = {p1_smul_58948_NarrowedMult__comb, p1_smul_57454_TrailingBits___117_comb};
  assign p1_concat_145783_comb = {p1_smul_58950_NarrowedMult__comb, p1_smul_57454_TrailingBits___118_comb};
  assign p1_concat_145784_comb = {p1_smul_58952_NarrowedMult__comb, p1_smul_57330_TrailingBits___342_comb};
  assign p1_concat_145785_comb = {p1_smul_58954_NarrowedMult__comb, p1_smul_57454_TrailingBits___119_comb};
  assign p1_concat_145786_comb = {p1_smul_58956_NarrowedMult__comb, p1_smul_57330_TrailingBits___343_comb};
  assign p1_concat_145787_comb = {p1_smul_58958_NarrowedMult__comb, p1_smul_57330_TrailingBits___344_comb};
  assign p1_concat_145788_comb = {p1_smul_58960_NarrowedMult__comb, p1_smul_57454_TrailingBits___120_comb};
  assign p1_concat_145789_comb = {p1_smul_58962_NarrowedMult__comb, p1_smul_57330_TrailingBits___345_comb};
  assign p1_concat_145790_comb = {p1_smul_58964_NarrowedMult__comb, p1_smul_57454_TrailingBits___121_comb};
  assign p1_concat_145791_comb = {p1_smul_58966_NarrowedMult__comb, p1_smul_57454_TrailingBits___122_comb};
  assign p1_concat_145792_comb = {p1_smul_58968_NarrowedMult__comb, p1_smul_57330_TrailingBits___346_comb};
  assign p1_concat_145793_comb = {p1_smul_58970_NarrowedMult__comb, p1_smul_57454_TrailingBits___123_comb};
  assign p1_concat_145794_comb = {p1_smul_58972_NarrowedMult__comb, p1_smul_57330_TrailingBits___347_comb};
  assign p1_concat_145795_comb = {p1_smul_58974_NarrowedMult__comb, p1_smul_57330_TrailingBits___348_comb};
  assign p1_concat_145796_comb = {p1_smul_58976_NarrowedMult__comb, p1_smul_57454_TrailingBits___124_comb};
  assign p1_concat_145797_comb = {p1_smul_58978_NarrowedMult__comb, p1_smul_57330_TrailingBits___349_comb};
  assign p1_concat_145798_comb = {p1_smul_58980_NarrowedMult__comb, p1_smul_57454_TrailingBits___125_comb};
  assign p1_concat_145799_comb = {p1_smul_58982_NarrowedMult__comb, p1_smul_57454_TrailingBits___126_comb};
  assign p1_concat_145800_comb = {p1_smul_58984_NarrowedMult__comb, p1_smul_57330_TrailingBits___350_comb};
  assign p1_concat_145801_comb = {p1_smul_58986_NarrowedMult__comb, p1_smul_57454_TrailingBits___127_comb};
  assign p1_concat_145802_comb = {p1_smul_58988_NarrowedMult__comb, p1_smul_57330_TrailingBits___351_comb};
  assign p1_smul_58990_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__64_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___352_comb = 9'h000;
  assign p1_concat_145805_comb = {p1_smul_58992_NarrowedMult__comb, p1_smul_57330_TrailingBits___353_comb};
  assign p1_concat_145806_comb = {p1_smul_59002_NarrowedMult__comb, p1_smul_57330_TrailingBits___354_comb};
  assign p1_smul_59004_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__71_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___355_comb = 9'h000;
  assign p1_smul_59006_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__72_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___356_comb = 9'h000;
  assign p1_concat_145811_comb = {p1_smul_59008_NarrowedMult__comb, p1_smul_57330_TrailingBits___357_comb};
  assign p1_concat_145812_comb = {p1_smul_59018_NarrowedMult__comb, p1_smul_57330_TrailingBits___358_comb};
  assign p1_smul_59020_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__79_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___359_comb = 9'h000;
  assign p1_smul_59022_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__80_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___360_comb = 9'h000;
  assign p1_concat_145817_comb = {p1_smul_59024_NarrowedMult__comb, p1_smul_57330_TrailingBits___361_comb};
  assign p1_concat_145818_comb = {p1_smul_59034_NarrowedMult__comb, p1_smul_57330_TrailingBits___362_comb};
  assign p1_smul_59036_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__87_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___363_comb = 9'h000;
  assign p1_smul_59038_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__88_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___364_comb = 9'h000;
  assign p1_concat_145823_comb = {p1_smul_59040_NarrowedMult__comb, p1_smul_57330_TrailingBits___365_comb};
  assign p1_concat_145824_comb = {p1_smul_59050_NarrowedMult__comb, p1_smul_57330_TrailingBits___366_comb};
  assign p1_smul_59052_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__95_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___367_comb = 9'h000;
  assign p1_smul_59054_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__96_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___368_comb = 9'h000;
  assign p1_concat_145829_comb = {p1_smul_59056_NarrowedMult__comb, p1_smul_57330_TrailingBits___369_comb};
  assign p1_concat_145830_comb = {p1_smul_59066_NarrowedMult__comb, p1_smul_57330_TrailingBits___370_comb};
  assign p1_smul_59068_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__103_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___371_comb = 9'h000;
  assign p1_smul_59070_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__104_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___372_comb = 9'h000;
  assign p1_concat_145835_comb = {p1_smul_59072_NarrowedMult__comb, p1_smul_57330_TrailingBits___373_comb};
  assign p1_concat_145836_comb = {p1_smul_59082_NarrowedMult__comb, p1_smul_57330_TrailingBits___374_comb};
  assign p1_smul_59084_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__111_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___375_comb = 9'h000;
  assign p1_smul_59086_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__112_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___376_comb = 9'h000;
  assign p1_concat_145841_comb = {p1_smul_59088_NarrowedMult__comb, p1_smul_57330_TrailingBits___377_comb};
  assign p1_concat_145842_comb = {p1_smul_59098_NarrowedMult__comb, p1_smul_57330_TrailingBits___378_comb};
  assign p1_smul_59100_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__119_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___379_comb = 9'h000;
  assign p1_smul_59102_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__120_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___380_comb = 9'h000;
  assign p1_concat_145847_comb = {p1_smul_59104_NarrowedMult__comb, p1_smul_57330_TrailingBits___381_comb};
  assign p1_concat_145848_comb = {p1_smul_59114_NarrowedMult__comb, p1_smul_57330_TrailingBits___382_comb};
  assign p1_smul_59116_NarrowedMult__comb = smul14b_8b_x_6b(p1_shifted__127_squeezed_comb, 6'h19);
  assign p1_smul_57330_TrailingBits___383_comb = 9'h000;
  assign p1_smul_57326_TrailingBits___192_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___193_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___194_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___195_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___196_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___197_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___198_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___199_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___200_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___201_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___202_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___203_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___204_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___205_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___206_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___207_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___208_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___209_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___210_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___211_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___212_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___213_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___214_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___215_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___216_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___217_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___218_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___219_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___220_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___221_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___222_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___223_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___224_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___225_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___226_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___227_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___228_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___229_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___230_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___231_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___232_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___233_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___234_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___235_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___236_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___237_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___238_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___239_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___240_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___241_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___242_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___243_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___244_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___245_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___246_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___247_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___248_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___249_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___250_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___251_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___252_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___253_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___254_comb = 8'h00;
  assign p1_smul_57326_TrailingBits___255_comb = 8'h00;
  assign p1_prod__519_comb = {{7{p1_concat_145531_comb[24]}}, p1_concat_145531_comb};
  assign p1_concat_146045_comb = {p1_smul_58228_NarrowedMult__comb, p1_smul_57330_TrailingBits___193_comb};
  assign p1_concat_146046_comb = {p1_smul_58230_NarrowedMult__comb, p1_smul_57330_TrailingBits___194_comb};
  assign p1_prod__534_comb = {{7{p1_concat_145536_comb[24]}}, p1_concat_145536_comb};
  assign p1_prod__583_comb = {{7{p1_concat_145537_comb[24]}}, p1_concat_145537_comb};
  assign p1_concat_146051_comb = {p1_smul_58244_NarrowedMult__comb, p1_smul_57330_TrailingBits___197_comb};
  assign p1_concat_146052_comb = {p1_smul_58246_NarrowedMult__comb, p1_smul_57330_TrailingBits___198_comb};
  assign p1_prod__598_comb = {{7{p1_concat_145542_comb[24]}}, p1_concat_145542_comb};
  assign p1_prod__647_comb = {{7{p1_concat_145543_comb[24]}}, p1_concat_145543_comb};
  assign p1_concat_146057_comb = {p1_smul_58260_NarrowedMult__comb, p1_smul_57330_TrailingBits___201_comb};
  assign p1_concat_146058_comb = {p1_smul_58262_NarrowedMult__comb, p1_smul_57330_TrailingBits___202_comb};
  assign p1_prod__662_comb = {{7{p1_concat_145548_comb[24]}}, p1_concat_145548_comb};
  assign p1_prod__711_comb = {{7{p1_concat_145549_comb[24]}}, p1_concat_145549_comb};
  assign p1_concat_146063_comb = {p1_smul_58276_NarrowedMult__comb, p1_smul_57330_TrailingBits___205_comb};
  assign p1_concat_146064_comb = {p1_smul_58278_NarrowedMult__comb, p1_smul_57330_TrailingBits___206_comb};
  assign p1_prod__726_comb = {{7{p1_concat_145554_comb[24]}}, p1_concat_145554_comb};
  assign p1_prod__775_comb = {{7{p1_concat_145555_comb[24]}}, p1_concat_145555_comb};
  assign p1_concat_146069_comb = {p1_smul_58292_NarrowedMult__comb, p1_smul_57330_TrailingBits___209_comb};
  assign p1_concat_146070_comb = {p1_smul_58294_NarrowedMult__comb, p1_smul_57330_TrailingBits___210_comb};
  assign p1_prod__790_comb = {{7{p1_concat_145560_comb[24]}}, p1_concat_145560_comb};
  assign p1_prod__839_comb = {{7{p1_concat_145561_comb[24]}}, p1_concat_145561_comb};
  assign p1_concat_146075_comb = {p1_smul_58308_NarrowedMult__comb, p1_smul_57330_TrailingBits___213_comb};
  assign p1_concat_146076_comb = {p1_smul_58310_NarrowedMult__comb, p1_smul_57330_TrailingBits___214_comb};
  assign p1_prod__854_comb = {{7{p1_concat_145566_comb[24]}}, p1_concat_145566_comb};
  assign p1_prod__903_comb = {{7{p1_concat_145567_comb[24]}}, p1_concat_145567_comb};
  assign p1_concat_146081_comb = {p1_smul_58324_NarrowedMult__comb, p1_smul_57330_TrailingBits___217_comb};
  assign p1_concat_146082_comb = {p1_smul_58326_NarrowedMult__comb, p1_smul_57330_TrailingBits___218_comb};
  assign p1_prod__918_comb = {{7{p1_concat_145572_comb[24]}}, p1_concat_145572_comb};
  assign p1_prod__967_comb = {{7{p1_concat_145573_comb[24]}}, p1_concat_145573_comb};
  assign p1_concat_146087_comb = {p1_smul_58340_NarrowedMult__comb, p1_smul_57330_TrailingBits___221_comb};
  assign p1_concat_146088_comb = {p1_smul_58342_NarrowedMult__comb, p1_smul_57330_TrailingBits___222_comb};
  assign p1_prod__982_comb = {{7{p1_concat_145578_comb[24]}}, p1_concat_145578_comb};
  assign p1_prod__517_comb = {{7{p1_concat_145579_comb[24]}}, p1_concat_145579_comb};
  assign p1_prod__520_comb = {{8{p1_concat_145580_comb[23]}}, p1_concat_145580_comb};
  assign p1_prod__524_comb = {{8{p1_concat_145581_comb[23]}}, p1_concat_145581_comb};
  assign p1_prod__529_comb = {{7{p1_concat_145582_comb[24]}}, p1_concat_145582_comb};
  assign p1_prod__535_comb = {{7{p1_concat_145583_comb[24]}}, p1_concat_145583_comb};
  assign p1_prod__542_comb = {{8{p1_concat_145584_comb[23]}}, p1_concat_145584_comb};
  assign p1_prod__549_comb = {{8{p1_concat_145585_comb[23]}}, p1_concat_145585_comb};
  assign p1_prod__555_comb = {{7{p1_concat_145586_comb[24]}}, p1_concat_145586_comb};
  assign p1_prod__581_comb = {{7{p1_concat_145587_comb[24]}}, p1_concat_145587_comb};
  assign p1_prod__584_comb = {{8{p1_concat_145588_comb[23]}}, p1_concat_145588_comb};
  assign p1_prod__588_comb = {{8{p1_concat_145589_comb[23]}}, p1_concat_145589_comb};
  assign p1_prod__593_comb = {{7{p1_concat_145590_comb[24]}}, p1_concat_145590_comb};
  assign p1_prod__599_comb = {{7{p1_concat_145591_comb[24]}}, p1_concat_145591_comb};
  assign p1_prod__606_comb = {{8{p1_concat_145592_comb[23]}}, p1_concat_145592_comb};
  assign p1_prod__613_comb = {{8{p1_concat_145593_comb[23]}}, p1_concat_145593_comb};
  assign p1_prod__619_comb = {{7{p1_concat_145594_comb[24]}}, p1_concat_145594_comb};
  assign p1_prod__645_comb = {{7{p1_concat_145595_comb[24]}}, p1_concat_145595_comb};
  assign p1_prod__648_comb = {{8{p1_concat_145596_comb[23]}}, p1_concat_145596_comb};
  assign p1_prod__652_comb = {{8{p1_concat_145597_comb[23]}}, p1_concat_145597_comb};
  assign p1_prod__657_comb = {{7{p1_concat_145598_comb[24]}}, p1_concat_145598_comb};
  assign p1_prod__663_comb = {{7{p1_concat_145599_comb[24]}}, p1_concat_145599_comb};
  assign p1_prod__670_comb = {{8{p1_concat_145600_comb[23]}}, p1_concat_145600_comb};
  assign p1_prod__677_comb = {{8{p1_concat_145601_comb[23]}}, p1_concat_145601_comb};
  assign p1_prod__683_comb = {{7{p1_concat_145602_comb[24]}}, p1_concat_145602_comb};
  assign p1_prod__709_comb = {{7{p1_concat_145603_comb[24]}}, p1_concat_145603_comb};
  assign p1_prod__712_comb = {{8{p1_concat_145604_comb[23]}}, p1_concat_145604_comb};
  assign p1_prod__716_comb = {{8{p1_concat_145605_comb[23]}}, p1_concat_145605_comb};
  assign p1_prod__721_comb = {{7{p1_concat_145606_comb[24]}}, p1_concat_145606_comb};
  assign p1_prod__727_comb = {{7{p1_concat_145607_comb[24]}}, p1_concat_145607_comb};
  assign p1_prod__734_comb = {{8{p1_concat_145608_comb[23]}}, p1_concat_145608_comb};
  assign p1_prod__741_comb = {{8{p1_concat_145609_comb[23]}}, p1_concat_145609_comb};
  assign p1_prod__747_comb = {{7{p1_concat_145610_comb[24]}}, p1_concat_145610_comb};
  assign p1_prod__773_comb = {{7{p1_concat_145611_comb[24]}}, p1_concat_145611_comb};
  assign p1_prod__776_comb = {{8{p1_concat_145612_comb[23]}}, p1_concat_145612_comb};
  assign p1_prod__780_comb = {{8{p1_concat_145613_comb[23]}}, p1_concat_145613_comb};
  assign p1_prod__785_comb = {{7{p1_concat_145614_comb[24]}}, p1_concat_145614_comb};
  assign p1_prod__791_comb = {{7{p1_concat_145615_comb[24]}}, p1_concat_145615_comb};
  assign p1_prod__798_comb = {{8{p1_concat_145616_comb[23]}}, p1_concat_145616_comb};
  assign p1_prod__805_comb = {{8{p1_concat_145617_comb[23]}}, p1_concat_145617_comb};
  assign p1_prod__811_comb = {{7{p1_concat_145618_comb[24]}}, p1_concat_145618_comb};
  assign p1_prod__837_comb = {{7{p1_concat_145619_comb[24]}}, p1_concat_145619_comb};
  assign p1_prod__840_comb = {{8{p1_concat_145620_comb[23]}}, p1_concat_145620_comb};
  assign p1_prod__844_comb = {{8{p1_concat_145621_comb[23]}}, p1_concat_145621_comb};
  assign p1_prod__849_comb = {{7{p1_concat_145622_comb[24]}}, p1_concat_145622_comb};
  assign p1_prod__855_comb = {{7{p1_concat_145623_comb[24]}}, p1_concat_145623_comb};
  assign p1_prod__862_comb = {{8{p1_concat_145624_comb[23]}}, p1_concat_145624_comb};
  assign p1_prod__869_comb = {{8{p1_concat_145625_comb[23]}}, p1_concat_145625_comb};
  assign p1_prod__875_comb = {{7{p1_concat_145626_comb[24]}}, p1_concat_145626_comb};
  assign p1_prod__901_comb = {{7{p1_concat_145627_comb[24]}}, p1_concat_145627_comb};
  assign p1_prod__904_comb = {{8{p1_concat_145628_comb[23]}}, p1_concat_145628_comb};
  assign p1_prod__908_comb = {{8{p1_concat_145629_comb[23]}}, p1_concat_145629_comb};
  assign p1_prod__913_comb = {{7{p1_concat_145630_comb[24]}}, p1_concat_145630_comb};
  assign p1_prod__919_comb = {{7{p1_concat_145631_comb[24]}}, p1_concat_145631_comb};
  assign p1_prod__926_comb = {{8{p1_concat_145632_comb[23]}}, p1_concat_145632_comb};
  assign p1_prod__933_comb = {{8{p1_concat_145633_comb[23]}}, p1_concat_145633_comb};
  assign p1_prod__939_comb = {{7{p1_concat_145634_comb[24]}}, p1_concat_145634_comb};
  assign p1_prod__965_comb = {{7{p1_concat_145635_comb[24]}}, p1_concat_145635_comb};
  assign p1_prod__968_comb = {{8{p1_concat_145636_comb[23]}}, p1_concat_145636_comb};
  assign p1_prod__972_comb = {{8{p1_concat_145637_comb[23]}}, p1_concat_145637_comb};
  assign p1_prod__977_comb = {{7{p1_concat_145638_comb[24]}}, p1_concat_145638_comb};
  assign p1_prod__983_comb = {{7{p1_concat_145639_comb[24]}}, p1_concat_145639_comb};
  assign p1_prod__990_comb = {{8{p1_concat_145640_comb[23]}}, p1_concat_145640_comb};
  assign p1_prod__997_comb = {{8{p1_concat_145641_comb[23]}}, p1_concat_145641_comb};
  assign p1_prod__1003_comb = {{7{p1_concat_145642_comb[24]}}, p1_concat_145642_comb};
  assign p1_concat_146187_comb = {p1_smul_58480_NarrowedMult__comb, p1_smul_57330_TrailingBits___256_comb};
  assign p1_prod__536_comb = {{7{p1_concat_145645_comb[24]}}, p1_concat_145645_comb};
  assign p1_prod__543_comb = {{7{p1_concat_145646_comb[24]}}, p1_concat_145646_comb};
  assign p1_concat_146192_comb = {p1_smul_58490_NarrowedMult__comb, p1_smul_57330_TrailingBits___259_comb};
  assign p1_concat_146193_comb = {p1_smul_58496_NarrowedMult__comb, p1_smul_57330_TrailingBits___260_comb};
  assign p1_prod__600_comb = {{7{p1_concat_145651_comb[24]}}, p1_concat_145651_comb};
  assign p1_prod__607_comb = {{7{p1_concat_145652_comb[24]}}, p1_concat_145652_comb};
  assign p1_concat_146198_comb = {p1_smul_58506_NarrowedMult__comb, p1_smul_57330_TrailingBits___263_comb};
  assign p1_concat_146199_comb = {p1_smul_58512_NarrowedMult__comb, p1_smul_57330_TrailingBits___264_comb};
  assign p1_prod__664_comb = {{7{p1_concat_145657_comb[24]}}, p1_concat_145657_comb};
  assign p1_prod__671_comb = {{7{p1_concat_145658_comb[24]}}, p1_concat_145658_comb};
  assign p1_concat_146204_comb = {p1_smul_58522_NarrowedMult__comb, p1_smul_57330_TrailingBits___267_comb};
  assign p1_concat_146205_comb = {p1_smul_58528_NarrowedMult__comb, p1_smul_57330_TrailingBits___268_comb};
  assign p1_prod__728_comb = {{7{p1_concat_145663_comb[24]}}, p1_concat_145663_comb};
  assign p1_prod__735_comb = {{7{p1_concat_145664_comb[24]}}, p1_concat_145664_comb};
  assign p1_concat_146210_comb = {p1_smul_58538_NarrowedMult__comb, p1_smul_57330_TrailingBits___271_comb};
  assign p1_concat_146211_comb = {p1_smul_58544_NarrowedMult__comb, p1_smul_57330_TrailingBits___272_comb};
  assign p1_prod__792_comb = {{7{p1_concat_145669_comb[24]}}, p1_concat_145669_comb};
  assign p1_prod__799_comb = {{7{p1_concat_145670_comb[24]}}, p1_concat_145670_comb};
  assign p1_concat_146216_comb = {p1_smul_58554_NarrowedMult__comb, p1_smul_57330_TrailingBits___275_comb};
  assign p1_concat_146217_comb = {p1_smul_58560_NarrowedMult__comb, p1_smul_57330_TrailingBits___276_comb};
  assign p1_prod__856_comb = {{7{p1_concat_145675_comb[24]}}, p1_concat_145675_comb};
  assign p1_prod__863_comb = {{7{p1_concat_145676_comb[24]}}, p1_concat_145676_comb};
  assign p1_concat_146222_comb = {p1_smul_58570_NarrowedMult__comb, p1_smul_57330_TrailingBits___279_comb};
  assign p1_concat_146223_comb = {p1_smul_58576_NarrowedMult__comb, p1_smul_57330_TrailingBits___280_comb};
  assign p1_prod__920_comb = {{7{p1_concat_145681_comb[24]}}, p1_concat_145681_comb};
  assign p1_prod__927_comb = {{7{p1_concat_145682_comb[24]}}, p1_concat_145682_comb};
  assign p1_concat_146228_comb = {p1_smul_58586_NarrowedMult__comb, p1_smul_57330_TrailingBits___283_comb};
  assign p1_concat_146229_comb = {p1_smul_58592_NarrowedMult__comb, p1_smul_57330_TrailingBits___284_comb};
  assign p1_prod__984_comb = {{7{p1_concat_145687_comb[24]}}, p1_concat_145687_comb};
  assign p1_prod__991_comb = {{7{p1_concat_145688_comb[24]}}, p1_concat_145688_comb};
  assign p1_concat_146234_comb = {p1_smul_58602_NarrowedMult__comb, p1_smul_57330_TrailingBits___287_comb};
  assign p1_prod__532_comb = {{7{p1_concat_145691_comb[24]}}, p1_concat_145691_comb};
  assign p1_concat_146237_comb = {p1_smul_58738_NarrowedMult__comb, p1_smul_57330_TrailingBits___289_comb};
  assign p1_concat_146238_comb = {p1_smul_58744_NarrowedMult__comb, p1_smul_57330_TrailingBits___290_comb};
  assign p1_prod__570_comb = {{7{p1_concat_145696_comb[24]}}, p1_concat_145696_comb};
  assign p1_prod__596_comb = {{7{p1_concat_145697_comb[24]}}, p1_concat_145697_comb};
  assign p1_concat_146243_comb = {p1_smul_58754_NarrowedMult__comb, p1_smul_57330_TrailingBits___293_comb};
  assign p1_concat_146244_comb = {p1_smul_58760_NarrowedMult__comb, p1_smul_57330_TrailingBits___294_comb};
  assign p1_prod__634_comb = {{7{p1_concat_145702_comb[24]}}, p1_concat_145702_comb};
  assign p1_prod__660_comb = {{7{p1_concat_145703_comb[24]}}, p1_concat_145703_comb};
  assign p1_concat_146249_comb = {p1_smul_58770_NarrowedMult__comb, p1_smul_57330_TrailingBits___297_comb};
  assign p1_concat_146250_comb = {p1_smul_58776_NarrowedMult__comb, p1_smul_57330_TrailingBits___298_comb};
  assign p1_prod__698_comb = {{7{p1_concat_145708_comb[24]}}, p1_concat_145708_comb};
  assign p1_prod__724_comb = {{7{p1_concat_145709_comb[24]}}, p1_concat_145709_comb};
  assign p1_concat_146255_comb = {p1_smul_58786_NarrowedMult__comb, p1_smul_57330_TrailingBits___301_comb};
  assign p1_concat_146256_comb = {p1_smul_58792_NarrowedMult__comb, p1_smul_57330_TrailingBits___302_comb};
  assign p1_prod__762_comb = {{7{p1_concat_145714_comb[24]}}, p1_concat_145714_comb};
  assign p1_prod__788_comb = {{7{p1_concat_145715_comb[24]}}, p1_concat_145715_comb};
  assign p1_concat_146261_comb = {p1_smul_58802_NarrowedMult__comb, p1_smul_57330_TrailingBits___305_comb};
  assign p1_concat_146262_comb = {p1_smul_58808_NarrowedMult__comb, p1_smul_57330_TrailingBits___306_comb};
  assign p1_prod__826_comb = {{7{p1_concat_145720_comb[24]}}, p1_concat_145720_comb};
  assign p1_prod__852_comb = {{7{p1_concat_145721_comb[24]}}, p1_concat_145721_comb};
  assign p1_concat_146267_comb = {p1_smul_58818_NarrowedMult__comb, p1_smul_57330_TrailingBits___309_comb};
  assign p1_concat_146268_comb = {p1_smul_58824_NarrowedMult__comb, p1_smul_57330_TrailingBits___310_comb};
  assign p1_prod__890_comb = {{7{p1_concat_145726_comb[24]}}, p1_concat_145726_comb};
  assign p1_prod__916_comb = {{7{p1_concat_145727_comb[24]}}, p1_concat_145727_comb};
  assign p1_concat_146273_comb = {p1_smul_58834_NarrowedMult__comb, p1_smul_57330_TrailingBits___313_comb};
  assign p1_concat_146274_comb = {p1_smul_58840_NarrowedMult__comb, p1_smul_57330_TrailingBits___314_comb};
  assign p1_prod__954_comb = {{7{p1_concat_145732_comb[24]}}, p1_concat_145732_comb};
  assign p1_prod__980_comb = {{7{p1_concat_145733_comb[24]}}, p1_concat_145733_comb};
  assign p1_concat_146279_comb = {p1_smul_58850_NarrowedMult__comb, p1_smul_57330_TrailingBits___317_comb};
  assign p1_concat_146280_comb = {p1_smul_58856_NarrowedMult__comb, p1_smul_57330_TrailingBits___318_comb};
  assign p1_prod__1018_comb = {{7{p1_concat_145738_comb[24]}}, p1_concat_145738_comb};
  assign p1_prod__539_comb = {{8{p1_concat_145739_comb[23]}}, p1_concat_145739_comb};
  assign p1_prod__546_comb = {{7{p1_concat_145740_comb[24]}}, p1_concat_145740_comb};
  assign p1_prod__553_comb = {{8{p1_concat_145741_comb[23]}}, p1_concat_145741_comb};
  assign p1_prod__559_comb = {{7{p1_concat_145742_comb[24]}}, p1_concat_145742_comb};
  assign p1_prod__564_comb = {{7{p1_concat_145743_comb[24]}}, p1_concat_145743_comb};
  assign p1_prod__568_comb = {{8{p1_concat_145744_comb[23]}}, p1_concat_145744_comb};
  assign p1_prod__571_comb = {{7{p1_concat_145745_comb[24]}}, p1_concat_145745_comb};
  assign p1_prod__573_comb = {{8{p1_concat_145746_comb[23]}}, p1_concat_145746_comb};
  assign p1_prod__603_comb = {{8{p1_concat_145747_comb[23]}}, p1_concat_145747_comb};
  assign p1_prod__610_comb = {{7{p1_concat_145748_comb[24]}}, p1_concat_145748_comb};
  assign p1_prod__617_comb = {{8{p1_concat_145749_comb[23]}}, p1_concat_145749_comb};
  assign p1_prod__623_comb = {{7{p1_concat_145750_comb[24]}}, p1_concat_145750_comb};
  assign p1_prod__628_comb = {{7{p1_concat_145751_comb[24]}}, p1_concat_145751_comb};
  assign p1_prod__632_comb = {{8{p1_concat_145752_comb[23]}}, p1_concat_145752_comb};
  assign p1_prod__635_comb = {{7{p1_concat_145753_comb[24]}}, p1_concat_145753_comb};
  assign p1_prod__637_comb = {{8{p1_concat_145754_comb[23]}}, p1_concat_145754_comb};
  assign p1_prod__667_comb = {{8{p1_concat_145755_comb[23]}}, p1_concat_145755_comb};
  assign p1_prod__674_comb = {{7{p1_concat_145756_comb[24]}}, p1_concat_145756_comb};
  assign p1_prod__681_comb = {{8{p1_concat_145757_comb[23]}}, p1_concat_145757_comb};
  assign p1_prod__687_comb = {{7{p1_concat_145758_comb[24]}}, p1_concat_145758_comb};
  assign p1_prod__692_comb = {{7{p1_concat_145759_comb[24]}}, p1_concat_145759_comb};
  assign p1_prod__696_comb = {{8{p1_concat_145760_comb[23]}}, p1_concat_145760_comb};
  assign p1_prod__699_comb = {{7{p1_concat_145761_comb[24]}}, p1_concat_145761_comb};
  assign p1_prod__701_comb = {{8{p1_concat_145762_comb[23]}}, p1_concat_145762_comb};
  assign p1_prod__731_comb = {{8{p1_concat_145763_comb[23]}}, p1_concat_145763_comb};
  assign p1_prod__738_comb = {{7{p1_concat_145764_comb[24]}}, p1_concat_145764_comb};
  assign p1_prod__745_comb = {{8{p1_concat_145765_comb[23]}}, p1_concat_145765_comb};
  assign p1_prod__751_comb = {{7{p1_concat_145766_comb[24]}}, p1_concat_145766_comb};
  assign p1_prod__756_comb = {{7{p1_concat_145767_comb[24]}}, p1_concat_145767_comb};
  assign p1_prod__760_comb = {{8{p1_concat_145768_comb[23]}}, p1_concat_145768_comb};
  assign p1_prod__763_comb = {{7{p1_concat_145769_comb[24]}}, p1_concat_145769_comb};
  assign p1_prod__765_comb = {{8{p1_concat_145770_comb[23]}}, p1_concat_145770_comb};
  assign p1_prod__795_comb = {{8{p1_concat_145771_comb[23]}}, p1_concat_145771_comb};
  assign p1_prod__802_comb = {{7{p1_concat_145772_comb[24]}}, p1_concat_145772_comb};
  assign p1_prod__809_comb = {{8{p1_concat_145773_comb[23]}}, p1_concat_145773_comb};
  assign p1_prod__815_comb = {{7{p1_concat_145774_comb[24]}}, p1_concat_145774_comb};
  assign p1_prod__820_comb = {{7{p1_concat_145775_comb[24]}}, p1_concat_145775_comb};
  assign p1_prod__824_comb = {{8{p1_concat_145776_comb[23]}}, p1_concat_145776_comb};
  assign p1_prod__827_comb = {{7{p1_concat_145777_comb[24]}}, p1_concat_145777_comb};
  assign p1_prod__829_comb = {{8{p1_concat_145778_comb[23]}}, p1_concat_145778_comb};
  assign p1_prod__859_comb = {{8{p1_concat_145779_comb[23]}}, p1_concat_145779_comb};
  assign p1_prod__866_comb = {{7{p1_concat_145780_comb[24]}}, p1_concat_145780_comb};
  assign p1_prod__873_comb = {{8{p1_concat_145781_comb[23]}}, p1_concat_145781_comb};
  assign p1_prod__879_comb = {{7{p1_concat_145782_comb[24]}}, p1_concat_145782_comb};
  assign p1_prod__884_comb = {{7{p1_concat_145783_comb[24]}}, p1_concat_145783_comb};
  assign p1_prod__888_comb = {{8{p1_concat_145784_comb[23]}}, p1_concat_145784_comb};
  assign p1_prod__891_comb = {{7{p1_concat_145785_comb[24]}}, p1_concat_145785_comb};
  assign p1_prod__893_comb = {{8{p1_concat_145786_comb[23]}}, p1_concat_145786_comb};
  assign p1_prod__923_comb = {{8{p1_concat_145787_comb[23]}}, p1_concat_145787_comb};
  assign p1_prod__930_comb = {{7{p1_concat_145788_comb[24]}}, p1_concat_145788_comb};
  assign p1_prod__937_comb = {{8{p1_concat_145789_comb[23]}}, p1_concat_145789_comb};
  assign p1_prod__943_comb = {{7{p1_concat_145790_comb[24]}}, p1_concat_145790_comb};
  assign p1_prod__948_comb = {{7{p1_concat_145791_comb[24]}}, p1_concat_145791_comb};
  assign p1_prod__952_comb = {{8{p1_concat_145792_comb[23]}}, p1_concat_145792_comb};
  assign p1_prod__955_comb = {{7{p1_concat_145793_comb[24]}}, p1_concat_145793_comb};
  assign p1_prod__957_comb = {{8{p1_concat_145794_comb[23]}}, p1_concat_145794_comb};
  assign p1_prod__987_comb = {{8{p1_concat_145795_comb[23]}}, p1_concat_145795_comb};
  assign p1_prod__994_comb = {{7{p1_concat_145796_comb[24]}}, p1_concat_145796_comb};
  assign p1_prod__1001_comb = {{8{p1_concat_145797_comb[23]}}, p1_concat_145797_comb};
  assign p1_prod__1007_comb = {{7{p1_concat_145798_comb[24]}}, p1_concat_145798_comb};
  assign p1_prod__1012_comb = {{7{p1_concat_145799_comb[24]}}, p1_concat_145799_comb};
  assign p1_prod__1016_comb = {{8{p1_concat_145800_comb[23]}}, p1_concat_145800_comb};
  assign p1_prod__1019_comb = {{7{p1_concat_145801_comb[24]}}, p1_concat_145801_comb};
  assign p1_prod__1021_comb = {{8{p1_concat_145802_comb[23]}}, p1_concat_145802_comb};
  assign p1_concat_146379_comb = {p1_smul_58990_NarrowedMult__comb, p1_smul_57330_TrailingBits___352_comb};
  assign p1_prod__554_comb = {{7{p1_concat_145805_comb[24]}}, p1_concat_145805_comb};
  assign p1_prod__574_comb = {{7{p1_concat_145806_comb[24]}}, p1_concat_145806_comb};
  assign p1_concat_146384_comb = {p1_smul_59004_NarrowedMult__comb, p1_smul_57330_TrailingBits___355_comb};
  assign p1_concat_146385_comb = {p1_smul_59006_NarrowedMult__comb, p1_smul_57330_TrailingBits___356_comb};
  assign p1_prod__618_comb = {{7{p1_concat_145811_comb[24]}}, p1_concat_145811_comb};
  assign p1_prod__638_comb = {{7{p1_concat_145812_comb[24]}}, p1_concat_145812_comb};
  assign p1_concat_146390_comb = {p1_smul_59020_NarrowedMult__comb, p1_smul_57330_TrailingBits___359_comb};
  assign p1_concat_146391_comb = {p1_smul_59022_NarrowedMult__comb, p1_smul_57330_TrailingBits___360_comb};
  assign p1_prod__682_comb = {{7{p1_concat_145817_comb[24]}}, p1_concat_145817_comb};
  assign p1_prod__702_comb = {{7{p1_concat_145818_comb[24]}}, p1_concat_145818_comb};
  assign p1_concat_146396_comb = {p1_smul_59036_NarrowedMult__comb, p1_smul_57330_TrailingBits___363_comb};
  assign p1_concat_146397_comb = {p1_smul_59038_NarrowedMult__comb, p1_smul_57330_TrailingBits___364_comb};
  assign p1_prod__746_comb = {{7{p1_concat_145823_comb[24]}}, p1_concat_145823_comb};
  assign p1_prod__766_comb = {{7{p1_concat_145824_comb[24]}}, p1_concat_145824_comb};
  assign p1_concat_146402_comb = {p1_smul_59052_NarrowedMult__comb, p1_smul_57330_TrailingBits___367_comb};
  assign p1_concat_146403_comb = {p1_smul_59054_NarrowedMult__comb, p1_smul_57330_TrailingBits___368_comb};
  assign p1_prod__810_comb = {{7{p1_concat_145829_comb[24]}}, p1_concat_145829_comb};
  assign p1_prod__830_comb = {{7{p1_concat_145830_comb[24]}}, p1_concat_145830_comb};
  assign p1_concat_146408_comb = {p1_smul_59068_NarrowedMult__comb, p1_smul_57330_TrailingBits___371_comb};
  assign p1_concat_146409_comb = {p1_smul_59070_NarrowedMult__comb, p1_smul_57330_TrailingBits___372_comb};
  assign p1_prod__874_comb = {{7{p1_concat_145835_comb[24]}}, p1_concat_145835_comb};
  assign p1_prod__894_comb = {{7{p1_concat_145836_comb[24]}}, p1_concat_145836_comb};
  assign p1_concat_146414_comb = {p1_smul_59084_NarrowedMult__comb, p1_smul_57330_TrailingBits___375_comb};
  assign p1_concat_146415_comb = {p1_smul_59086_NarrowedMult__comb, p1_smul_57330_TrailingBits___376_comb};
  assign p1_prod__938_comb = {{7{p1_concat_145841_comb[24]}}, p1_concat_145841_comb};
  assign p1_prod__958_comb = {{7{p1_concat_145842_comb[24]}}, p1_concat_145842_comb};
  assign p1_concat_146420_comb = {p1_smul_59100_NarrowedMult__comb, p1_smul_57330_TrailingBits___379_comb};
  assign p1_concat_146421_comb = {p1_smul_59102_NarrowedMult__comb, p1_smul_57330_TrailingBits___380_comb};
  assign p1_prod__1002_comb = {{7{p1_concat_145847_comb[24]}}, p1_concat_145847_comb};
  assign p1_prod__1022_comb = {{7{p1_concat_145848_comb[24]}}, p1_concat_145848_comb};
  assign p1_concat_146426_comb = {p1_smul_59116_NarrowedMult__comb, p1_smul_57330_TrailingBits___383_comb};
  assign p1_shifted__64_comb = {~p1_clipped__8_comb[7], p1_clipped__8_comb[6:0], p1_smul_57326_TrailingBits___192_comb};
  assign p1_smul_57326_TrailingBits___64_comb = 8'h00;
  assign p1_shifted__65_comb = {~p1_clipped__24_comb[7], p1_clipped__24_comb[6:0], p1_smul_57326_TrailingBits___193_comb};
  assign p1_smul_57326_TrailingBits___65_comb = 8'h00;
  assign p1_shifted__66_comb = {~p1_clipped__40_comb[7], p1_clipped__40_comb[6:0], p1_smul_57326_TrailingBits___194_comb};
  assign p1_smul_57326_TrailingBits___66_comb = 8'h00;
  assign p1_shifted__67_comb = {~p1_clipped__56_comb[7], p1_clipped__56_comb[6:0], p1_smul_57326_TrailingBits___195_comb};
  assign p1_smul_57326_TrailingBits___67_comb = 8'h00;
  assign p1_shifted__68_comb = {~p1_clipped__72_comb[7], p1_clipped__72_comb[6:0], p1_smul_57326_TrailingBits___196_comb};
  assign p1_smul_57326_TrailingBits___68_comb = 8'h00;
  assign p1_shifted__69_comb = {~p1_clipped__88_comb[7], p1_clipped__88_comb[6:0], p1_smul_57326_TrailingBits___197_comb};
  assign p1_smul_57326_TrailingBits___69_comb = 8'h00;
  assign p1_shifted__70_comb = {~p1_clipped__104_comb[7], p1_clipped__104_comb[6:0], p1_smul_57326_TrailingBits___198_comb};
  assign p1_smul_57326_TrailingBits___70_comb = 8'h00;
  assign p1_shifted__71_comb = {~p1_clipped__120_comb[7], p1_clipped__120_comb[6:0], p1_smul_57326_TrailingBits___199_comb};
  assign p1_smul_57326_TrailingBits___71_comb = 8'h00;
  assign p1_shifted__72_comb = {~p1_clipped__9_comb[7], p1_clipped__9_comb[6:0], p1_smul_57326_TrailingBits___200_comb};
  assign p1_smul_57326_TrailingBits___72_comb = 8'h00;
  assign p1_shifted__73_comb = {~p1_clipped__25_comb[7], p1_clipped__25_comb[6:0], p1_smul_57326_TrailingBits___201_comb};
  assign p1_smul_57326_TrailingBits___73_comb = 8'h00;
  assign p1_shifted__74_comb = {~p1_clipped__41_comb[7], p1_clipped__41_comb[6:0], p1_smul_57326_TrailingBits___202_comb};
  assign p1_smul_57326_TrailingBits___74_comb = 8'h00;
  assign p1_shifted__75_comb = {~p1_clipped__57_comb[7], p1_clipped__57_comb[6:0], p1_smul_57326_TrailingBits___203_comb};
  assign p1_smul_57326_TrailingBits___75_comb = 8'h00;
  assign p1_shifted__76_comb = {~p1_clipped__73_comb[7], p1_clipped__73_comb[6:0], p1_smul_57326_TrailingBits___204_comb};
  assign p1_smul_57326_TrailingBits___76_comb = 8'h00;
  assign p1_shifted__77_comb = {~p1_clipped__89_comb[7], p1_clipped__89_comb[6:0], p1_smul_57326_TrailingBits___205_comb};
  assign p1_smul_57326_TrailingBits___77_comb = 8'h00;
  assign p1_shifted__78_comb = {~p1_clipped__105_comb[7], p1_clipped__105_comb[6:0], p1_smul_57326_TrailingBits___206_comb};
  assign p1_smul_57326_TrailingBits___78_comb = 8'h00;
  assign p1_shifted__79_comb = {~p1_clipped__121_comb[7], p1_clipped__121_comb[6:0], p1_smul_57326_TrailingBits___207_comb};
  assign p1_smul_57326_TrailingBits___79_comb = 8'h00;
  assign p1_shifted__80_comb = {~p1_clipped__10_comb[7], p1_clipped__10_comb[6:0], p1_smul_57326_TrailingBits___208_comb};
  assign p1_smul_57326_TrailingBits___80_comb = 8'h00;
  assign p1_shifted__81_comb = {~p1_clipped__26_comb[7], p1_clipped__26_comb[6:0], p1_smul_57326_TrailingBits___209_comb};
  assign p1_smul_57326_TrailingBits___81_comb = 8'h00;
  assign p1_shifted__82_comb = {~p1_clipped__42_comb[7], p1_clipped__42_comb[6:0], p1_smul_57326_TrailingBits___210_comb};
  assign p1_smul_57326_TrailingBits___82_comb = 8'h00;
  assign p1_shifted__83_comb = {~p1_clipped__58_comb[7], p1_clipped__58_comb[6:0], p1_smul_57326_TrailingBits___211_comb};
  assign p1_smul_57326_TrailingBits___83_comb = 8'h00;
  assign p1_shifted__84_comb = {~p1_clipped__74_comb[7], p1_clipped__74_comb[6:0], p1_smul_57326_TrailingBits___212_comb};
  assign p1_smul_57326_TrailingBits___84_comb = 8'h00;
  assign p1_shifted__85_comb = {~p1_clipped__90_comb[7], p1_clipped__90_comb[6:0], p1_smul_57326_TrailingBits___213_comb};
  assign p1_smul_57326_TrailingBits___85_comb = 8'h00;
  assign p1_shifted__86_comb = {~p1_clipped__106_comb[7], p1_clipped__106_comb[6:0], p1_smul_57326_TrailingBits___214_comb};
  assign p1_smul_57326_TrailingBits___86_comb = 8'h00;
  assign p1_shifted__87_comb = {~p1_clipped__122_comb[7], p1_clipped__122_comb[6:0], p1_smul_57326_TrailingBits___215_comb};
  assign p1_smul_57326_TrailingBits___87_comb = 8'h00;
  assign p1_shifted__88_comb = {~p1_clipped__11_comb[7], p1_clipped__11_comb[6:0], p1_smul_57326_TrailingBits___216_comb};
  assign p1_smul_57326_TrailingBits___88_comb = 8'h00;
  assign p1_shifted__89_comb = {~p1_clipped__27_comb[7], p1_clipped__27_comb[6:0], p1_smul_57326_TrailingBits___217_comb};
  assign p1_smul_57326_TrailingBits___89_comb = 8'h00;
  assign p1_shifted__90_comb = {~p1_clipped__43_comb[7], p1_clipped__43_comb[6:0], p1_smul_57326_TrailingBits___218_comb};
  assign p1_smul_57326_TrailingBits___90_comb = 8'h00;
  assign p1_shifted__91_comb = {~p1_clipped__59_comb[7], p1_clipped__59_comb[6:0], p1_smul_57326_TrailingBits___219_comb};
  assign p1_smul_57326_TrailingBits___91_comb = 8'h00;
  assign p1_shifted__92_comb = {~p1_clipped__75_comb[7], p1_clipped__75_comb[6:0], p1_smul_57326_TrailingBits___220_comb};
  assign p1_smul_57326_TrailingBits___92_comb = 8'h00;
  assign p1_shifted__93_comb = {~p1_clipped__91_comb[7], p1_clipped__91_comb[6:0], p1_smul_57326_TrailingBits___221_comb};
  assign p1_smul_57326_TrailingBits___93_comb = 8'h00;
  assign p1_shifted__94_comb = {~p1_clipped__107_comb[7], p1_clipped__107_comb[6:0], p1_smul_57326_TrailingBits___222_comb};
  assign p1_smul_57326_TrailingBits___94_comb = 8'h00;
  assign p1_shifted__95_comb = {~p1_clipped__123_comb[7], p1_clipped__123_comb[6:0], p1_smul_57326_TrailingBits___223_comb};
  assign p1_smul_57326_TrailingBits___95_comb = 8'h00;
  assign p1_shifted__96_comb = {~p1_clipped__12_comb[7], p1_clipped__12_comb[6:0], p1_smul_57326_TrailingBits___224_comb};
  assign p1_smul_57326_TrailingBits___96_comb = 8'h00;
  assign p1_shifted__97_comb = {~p1_clipped__28_comb[7], p1_clipped__28_comb[6:0], p1_smul_57326_TrailingBits___225_comb};
  assign p1_smul_57326_TrailingBits___97_comb = 8'h00;
  assign p1_shifted__98_comb = {~p1_clipped__44_comb[7], p1_clipped__44_comb[6:0], p1_smul_57326_TrailingBits___226_comb};
  assign p1_smul_57326_TrailingBits___98_comb = 8'h00;
  assign p1_shifted__99_comb = {~p1_clipped__60_comb[7], p1_clipped__60_comb[6:0], p1_smul_57326_TrailingBits___227_comb};
  assign p1_smul_57326_TrailingBits___99_comb = 8'h00;
  assign p1_shifted__100_comb = {~p1_clipped__76_comb[7], p1_clipped__76_comb[6:0], p1_smul_57326_TrailingBits___228_comb};
  assign p1_smul_57326_TrailingBits___100_comb = 8'h00;
  assign p1_shifted__101_comb = {~p1_clipped__92_comb[7], p1_clipped__92_comb[6:0], p1_smul_57326_TrailingBits___229_comb};
  assign p1_smul_57326_TrailingBits___101_comb = 8'h00;
  assign p1_shifted__102_comb = {~p1_clipped__108_comb[7], p1_clipped__108_comb[6:0], p1_smul_57326_TrailingBits___230_comb};
  assign p1_smul_57326_TrailingBits___102_comb = 8'h00;
  assign p1_shifted__103_comb = {~p1_clipped__124_comb[7], p1_clipped__124_comb[6:0], p1_smul_57326_TrailingBits___231_comb};
  assign p1_smul_57326_TrailingBits___103_comb = 8'h00;
  assign p1_shifted__104_comb = {~p1_clipped__13_comb[7], p1_clipped__13_comb[6:0], p1_smul_57326_TrailingBits___232_comb};
  assign p1_smul_57326_TrailingBits___104_comb = 8'h00;
  assign p1_shifted__105_comb = {~p1_clipped__29_comb[7], p1_clipped__29_comb[6:0], p1_smul_57326_TrailingBits___233_comb};
  assign p1_smul_57326_TrailingBits___105_comb = 8'h00;
  assign p1_shifted__106_comb = {~p1_clipped__45_comb[7], p1_clipped__45_comb[6:0], p1_smul_57326_TrailingBits___234_comb};
  assign p1_smul_57326_TrailingBits___106_comb = 8'h00;
  assign p1_shifted__107_comb = {~p1_clipped__61_comb[7], p1_clipped__61_comb[6:0], p1_smul_57326_TrailingBits___235_comb};
  assign p1_smul_57326_TrailingBits___107_comb = 8'h00;
  assign p1_shifted__108_comb = {~p1_clipped__77_comb[7], p1_clipped__77_comb[6:0], p1_smul_57326_TrailingBits___236_comb};
  assign p1_smul_57326_TrailingBits___108_comb = 8'h00;
  assign p1_shifted__109_comb = {~p1_clipped__93_comb[7], p1_clipped__93_comb[6:0], p1_smul_57326_TrailingBits___237_comb};
  assign p1_smul_57326_TrailingBits___109_comb = 8'h00;
  assign p1_shifted__110_comb = {~p1_clipped__109_comb[7], p1_clipped__109_comb[6:0], p1_smul_57326_TrailingBits___238_comb};
  assign p1_smul_57326_TrailingBits___110_comb = 8'h00;
  assign p1_shifted__111_comb = {~p1_clipped__125_comb[7], p1_clipped__125_comb[6:0], p1_smul_57326_TrailingBits___239_comb};
  assign p1_smul_57326_TrailingBits___111_comb = 8'h00;
  assign p1_shifted__112_comb = {~p1_clipped__14_comb[7], p1_clipped__14_comb[6:0], p1_smul_57326_TrailingBits___240_comb};
  assign p1_smul_57326_TrailingBits___112_comb = 8'h00;
  assign p1_shifted__113_comb = {~p1_clipped__30_comb[7], p1_clipped__30_comb[6:0], p1_smul_57326_TrailingBits___241_comb};
  assign p1_smul_57326_TrailingBits___113_comb = 8'h00;
  assign p1_shifted__114_comb = {~p1_clipped__46_comb[7], p1_clipped__46_comb[6:0], p1_smul_57326_TrailingBits___242_comb};
  assign p1_smul_57326_TrailingBits___114_comb = 8'h00;
  assign p1_shifted__115_comb = {~p1_clipped__62_comb[7], p1_clipped__62_comb[6:0], p1_smul_57326_TrailingBits___243_comb};
  assign p1_smul_57326_TrailingBits___115_comb = 8'h00;
  assign p1_shifted__116_comb = {~p1_clipped__78_comb[7], p1_clipped__78_comb[6:0], p1_smul_57326_TrailingBits___244_comb};
  assign p1_smul_57326_TrailingBits___116_comb = 8'h00;
  assign p1_shifted__117_comb = {~p1_clipped__94_comb[7], p1_clipped__94_comb[6:0], p1_smul_57326_TrailingBits___245_comb};
  assign p1_smul_57326_TrailingBits___117_comb = 8'h00;
  assign p1_shifted__118_comb = {~p1_clipped__110_comb[7], p1_clipped__110_comb[6:0], p1_smul_57326_TrailingBits___246_comb};
  assign p1_smul_57326_TrailingBits___118_comb = 8'h00;
  assign p1_shifted__119_comb = {~p1_clipped__126_comb[7], p1_clipped__126_comb[6:0], p1_smul_57326_TrailingBits___247_comb};
  assign p1_smul_57326_TrailingBits___119_comb = 8'h00;
  assign p1_shifted__120_comb = {~p1_clipped__15_comb[7], p1_clipped__15_comb[6:0], p1_smul_57326_TrailingBits___248_comb};
  assign p1_smul_57326_TrailingBits___120_comb = 8'h00;
  assign p1_shifted__121_comb = {~p1_clipped__31_comb[7], p1_clipped__31_comb[6:0], p1_smul_57326_TrailingBits___249_comb};
  assign p1_smul_57326_TrailingBits___121_comb = 8'h00;
  assign p1_shifted__122_comb = {~p1_clipped__47_comb[7], p1_clipped__47_comb[6:0], p1_smul_57326_TrailingBits___250_comb};
  assign p1_smul_57326_TrailingBits___122_comb = 8'h00;
  assign p1_shifted__123_comb = {~p1_clipped__63_comb[7], p1_clipped__63_comb[6:0], p1_smul_57326_TrailingBits___251_comb};
  assign p1_smul_57326_TrailingBits___123_comb = 8'h00;
  assign p1_shifted__124_comb = {~p1_clipped__79_comb[7], p1_clipped__79_comb[6:0], p1_smul_57326_TrailingBits___252_comb};
  assign p1_smul_57326_TrailingBits___124_comb = 8'h00;
  assign p1_shifted__125_comb = {~p1_clipped__95_comb[7], p1_clipped__95_comb[6:0], p1_smul_57326_TrailingBits___253_comb};
  assign p1_smul_57326_TrailingBits___125_comb = 8'h00;
  assign p1_shifted__126_comb = {~p1_clipped__111_comb[7], p1_clipped__111_comb[6:0], p1_smul_57326_TrailingBits___254_comb};
  assign p1_smul_57326_TrailingBits___126_comb = 8'h00;
  assign p1_shifted__127_comb = {~p1_clipped__127_comb[7], p1_clipped__127_comb[6:0], p1_smul_57326_TrailingBits___255_comb};
  assign p1_smul_57326_TrailingBits___127_comb = 8'h00;
  assign p1_or_146687_comb = p1_prod__519_comb | 32'h0000_0080;
  assign p1_prod__523_comb = {{9{p1_concat_146045_comb[22]}}, p1_concat_146045_comb};
  assign p1_prod__528_comb = {{9{p1_concat_146046_comb[22]}}, p1_concat_146046_comb};
  assign p1_or_146694_comb = p1_prod__534_comb | 32'h0000_0080;
  assign p1_or_146701_comb = p1_prod__583_comb | 32'h0000_0080;
  assign p1_prod__587_comb = {{9{p1_concat_146051_comb[22]}}, p1_concat_146051_comb};
  assign p1_prod__592_comb = {{9{p1_concat_146052_comb[22]}}, p1_concat_146052_comb};
  assign p1_or_146708_comb = p1_prod__598_comb | 32'h0000_0080;
  assign p1_or_146715_comb = p1_prod__647_comb | 32'h0000_0080;
  assign p1_prod__651_comb = {{9{p1_concat_146057_comb[22]}}, p1_concat_146057_comb};
  assign p1_prod__656_comb = {{9{p1_concat_146058_comb[22]}}, p1_concat_146058_comb};
  assign p1_or_146722_comb = p1_prod__662_comb | 32'h0000_0080;
  assign p1_or_146729_comb = p1_prod__711_comb | 32'h0000_0080;
  assign p1_prod__715_comb = {{9{p1_concat_146063_comb[22]}}, p1_concat_146063_comb};
  assign p1_prod__720_comb = {{9{p1_concat_146064_comb[22]}}, p1_concat_146064_comb};
  assign p1_or_146736_comb = p1_prod__726_comb | 32'h0000_0080;
  assign p1_or_146743_comb = p1_prod__775_comb | 32'h0000_0080;
  assign p1_prod__779_comb = {{9{p1_concat_146069_comb[22]}}, p1_concat_146069_comb};
  assign p1_prod__784_comb = {{9{p1_concat_146070_comb[22]}}, p1_concat_146070_comb};
  assign p1_or_146750_comb = p1_prod__790_comb | 32'h0000_0080;
  assign p1_or_146757_comb = p1_prod__839_comb | 32'h0000_0080;
  assign p1_prod__843_comb = {{9{p1_concat_146075_comb[22]}}, p1_concat_146075_comb};
  assign p1_prod__848_comb = {{9{p1_concat_146076_comb[22]}}, p1_concat_146076_comb};
  assign p1_or_146764_comb = p1_prod__854_comb | 32'h0000_0080;
  assign p1_or_146771_comb = p1_prod__903_comb | 32'h0000_0080;
  assign p1_prod__907_comb = {{9{p1_concat_146081_comb[22]}}, p1_concat_146081_comb};
  assign p1_prod__912_comb = {{9{p1_concat_146082_comb[22]}}, p1_concat_146082_comb};
  assign p1_or_146778_comb = p1_prod__918_comb | 32'h0000_0080;
  assign p1_or_146785_comb = p1_prod__967_comb | 32'h0000_0080;
  assign p1_prod__971_comb = {{9{p1_concat_146087_comb[22]}}, p1_concat_146087_comb};
  assign p1_prod__976_comb = {{9{p1_concat_146088_comb[22]}}, p1_concat_146088_comb};
  assign p1_or_146792_comb = p1_prod__982_comb | 32'h0000_0080;
  assign p1_or_146797_comb = p1_prod__517_comb | 32'h0000_0080;
  assign p1_or_146804_comb = p1_prod__529_comb | 32'h0000_0080;
  assign p1_or_146807_comb = p1_prod__535_comb | 32'h0000_0080;
  assign p1_or_146814_comb = p1_prod__555_comb | 32'h0000_0080;
  assign p1_or_146817_comb = p1_prod__581_comb | 32'h0000_0080;
  assign p1_or_146824_comb = p1_prod__593_comb | 32'h0000_0080;
  assign p1_or_146827_comb = p1_prod__599_comb | 32'h0000_0080;
  assign p1_or_146834_comb = p1_prod__619_comb | 32'h0000_0080;
  assign p1_or_146837_comb = p1_prod__645_comb | 32'h0000_0080;
  assign p1_or_146844_comb = p1_prod__657_comb | 32'h0000_0080;
  assign p1_or_146847_comb = p1_prod__663_comb | 32'h0000_0080;
  assign p1_or_146854_comb = p1_prod__683_comb | 32'h0000_0080;
  assign p1_or_146857_comb = p1_prod__709_comb | 32'h0000_0080;
  assign p1_or_146864_comb = p1_prod__721_comb | 32'h0000_0080;
  assign p1_or_146867_comb = p1_prod__727_comb | 32'h0000_0080;
  assign p1_or_146874_comb = p1_prod__747_comb | 32'h0000_0080;
  assign p1_or_146877_comb = p1_prod__773_comb | 32'h0000_0080;
  assign p1_or_146884_comb = p1_prod__785_comb | 32'h0000_0080;
  assign p1_or_146887_comb = p1_prod__791_comb | 32'h0000_0080;
  assign p1_or_146894_comb = p1_prod__811_comb | 32'h0000_0080;
  assign p1_or_146897_comb = p1_prod__837_comb | 32'h0000_0080;
  assign p1_or_146904_comb = p1_prod__849_comb | 32'h0000_0080;
  assign p1_or_146907_comb = p1_prod__855_comb | 32'h0000_0080;
  assign p1_or_146914_comb = p1_prod__875_comb | 32'h0000_0080;
  assign p1_or_146917_comb = p1_prod__901_comb | 32'h0000_0080;
  assign p1_or_146924_comb = p1_prod__913_comb | 32'h0000_0080;
  assign p1_or_146927_comb = p1_prod__919_comb | 32'h0000_0080;
  assign p1_or_146934_comb = p1_prod__939_comb | 32'h0000_0080;
  assign p1_or_146937_comb = p1_prod__965_comb | 32'h0000_0080;
  assign p1_or_146944_comb = p1_prod__977_comb | 32'h0000_0080;
  assign p1_or_146947_comb = p1_prod__983_comb | 32'h0000_0080;
  assign p1_or_146954_comb = p1_prod__1003_comb | 32'h0000_0080;
  assign p1_prod__525_comb = {{9{p1_concat_146187_comb[22]}}, p1_concat_146187_comb};
  assign p1_or_146961_comb = p1_prod__536_comb | 32'h0000_0080;
  assign p1_or_146964_comb = p1_prod__543_comb | 32'h0000_0080;
  assign p1_prod__556_comb = {{9{p1_concat_146192_comb[22]}}, p1_concat_146192_comb};
  assign p1_prod__589_comb = {{9{p1_concat_146193_comb[22]}}, p1_concat_146193_comb};
  assign p1_or_146975_comb = p1_prod__600_comb | 32'h0000_0080;
  assign p1_or_146978_comb = p1_prod__607_comb | 32'h0000_0080;
  assign p1_prod__620_comb = {{9{p1_concat_146198_comb[22]}}, p1_concat_146198_comb};
  assign p1_prod__653_comb = {{9{p1_concat_146199_comb[22]}}, p1_concat_146199_comb};
  assign p1_or_146989_comb = p1_prod__664_comb | 32'h0000_0080;
  assign p1_or_146992_comb = p1_prod__671_comb | 32'h0000_0080;
  assign p1_prod__684_comb = {{9{p1_concat_146204_comb[22]}}, p1_concat_146204_comb};
  assign p1_prod__717_comb = {{9{p1_concat_146205_comb[22]}}, p1_concat_146205_comb};
  assign p1_or_147003_comb = p1_prod__728_comb | 32'h0000_0080;
  assign p1_or_147006_comb = p1_prod__735_comb | 32'h0000_0080;
  assign p1_prod__748_comb = {{9{p1_concat_146210_comb[22]}}, p1_concat_146210_comb};
  assign p1_prod__781_comb = {{9{p1_concat_146211_comb[22]}}, p1_concat_146211_comb};
  assign p1_or_147017_comb = p1_prod__792_comb | 32'h0000_0080;
  assign p1_or_147020_comb = p1_prod__799_comb | 32'h0000_0080;
  assign p1_prod__812_comb = {{9{p1_concat_146216_comb[22]}}, p1_concat_146216_comb};
  assign p1_prod__845_comb = {{9{p1_concat_146217_comb[22]}}, p1_concat_146217_comb};
  assign p1_or_147031_comb = p1_prod__856_comb | 32'h0000_0080;
  assign p1_or_147034_comb = p1_prod__863_comb | 32'h0000_0080;
  assign p1_prod__876_comb = {{9{p1_concat_146222_comb[22]}}, p1_concat_146222_comb};
  assign p1_prod__909_comb = {{9{p1_concat_146223_comb[22]}}, p1_concat_146223_comb};
  assign p1_or_147045_comb = p1_prod__920_comb | 32'h0000_0080;
  assign p1_or_147048_comb = p1_prod__927_comb | 32'h0000_0080;
  assign p1_prod__940_comb = {{9{p1_concat_146228_comb[22]}}, p1_concat_146228_comb};
  assign p1_prod__973_comb = {{9{p1_concat_146229_comb[22]}}, p1_concat_146229_comb};
  assign p1_or_147059_comb = p1_prod__984_comb | 32'h0000_0080;
  assign p1_or_147062_comb = p1_prod__991_comb | 32'h0000_0080;
  assign p1_prod__1004_comb = {{9{p1_concat_146234_comb[22]}}, p1_concat_146234_comb};
  assign p1_or_147133_comb = p1_prod__532_comb | 32'h0000_0080;
  assign p1_prod__545_comb = {{9{p1_concat_146237_comb[22]}}, p1_concat_146237_comb};
  assign p1_prod__563_comb = {{9{p1_concat_146238_comb[22]}}, p1_concat_146238_comb};
  assign p1_or_147144_comb = p1_prod__570_comb | 32'h0000_0080;
  assign p1_or_147147_comb = p1_prod__596_comb | 32'h0000_0080;
  assign p1_prod__609_comb = {{9{p1_concat_146243_comb[22]}}, p1_concat_146243_comb};
  assign p1_prod__627_comb = {{9{p1_concat_146244_comb[22]}}, p1_concat_146244_comb};
  assign p1_or_147158_comb = p1_prod__634_comb | 32'h0000_0080;
  assign p1_or_147161_comb = p1_prod__660_comb | 32'h0000_0080;
  assign p1_prod__673_comb = {{9{p1_concat_146249_comb[22]}}, p1_concat_146249_comb};
  assign p1_prod__691_comb = {{9{p1_concat_146250_comb[22]}}, p1_concat_146250_comb};
  assign p1_or_147172_comb = p1_prod__698_comb | 32'h0000_0080;
  assign p1_or_147175_comb = p1_prod__724_comb | 32'h0000_0080;
  assign p1_prod__737_comb = {{9{p1_concat_146255_comb[22]}}, p1_concat_146255_comb};
  assign p1_prod__755_comb = {{9{p1_concat_146256_comb[22]}}, p1_concat_146256_comb};
  assign p1_or_147186_comb = p1_prod__762_comb | 32'h0000_0080;
  assign p1_or_147189_comb = p1_prod__788_comb | 32'h0000_0080;
  assign p1_prod__801_comb = {{9{p1_concat_146261_comb[22]}}, p1_concat_146261_comb};
  assign p1_prod__819_comb = {{9{p1_concat_146262_comb[22]}}, p1_concat_146262_comb};
  assign p1_or_147200_comb = p1_prod__826_comb | 32'h0000_0080;
  assign p1_or_147203_comb = p1_prod__852_comb | 32'h0000_0080;
  assign p1_prod__865_comb = {{9{p1_concat_146267_comb[22]}}, p1_concat_146267_comb};
  assign p1_prod__883_comb = {{9{p1_concat_146268_comb[22]}}, p1_concat_146268_comb};
  assign p1_or_147214_comb = p1_prod__890_comb | 32'h0000_0080;
  assign p1_or_147217_comb = p1_prod__916_comb | 32'h0000_0080;
  assign p1_prod__929_comb = {{9{p1_concat_146273_comb[22]}}, p1_concat_146273_comb};
  assign p1_prod__947_comb = {{9{p1_concat_146274_comb[22]}}, p1_concat_146274_comb};
  assign p1_or_147228_comb = p1_prod__954_comb | 32'h0000_0080;
  assign p1_or_147231_comb = p1_prod__980_comb | 32'h0000_0080;
  assign p1_prod__993_comb = {{9{p1_concat_146279_comb[22]}}, p1_concat_146279_comb};
  assign p1_prod__1011_comb = {{9{p1_concat_146280_comb[22]}}, p1_concat_146280_comb};
  assign p1_or_147242_comb = p1_prod__1018_comb | 32'h0000_0080;
  assign p1_or_147247_comb = p1_prod__546_comb | 32'h0000_0080;
  assign p1_or_147252_comb = p1_prod__559_comb | 32'h0000_0080;
  assign p1_or_147255_comb = p1_prod__564_comb | 32'h0000_0080;
  assign p1_or_147260_comb = p1_prod__571_comb | 32'h0000_0080;
  assign p1_or_147267_comb = p1_prod__610_comb | 32'h0000_0080;
  assign p1_or_147272_comb = p1_prod__623_comb | 32'h0000_0080;
  assign p1_or_147275_comb = p1_prod__628_comb | 32'h0000_0080;
  assign p1_or_147280_comb = p1_prod__635_comb | 32'h0000_0080;
  assign p1_or_147287_comb = p1_prod__674_comb | 32'h0000_0080;
  assign p1_or_147292_comb = p1_prod__687_comb | 32'h0000_0080;
  assign p1_or_147295_comb = p1_prod__692_comb | 32'h0000_0080;
  assign p1_or_147300_comb = p1_prod__699_comb | 32'h0000_0080;
  assign p1_or_147307_comb = p1_prod__738_comb | 32'h0000_0080;
  assign p1_or_147312_comb = p1_prod__751_comb | 32'h0000_0080;
  assign p1_or_147315_comb = p1_prod__756_comb | 32'h0000_0080;
  assign p1_or_147320_comb = p1_prod__763_comb | 32'h0000_0080;
  assign p1_or_147327_comb = p1_prod__802_comb | 32'h0000_0080;
  assign p1_or_147332_comb = p1_prod__815_comb | 32'h0000_0080;
  assign p1_or_147335_comb = p1_prod__820_comb | 32'h0000_0080;
  assign p1_or_147340_comb = p1_prod__827_comb | 32'h0000_0080;
  assign p1_or_147347_comb = p1_prod__866_comb | 32'h0000_0080;
  assign p1_or_147352_comb = p1_prod__879_comb | 32'h0000_0080;
  assign p1_or_147355_comb = p1_prod__884_comb | 32'h0000_0080;
  assign p1_or_147360_comb = p1_prod__891_comb | 32'h0000_0080;
  assign p1_or_147367_comb = p1_prod__930_comb | 32'h0000_0080;
  assign p1_or_147372_comb = p1_prod__943_comb | 32'h0000_0080;
  assign p1_or_147375_comb = p1_prod__948_comb | 32'h0000_0080;
  assign p1_or_147380_comb = p1_prod__955_comb | 32'h0000_0080;
  assign p1_or_147387_comb = p1_prod__994_comb | 32'h0000_0080;
  assign p1_or_147392_comb = p1_prod__1007_comb | 32'h0000_0080;
  assign p1_or_147395_comb = p1_prod__1012_comb | 32'h0000_0080;
  assign p1_or_147400_comb = p1_prod__1019_comb | 32'h0000_0080;
  assign p1_prod__547_comb = {{9{p1_concat_146379_comb[22]}}, p1_concat_146379_comb};
  assign p1_or_147407_comb = p1_prod__554_comb | 32'h0000_0080;
  assign p1_or_147414_comb = p1_prod__574_comb | 32'h0000_0080;
  assign p1_prod__575_comb = {{9{p1_concat_146384_comb[22]}}, p1_concat_146384_comb};
  assign p1_prod__611_comb = {{9{p1_concat_146385_comb[22]}}, p1_concat_146385_comb};
  assign p1_or_147421_comb = p1_prod__618_comb | 32'h0000_0080;
  assign p1_or_147428_comb = p1_prod__638_comb | 32'h0000_0080;
  assign p1_prod__639_comb = {{9{p1_concat_146390_comb[22]}}, p1_concat_146390_comb};
  assign p1_prod__675_comb = {{9{p1_concat_146391_comb[22]}}, p1_concat_146391_comb};
  assign p1_or_147435_comb = p1_prod__682_comb | 32'h0000_0080;
  assign p1_or_147442_comb = p1_prod__702_comb | 32'h0000_0080;
  assign p1_prod__703_comb = {{9{p1_concat_146396_comb[22]}}, p1_concat_146396_comb};
  assign p1_prod__739_comb = {{9{p1_concat_146397_comb[22]}}, p1_concat_146397_comb};
  assign p1_or_147449_comb = p1_prod__746_comb | 32'h0000_0080;
  assign p1_or_147456_comb = p1_prod__766_comb | 32'h0000_0080;
  assign p1_prod__767_comb = {{9{p1_concat_146402_comb[22]}}, p1_concat_146402_comb};
  assign p1_prod__803_comb = {{9{p1_concat_146403_comb[22]}}, p1_concat_146403_comb};
  assign p1_or_147463_comb = p1_prod__810_comb | 32'h0000_0080;
  assign p1_or_147470_comb = p1_prod__830_comb | 32'h0000_0080;
  assign p1_prod__831_comb = {{9{p1_concat_146408_comb[22]}}, p1_concat_146408_comb};
  assign p1_prod__867_comb = {{9{p1_concat_146409_comb[22]}}, p1_concat_146409_comb};
  assign p1_or_147477_comb = p1_prod__874_comb | 32'h0000_0080;
  assign p1_or_147484_comb = p1_prod__894_comb | 32'h0000_0080;
  assign p1_prod__895_comb = {{9{p1_concat_146414_comb[22]}}, p1_concat_146414_comb};
  assign p1_prod__931_comb = {{9{p1_concat_146415_comb[22]}}, p1_concat_146415_comb};
  assign p1_or_147491_comb = p1_prod__938_comb | 32'h0000_0080;
  assign p1_or_147498_comb = p1_prod__958_comb | 32'h0000_0080;
  assign p1_prod__959_comb = {{9{p1_concat_146420_comb[22]}}, p1_concat_146420_comb};
  assign p1_prod__995_comb = {{9{p1_concat_146421_comb[22]}}, p1_concat_146421_comb};
  assign p1_or_147505_comb = p1_prod__1002_comb | 32'h0000_0080;
  assign p1_or_147512_comb = p1_prod__1022_comb | 32'h0000_0080;
  assign p1_prod__1023_comb = {{9{p1_concat_146426_comb[22]}}, p1_concat_146426_comb};
  assign p1_smul_58222_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__64_squeezed_comb, 9'h0fb);
  assign p1_smul_58224_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__65_squeezed_comb, 9'h0d5);
  assign p1_or_147714_comb = p1_prod__523_comb | 32'h0000_0080;
  assign p1_or_147715_comb = p1_prod__528_comb | 32'h0000_0080;
  assign p1_smul_58234_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__70_squeezed_comb, 9'h12b);
  assign p1_smul_58236_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__71_squeezed_comb, 9'h105);
  assign p1_smul_58238_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__72_squeezed_comb, 9'h0fb);
  assign p1_smul_58240_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__73_squeezed_comb, 9'h0d5);
  assign p1_or_147730_comb = p1_prod__587_comb | 32'h0000_0080;
  assign p1_or_147731_comb = p1_prod__592_comb | 32'h0000_0080;
  assign p1_smul_58250_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__78_squeezed_comb, 9'h12b);
  assign p1_smul_58252_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__79_squeezed_comb, 9'h105);
  assign p1_smul_58254_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__80_squeezed_comb, 9'h0fb);
  assign p1_smul_58256_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__81_squeezed_comb, 9'h0d5);
  assign p1_or_147746_comb = p1_prod__651_comb | 32'h0000_0080;
  assign p1_or_147747_comb = p1_prod__656_comb | 32'h0000_0080;
  assign p1_smul_58266_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__86_squeezed_comb, 9'h12b);
  assign p1_smul_58268_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__87_squeezed_comb, 9'h105);
  assign p1_smul_58270_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__88_squeezed_comb, 9'h0fb);
  assign p1_smul_58272_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__89_squeezed_comb, 9'h0d5);
  assign p1_or_147762_comb = p1_prod__715_comb | 32'h0000_0080;
  assign p1_or_147763_comb = p1_prod__720_comb | 32'h0000_0080;
  assign p1_smul_58282_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__94_squeezed_comb, 9'h12b);
  assign p1_smul_58284_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__95_squeezed_comb, 9'h105);
  assign p1_smul_58286_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__96_squeezed_comb, 9'h0fb);
  assign p1_smul_58288_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__97_squeezed_comb, 9'h0d5);
  assign p1_or_147778_comb = p1_prod__779_comb | 32'h0000_0080;
  assign p1_or_147779_comb = p1_prod__784_comb | 32'h0000_0080;
  assign p1_smul_58298_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__102_squeezed_comb, 9'h12b);
  assign p1_smul_58300_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__103_squeezed_comb, 9'h105);
  assign p1_smul_58302_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__104_squeezed_comb, 9'h0fb);
  assign p1_smul_58304_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__105_squeezed_comb, 9'h0d5);
  assign p1_or_147794_comb = p1_prod__843_comb | 32'h0000_0080;
  assign p1_or_147795_comb = p1_prod__848_comb | 32'h0000_0080;
  assign p1_smul_58314_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__110_squeezed_comb, 9'h12b);
  assign p1_smul_58316_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__111_squeezed_comb, 9'h105);
  assign p1_smul_58318_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__112_squeezed_comb, 9'h0fb);
  assign p1_smul_58320_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__113_squeezed_comb, 9'h0d5);
  assign p1_or_147810_comb = p1_prod__907_comb | 32'h0000_0080;
  assign p1_or_147811_comb = p1_prod__912_comb | 32'h0000_0080;
  assign p1_smul_58330_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__118_squeezed_comb, 9'h12b);
  assign p1_smul_58332_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__119_squeezed_comb, 9'h105);
  assign p1_smul_58334_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__120_squeezed_comb, 9'h0fb);
  assign p1_smul_58336_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__121_squeezed_comb, 9'h0d5);
  assign p1_or_147826_comb = p1_prod__971_comb | 32'h0000_0080;
  assign p1_or_147827_comb = p1_prod__976_comb | 32'h0000_0080;
  assign p1_smul_58346_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__126_squeezed_comb, 9'h12b);
  assign p1_smul_58348_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__127_squeezed_comb, 9'h105);
  assign p1_smul_58478_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__64_squeezed_comb, 9'h0d5);
  assign p1_or_147997_comb = p1_prod__525_comb | 32'h0000_0080;
  assign p1_smul_58482_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__66_squeezed_comb, 9'h105);
  assign p1_smul_58488_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__69_squeezed_comb, 9'h0fb);
  assign p1_or_148008_comb = p1_prod__556_comb | 32'h0000_0080;
  assign p1_smul_58492_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__71_squeezed_comb, 9'h12b);
  assign p1_smul_58494_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__72_squeezed_comb, 9'h0d5);
  assign p1_or_148013_comb = p1_prod__589_comb | 32'h0000_0080;
  assign p1_smul_58498_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__74_squeezed_comb, 9'h105);
  assign p1_smul_58504_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__77_squeezed_comb, 9'h0fb);
  assign p1_or_148024_comb = p1_prod__620_comb | 32'h0000_0080;
  assign p1_smul_58508_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__79_squeezed_comb, 9'h12b);
  assign p1_smul_58510_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__80_squeezed_comb, 9'h0d5);
  assign p1_or_148029_comb = p1_prod__653_comb | 32'h0000_0080;
  assign p1_smul_58514_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__82_squeezed_comb, 9'h105);
  assign p1_smul_58520_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__85_squeezed_comb, 9'h0fb);
  assign p1_or_148040_comb = p1_prod__684_comb | 32'h0000_0080;
  assign p1_smul_58524_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__87_squeezed_comb, 9'h12b);
  assign p1_smul_58526_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__88_squeezed_comb, 9'h0d5);
  assign p1_or_148045_comb = p1_prod__717_comb | 32'h0000_0080;
  assign p1_smul_58530_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__90_squeezed_comb, 9'h105);
  assign p1_smul_58536_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__93_squeezed_comb, 9'h0fb);
  assign p1_or_148056_comb = p1_prod__748_comb | 32'h0000_0080;
  assign p1_smul_58540_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__95_squeezed_comb, 9'h12b);
  assign p1_smul_58542_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__96_squeezed_comb, 9'h0d5);
  assign p1_or_148061_comb = p1_prod__781_comb | 32'h0000_0080;
  assign p1_smul_58546_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__98_squeezed_comb, 9'h105);
  assign p1_smul_58552_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__101_squeezed_comb, 9'h0fb);
  assign p1_or_148072_comb = p1_prod__812_comb | 32'h0000_0080;
  assign p1_smul_58556_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__103_squeezed_comb, 9'h12b);
  assign p1_smul_58558_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__104_squeezed_comb, 9'h0d5);
  assign p1_or_148077_comb = p1_prod__845_comb | 32'h0000_0080;
  assign p1_smul_58562_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__106_squeezed_comb, 9'h105);
  assign p1_smul_58568_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__109_squeezed_comb, 9'h0fb);
  assign p1_or_148088_comb = p1_prod__876_comb | 32'h0000_0080;
  assign p1_smul_58572_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__111_squeezed_comb, 9'h12b);
  assign p1_smul_58574_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__112_squeezed_comb, 9'h0d5);
  assign p1_or_148093_comb = p1_prod__909_comb | 32'h0000_0080;
  assign p1_smul_58578_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__114_squeezed_comb, 9'h105);
  assign p1_smul_58584_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__117_squeezed_comb, 9'h0fb);
  assign p1_or_148104_comb = p1_prod__940_comb | 32'h0000_0080;
  assign p1_smul_58588_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__119_squeezed_comb, 9'h12b);
  assign p1_smul_58590_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__120_squeezed_comb, 9'h0d5);
  assign p1_or_148109_comb = p1_prod__973_comb | 32'h0000_0080;
  assign p1_smul_58594_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__122_squeezed_comb, 9'h105);
  assign p1_smul_58600_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__125_squeezed_comb, 9'h0fb);
  assign p1_or_148120_comb = p1_prod__1004_comb | 32'h0000_0080;
  assign p1_smul_58604_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__127_squeezed_comb, 9'h12b);
  assign p1_smul_58606_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__64_squeezed_comb, 9'h0b5);
  assign p1_smul_58608_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__65_squeezed_comb, 9'h14b);
  assign p1_smul_58610_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__66_squeezed_comb, 9'h14b);
  assign p1_smul_58612_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__67_squeezed_comb, 9'h0b5);
  assign p1_smul_58614_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__68_squeezed_comb, 9'h0b5);
  assign p1_smul_58616_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__69_squeezed_comb, 9'h14b);
  assign p1_smul_58618_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__70_squeezed_comb, 9'h14b);
  assign p1_smul_58620_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__71_squeezed_comb, 9'h0b5);
  assign p1_smul_58622_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__72_squeezed_comb, 9'h0b5);
  assign p1_smul_58624_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__73_squeezed_comb, 9'h14b);
  assign p1_smul_58626_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__74_squeezed_comb, 9'h14b);
  assign p1_smul_58628_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__75_squeezed_comb, 9'h0b5);
  assign p1_smul_58630_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__76_squeezed_comb, 9'h0b5);
  assign p1_smul_58632_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__77_squeezed_comb, 9'h14b);
  assign p1_smul_58634_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__78_squeezed_comb, 9'h14b);
  assign p1_smul_58636_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__79_squeezed_comb, 9'h0b5);
  assign p1_smul_58638_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__80_squeezed_comb, 9'h0b5);
  assign p1_smul_58640_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__81_squeezed_comb, 9'h14b);
  assign p1_smul_58642_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__82_squeezed_comb, 9'h14b);
  assign p1_smul_58644_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__83_squeezed_comb, 9'h0b5);
  assign p1_smul_58646_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__84_squeezed_comb, 9'h0b5);
  assign p1_smul_58648_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__85_squeezed_comb, 9'h14b);
  assign p1_smul_58650_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__86_squeezed_comb, 9'h14b);
  assign p1_smul_58652_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__87_squeezed_comb, 9'h0b5);
  assign p1_smul_58654_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__88_squeezed_comb, 9'h0b5);
  assign p1_smul_58656_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__89_squeezed_comb, 9'h14b);
  assign p1_smul_58658_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__90_squeezed_comb, 9'h14b);
  assign p1_smul_58660_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__91_squeezed_comb, 9'h0b5);
  assign p1_smul_58662_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__92_squeezed_comb, 9'h0b5);
  assign p1_smul_58664_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__93_squeezed_comb, 9'h14b);
  assign p1_smul_58666_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__94_squeezed_comb, 9'h14b);
  assign p1_smul_58668_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__95_squeezed_comb, 9'h0b5);
  assign p1_smul_58670_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__96_squeezed_comb, 9'h0b5);
  assign p1_smul_58672_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__97_squeezed_comb, 9'h14b);
  assign p1_smul_58674_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__98_squeezed_comb, 9'h14b);
  assign p1_smul_58676_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__99_squeezed_comb, 9'h0b5);
  assign p1_smul_58678_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__100_squeezed_comb, 9'h0b5);
  assign p1_smul_58680_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__101_squeezed_comb, 9'h14b);
  assign p1_smul_58682_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__102_squeezed_comb, 9'h14b);
  assign p1_smul_58684_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__103_squeezed_comb, 9'h0b5);
  assign p1_smul_58686_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__104_squeezed_comb, 9'h0b5);
  assign p1_smul_58688_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__105_squeezed_comb, 9'h14b);
  assign p1_smul_58690_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__106_squeezed_comb, 9'h14b);
  assign p1_smul_58692_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__107_squeezed_comb, 9'h0b5);
  assign p1_smul_58694_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__108_squeezed_comb, 9'h0b5);
  assign p1_smul_58696_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__109_squeezed_comb, 9'h14b);
  assign p1_smul_58698_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__110_squeezed_comb, 9'h14b);
  assign p1_smul_58700_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__111_squeezed_comb, 9'h0b5);
  assign p1_smul_58702_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__112_squeezed_comb, 9'h0b5);
  assign p1_smul_58704_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__113_squeezed_comb, 9'h14b);
  assign p1_smul_58706_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__114_squeezed_comb, 9'h14b);
  assign p1_smul_58708_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__115_squeezed_comb, 9'h0b5);
  assign p1_smul_58710_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__116_squeezed_comb, 9'h0b5);
  assign p1_smul_58712_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__117_squeezed_comb, 9'h14b);
  assign p1_smul_58714_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__118_squeezed_comb, 9'h14b);
  assign p1_smul_58716_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__119_squeezed_comb, 9'h0b5);
  assign p1_smul_58718_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__120_squeezed_comb, 9'h0b5);
  assign p1_smul_58720_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__121_squeezed_comb, 9'h14b);
  assign p1_smul_58722_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__122_squeezed_comb, 9'h14b);
  assign p1_smul_58724_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__123_squeezed_comb, 9'h0b5);
  assign p1_smul_58726_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__124_squeezed_comb, 9'h0b5);
  assign p1_smul_58728_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__125_squeezed_comb, 9'h14b);
  assign p1_smul_58730_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__126_squeezed_comb, 9'h14b);
  assign p1_smul_58732_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__127_squeezed_comb, 9'h0b5);
  assign p1_smul_58736_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__65_squeezed_comb, 9'h105);
  assign p1_or_148256_comb = p1_prod__545_comb | 32'h0000_0080;
  assign p1_smul_58740_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__67_squeezed_comb, 9'h0d5);
  assign p1_smul_58742_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__68_squeezed_comb, 9'h0d5);
  assign p1_or_148261_comb = p1_prod__563_comb | 32'h0000_0080;
  assign p1_smul_58746_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__70_squeezed_comb, 9'h105);
  assign p1_smul_58752_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__73_squeezed_comb, 9'h105);
  assign p1_or_148272_comb = p1_prod__609_comb | 32'h0000_0080;
  assign p1_smul_58756_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__75_squeezed_comb, 9'h0d5);
  assign p1_smul_58758_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__76_squeezed_comb, 9'h0d5);
  assign p1_or_148277_comb = p1_prod__627_comb | 32'h0000_0080;
  assign p1_smul_58762_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__78_squeezed_comb, 9'h105);
  assign p1_smul_58768_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__81_squeezed_comb, 9'h105);
  assign p1_or_148288_comb = p1_prod__673_comb | 32'h0000_0080;
  assign p1_smul_58772_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__83_squeezed_comb, 9'h0d5);
  assign p1_smul_58774_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__84_squeezed_comb, 9'h0d5);
  assign p1_or_148293_comb = p1_prod__691_comb | 32'h0000_0080;
  assign p1_smul_58778_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__86_squeezed_comb, 9'h105);
  assign p1_smul_58784_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__89_squeezed_comb, 9'h105);
  assign p1_or_148304_comb = p1_prod__737_comb | 32'h0000_0080;
  assign p1_smul_58788_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__91_squeezed_comb, 9'h0d5);
  assign p1_smul_58790_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__92_squeezed_comb, 9'h0d5);
  assign p1_or_148309_comb = p1_prod__755_comb | 32'h0000_0080;
  assign p1_smul_58794_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__94_squeezed_comb, 9'h105);
  assign p1_smul_58800_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__97_squeezed_comb, 9'h105);
  assign p1_or_148320_comb = p1_prod__801_comb | 32'h0000_0080;
  assign p1_smul_58804_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__99_squeezed_comb, 9'h0d5);
  assign p1_smul_58806_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__100_squeezed_comb, 9'h0d5);
  assign p1_or_148325_comb = p1_prod__819_comb | 32'h0000_0080;
  assign p1_smul_58810_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__102_squeezed_comb, 9'h105);
  assign p1_smul_58816_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__105_squeezed_comb, 9'h105);
  assign p1_or_148336_comb = p1_prod__865_comb | 32'h0000_0080;
  assign p1_smul_58820_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__107_squeezed_comb, 9'h0d5);
  assign p1_smul_58822_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__108_squeezed_comb, 9'h0d5);
  assign p1_or_148341_comb = p1_prod__883_comb | 32'h0000_0080;
  assign p1_smul_58826_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__110_squeezed_comb, 9'h105);
  assign p1_smul_58832_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__113_squeezed_comb, 9'h105);
  assign p1_or_148352_comb = p1_prod__929_comb | 32'h0000_0080;
  assign p1_smul_58836_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__115_squeezed_comb, 9'h0d5);
  assign p1_smul_58838_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__116_squeezed_comb, 9'h0d5);
  assign p1_or_148357_comb = p1_prod__947_comb | 32'h0000_0080;
  assign p1_smul_58842_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__118_squeezed_comb, 9'h105);
  assign p1_smul_58848_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__121_squeezed_comb, 9'h105);
  assign p1_or_148368_comb = p1_prod__993_comb | 32'h0000_0080;
  assign p1_smul_58852_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__123_squeezed_comb, 9'h0d5);
  assign p1_smul_58854_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__124_squeezed_comb, 9'h0d5);
  assign p1_or_148373_comb = p1_prod__1011_comb | 32'h0000_0080;
  assign p1_smul_58858_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__126_squeezed_comb, 9'h105);
  assign p1_or_148539_comb = p1_prod__547_comb | 32'h0000_0080;
  assign p1_smul_58994_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__66_squeezed_comb, 9'h0d5);
  assign p1_smul_58996_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__67_squeezed_comb, 9'h105);
  assign p1_smul_58998_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__68_squeezed_comb, 9'h105);
  assign p1_smul_59000_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__69_squeezed_comb, 9'h0d5);
  assign p1_or_148554_comb = p1_prod__575_comb | 32'h0000_0080;
  assign p1_or_148555_comb = p1_prod__611_comb | 32'h0000_0080;
  assign p1_smul_59010_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__74_squeezed_comb, 9'h0d5);
  assign p1_smul_59012_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__75_squeezed_comb, 9'h105);
  assign p1_smul_59014_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__76_squeezed_comb, 9'h105);
  assign p1_smul_59016_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__77_squeezed_comb, 9'h0d5);
  assign p1_or_148570_comb = p1_prod__639_comb | 32'h0000_0080;
  assign p1_or_148571_comb = p1_prod__675_comb | 32'h0000_0080;
  assign p1_smul_59026_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__82_squeezed_comb, 9'h0d5);
  assign p1_smul_59028_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__83_squeezed_comb, 9'h105);
  assign p1_smul_59030_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__84_squeezed_comb, 9'h105);
  assign p1_smul_59032_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__85_squeezed_comb, 9'h0d5);
  assign p1_or_148586_comb = p1_prod__703_comb | 32'h0000_0080;
  assign p1_or_148587_comb = p1_prod__739_comb | 32'h0000_0080;
  assign p1_smul_59042_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__90_squeezed_comb, 9'h0d5);
  assign p1_smul_59044_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__91_squeezed_comb, 9'h105);
  assign p1_smul_59046_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__92_squeezed_comb, 9'h105);
  assign p1_smul_59048_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__93_squeezed_comb, 9'h0d5);
  assign p1_or_148602_comb = p1_prod__767_comb | 32'h0000_0080;
  assign p1_or_148603_comb = p1_prod__803_comb | 32'h0000_0080;
  assign p1_smul_59058_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__98_squeezed_comb, 9'h0d5);
  assign p1_smul_59060_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__99_squeezed_comb, 9'h105);
  assign p1_smul_59062_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__100_squeezed_comb, 9'h105);
  assign p1_smul_59064_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__101_squeezed_comb, 9'h0d5);
  assign p1_or_148618_comb = p1_prod__831_comb | 32'h0000_0080;
  assign p1_or_148619_comb = p1_prod__867_comb | 32'h0000_0080;
  assign p1_smul_59074_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__106_squeezed_comb, 9'h0d5);
  assign p1_smul_59076_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__107_squeezed_comb, 9'h105);
  assign p1_smul_59078_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__108_squeezed_comb, 9'h105);
  assign p1_smul_59080_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__109_squeezed_comb, 9'h0d5);
  assign p1_or_148634_comb = p1_prod__895_comb | 32'h0000_0080;
  assign p1_or_148635_comb = p1_prod__931_comb | 32'h0000_0080;
  assign p1_smul_59090_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__114_squeezed_comb, 9'h0d5);
  assign p1_smul_59092_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__115_squeezed_comb, 9'h105);
  assign p1_smul_59094_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__116_squeezed_comb, 9'h105);
  assign p1_smul_59096_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__117_squeezed_comb, 9'h0d5);
  assign p1_or_148650_comb = p1_prod__959_comb | 32'h0000_0080;
  assign p1_or_148651_comb = p1_prod__995_comb | 32'h0000_0080;
  assign p1_smul_59106_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__122_squeezed_comb, 9'h0d5);
  assign p1_smul_59108_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__123_squeezed_comb, 9'h105);
  assign p1_smul_59110_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__124_squeezed_comb, 9'h105);
  assign p1_smul_59112_NarrowedMult__comb = smul17b_8b_x_9b(p1_shifted__125_squeezed_comb, 9'h0d5);
  assign p1_or_148666_comb = p1_prod__1023_comb | 32'h0000_0080;
  assign p1_sel_148667_comb = $signed(p1_shifted__64_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__64_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__64_squeezed_comb, p1_smul_57326_TrailingBits___64_comb};
  assign p1_sel_148668_comb = $signed(p1_shifted__65_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__65_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__65_squeezed_comb, p1_smul_57326_TrailingBits___65_comb};
  assign p1_sel_148669_comb = $signed(p1_shifted__66_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__66_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__66_squeezed_comb, p1_smul_57326_TrailingBits___66_comb};
  assign p1_sel_148670_comb = $signed(p1_shifted__67_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__67_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__67_squeezed_comb, p1_smul_57326_TrailingBits___67_comb};
  assign p1_sel_148671_comb = $signed(p1_shifted__68_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__68_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__68_squeezed_comb, p1_smul_57326_TrailingBits___68_comb};
  assign p1_sel_148672_comb = $signed(p1_shifted__69_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__69_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__69_squeezed_comb, p1_smul_57326_TrailingBits___69_comb};
  assign p1_sel_148673_comb = $signed(p1_shifted__70_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__70_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__70_squeezed_comb, p1_smul_57326_TrailingBits___70_comb};
  assign p1_sel_148674_comb = $signed(p1_shifted__71_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__71_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__71_squeezed_comb, p1_smul_57326_TrailingBits___71_comb};
  assign p1_sel_148675_comb = $signed(p1_shifted__72_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__72_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__72_squeezed_comb, p1_smul_57326_TrailingBits___72_comb};
  assign p1_sel_148676_comb = $signed(p1_shifted__73_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__73_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__73_squeezed_comb, p1_smul_57326_TrailingBits___73_comb};
  assign p1_sel_148677_comb = $signed(p1_shifted__74_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__74_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__74_squeezed_comb, p1_smul_57326_TrailingBits___74_comb};
  assign p1_sel_148678_comb = $signed(p1_shifted__75_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__75_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__75_squeezed_comb, p1_smul_57326_TrailingBits___75_comb};
  assign p1_sel_148679_comb = $signed(p1_shifted__76_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__76_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__76_squeezed_comb, p1_smul_57326_TrailingBits___76_comb};
  assign p1_sel_148680_comb = $signed(p1_shifted__77_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__77_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__77_squeezed_comb, p1_smul_57326_TrailingBits___77_comb};
  assign p1_sel_148681_comb = $signed(p1_shifted__78_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__78_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__78_squeezed_comb, p1_smul_57326_TrailingBits___78_comb};
  assign p1_sel_148682_comb = $signed(p1_shifted__79_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__79_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__79_squeezed_comb, p1_smul_57326_TrailingBits___79_comb};
  assign p1_sel_148683_comb = $signed(p1_shifted__80_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__80_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__80_squeezed_comb, p1_smul_57326_TrailingBits___80_comb};
  assign p1_sel_148684_comb = $signed(p1_shifted__81_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__81_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__81_squeezed_comb, p1_smul_57326_TrailingBits___81_comb};
  assign p1_sel_148685_comb = $signed(p1_shifted__82_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__82_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__82_squeezed_comb, p1_smul_57326_TrailingBits___82_comb};
  assign p1_sel_148686_comb = $signed(p1_shifted__83_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__83_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__83_squeezed_comb, p1_smul_57326_TrailingBits___83_comb};
  assign p1_sel_148687_comb = $signed(p1_shifted__84_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__84_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__84_squeezed_comb, p1_smul_57326_TrailingBits___84_comb};
  assign p1_sel_148688_comb = $signed(p1_shifted__85_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__85_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__85_squeezed_comb, p1_smul_57326_TrailingBits___85_comb};
  assign p1_sel_148689_comb = $signed(p1_shifted__86_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__86_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__86_squeezed_comb, p1_smul_57326_TrailingBits___86_comb};
  assign p1_sel_148690_comb = $signed(p1_shifted__87_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__87_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__87_squeezed_comb, p1_smul_57326_TrailingBits___87_comb};
  assign p1_sel_148691_comb = $signed(p1_shifted__88_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__88_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__88_squeezed_comb, p1_smul_57326_TrailingBits___88_comb};
  assign p1_sel_148692_comb = $signed(p1_shifted__89_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__89_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__89_squeezed_comb, p1_smul_57326_TrailingBits___89_comb};
  assign p1_sel_148693_comb = $signed(p1_shifted__90_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__90_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__90_squeezed_comb, p1_smul_57326_TrailingBits___90_comb};
  assign p1_sel_148694_comb = $signed(p1_shifted__91_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__91_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__91_squeezed_comb, p1_smul_57326_TrailingBits___91_comb};
  assign p1_sel_148695_comb = $signed(p1_shifted__92_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__92_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__92_squeezed_comb, p1_smul_57326_TrailingBits___92_comb};
  assign p1_sel_148696_comb = $signed(p1_shifted__93_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__93_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__93_squeezed_comb, p1_smul_57326_TrailingBits___93_comb};
  assign p1_sel_148697_comb = $signed(p1_shifted__94_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__94_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__94_squeezed_comb, p1_smul_57326_TrailingBits___94_comb};
  assign p1_sel_148698_comb = $signed(p1_shifted__95_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__95_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__95_squeezed_comb, p1_smul_57326_TrailingBits___95_comb};
  assign p1_sel_148699_comb = $signed(p1_shifted__96_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__96_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__96_squeezed_comb, p1_smul_57326_TrailingBits___96_comb};
  assign p1_sel_148700_comb = $signed(p1_shifted__97_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__97_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__97_squeezed_comb, p1_smul_57326_TrailingBits___97_comb};
  assign p1_sel_148701_comb = $signed(p1_shifted__98_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__98_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__98_squeezed_comb, p1_smul_57326_TrailingBits___98_comb};
  assign p1_sel_148702_comb = $signed(p1_shifted__99_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__99_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__99_squeezed_comb, p1_smul_57326_TrailingBits___99_comb};
  assign p1_sel_148703_comb = $signed(p1_shifted__100_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__100_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__100_squeezed_comb, p1_smul_57326_TrailingBits___100_comb};
  assign p1_sel_148704_comb = $signed(p1_shifted__101_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__101_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__101_squeezed_comb, p1_smul_57326_TrailingBits___101_comb};
  assign p1_sel_148705_comb = $signed(p1_shifted__102_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__102_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__102_squeezed_comb, p1_smul_57326_TrailingBits___102_comb};
  assign p1_sel_148706_comb = $signed(p1_shifted__103_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__103_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__103_squeezed_comb, p1_smul_57326_TrailingBits___103_comb};
  assign p1_sel_148707_comb = $signed(p1_shifted__104_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__104_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__104_squeezed_comb, p1_smul_57326_TrailingBits___104_comb};
  assign p1_sel_148708_comb = $signed(p1_shifted__105_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__105_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__105_squeezed_comb, p1_smul_57326_TrailingBits___105_comb};
  assign p1_sel_148709_comb = $signed(p1_shifted__106_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__106_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__106_squeezed_comb, p1_smul_57326_TrailingBits___106_comb};
  assign p1_sel_148710_comb = $signed(p1_shifted__107_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__107_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__107_squeezed_comb, p1_smul_57326_TrailingBits___107_comb};
  assign p1_sel_148711_comb = $signed(p1_shifted__108_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__108_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__108_squeezed_comb, p1_smul_57326_TrailingBits___108_comb};
  assign p1_sel_148712_comb = $signed(p1_shifted__109_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__109_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__109_squeezed_comb, p1_smul_57326_TrailingBits___109_comb};
  assign p1_sel_148713_comb = $signed(p1_shifted__110_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__110_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__110_squeezed_comb, p1_smul_57326_TrailingBits___110_comb};
  assign p1_sel_148714_comb = $signed(p1_shifted__111_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__111_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__111_squeezed_comb, p1_smul_57326_TrailingBits___111_comb};
  assign p1_sel_148715_comb = $signed(p1_shifted__112_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__112_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__112_squeezed_comb, p1_smul_57326_TrailingBits___112_comb};
  assign p1_sel_148716_comb = $signed(p1_shifted__113_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__113_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__113_squeezed_comb, p1_smul_57326_TrailingBits___113_comb};
  assign p1_sel_148717_comb = $signed(p1_shifted__114_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__114_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__114_squeezed_comb, p1_smul_57326_TrailingBits___114_comb};
  assign p1_sel_148718_comb = $signed(p1_shifted__115_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__115_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__115_squeezed_comb, p1_smul_57326_TrailingBits___115_comb};
  assign p1_sel_148719_comb = $signed(p1_shifted__116_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__116_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__116_squeezed_comb, p1_smul_57326_TrailingBits___116_comb};
  assign p1_sel_148720_comb = $signed(p1_shifted__117_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__117_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__117_squeezed_comb, p1_smul_57326_TrailingBits___117_comb};
  assign p1_sel_148721_comb = $signed(p1_shifted__118_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__118_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__118_squeezed_comb, p1_smul_57326_TrailingBits___118_comb};
  assign p1_sel_148722_comb = $signed(p1_shifted__119_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__119_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__119_squeezed_comb, p1_smul_57326_TrailingBits___119_comb};
  assign p1_sel_148723_comb = $signed(p1_shifted__120_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__120_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__120_squeezed_comb, p1_smul_57326_TrailingBits___120_comb};
  assign p1_sel_148724_comb = $signed(p1_shifted__121_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__121_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__121_squeezed_comb, p1_smul_57326_TrailingBits___121_comb};
  assign p1_sel_148725_comb = $signed(p1_shifted__122_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__122_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__122_squeezed_comb, p1_smul_57326_TrailingBits___122_comb};
  assign p1_sel_148726_comb = $signed(p1_shifted__123_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__123_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__123_squeezed_comb, p1_smul_57326_TrailingBits___123_comb};
  assign p1_sel_148727_comb = $signed(p1_shifted__124_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__124_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__124_squeezed_comb, p1_smul_57326_TrailingBits___124_comb};
  assign p1_sel_148728_comb = $signed(p1_shifted__125_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__125_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__125_squeezed_comb, p1_smul_57326_TrailingBits___125_comb};
  assign p1_sel_148729_comb = $signed(p1_shifted__126_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__126_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__126_squeezed_comb, p1_smul_57326_TrailingBits___126_comb};
  assign p1_sel_148730_comb = $signed(p1_shifted__127_comb) > $signed(16'h7fff) ? 16'h7fff : {$signed(p1_shifted__127_squeezed_comb) < $signed(8'h80) ? 8'h80 : p1_shifted__127_squeezed_comb, p1_smul_57326_TrailingBits___127_comb};
  assign p1_add_151931_comb = {{1{p1_sel_148667_comb[15]}}, p1_sel_148667_comb} + {{1{p1_sel_148668_comb[15]}}, p1_sel_148668_comb};
  assign p1_add_151932_comb = {{1{p1_sel_148669_comb[15]}}, p1_sel_148669_comb} + {{1{p1_sel_148670_comb[15]}}, p1_sel_148670_comb};
  assign p1_add_151933_comb = {{1{p1_sel_148671_comb[15]}}, p1_sel_148671_comb} + {{1{p1_sel_148672_comb[15]}}, p1_sel_148672_comb};
  assign p1_add_151934_comb = {{1{p1_sel_148673_comb[15]}}, p1_sel_148673_comb} + {{1{p1_sel_148674_comb[15]}}, p1_sel_148674_comb};
  assign p1_add_151935_comb = {{1{p1_sel_148675_comb[15]}}, p1_sel_148675_comb} + {{1{p1_sel_148676_comb[15]}}, p1_sel_148676_comb};
  assign p1_add_151936_comb = {{1{p1_sel_148677_comb[15]}}, p1_sel_148677_comb} + {{1{p1_sel_148678_comb[15]}}, p1_sel_148678_comb};
  assign p1_add_151937_comb = {{1{p1_sel_148679_comb[15]}}, p1_sel_148679_comb} + {{1{p1_sel_148680_comb[15]}}, p1_sel_148680_comb};
  assign p1_add_151938_comb = {{1{p1_sel_148681_comb[15]}}, p1_sel_148681_comb} + {{1{p1_sel_148682_comb[15]}}, p1_sel_148682_comb};
  assign p1_add_151939_comb = {{1{p1_sel_148683_comb[15]}}, p1_sel_148683_comb} + {{1{p1_sel_148684_comb[15]}}, p1_sel_148684_comb};
  assign p1_add_151940_comb = {{1{p1_sel_148685_comb[15]}}, p1_sel_148685_comb} + {{1{p1_sel_148686_comb[15]}}, p1_sel_148686_comb};
  assign p1_add_151941_comb = {{1{p1_sel_148687_comb[15]}}, p1_sel_148687_comb} + {{1{p1_sel_148688_comb[15]}}, p1_sel_148688_comb};
  assign p1_add_151942_comb = {{1{p1_sel_148689_comb[15]}}, p1_sel_148689_comb} + {{1{p1_sel_148690_comb[15]}}, p1_sel_148690_comb};
  assign p1_add_151943_comb = {{1{p1_sel_148691_comb[15]}}, p1_sel_148691_comb} + {{1{p1_sel_148692_comb[15]}}, p1_sel_148692_comb};
  assign p1_add_151944_comb = {{1{p1_sel_148693_comb[15]}}, p1_sel_148693_comb} + {{1{p1_sel_148694_comb[15]}}, p1_sel_148694_comb};
  assign p1_add_151945_comb = {{1{p1_sel_148695_comb[15]}}, p1_sel_148695_comb} + {{1{p1_sel_148696_comb[15]}}, p1_sel_148696_comb};
  assign p1_add_151946_comb = {{1{p1_sel_148697_comb[15]}}, p1_sel_148697_comb} + {{1{p1_sel_148698_comb[15]}}, p1_sel_148698_comb};
  assign p1_add_151947_comb = {{1{p1_sel_148699_comb[15]}}, p1_sel_148699_comb} + {{1{p1_sel_148700_comb[15]}}, p1_sel_148700_comb};
  assign p1_add_151948_comb = {{1{p1_sel_148701_comb[15]}}, p1_sel_148701_comb} + {{1{p1_sel_148702_comb[15]}}, p1_sel_148702_comb};
  assign p1_add_151949_comb = {{1{p1_sel_148703_comb[15]}}, p1_sel_148703_comb} + {{1{p1_sel_148704_comb[15]}}, p1_sel_148704_comb};
  assign p1_add_151950_comb = {{1{p1_sel_148705_comb[15]}}, p1_sel_148705_comb} + {{1{p1_sel_148706_comb[15]}}, p1_sel_148706_comb};
  assign p1_add_151951_comb = {{1{p1_sel_148707_comb[15]}}, p1_sel_148707_comb} + {{1{p1_sel_148708_comb[15]}}, p1_sel_148708_comb};
  assign p1_add_151952_comb = {{1{p1_sel_148709_comb[15]}}, p1_sel_148709_comb} + {{1{p1_sel_148710_comb[15]}}, p1_sel_148710_comb};
  assign p1_add_151953_comb = {{1{p1_sel_148711_comb[15]}}, p1_sel_148711_comb} + {{1{p1_sel_148712_comb[15]}}, p1_sel_148712_comb};
  assign p1_add_151954_comb = {{1{p1_sel_148713_comb[15]}}, p1_sel_148713_comb} + {{1{p1_sel_148714_comb[15]}}, p1_sel_148714_comb};
  assign p1_add_151955_comb = {{1{p1_sel_148715_comb[15]}}, p1_sel_148715_comb} + {{1{p1_sel_148716_comb[15]}}, p1_sel_148716_comb};
  assign p1_add_151956_comb = {{1{p1_sel_148717_comb[15]}}, p1_sel_148717_comb} + {{1{p1_sel_148718_comb[15]}}, p1_sel_148718_comb};
  assign p1_add_151957_comb = {{1{p1_sel_148719_comb[15]}}, p1_sel_148719_comb} + {{1{p1_sel_148720_comb[15]}}, p1_sel_148720_comb};
  assign p1_add_151958_comb = {{1{p1_sel_148721_comb[15]}}, p1_sel_148721_comb} + {{1{p1_sel_148722_comb[15]}}, p1_sel_148722_comb};
  assign p1_add_151959_comb = {{1{p1_sel_148723_comb[15]}}, p1_sel_148723_comb} + {{1{p1_sel_148724_comb[15]}}, p1_sel_148724_comb};
  assign p1_add_151960_comb = {{1{p1_sel_148725_comb[15]}}, p1_sel_148725_comb} + {{1{p1_sel_148726_comb[15]}}, p1_sel_148726_comb};
  assign p1_add_151961_comb = {{1{p1_sel_148727_comb[15]}}, p1_sel_148727_comb} + {{1{p1_sel_148728_comb[15]}}, p1_sel_148728_comb};
  assign p1_add_151962_comb = {{1{p1_sel_148729_comb[15]}}, p1_sel_148729_comb} + {{1{p1_sel_148730_comb[15]}}, p1_sel_148730_comb};
  assign p1_sel_151963_comb = $signed(p1_smul_58222_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58222_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58222_NarrowedMult__comb[15:0]);
  assign p1_sel_151964_comb = $signed(p1_smul_58224_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58224_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58224_NarrowedMult__comb[15:0]);
  assign p1_sel_151965_comb = $signed(p1_or_146687_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__519_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146687_comb[23:9], 1'h0};
  assign p1_sel_151966_comb = $signed(p1_or_147714_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147714_comb[23:9], 1'h0};
  assign p1_sel_151967_comb = $signed(p1_or_147715_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147715_comb[23:9], 1'h0};
  assign p1_sel_151968_comb = $signed(p1_or_146694_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__534_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146694_comb[23:9], 1'h0};
  assign p1_sel_151969_comb = $signed(p1_smul_58234_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58234_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58234_NarrowedMult__comb[15:0]);
  assign p1_sel_151970_comb = $signed(p1_smul_58236_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58236_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58236_NarrowedMult__comb[15:0]);
  assign p1_sel_151971_comb = $signed(p1_smul_58238_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58238_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58238_NarrowedMult__comb[15:0]);
  assign p1_sel_151972_comb = $signed(p1_smul_58240_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58240_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58240_NarrowedMult__comb[15:0]);
  assign p1_sel_151973_comb = $signed(p1_or_146701_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__583_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146701_comb[23:9], 1'h0};
  assign p1_sel_151974_comb = $signed(p1_or_147730_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147730_comb[23:9], 1'h0};
  assign p1_sel_151975_comb = $signed(p1_or_147731_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147731_comb[23:9], 1'h0};
  assign p1_sel_151976_comb = $signed(p1_or_146708_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__598_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146708_comb[23:9], 1'h0};
  assign p1_sel_151977_comb = $signed(p1_smul_58250_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58250_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58250_NarrowedMult__comb[15:0]);
  assign p1_sel_151978_comb = $signed(p1_smul_58252_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58252_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58252_NarrowedMult__comb[15:0]);
  assign p1_sel_151979_comb = $signed(p1_smul_58254_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58254_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58254_NarrowedMult__comb[15:0]);
  assign p1_sel_151980_comb = $signed(p1_smul_58256_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58256_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58256_NarrowedMult__comb[15:0]);
  assign p1_sel_151981_comb = $signed(p1_or_146715_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__647_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146715_comb[23:9], 1'h0};
  assign p1_sel_151982_comb = $signed(p1_or_147746_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147746_comb[23:9], 1'h0};
  assign p1_sel_151983_comb = $signed(p1_or_147747_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147747_comb[23:9], 1'h0};
  assign p1_sel_151984_comb = $signed(p1_or_146722_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__662_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146722_comb[23:9], 1'h0};
  assign p1_sel_151985_comb = $signed(p1_smul_58266_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58266_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58266_NarrowedMult__comb[15:0]);
  assign p1_sel_151986_comb = $signed(p1_smul_58268_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58268_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58268_NarrowedMult__comb[15:0]);
  assign p1_sel_151987_comb = $signed(p1_smul_58270_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58270_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58270_NarrowedMult__comb[15:0]);
  assign p1_sel_151988_comb = $signed(p1_smul_58272_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58272_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58272_NarrowedMult__comb[15:0]);
  assign p1_sel_151989_comb = $signed(p1_or_146729_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__711_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146729_comb[23:9], 1'h0};
  assign p1_sel_151990_comb = $signed(p1_or_147762_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147762_comb[23:9], 1'h0};
  assign p1_sel_151991_comb = $signed(p1_or_147763_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147763_comb[23:9], 1'h0};
  assign p1_sel_151992_comb = $signed(p1_or_146736_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__726_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146736_comb[23:9], 1'h0};
  assign p1_sel_151993_comb = $signed(p1_smul_58282_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58282_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58282_NarrowedMult__comb[15:0]);
  assign p1_sel_151994_comb = $signed(p1_smul_58284_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58284_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58284_NarrowedMult__comb[15:0]);
  assign p1_sel_151995_comb = $signed(p1_smul_58286_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58286_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58286_NarrowedMult__comb[15:0]);
  assign p1_sel_151996_comb = $signed(p1_smul_58288_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58288_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58288_NarrowedMult__comb[15:0]);
  assign p1_sel_151997_comb = $signed(p1_or_146743_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__775_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146743_comb[23:9], 1'h0};
  assign p1_sel_151998_comb = $signed(p1_or_147778_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147778_comb[23:9], 1'h0};
  assign p1_sel_151999_comb = $signed(p1_or_147779_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147779_comb[23:9], 1'h0};
  assign p1_sel_152000_comb = $signed(p1_or_146750_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__790_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146750_comb[23:9], 1'h0};
  assign p1_sel_152001_comb = $signed(p1_smul_58298_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58298_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58298_NarrowedMult__comb[15:0]);
  assign p1_sel_152002_comb = $signed(p1_smul_58300_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58300_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58300_NarrowedMult__comb[15:0]);
  assign p1_sel_152003_comb = $signed(p1_smul_58302_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58302_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58302_NarrowedMult__comb[15:0]);
  assign p1_sel_152004_comb = $signed(p1_smul_58304_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58304_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58304_NarrowedMult__comb[15:0]);
  assign p1_sel_152005_comb = $signed(p1_or_146757_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__839_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146757_comb[23:9], 1'h0};
  assign p1_sel_152006_comb = $signed(p1_or_147794_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147794_comb[23:9], 1'h0};
  assign p1_sel_152007_comb = $signed(p1_or_147795_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147795_comb[23:9], 1'h0};
  assign p1_sel_152008_comb = $signed(p1_or_146764_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__854_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146764_comb[23:9], 1'h0};
  assign p1_sel_152009_comb = $signed(p1_smul_58314_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58314_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58314_NarrowedMult__comb[15:0]);
  assign p1_sel_152010_comb = $signed(p1_smul_58316_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58316_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58316_NarrowedMult__comb[15:0]);
  assign p1_sel_152011_comb = $signed(p1_smul_58318_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58318_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58318_NarrowedMult__comb[15:0]);
  assign p1_sel_152012_comb = $signed(p1_smul_58320_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58320_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58320_NarrowedMult__comb[15:0]);
  assign p1_sel_152013_comb = $signed(p1_or_146771_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__903_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146771_comb[23:9], 1'h0};
  assign p1_sel_152014_comb = $signed(p1_or_147810_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147810_comb[23:9], 1'h0};
  assign p1_sel_152015_comb = $signed(p1_or_147811_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147811_comb[23:9], 1'h0};
  assign p1_sel_152016_comb = $signed(p1_or_146778_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__918_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146778_comb[23:9], 1'h0};
  assign p1_sel_152017_comb = $signed(p1_smul_58330_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58330_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58330_NarrowedMult__comb[15:0]);
  assign p1_sel_152018_comb = $signed(p1_smul_58332_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58332_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58332_NarrowedMult__comb[15:0]);
  assign p1_sel_152019_comb = $signed(p1_smul_58334_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58334_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58334_NarrowedMult__comb[15:0]);
  assign p1_sel_152020_comb = $signed(p1_smul_58336_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58336_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58336_NarrowedMult__comb[15:0]);
  assign p1_sel_152021_comb = $signed(p1_or_146785_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__967_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146785_comb[23:9], 1'h0};
  assign p1_sel_152022_comb = $signed(p1_or_147826_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147826_comb[23:9], 1'h0};
  assign p1_sel_152023_comb = $signed(p1_or_147827_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147827_comb[23:9], 1'h0};
  assign p1_sel_152024_comb = $signed(p1_or_146792_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__982_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146792_comb[23:9], 1'h0};
  assign p1_sel_152025_comb = $signed(p1_smul_58346_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58346_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58346_NarrowedMult__comb[15:0]);
  assign p1_sel_152026_comb = $signed(p1_smul_58348_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58348_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58348_NarrowedMult__comb[15:0]);
  assign p1_sel_152027_comb = $signed(p1_or_146797_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__517_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146797_comb[23:10], 2'h0};
  assign p1_sel_152028_comb = $signed(p1_prod__520_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__520_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58352_NarrowedMult__comb, 1'h0};
  assign p1_sel_152029_comb = $signed(p1_prod__524_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__524_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58354_NarrowedMult__comb, 1'h0};
  assign p1_sel_152030_comb = $signed(p1_or_146804_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__529_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146804_comb[23:10], 2'h0};
  assign p1_sel_152031_comb = $signed(p1_or_146807_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__535_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146807_comb[23:10], 2'h0};
  assign p1_sel_152032_comb = $signed(p1_prod__542_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__542_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58360_NarrowedMult__comb, 1'h0};
  assign p1_sel_152033_comb = $signed(p1_prod__549_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__549_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58362_NarrowedMult__comb, 1'h0};
  assign p1_sel_152034_comb = $signed(p1_or_146814_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__555_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146814_comb[23:10], 2'h0};
  assign p1_sel_152035_comb = $signed(p1_or_146817_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__581_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146817_comb[23:10], 2'h0};
  assign p1_sel_152036_comb = $signed(p1_prod__584_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__584_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58368_NarrowedMult__comb, 1'h0};
  assign p1_sel_152037_comb = $signed(p1_prod__588_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__588_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58370_NarrowedMult__comb, 1'h0};
  assign p1_sel_152038_comb = $signed(p1_or_146824_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__593_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146824_comb[23:10], 2'h0};
  assign p1_sel_152039_comb = $signed(p1_or_146827_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__599_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146827_comb[23:10], 2'h0};
  assign p1_sel_152040_comb = $signed(p1_prod__606_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__606_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58376_NarrowedMult__comb, 1'h0};
  assign p1_sel_152041_comb = $signed(p1_prod__613_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__613_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58378_NarrowedMult__comb, 1'h0};
  assign p1_sel_152042_comb = $signed(p1_or_146834_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__619_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146834_comb[23:10], 2'h0};
  assign p1_sel_152043_comb = $signed(p1_or_146837_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__645_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146837_comb[23:10], 2'h0};
  assign p1_sel_152044_comb = $signed(p1_prod__648_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__648_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58384_NarrowedMult__comb, 1'h0};
  assign p1_sel_152045_comb = $signed(p1_prod__652_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__652_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58386_NarrowedMult__comb, 1'h0};
  assign p1_sel_152046_comb = $signed(p1_or_146844_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__657_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146844_comb[23:10], 2'h0};
  assign p1_sel_152047_comb = $signed(p1_or_146847_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__663_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146847_comb[23:10], 2'h0};
  assign p1_sel_152048_comb = $signed(p1_prod__670_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__670_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58392_NarrowedMult__comb, 1'h0};
  assign p1_sel_152049_comb = $signed(p1_prod__677_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__677_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58394_NarrowedMult__comb, 1'h0};
  assign p1_sel_152050_comb = $signed(p1_or_146854_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__683_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146854_comb[23:10], 2'h0};
  assign p1_sel_152051_comb = $signed(p1_or_146857_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__709_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146857_comb[23:10], 2'h0};
  assign p1_sel_152052_comb = $signed(p1_prod__712_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__712_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58400_NarrowedMult__comb, 1'h0};
  assign p1_sel_152053_comb = $signed(p1_prod__716_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__716_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58402_NarrowedMult__comb, 1'h0};
  assign p1_sel_152054_comb = $signed(p1_or_146864_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__721_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146864_comb[23:10], 2'h0};
  assign p1_sel_152055_comb = $signed(p1_or_146867_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__727_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146867_comb[23:10], 2'h0};
  assign p1_sel_152056_comb = $signed(p1_prod__734_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__734_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58408_NarrowedMult__comb, 1'h0};
  assign p1_sel_152057_comb = $signed(p1_prod__741_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__741_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58410_NarrowedMult__comb, 1'h0};
  assign p1_sel_152058_comb = $signed(p1_or_146874_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__747_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146874_comb[23:10], 2'h0};
  assign p1_sel_152059_comb = $signed(p1_or_146877_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__773_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146877_comb[23:10], 2'h0};
  assign p1_sel_152060_comb = $signed(p1_prod__776_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__776_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58416_NarrowedMult__comb, 1'h0};
  assign p1_sel_152061_comb = $signed(p1_prod__780_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__780_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58418_NarrowedMult__comb, 1'h0};
  assign p1_sel_152062_comb = $signed(p1_or_146884_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__785_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146884_comb[23:10], 2'h0};
  assign p1_sel_152063_comb = $signed(p1_or_146887_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__791_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146887_comb[23:10], 2'h0};
  assign p1_sel_152064_comb = $signed(p1_prod__798_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__798_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58424_NarrowedMult__comb, 1'h0};
  assign p1_sel_152065_comb = $signed(p1_prod__805_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__805_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58426_NarrowedMult__comb, 1'h0};
  assign p1_sel_152066_comb = $signed(p1_or_146894_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__811_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146894_comb[23:10], 2'h0};
  assign p1_sel_152067_comb = $signed(p1_or_146897_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__837_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146897_comb[23:10], 2'h0};
  assign p1_sel_152068_comb = $signed(p1_prod__840_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__840_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58432_NarrowedMult__comb, 1'h0};
  assign p1_sel_152069_comb = $signed(p1_prod__844_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__844_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58434_NarrowedMult__comb, 1'h0};
  assign p1_sel_152070_comb = $signed(p1_or_146904_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__849_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146904_comb[23:10], 2'h0};
  assign p1_sel_152071_comb = $signed(p1_or_146907_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__855_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146907_comb[23:10], 2'h0};
  assign p1_sel_152072_comb = $signed(p1_prod__862_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__862_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58440_NarrowedMult__comb, 1'h0};
  assign p1_sel_152073_comb = $signed(p1_prod__869_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__869_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58442_NarrowedMult__comb, 1'h0};
  assign p1_sel_152074_comb = $signed(p1_or_146914_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__875_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146914_comb[23:10], 2'h0};
  assign p1_sel_152075_comb = $signed(p1_or_146917_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__901_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146917_comb[23:10], 2'h0};
  assign p1_sel_152076_comb = $signed(p1_prod__904_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__904_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58448_NarrowedMult__comb, 1'h0};
  assign p1_sel_152077_comb = $signed(p1_prod__908_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__908_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58450_NarrowedMult__comb, 1'h0};
  assign p1_sel_152078_comb = $signed(p1_or_146924_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__913_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146924_comb[23:10], 2'h0};
  assign p1_sel_152079_comb = $signed(p1_or_146927_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__919_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146927_comb[23:10], 2'h0};
  assign p1_sel_152080_comb = $signed(p1_prod__926_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__926_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58456_NarrowedMult__comb, 1'h0};
  assign p1_sel_152081_comb = $signed(p1_prod__933_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__933_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58458_NarrowedMult__comb, 1'h0};
  assign p1_sel_152082_comb = $signed(p1_or_146934_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__939_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146934_comb[23:10], 2'h0};
  assign p1_sel_152083_comb = $signed(p1_or_146937_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__965_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146937_comb[23:10], 2'h0};
  assign p1_sel_152084_comb = $signed(p1_prod__968_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__968_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58464_NarrowedMult__comb, 1'h0};
  assign p1_sel_152085_comb = $signed(p1_prod__972_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__972_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58466_NarrowedMult__comb, 1'h0};
  assign p1_sel_152086_comb = $signed(p1_or_146944_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__977_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146944_comb[23:10], 2'h0};
  assign p1_sel_152087_comb = $signed(p1_or_146947_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__983_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146947_comb[23:10], 2'h0};
  assign p1_sel_152088_comb = $signed(p1_prod__990_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__990_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58472_NarrowedMult__comb, 1'h0};
  assign p1_sel_152089_comb = $signed(p1_prod__997_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__997_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58474_NarrowedMult__comb, 1'h0};
  assign p1_sel_152090_comb = $signed(p1_or_146954_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1003_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_146954_comb[23:10], 2'h0};
  assign p1_sel_152091_comb = $signed(p1_smul_58478_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58478_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58478_NarrowedMult__comb[15:0]);
  assign p1_sel_152092_comb = $signed(p1_or_147997_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_147997_comb[23:9], 1'h0};
  assign p1_sel_152093_comb = $signed(p1_smul_58482_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58482_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58482_NarrowedMult__comb[15:0]);
  assign p1_sel_152094_comb = $signed(p1_or_146961_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__536_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146961_comb[23:9], 1'h0};
  assign p1_sel_152095_comb = $signed(p1_or_146964_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__543_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146964_comb[23:9], 1'h0};
  assign p1_sel_152096_comb = $signed(p1_smul_58488_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58488_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58488_NarrowedMult__comb[15:0]);
  assign p1_sel_152097_comb = $signed(p1_or_148008_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148008_comb[23:9], 1'h0};
  assign p1_sel_152098_comb = $signed(p1_smul_58492_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58492_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58492_NarrowedMult__comb[15:0]);
  assign p1_sel_152099_comb = $signed(p1_smul_58494_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58494_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58494_NarrowedMult__comb[15:0]);
  assign p1_sel_152100_comb = $signed(p1_or_148013_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148013_comb[23:9], 1'h0};
  assign p1_sel_152101_comb = $signed(p1_smul_58498_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58498_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58498_NarrowedMult__comb[15:0]);
  assign p1_sel_152102_comb = $signed(p1_or_146975_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__600_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146975_comb[23:9], 1'h0};
  assign p1_sel_152103_comb = $signed(p1_or_146978_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__607_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146978_comb[23:9], 1'h0};
  assign p1_sel_152104_comb = $signed(p1_smul_58504_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58504_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58504_NarrowedMult__comb[15:0]);
  assign p1_sel_152105_comb = $signed(p1_or_148024_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148024_comb[23:9], 1'h0};
  assign p1_sel_152106_comb = $signed(p1_smul_58508_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58508_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58508_NarrowedMult__comb[15:0]);
  assign p1_sel_152107_comb = $signed(p1_smul_58510_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58510_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58510_NarrowedMult__comb[15:0]);
  assign p1_sel_152108_comb = $signed(p1_or_148029_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148029_comb[23:9], 1'h0};
  assign p1_sel_152109_comb = $signed(p1_smul_58514_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58514_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58514_NarrowedMult__comb[15:0]);
  assign p1_sel_152110_comb = $signed(p1_or_146989_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__664_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146989_comb[23:9], 1'h0};
  assign p1_sel_152111_comb = $signed(p1_or_146992_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__671_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_146992_comb[23:9], 1'h0};
  assign p1_sel_152112_comb = $signed(p1_smul_58520_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58520_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58520_NarrowedMult__comb[15:0]);
  assign p1_sel_152113_comb = $signed(p1_or_148040_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148040_comb[23:9], 1'h0};
  assign p1_sel_152114_comb = $signed(p1_smul_58524_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58524_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58524_NarrowedMult__comb[15:0]);
  assign p1_sel_152115_comb = $signed(p1_smul_58526_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58526_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58526_NarrowedMult__comb[15:0]);
  assign p1_sel_152116_comb = $signed(p1_or_148045_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148045_comb[23:9], 1'h0};
  assign p1_sel_152117_comb = $signed(p1_smul_58530_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58530_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58530_NarrowedMult__comb[15:0]);
  assign p1_sel_152118_comb = $signed(p1_or_147003_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__728_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147003_comb[23:9], 1'h0};
  assign p1_sel_152119_comb = $signed(p1_or_147006_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__735_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147006_comb[23:9], 1'h0};
  assign p1_sel_152120_comb = $signed(p1_smul_58536_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58536_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58536_NarrowedMult__comb[15:0]);
  assign p1_sel_152121_comb = $signed(p1_or_148056_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148056_comb[23:9], 1'h0};
  assign p1_sel_152122_comb = $signed(p1_smul_58540_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58540_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58540_NarrowedMult__comb[15:0]);
  assign p1_sel_152123_comb = $signed(p1_smul_58542_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58542_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58542_NarrowedMult__comb[15:0]);
  assign p1_sel_152124_comb = $signed(p1_or_148061_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148061_comb[23:9], 1'h0};
  assign p1_sel_152125_comb = $signed(p1_smul_58546_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58546_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58546_NarrowedMult__comb[15:0]);
  assign p1_sel_152126_comb = $signed(p1_or_147017_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__792_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147017_comb[23:9], 1'h0};
  assign p1_sel_152127_comb = $signed(p1_or_147020_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__799_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147020_comb[23:9], 1'h0};
  assign p1_sel_152128_comb = $signed(p1_smul_58552_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58552_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58552_NarrowedMult__comb[15:0]);
  assign p1_sel_152129_comb = $signed(p1_or_148072_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148072_comb[23:9], 1'h0};
  assign p1_sel_152130_comb = $signed(p1_smul_58556_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58556_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58556_NarrowedMult__comb[15:0]);
  assign p1_sel_152131_comb = $signed(p1_smul_58558_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58558_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58558_NarrowedMult__comb[15:0]);
  assign p1_sel_152132_comb = $signed(p1_or_148077_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148077_comb[23:9], 1'h0};
  assign p1_sel_152133_comb = $signed(p1_smul_58562_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58562_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58562_NarrowedMult__comb[15:0]);
  assign p1_sel_152134_comb = $signed(p1_or_147031_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__856_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147031_comb[23:9], 1'h0};
  assign p1_sel_152135_comb = $signed(p1_or_147034_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__863_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147034_comb[23:9], 1'h0};
  assign p1_sel_152136_comb = $signed(p1_smul_58568_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58568_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58568_NarrowedMult__comb[15:0]);
  assign p1_sel_152137_comb = $signed(p1_or_148088_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148088_comb[23:9], 1'h0};
  assign p1_sel_152138_comb = $signed(p1_smul_58572_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58572_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58572_NarrowedMult__comb[15:0]);
  assign p1_sel_152139_comb = $signed(p1_smul_58574_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58574_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58574_NarrowedMult__comb[15:0]);
  assign p1_sel_152140_comb = $signed(p1_or_148093_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148093_comb[23:9], 1'h0};
  assign p1_sel_152141_comb = $signed(p1_smul_58578_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58578_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58578_NarrowedMult__comb[15:0]);
  assign p1_sel_152142_comb = $signed(p1_or_147045_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__920_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147045_comb[23:9], 1'h0};
  assign p1_sel_152143_comb = $signed(p1_or_147048_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__927_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147048_comb[23:9], 1'h0};
  assign p1_sel_152144_comb = $signed(p1_smul_58584_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58584_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58584_NarrowedMult__comb[15:0]);
  assign p1_sel_152145_comb = $signed(p1_or_148104_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148104_comb[23:9], 1'h0};
  assign p1_sel_152146_comb = $signed(p1_smul_58588_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58588_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58588_NarrowedMult__comb[15:0]);
  assign p1_sel_152147_comb = $signed(p1_smul_58590_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58590_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58590_NarrowedMult__comb[15:0]);
  assign p1_sel_152148_comb = $signed(p1_or_148109_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148109_comb[23:9], 1'h0};
  assign p1_sel_152149_comb = $signed(p1_smul_58594_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58594_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58594_NarrowedMult__comb[15:0]);
  assign p1_sel_152150_comb = $signed(p1_or_147059_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__984_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147059_comb[23:9], 1'h0};
  assign p1_sel_152151_comb = $signed(p1_or_147062_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__991_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147062_comb[23:9], 1'h0};
  assign p1_sel_152152_comb = $signed(p1_smul_58600_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58600_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58600_NarrowedMult__comb[15:0]);
  assign p1_sel_152153_comb = $signed(p1_or_148120_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148120_comb[23:9], 1'h0};
  assign p1_sel_152154_comb = $signed(p1_smul_58604_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58604_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58604_NarrowedMult__comb[15:0]);
  assign p1_sel_152155_comb = $signed(p1_smul_58606_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58606_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58606_NarrowedMult__comb[15:0]);
  assign p1_sel_152156_comb = $signed(p1_smul_58608_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58608_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58608_NarrowedMult__comb[15:0]);
  assign p1_sel_152157_comb = $signed(p1_smul_58610_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58610_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58610_NarrowedMult__comb[15:0]);
  assign p1_sel_152158_comb = $signed(p1_smul_58612_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58612_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58612_NarrowedMult__comb[15:0]);
  assign p1_sel_152159_comb = $signed(p1_smul_58614_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58614_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58614_NarrowedMult__comb[15:0]);
  assign p1_sel_152160_comb = $signed(p1_smul_58616_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58616_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58616_NarrowedMult__comb[15:0]);
  assign p1_sel_152161_comb = $signed(p1_smul_58618_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58618_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58618_NarrowedMult__comb[15:0]);
  assign p1_sel_152162_comb = $signed(p1_smul_58620_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58620_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58620_NarrowedMult__comb[15:0]);
  assign p1_sel_152163_comb = $signed(p1_smul_58622_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58622_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58622_NarrowedMult__comb[15:0]);
  assign p1_sel_152164_comb = $signed(p1_smul_58624_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58624_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58624_NarrowedMult__comb[15:0]);
  assign p1_sel_152165_comb = $signed(p1_smul_58626_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58626_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58626_NarrowedMult__comb[15:0]);
  assign p1_sel_152166_comb = $signed(p1_smul_58628_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58628_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58628_NarrowedMult__comb[15:0]);
  assign p1_sel_152167_comb = $signed(p1_smul_58630_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58630_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58630_NarrowedMult__comb[15:0]);
  assign p1_sel_152168_comb = $signed(p1_smul_58632_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58632_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58632_NarrowedMult__comb[15:0]);
  assign p1_sel_152169_comb = $signed(p1_smul_58634_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58634_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58634_NarrowedMult__comb[15:0]);
  assign p1_sel_152170_comb = $signed(p1_smul_58636_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58636_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58636_NarrowedMult__comb[15:0]);
  assign p1_sel_152171_comb = $signed(p1_smul_58638_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58638_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58638_NarrowedMult__comb[15:0]);
  assign p1_sel_152172_comb = $signed(p1_smul_58640_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58640_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58640_NarrowedMult__comb[15:0]);
  assign p1_sel_152173_comb = $signed(p1_smul_58642_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58642_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58642_NarrowedMult__comb[15:0]);
  assign p1_sel_152174_comb = $signed(p1_smul_58644_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58644_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58644_NarrowedMult__comb[15:0]);
  assign p1_sel_152175_comb = $signed(p1_smul_58646_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58646_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58646_NarrowedMult__comb[15:0]);
  assign p1_sel_152176_comb = $signed(p1_smul_58648_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58648_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58648_NarrowedMult__comb[15:0]);
  assign p1_sel_152177_comb = $signed(p1_smul_58650_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58650_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58650_NarrowedMult__comb[15:0]);
  assign p1_sel_152178_comb = $signed(p1_smul_58652_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58652_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58652_NarrowedMult__comb[15:0]);
  assign p1_sel_152179_comb = $signed(p1_smul_58654_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58654_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58654_NarrowedMult__comb[15:0]);
  assign p1_sel_152180_comb = $signed(p1_smul_58656_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58656_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58656_NarrowedMult__comb[15:0]);
  assign p1_sel_152181_comb = $signed(p1_smul_58658_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58658_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58658_NarrowedMult__comb[15:0]);
  assign p1_sel_152182_comb = $signed(p1_smul_58660_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58660_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58660_NarrowedMult__comb[15:0]);
  assign p1_sel_152183_comb = $signed(p1_smul_58662_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58662_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58662_NarrowedMult__comb[15:0]);
  assign p1_sel_152184_comb = $signed(p1_smul_58664_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58664_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58664_NarrowedMult__comb[15:0]);
  assign p1_sel_152185_comb = $signed(p1_smul_58666_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58666_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58666_NarrowedMult__comb[15:0]);
  assign p1_sel_152186_comb = $signed(p1_smul_58668_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58668_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58668_NarrowedMult__comb[15:0]);
  assign p1_sel_152187_comb = $signed(p1_smul_58670_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58670_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58670_NarrowedMult__comb[15:0]);
  assign p1_sel_152188_comb = $signed(p1_smul_58672_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58672_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58672_NarrowedMult__comb[15:0]);
  assign p1_sel_152189_comb = $signed(p1_smul_58674_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58674_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58674_NarrowedMult__comb[15:0]);
  assign p1_sel_152190_comb = $signed(p1_smul_58676_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58676_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58676_NarrowedMult__comb[15:0]);
  assign p1_sel_152191_comb = $signed(p1_smul_58678_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58678_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58678_NarrowedMult__comb[15:0]);
  assign p1_sel_152192_comb = $signed(p1_smul_58680_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58680_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58680_NarrowedMult__comb[15:0]);
  assign p1_sel_152193_comb = $signed(p1_smul_58682_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58682_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58682_NarrowedMult__comb[15:0]);
  assign p1_sel_152194_comb = $signed(p1_smul_58684_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58684_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58684_NarrowedMult__comb[15:0]);
  assign p1_sel_152195_comb = $signed(p1_smul_58686_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58686_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58686_NarrowedMult__comb[15:0]);
  assign p1_sel_152196_comb = $signed(p1_smul_58688_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58688_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58688_NarrowedMult__comb[15:0]);
  assign p1_sel_152197_comb = $signed(p1_smul_58690_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58690_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58690_NarrowedMult__comb[15:0]);
  assign p1_sel_152198_comb = $signed(p1_smul_58692_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58692_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58692_NarrowedMult__comb[15:0]);
  assign p1_sel_152199_comb = $signed(p1_smul_58694_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58694_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58694_NarrowedMult__comb[15:0]);
  assign p1_sel_152200_comb = $signed(p1_smul_58696_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58696_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58696_NarrowedMult__comb[15:0]);
  assign p1_sel_152201_comb = $signed(p1_smul_58698_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58698_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58698_NarrowedMult__comb[15:0]);
  assign p1_sel_152202_comb = $signed(p1_smul_58700_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58700_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58700_NarrowedMult__comb[15:0]);
  assign p1_sel_152203_comb = $signed(p1_smul_58702_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58702_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58702_NarrowedMult__comb[15:0]);
  assign p1_sel_152204_comb = $signed(p1_smul_58704_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58704_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58704_NarrowedMult__comb[15:0]);
  assign p1_sel_152205_comb = $signed(p1_smul_58706_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58706_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58706_NarrowedMult__comb[15:0]);
  assign p1_sel_152206_comb = $signed(p1_smul_58708_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58708_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58708_NarrowedMult__comb[15:0]);
  assign p1_sel_152207_comb = $signed(p1_smul_58710_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58710_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58710_NarrowedMult__comb[15:0]);
  assign p1_sel_152208_comb = $signed(p1_smul_58712_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58712_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58712_NarrowedMult__comb[15:0]);
  assign p1_sel_152209_comb = $signed(p1_smul_58714_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58714_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58714_NarrowedMult__comb[15:0]);
  assign p1_sel_152210_comb = $signed(p1_smul_58716_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58716_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58716_NarrowedMult__comb[15:0]);
  assign p1_sel_152211_comb = $signed(p1_smul_58718_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58718_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58718_NarrowedMult__comb[15:0]);
  assign p1_sel_152212_comb = $signed(p1_smul_58720_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58720_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58720_NarrowedMult__comb[15:0]);
  assign p1_sel_152213_comb = $signed(p1_smul_58722_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58722_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58722_NarrowedMult__comb[15:0]);
  assign p1_sel_152214_comb = $signed(p1_smul_58724_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58724_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58724_NarrowedMult__comb[15:0]);
  assign p1_sel_152215_comb = $signed(p1_smul_58726_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58726_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58726_NarrowedMult__comb[15:0]);
  assign p1_sel_152216_comb = $signed(p1_smul_58728_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58728_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58728_NarrowedMult__comb[15:0]);
  assign p1_sel_152217_comb = $signed(p1_smul_58730_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58730_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58730_NarrowedMult__comb[15:0]);
  assign p1_sel_152218_comb = $signed(p1_smul_58732_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58732_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58732_NarrowedMult__comb[15:0]);
  assign p1_sel_152219_comb = $signed(p1_or_147133_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__532_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147133_comb[23:9], 1'h0};
  assign p1_sel_152220_comb = $signed(p1_smul_58736_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58736_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58736_NarrowedMult__comb[15:0]);
  assign p1_sel_152221_comb = $signed(p1_or_148256_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148256_comb[23:9], 1'h0};
  assign p1_sel_152222_comb = $signed(p1_smul_58740_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58740_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58740_NarrowedMult__comb[15:0]);
  assign p1_sel_152223_comb = $signed(p1_smul_58742_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58742_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58742_NarrowedMult__comb[15:0]);
  assign p1_sel_152224_comb = $signed(p1_or_148261_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148261_comb[23:9], 1'h0};
  assign p1_sel_152225_comb = $signed(p1_smul_58746_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58746_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58746_NarrowedMult__comb[15:0]);
  assign p1_sel_152226_comb = $signed(p1_or_147144_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__570_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147144_comb[23:9], 1'h0};
  assign p1_sel_152227_comb = $signed(p1_or_147147_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__596_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147147_comb[23:9], 1'h0};
  assign p1_sel_152228_comb = $signed(p1_smul_58752_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58752_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58752_NarrowedMult__comb[15:0]);
  assign p1_sel_152229_comb = $signed(p1_or_148272_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148272_comb[23:9], 1'h0};
  assign p1_sel_152230_comb = $signed(p1_smul_58756_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58756_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58756_NarrowedMult__comb[15:0]);
  assign p1_sel_152231_comb = $signed(p1_smul_58758_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58758_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58758_NarrowedMult__comb[15:0]);
  assign p1_sel_152232_comb = $signed(p1_or_148277_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148277_comb[23:9], 1'h0};
  assign p1_sel_152233_comb = $signed(p1_smul_58762_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58762_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58762_NarrowedMult__comb[15:0]);
  assign p1_sel_152234_comb = $signed(p1_or_147158_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__634_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147158_comb[23:9], 1'h0};
  assign p1_sel_152235_comb = $signed(p1_or_147161_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__660_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147161_comb[23:9], 1'h0};
  assign p1_sel_152236_comb = $signed(p1_smul_58768_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58768_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58768_NarrowedMult__comb[15:0]);
  assign p1_sel_152237_comb = $signed(p1_or_148288_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148288_comb[23:9], 1'h0};
  assign p1_sel_152238_comb = $signed(p1_smul_58772_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58772_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58772_NarrowedMult__comb[15:0]);
  assign p1_sel_152239_comb = $signed(p1_smul_58774_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58774_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58774_NarrowedMult__comb[15:0]);
  assign p1_sel_152240_comb = $signed(p1_or_148293_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148293_comb[23:9], 1'h0};
  assign p1_sel_152241_comb = $signed(p1_smul_58778_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58778_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58778_NarrowedMult__comb[15:0]);
  assign p1_sel_152242_comb = $signed(p1_or_147172_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__698_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147172_comb[23:9], 1'h0};
  assign p1_sel_152243_comb = $signed(p1_or_147175_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__724_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147175_comb[23:9], 1'h0};
  assign p1_sel_152244_comb = $signed(p1_smul_58784_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58784_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58784_NarrowedMult__comb[15:0]);
  assign p1_sel_152245_comb = $signed(p1_or_148304_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148304_comb[23:9], 1'h0};
  assign p1_sel_152246_comb = $signed(p1_smul_58788_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58788_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58788_NarrowedMult__comb[15:0]);
  assign p1_sel_152247_comb = $signed(p1_smul_58790_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58790_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58790_NarrowedMult__comb[15:0]);
  assign p1_sel_152248_comb = $signed(p1_or_148309_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148309_comb[23:9], 1'h0};
  assign p1_sel_152249_comb = $signed(p1_smul_58794_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58794_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58794_NarrowedMult__comb[15:0]);
  assign p1_sel_152250_comb = $signed(p1_or_147186_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__762_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147186_comb[23:9], 1'h0};
  assign p1_sel_152251_comb = $signed(p1_or_147189_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__788_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147189_comb[23:9], 1'h0};
  assign p1_sel_152252_comb = $signed(p1_smul_58800_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58800_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58800_NarrowedMult__comb[15:0]);
  assign p1_sel_152253_comb = $signed(p1_or_148320_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148320_comb[23:9], 1'h0};
  assign p1_sel_152254_comb = $signed(p1_smul_58804_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58804_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58804_NarrowedMult__comb[15:0]);
  assign p1_sel_152255_comb = $signed(p1_smul_58806_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58806_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58806_NarrowedMult__comb[15:0]);
  assign p1_sel_152256_comb = $signed(p1_or_148325_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148325_comb[23:9], 1'h0};
  assign p1_sel_152257_comb = $signed(p1_smul_58810_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58810_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58810_NarrowedMult__comb[15:0]);
  assign p1_sel_152258_comb = $signed(p1_or_147200_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__826_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147200_comb[23:9], 1'h0};
  assign p1_sel_152259_comb = $signed(p1_or_147203_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__852_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147203_comb[23:9], 1'h0};
  assign p1_sel_152260_comb = $signed(p1_smul_58816_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58816_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58816_NarrowedMult__comb[15:0]);
  assign p1_sel_152261_comb = $signed(p1_or_148336_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148336_comb[23:9], 1'h0};
  assign p1_sel_152262_comb = $signed(p1_smul_58820_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58820_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58820_NarrowedMult__comb[15:0]);
  assign p1_sel_152263_comb = $signed(p1_smul_58822_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58822_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58822_NarrowedMult__comb[15:0]);
  assign p1_sel_152264_comb = $signed(p1_or_148341_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148341_comb[23:9], 1'h0};
  assign p1_sel_152265_comb = $signed(p1_smul_58826_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58826_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58826_NarrowedMult__comb[15:0]);
  assign p1_sel_152266_comb = $signed(p1_or_147214_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__890_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147214_comb[23:9], 1'h0};
  assign p1_sel_152267_comb = $signed(p1_or_147217_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__916_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147217_comb[23:9], 1'h0};
  assign p1_sel_152268_comb = $signed(p1_smul_58832_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58832_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58832_NarrowedMult__comb[15:0]);
  assign p1_sel_152269_comb = $signed(p1_or_148352_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148352_comb[23:9], 1'h0};
  assign p1_sel_152270_comb = $signed(p1_smul_58836_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58836_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58836_NarrowedMult__comb[15:0]);
  assign p1_sel_152271_comb = $signed(p1_smul_58838_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58838_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58838_NarrowedMult__comb[15:0]);
  assign p1_sel_152272_comb = $signed(p1_or_148357_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148357_comb[23:9], 1'h0};
  assign p1_sel_152273_comb = $signed(p1_smul_58842_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58842_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58842_NarrowedMult__comb[15:0]);
  assign p1_sel_152274_comb = $signed(p1_or_147228_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__954_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147228_comb[23:9], 1'h0};
  assign p1_sel_152275_comb = $signed(p1_or_147231_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__980_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147231_comb[23:9], 1'h0};
  assign p1_sel_152276_comb = $signed(p1_smul_58848_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58848_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58848_NarrowedMult__comb[15:0]);
  assign p1_sel_152277_comb = $signed(p1_or_148368_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148368_comb[23:9], 1'h0};
  assign p1_sel_152278_comb = $signed(p1_smul_58852_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58852_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58852_NarrowedMult__comb[15:0]);
  assign p1_sel_152279_comb = $signed(p1_smul_58854_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58854_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58854_NarrowedMult__comb[15:0]);
  assign p1_sel_152280_comb = $signed(p1_or_148373_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148373_comb[23:9], 1'h0};
  assign p1_sel_152281_comb = $signed(p1_smul_58858_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58858_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58858_NarrowedMult__comb[15:0]);
  assign p1_sel_152282_comb = $signed(p1_or_147242_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1018_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147242_comb[23:9], 1'h0};
  assign p1_sel_152283_comb = $signed(p1_prod__539_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__539_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58862_NarrowedMult__comb, 1'h0};
  assign p1_sel_152284_comb = $signed(p1_or_147247_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__546_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147247_comb[23:10], 2'h0};
  assign p1_sel_152285_comb = $signed(p1_prod__553_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__553_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58866_NarrowedMult__comb, 1'h0};
  assign p1_sel_152286_comb = $signed(p1_or_147252_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__559_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147252_comb[23:10], 2'h0};
  assign p1_sel_152287_comb = $signed(p1_or_147255_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__564_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147255_comb[23:10], 2'h0};
  assign p1_sel_152288_comb = $signed(p1_prod__568_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__568_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58872_NarrowedMult__comb, 1'h0};
  assign p1_sel_152289_comb = $signed(p1_or_147260_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__571_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147260_comb[23:10], 2'h0};
  assign p1_sel_152290_comb = $signed(p1_prod__573_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__573_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58876_NarrowedMult__comb, 1'h0};
  assign p1_sel_152291_comb = $signed(p1_prod__603_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__603_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58878_NarrowedMult__comb, 1'h0};
  assign p1_sel_152292_comb = $signed(p1_or_147267_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__610_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147267_comb[23:10], 2'h0};
  assign p1_sel_152293_comb = $signed(p1_prod__617_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__617_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58882_NarrowedMult__comb, 1'h0};
  assign p1_sel_152294_comb = $signed(p1_or_147272_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__623_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147272_comb[23:10], 2'h0};
  assign p1_sel_152295_comb = $signed(p1_or_147275_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__628_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147275_comb[23:10], 2'h0};
  assign p1_sel_152296_comb = $signed(p1_prod__632_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__632_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58888_NarrowedMult__comb, 1'h0};
  assign p1_sel_152297_comb = $signed(p1_or_147280_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__635_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147280_comb[23:10], 2'h0};
  assign p1_sel_152298_comb = $signed(p1_prod__637_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__637_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58892_NarrowedMult__comb, 1'h0};
  assign p1_sel_152299_comb = $signed(p1_prod__667_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__667_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58894_NarrowedMult__comb, 1'h0};
  assign p1_sel_152300_comb = $signed(p1_or_147287_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__674_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147287_comb[23:10], 2'h0};
  assign p1_sel_152301_comb = $signed(p1_prod__681_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__681_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58898_NarrowedMult__comb, 1'h0};
  assign p1_sel_152302_comb = $signed(p1_or_147292_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__687_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147292_comb[23:10], 2'h0};
  assign p1_sel_152303_comb = $signed(p1_or_147295_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__692_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147295_comb[23:10], 2'h0};
  assign p1_sel_152304_comb = $signed(p1_prod__696_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__696_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58904_NarrowedMult__comb, 1'h0};
  assign p1_sel_152305_comb = $signed(p1_or_147300_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__699_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147300_comb[23:10], 2'h0};
  assign p1_sel_152306_comb = $signed(p1_prod__701_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__701_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58908_NarrowedMult__comb, 1'h0};
  assign p1_sel_152307_comb = $signed(p1_prod__731_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__731_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58910_NarrowedMult__comb, 1'h0};
  assign p1_sel_152308_comb = $signed(p1_or_147307_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__738_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147307_comb[23:10], 2'h0};
  assign p1_sel_152309_comb = $signed(p1_prod__745_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__745_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58914_NarrowedMult__comb, 1'h0};
  assign p1_sel_152310_comb = $signed(p1_or_147312_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__751_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147312_comb[23:10], 2'h0};
  assign p1_sel_152311_comb = $signed(p1_or_147315_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__756_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147315_comb[23:10], 2'h0};
  assign p1_sel_152312_comb = $signed(p1_prod__760_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__760_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58920_NarrowedMult__comb, 1'h0};
  assign p1_sel_152313_comb = $signed(p1_or_147320_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__763_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147320_comb[23:10], 2'h0};
  assign p1_sel_152314_comb = $signed(p1_prod__765_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__765_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58924_NarrowedMult__comb, 1'h0};
  assign p1_sel_152315_comb = $signed(p1_prod__795_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__795_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58926_NarrowedMult__comb, 1'h0};
  assign p1_sel_152316_comb = $signed(p1_or_147327_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__802_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147327_comb[23:10], 2'h0};
  assign p1_sel_152317_comb = $signed(p1_prod__809_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__809_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58930_NarrowedMult__comb, 1'h0};
  assign p1_sel_152318_comb = $signed(p1_or_147332_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__815_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147332_comb[23:10], 2'h0};
  assign p1_sel_152319_comb = $signed(p1_or_147335_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__820_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147335_comb[23:10], 2'h0};
  assign p1_sel_152320_comb = $signed(p1_prod__824_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__824_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58936_NarrowedMult__comb, 1'h0};
  assign p1_sel_152321_comb = $signed(p1_or_147340_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__827_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147340_comb[23:10], 2'h0};
  assign p1_sel_152322_comb = $signed(p1_prod__829_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__829_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58940_NarrowedMult__comb, 1'h0};
  assign p1_sel_152323_comb = $signed(p1_prod__859_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__859_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58942_NarrowedMult__comb, 1'h0};
  assign p1_sel_152324_comb = $signed(p1_or_147347_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__866_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147347_comb[23:10], 2'h0};
  assign p1_sel_152325_comb = $signed(p1_prod__873_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__873_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58946_NarrowedMult__comb, 1'h0};
  assign p1_sel_152326_comb = $signed(p1_or_147352_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__879_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147352_comb[23:10], 2'h0};
  assign p1_sel_152327_comb = $signed(p1_or_147355_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__884_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147355_comb[23:10], 2'h0};
  assign p1_sel_152328_comb = $signed(p1_prod__888_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__888_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58952_NarrowedMult__comb, 1'h0};
  assign p1_sel_152329_comb = $signed(p1_or_147360_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__891_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147360_comb[23:10], 2'h0};
  assign p1_sel_152330_comb = $signed(p1_prod__893_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__893_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58956_NarrowedMult__comb, 1'h0};
  assign p1_sel_152331_comb = $signed(p1_prod__923_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__923_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58958_NarrowedMult__comb, 1'h0};
  assign p1_sel_152332_comb = $signed(p1_or_147367_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__930_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147367_comb[23:10], 2'h0};
  assign p1_sel_152333_comb = $signed(p1_prod__937_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__937_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58962_NarrowedMult__comb, 1'h0};
  assign p1_sel_152334_comb = $signed(p1_or_147372_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__943_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147372_comb[23:10], 2'h0};
  assign p1_sel_152335_comb = $signed(p1_or_147375_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__948_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147375_comb[23:10], 2'h0};
  assign p1_sel_152336_comb = $signed(p1_prod__952_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__952_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58968_NarrowedMult__comb, 1'h0};
  assign p1_sel_152337_comb = $signed(p1_or_147380_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__955_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147380_comb[23:10], 2'h0};
  assign p1_sel_152338_comb = $signed(p1_prod__957_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__957_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58972_NarrowedMult__comb, 1'h0};
  assign p1_sel_152339_comb = $signed(p1_prod__987_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__987_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58974_NarrowedMult__comb, 1'h0};
  assign p1_sel_152340_comb = $signed(p1_or_147387_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__994_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147387_comb[23:10], 2'h0};
  assign p1_sel_152341_comb = $signed(p1_prod__1001_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1001_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58978_NarrowedMult__comb, 1'h0};
  assign p1_sel_152342_comb = $signed(p1_or_147392_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1007_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147392_comb[23:10], 2'h0};
  assign p1_sel_152343_comb = $signed(p1_or_147395_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1012_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147395_comb[23:10], 2'h0};
  assign p1_sel_152344_comb = $signed(p1_prod__1016_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1016_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58984_NarrowedMult__comb, 1'h0};
  assign p1_sel_152345_comb = $signed(p1_or_147400_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1019_comb[31:10]) < $signed(22'h3f_e000) ? 14'h2000 : p1_or_147400_comb[23:10], 2'h0};
  assign p1_sel_152346_comb = $signed(p1_prod__1021_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1021_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_smul_58988_NarrowedMult__comb, 1'h0};
  assign p1_sel_152347_comb = $signed(p1_or_148539_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148539_comb[23:9], 1'h0};
  assign p1_sel_152348_comb = $signed(p1_or_147407_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__554_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147407_comb[23:9], 1'h0};
  assign p1_sel_152349_comb = $signed(p1_smul_58994_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58994_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58994_NarrowedMult__comb[15:0]);
  assign p1_sel_152350_comb = $signed(p1_smul_58996_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58996_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58996_NarrowedMult__comb[15:0]);
  assign p1_sel_152351_comb = $signed(p1_smul_58998_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_58998_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_58998_NarrowedMult__comb[15:0]);
  assign p1_sel_152352_comb = $signed(p1_smul_59000_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59000_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59000_NarrowedMult__comb[15:0]);
  assign p1_sel_152353_comb = $signed(p1_or_147414_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__574_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147414_comb[23:9], 1'h0};
  assign p1_sel_152354_comb = $signed(p1_or_148554_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148554_comb[23:9], 1'h0};
  assign p1_sel_152355_comb = $signed(p1_or_148555_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148555_comb[23:9], 1'h0};
  assign p1_sel_152356_comb = $signed(p1_or_147421_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__618_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147421_comb[23:9], 1'h0};
  assign p1_sel_152357_comb = $signed(p1_smul_59010_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59010_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59010_NarrowedMult__comb[15:0]);
  assign p1_sel_152358_comb = $signed(p1_smul_59012_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59012_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59012_NarrowedMult__comb[15:0]);
  assign p1_sel_152359_comb = $signed(p1_smul_59014_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59014_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59014_NarrowedMult__comb[15:0]);
  assign p1_sel_152360_comb = $signed(p1_smul_59016_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59016_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59016_NarrowedMult__comb[15:0]);
  assign p1_sel_152361_comb = $signed(p1_or_147428_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__638_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147428_comb[23:9], 1'h0};
  assign p1_sel_152362_comb = $signed(p1_or_148570_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148570_comb[23:9], 1'h0};
  assign p1_sel_152363_comb = $signed(p1_or_148571_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148571_comb[23:9], 1'h0};
  assign p1_sel_152364_comb = $signed(p1_or_147435_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__682_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147435_comb[23:9], 1'h0};
  assign p1_sel_152365_comb = $signed(p1_smul_59026_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59026_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59026_NarrowedMult__comb[15:0]);
  assign p1_sel_152366_comb = $signed(p1_smul_59028_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59028_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59028_NarrowedMult__comb[15:0]);
  assign p1_sel_152367_comb = $signed(p1_smul_59030_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59030_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59030_NarrowedMult__comb[15:0]);
  assign p1_sel_152368_comb = $signed(p1_smul_59032_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59032_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59032_NarrowedMult__comb[15:0]);
  assign p1_sel_152369_comb = $signed(p1_or_147442_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__702_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147442_comb[23:9], 1'h0};
  assign p1_sel_152370_comb = $signed(p1_or_148586_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148586_comb[23:9], 1'h0};
  assign p1_sel_152371_comb = $signed(p1_or_148587_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148587_comb[23:9], 1'h0};
  assign p1_sel_152372_comb = $signed(p1_or_147449_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__746_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147449_comb[23:9], 1'h0};
  assign p1_sel_152373_comb = $signed(p1_smul_59042_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59042_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59042_NarrowedMult__comb[15:0]);
  assign p1_sel_152374_comb = $signed(p1_smul_59044_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59044_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59044_NarrowedMult__comb[15:0]);
  assign p1_sel_152375_comb = $signed(p1_smul_59046_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59046_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59046_NarrowedMult__comb[15:0]);
  assign p1_sel_152376_comb = $signed(p1_smul_59048_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59048_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59048_NarrowedMult__comb[15:0]);
  assign p1_sel_152377_comb = $signed(p1_or_147456_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__766_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147456_comb[23:9], 1'h0};
  assign p1_sel_152378_comb = $signed(p1_or_148602_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148602_comb[23:9], 1'h0};
  assign p1_sel_152379_comb = $signed(p1_or_148603_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148603_comb[23:9], 1'h0};
  assign p1_sel_152380_comb = $signed(p1_or_147463_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__810_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147463_comb[23:9], 1'h0};
  assign p1_sel_152381_comb = $signed(p1_smul_59058_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59058_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59058_NarrowedMult__comb[15:0]);
  assign p1_sel_152382_comb = $signed(p1_smul_59060_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59060_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59060_NarrowedMult__comb[15:0]);
  assign p1_sel_152383_comb = $signed(p1_smul_59062_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59062_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59062_NarrowedMult__comb[15:0]);
  assign p1_sel_152384_comb = $signed(p1_smul_59064_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59064_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59064_NarrowedMult__comb[15:0]);
  assign p1_sel_152385_comb = $signed(p1_or_147470_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__830_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147470_comb[23:9], 1'h0};
  assign p1_sel_152386_comb = $signed(p1_or_148618_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148618_comb[23:9], 1'h0};
  assign p1_sel_152387_comb = $signed(p1_or_148619_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148619_comb[23:9], 1'h0};
  assign p1_sel_152388_comb = $signed(p1_or_147477_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__874_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147477_comb[23:9], 1'h0};
  assign p1_sel_152389_comb = $signed(p1_smul_59074_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59074_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59074_NarrowedMult__comb[15:0]);
  assign p1_sel_152390_comb = $signed(p1_smul_59076_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59076_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59076_NarrowedMult__comb[15:0]);
  assign p1_sel_152391_comb = $signed(p1_smul_59078_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59078_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59078_NarrowedMult__comb[15:0]);
  assign p1_sel_152392_comb = $signed(p1_smul_59080_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59080_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59080_NarrowedMult__comb[15:0]);
  assign p1_sel_152393_comb = $signed(p1_or_147484_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__894_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147484_comb[23:9], 1'h0};
  assign p1_sel_152394_comb = $signed(p1_or_148634_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148634_comb[23:9], 1'h0};
  assign p1_sel_152395_comb = $signed(p1_or_148635_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148635_comb[23:9], 1'h0};
  assign p1_sel_152396_comb = $signed(p1_or_147491_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__938_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147491_comb[23:9], 1'h0};
  assign p1_sel_152397_comb = $signed(p1_smul_59090_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59090_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59090_NarrowedMult__comb[15:0]);
  assign p1_sel_152398_comb = $signed(p1_smul_59092_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59092_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59092_NarrowedMult__comb[15:0]);
  assign p1_sel_152399_comb = $signed(p1_smul_59094_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59094_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59094_NarrowedMult__comb[15:0]);
  assign p1_sel_152400_comb = $signed(p1_smul_59096_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59096_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59096_NarrowedMult__comb[15:0]);
  assign p1_sel_152401_comb = $signed(p1_or_147498_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__958_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147498_comb[23:9], 1'h0};
  assign p1_sel_152402_comb = $signed(p1_or_148650_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148650_comb[23:9], 1'h0};
  assign p1_sel_152403_comb = $signed(p1_or_148651_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148651_comb[23:9], 1'h0};
  assign p1_sel_152404_comb = $signed(p1_or_147505_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1002_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147505_comb[23:9], 1'h0};
  assign p1_sel_152405_comb = $signed(p1_smul_59106_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59106_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59106_NarrowedMult__comb[15:0]);
  assign p1_sel_152406_comb = $signed(p1_smul_59108_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59108_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59108_NarrowedMult__comb[15:0]);
  assign p1_sel_152407_comb = $signed(p1_smul_59110_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59110_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59110_NarrowedMult__comb[15:0]);
  assign p1_sel_152408_comb = $signed(p1_smul_59112_NarrowedMult__comb) > $signed(17'h0_7fff) ? 16'h7fff : ($signed(p1_smul_59112_NarrowedMult__comb) < $signed(17'h1_8000) ? 16'h8000 : p1_smul_59112_NarrowedMult__comb[15:0]);
  assign p1_sel_152409_comb = $signed(p1_or_147512_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {$signed(p1_prod__1022_comb[31:9]) < $signed(23'h7f_c000) ? 15'h4000 : p1_or_147512_comb[23:9], 1'h0};
  assign p1_sel_152410_comb = $signed(p1_or_148666_comb[31:8]) > $signed(24'h00_7fff) ? 16'h7fff : {p1_or_148666_comb[23:9], 1'h0};
  assign p1_sum__520_comb = {{15{p1_add_151931_comb[16]}}, p1_add_151931_comb};
  assign p1_sum__521_comb = {{15{p1_add_151932_comb[16]}}, p1_add_151932_comb};
  assign p1_sum__522_comb = {{15{p1_add_151933_comb[16]}}, p1_add_151933_comb};
  assign p1_sum__523_comb = {{15{p1_add_151934_comb[16]}}, p1_add_151934_comb};
  assign p1_sum__464_comb = {{15{p1_add_151935_comb[16]}}, p1_add_151935_comb};
  assign p1_sum__465_comb = {{15{p1_add_151936_comb[16]}}, p1_add_151936_comb};
  assign p1_sum__466_comb = {{15{p1_add_151937_comb[16]}}, p1_add_151937_comb};
  assign p1_sum__467_comb = {{15{p1_add_151938_comb[16]}}, p1_add_151938_comb};
  assign p1_sum__408_comb = {{15{p1_add_151939_comb[16]}}, p1_add_151939_comb};
  assign p1_sum__409_comb = {{15{p1_add_151940_comb[16]}}, p1_add_151940_comb};
  assign p1_sum__410_comb = {{15{p1_add_151941_comb[16]}}, p1_add_151941_comb};
  assign p1_sum__411_comb = {{15{p1_add_151942_comb[16]}}, p1_add_151942_comb};
  assign p1_sum__352_comb = {{15{p1_add_151943_comb[16]}}, p1_add_151943_comb};
  assign p1_sum__353_comb = {{15{p1_add_151944_comb[16]}}, p1_add_151944_comb};
  assign p1_sum__354_comb = {{15{p1_add_151945_comb[16]}}, p1_add_151945_comb};
  assign p1_sum__355_comb = {{15{p1_add_151946_comb[16]}}, p1_add_151946_comb};
  assign p1_sum__296_comb = {{15{p1_add_151947_comb[16]}}, p1_add_151947_comb};
  assign p1_sum__297_comb = {{15{p1_add_151948_comb[16]}}, p1_add_151948_comb};
  assign p1_sum__298_comb = {{15{p1_add_151949_comb[16]}}, p1_add_151949_comb};
  assign p1_sum__299_comb = {{15{p1_add_151950_comb[16]}}, p1_add_151950_comb};
  assign p1_sum__240_comb = {{15{p1_add_151951_comb[16]}}, p1_add_151951_comb};
  assign p1_sum__241_comb = {{15{p1_add_151952_comb[16]}}, p1_add_151952_comb};
  assign p1_sum__242_comb = {{15{p1_add_151953_comb[16]}}, p1_add_151953_comb};
  assign p1_sum__243_comb = {{15{p1_add_151954_comb[16]}}, p1_add_151954_comb};
  assign p1_sum__184_comb = {{15{p1_add_151955_comb[16]}}, p1_add_151955_comb};
  assign p1_sum__185_comb = {{15{p1_add_151956_comb[16]}}, p1_add_151956_comb};
  assign p1_sum__186_comb = {{15{p1_add_151957_comb[16]}}, p1_add_151957_comb};
  assign p1_sum__187_comb = {{15{p1_add_151958_comb[16]}}, p1_add_151958_comb};
  assign p1_sum__128_comb = {{15{p1_add_151959_comb[16]}}, p1_add_151959_comb};
  assign p1_sum__129_comb = {{15{p1_add_151960_comb[16]}}, p1_add_151960_comb};
  assign p1_sum__130_comb = {{15{p1_add_151961_comb[16]}}, p1_add_151961_comb};
  assign p1_sum__131_comb = {{15{p1_add_151962_comb[16]}}, p1_add_151962_comb};
  assign p1_sum__524_comb = p1_sum__520_comb + p1_sum__521_comb;
  assign p1_sum__525_comb = p1_sum__522_comb + p1_sum__523_comb;
  assign p1_sum__468_comb = p1_sum__464_comb + p1_sum__465_comb;
  assign p1_sum__469_comb = p1_sum__466_comb + p1_sum__467_comb;
  assign p1_sum__412_comb = p1_sum__408_comb + p1_sum__409_comb;
  assign p1_sum__413_comb = p1_sum__410_comb + p1_sum__411_comb;
  assign p1_sum__356_comb = p1_sum__352_comb + p1_sum__353_comb;
  assign p1_sum__357_comb = p1_sum__354_comb + p1_sum__355_comb;
  assign p1_sum__300_comb = p1_sum__296_comb + p1_sum__297_comb;
  assign p1_sum__301_comb = p1_sum__298_comb + p1_sum__299_comb;
  assign p1_sum__244_comb = p1_sum__240_comb + p1_sum__241_comb;
  assign p1_sum__245_comb = p1_sum__242_comb + p1_sum__243_comb;
  assign p1_sum__188_comb = p1_sum__184_comb + p1_sum__185_comb;
  assign p1_sum__189_comb = p1_sum__186_comb + p1_sum__187_comb;
  assign p1_sum__132_comb = p1_sum__128_comb + p1_sum__129_comb;
  assign p1_sum__133_comb = p1_sum__130_comb + p1_sum__131_comb;
  assign p1_add_152907_comb = {{1{p1_sel_151963_comb[15]}}, p1_sel_151963_comb} + {{1{p1_sel_151964_comb[15]}}, p1_sel_151964_comb};
  assign p1_add_152908_comb = {{1{p1_sel_151965_comb[15]}}, p1_sel_151965_comb} + {{1{p1_sel_151966_comb[15]}}, p1_sel_151966_comb};
  assign p1_add_152909_comb = {{1{p1_sel_151967_comb[15]}}, p1_sel_151967_comb} + {{1{p1_sel_151968_comb[15]}}, p1_sel_151968_comb};
  assign p1_add_152910_comb = {{1{p1_sel_151969_comb[15]}}, p1_sel_151969_comb} + {{1{p1_sel_151970_comb[15]}}, p1_sel_151970_comb};
  assign p1_add_152911_comb = {{1{p1_sel_151971_comb[15]}}, p1_sel_151971_comb} + {{1{p1_sel_151972_comb[15]}}, p1_sel_151972_comb};
  assign p1_add_152912_comb = {{1{p1_sel_151973_comb[15]}}, p1_sel_151973_comb} + {{1{p1_sel_151974_comb[15]}}, p1_sel_151974_comb};
  assign p1_add_152913_comb = {{1{p1_sel_151975_comb[15]}}, p1_sel_151975_comb} + {{1{p1_sel_151976_comb[15]}}, p1_sel_151976_comb};
  assign p1_add_152914_comb = {{1{p1_sel_151977_comb[15]}}, p1_sel_151977_comb} + {{1{p1_sel_151978_comb[15]}}, p1_sel_151978_comb};
  assign p1_add_152915_comb = {{1{p1_sel_151979_comb[15]}}, p1_sel_151979_comb} + {{1{p1_sel_151980_comb[15]}}, p1_sel_151980_comb};
  assign p1_add_152916_comb = {{1{p1_sel_151981_comb[15]}}, p1_sel_151981_comb} + {{1{p1_sel_151982_comb[15]}}, p1_sel_151982_comb};
  assign p1_add_152917_comb = {{1{p1_sel_151983_comb[15]}}, p1_sel_151983_comb} + {{1{p1_sel_151984_comb[15]}}, p1_sel_151984_comb};
  assign p1_add_152918_comb = {{1{p1_sel_151985_comb[15]}}, p1_sel_151985_comb} + {{1{p1_sel_151986_comb[15]}}, p1_sel_151986_comb};
  assign p1_add_152919_comb = {{1{p1_sel_151987_comb[15]}}, p1_sel_151987_comb} + {{1{p1_sel_151988_comb[15]}}, p1_sel_151988_comb};
  assign p1_add_152920_comb = {{1{p1_sel_151989_comb[15]}}, p1_sel_151989_comb} + {{1{p1_sel_151990_comb[15]}}, p1_sel_151990_comb};
  assign p1_add_152921_comb = {{1{p1_sel_151991_comb[15]}}, p1_sel_151991_comb} + {{1{p1_sel_151992_comb[15]}}, p1_sel_151992_comb};
  assign p1_add_152922_comb = {{1{p1_sel_151993_comb[15]}}, p1_sel_151993_comb} + {{1{p1_sel_151994_comb[15]}}, p1_sel_151994_comb};
  assign p1_add_152923_comb = {{1{p1_sel_151995_comb[15]}}, p1_sel_151995_comb} + {{1{p1_sel_151996_comb[15]}}, p1_sel_151996_comb};
  assign p1_add_152924_comb = {{1{p1_sel_151997_comb[15]}}, p1_sel_151997_comb} + {{1{p1_sel_151998_comb[15]}}, p1_sel_151998_comb};
  assign p1_add_152925_comb = {{1{p1_sel_151999_comb[15]}}, p1_sel_151999_comb} + {{1{p1_sel_152000_comb[15]}}, p1_sel_152000_comb};
  assign p1_add_152926_comb = {{1{p1_sel_152001_comb[15]}}, p1_sel_152001_comb} + {{1{p1_sel_152002_comb[15]}}, p1_sel_152002_comb};
  assign p1_add_152927_comb = {{1{p1_sel_152003_comb[15]}}, p1_sel_152003_comb} + {{1{p1_sel_152004_comb[15]}}, p1_sel_152004_comb};
  assign p1_add_152928_comb = {{1{p1_sel_152005_comb[15]}}, p1_sel_152005_comb} + {{1{p1_sel_152006_comb[15]}}, p1_sel_152006_comb};
  assign p1_add_152929_comb = {{1{p1_sel_152007_comb[15]}}, p1_sel_152007_comb} + {{1{p1_sel_152008_comb[15]}}, p1_sel_152008_comb};
  assign p1_add_152930_comb = {{1{p1_sel_152009_comb[15]}}, p1_sel_152009_comb} + {{1{p1_sel_152010_comb[15]}}, p1_sel_152010_comb};
  assign p1_add_152931_comb = {{1{p1_sel_152011_comb[15]}}, p1_sel_152011_comb} + {{1{p1_sel_152012_comb[15]}}, p1_sel_152012_comb};
  assign p1_add_152932_comb = {{1{p1_sel_152013_comb[15]}}, p1_sel_152013_comb} + {{1{p1_sel_152014_comb[15]}}, p1_sel_152014_comb};
  assign p1_add_152933_comb = {{1{p1_sel_152015_comb[15]}}, p1_sel_152015_comb} + {{1{p1_sel_152016_comb[15]}}, p1_sel_152016_comb};
  assign p1_add_152934_comb = {{1{p1_sel_152017_comb[15]}}, p1_sel_152017_comb} + {{1{p1_sel_152018_comb[15]}}, p1_sel_152018_comb};
  assign p1_add_152935_comb = {{1{p1_sel_152019_comb[15]}}, p1_sel_152019_comb} + {{1{p1_sel_152020_comb[15]}}, p1_sel_152020_comb};
  assign p1_add_152936_comb = {{1{p1_sel_152021_comb[15]}}, p1_sel_152021_comb} + {{1{p1_sel_152022_comb[15]}}, p1_sel_152022_comb};
  assign p1_add_152937_comb = {{1{p1_sel_152023_comb[15]}}, p1_sel_152023_comb} + {{1{p1_sel_152024_comb[15]}}, p1_sel_152024_comb};
  assign p1_add_152938_comb = {{1{p1_sel_152025_comb[15]}}, p1_sel_152025_comb} + {{1{p1_sel_152026_comb[15]}}, p1_sel_152026_comb};
  assign p1_add_152939_comb = {{1{p1_sel_152027_comb[15]}}, p1_sel_152027_comb} + {{1{p1_sel_152028_comb[15]}}, p1_sel_152028_comb};
  assign p1_add_152940_comb = {{1{p1_sel_152029_comb[15]}}, p1_sel_152029_comb} + {{1{p1_sel_152030_comb[15]}}, p1_sel_152030_comb};
  assign p1_add_152941_comb = {{1{p1_sel_152031_comb[15]}}, p1_sel_152031_comb} + {{1{p1_sel_152032_comb[15]}}, p1_sel_152032_comb};
  assign p1_add_152942_comb = {{1{p1_sel_152033_comb[15]}}, p1_sel_152033_comb} + {{1{p1_sel_152034_comb[15]}}, p1_sel_152034_comb};
  assign p1_add_152943_comb = {{1{p1_sel_152035_comb[15]}}, p1_sel_152035_comb} + {{1{p1_sel_152036_comb[15]}}, p1_sel_152036_comb};
  assign p1_add_152944_comb = {{1{p1_sel_152037_comb[15]}}, p1_sel_152037_comb} + {{1{p1_sel_152038_comb[15]}}, p1_sel_152038_comb};
  assign p1_add_152945_comb = {{1{p1_sel_152039_comb[15]}}, p1_sel_152039_comb} + {{1{p1_sel_152040_comb[15]}}, p1_sel_152040_comb};
  assign p1_add_152946_comb = {{1{p1_sel_152041_comb[15]}}, p1_sel_152041_comb} + {{1{p1_sel_152042_comb[15]}}, p1_sel_152042_comb};
  assign p1_add_152947_comb = {{1{p1_sel_152043_comb[15]}}, p1_sel_152043_comb} + {{1{p1_sel_152044_comb[15]}}, p1_sel_152044_comb};
  assign p1_add_152948_comb = {{1{p1_sel_152045_comb[15]}}, p1_sel_152045_comb} + {{1{p1_sel_152046_comb[15]}}, p1_sel_152046_comb};
  assign p1_add_152949_comb = {{1{p1_sel_152047_comb[15]}}, p1_sel_152047_comb} + {{1{p1_sel_152048_comb[15]}}, p1_sel_152048_comb};
  assign p1_add_152950_comb = {{1{p1_sel_152049_comb[15]}}, p1_sel_152049_comb} + {{1{p1_sel_152050_comb[15]}}, p1_sel_152050_comb};
  assign p1_add_152951_comb = {{1{p1_sel_152051_comb[15]}}, p1_sel_152051_comb} + {{1{p1_sel_152052_comb[15]}}, p1_sel_152052_comb};
  assign p1_add_152952_comb = {{1{p1_sel_152053_comb[15]}}, p1_sel_152053_comb} + {{1{p1_sel_152054_comb[15]}}, p1_sel_152054_comb};
  assign p1_add_152953_comb = {{1{p1_sel_152055_comb[15]}}, p1_sel_152055_comb} + {{1{p1_sel_152056_comb[15]}}, p1_sel_152056_comb};
  assign p1_add_152954_comb = {{1{p1_sel_152057_comb[15]}}, p1_sel_152057_comb} + {{1{p1_sel_152058_comb[15]}}, p1_sel_152058_comb};
  assign p1_add_152955_comb = {{1{p1_sel_152059_comb[15]}}, p1_sel_152059_comb} + {{1{p1_sel_152060_comb[15]}}, p1_sel_152060_comb};
  assign p1_add_152956_comb = {{1{p1_sel_152061_comb[15]}}, p1_sel_152061_comb} + {{1{p1_sel_152062_comb[15]}}, p1_sel_152062_comb};
  assign p1_add_152957_comb = {{1{p1_sel_152063_comb[15]}}, p1_sel_152063_comb} + {{1{p1_sel_152064_comb[15]}}, p1_sel_152064_comb};
  assign p1_add_152958_comb = {{1{p1_sel_152065_comb[15]}}, p1_sel_152065_comb} + {{1{p1_sel_152066_comb[15]}}, p1_sel_152066_comb};
  assign p1_add_152959_comb = {{1{p1_sel_152067_comb[15]}}, p1_sel_152067_comb} + {{1{p1_sel_152068_comb[15]}}, p1_sel_152068_comb};
  assign p1_add_152960_comb = {{1{p1_sel_152069_comb[15]}}, p1_sel_152069_comb} + {{1{p1_sel_152070_comb[15]}}, p1_sel_152070_comb};
  assign p1_add_152961_comb = {{1{p1_sel_152071_comb[15]}}, p1_sel_152071_comb} + {{1{p1_sel_152072_comb[15]}}, p1_sel_152072_comb};
  assign p1_add_152962_comb = {{1{p1_sel_152073_comb[15]}}, p1_sel_152073_comb} + {{1{p1_sel_152074_comb[15]}}, p1_sel_152074_comb};
  assign p1_add_152963_comb = {{1{p1_sel_152075_comb[15]}}, p1_sel_152075_comb} + {{1{p1_sel_152076_comb[15]}}, p1_sel_152076_comb};
  assign p1_add_152964_comb = {{1{p1_sel_152077_comb[15]}}, p1_sel_152077_comb} + {{1{p1_sel_152078_comb[15]}}, p1_sel_152078_comb};
  assign p1_add_152965_comb = {{1{p1_sel_152079_comb[15]}}, p1_sel_152079_comb} + {{1{p1_sel_152080_comb[15]}}, p1_sel_152080_comb};
  assign p1_add_152966_comb = {{1{p1_sel_152081_comb[15]}}, p1_sel_152081_comb} + {{1{p1_sel_152082_comb[15]}}, p1_sel_152082_comb};
  assign p1_add_152967_comb = {{1{p1_sel_152083_comb[15]}}, p1_sel_152083_comb} + {{1{p1_sel_152084_comb[15]}}, p1_sel_152084_comb};
  assign p1_add_152968_comb = {{1{p1_sel_152085_comb[15]}}, p1_sel_152085_comb} + {{1{p1_sel_152086_comb[15]}}, p1_sel_152086_comb};
  assign p1_add_152969_comb = {{1{p1_sel_152087_comb[15]}}, p1_sel_152087_comb} + {{1{p1_sel_152088_comb[15]}}, p1_sel_152088_comb};
  assign p1_add_152970_comb = {{1{p1_sel_152089_comb[15]}}, p1_sel_152089_comb} + {{1{p1_sel_152090_comb[15]}}, p1_sel_152090_comb};
  assign p1_add_152971_comb = {{1{p1_sel_152091_comb[15]}}, p1_sel_152091_comb} + {{1{p1_sel_152092_comb[15]}}, p1_sel_152092_comb};
  assign p1_add_152972_comb = {{1{p1_sel_152093_comb[15]}}, p1_sel_152093_comb} + {{1{p1_sel_152094_comb[15]}}, p1_sel_152094_comb};
  assign p1_add_152973_comb = {{1{p1_sel_152095_comb[15]}}, p1_sel_152095_comb} + {{1{p1_sel_152096_comb[15]}}, p1_sel_152096_comb};
  assign p1_add_152974_comb = {{1{p1_sel_152097_comb[15]}}, p1_sel_152097_comb} + {{1{p1_sel_152098_comb[15]}}, p1_sel_152098_comb};
  assign p1_add_152975_comb = {{1{p1_sel_152099_comb[15]}}, p1_sel_152099_comb} + {{1{p1_sel_152100_comb[15]}}, p1_sel_152100_comb};
  assign p1_add_152976_comb = {{1{p1_sel_152101_comb[15]}}, p1_sel_152101_comb} + {{1{p1_sel_152102_comb[15]}}, p1_sel_152102_comb};
  assign p1_add_152977_comb = {{1{p1_sel_152103_comb[15]}}, p1_sel_152103_comb} + {{1{p1_sel_152104_comb[15]}}, p1_sel_152104_comb};
  assign p1_add_152978_comb = {{1{p1_sel_152105_comb[15]}}, p1_sel_152105_comb} + {{1{p1_sel_152106_comb[15]}}, p1_sel_152106_comb};
  assign p1_add_152979_comb = {{1{p1_sel_152107_comb[15]}}, p1_sel_152107_comb} + {{1{p1_sel_152108_comb[15]}}, p1_sel_152108_comb};
  assign p1_add_152980_comb = {{1{p1_sel_152109_comb[15]}}, p1_sel_152109_comb} + {{1{p1_sel_152110_comb[15]}}, p1_sel_152110_comb};
  assign p1_add_152981_comb = {{1{p1_sel_152111_comb[15]}}, p1_sel_152111_comb} + {{1{p1_sel_152112_comb[15]}}, p1_sel_152112_comb};
  assign p1_add_152982_comb = {{1{p1_sel_152113_comb[15]}}, p1_sel_152113_comb} + {{1{p1_sel_152114_comb[15]}}, p1_sel_152114_comb};
  assign p1_add_152983_comb = {{1{p1_sel_152115_comb[15]}}, p1_sel_152115_comb} + {{1{p1_sel_152116_comb[15]}}, p1_sel_152116_comb};
  assign p1_add_152984_comb = {{1{p1_sel_152117_comb[15]}}, p1_sel_152117_comb} + {{1{p1_sel_152118_comb[15]}}, p1_sel_152118_comb};
  assign p1_add_152985_comb = {{1{p1_sel_152119_comb[15]}}, p1_sel_152119_comb} + {{1{p1_sel_152120_comb[15]}}, p1_sel_152120_comb};
  assign p1_add_152986_comb = {{1{p1_sel_152121_comb[15]}}, p1_sel_152121_comb} + {{1{p1_sel_152122_comb[15]}}, p1_sel_152122_comb};
  assign p1_add_152987_comb = {{1{p1_sel_152123_comb[15]}}, p1_sel_152123_comb} + {{1{p1_sel_152124_comb[15]}}, p1_sel_152124_comb};
  assign p1_add_152988_comb = {{1{p1_sel_152125_comb[15]}}, p1_sel_152125_comb} + {{1{p1_sel_152126_comb[15]}}, p1_sel_152126_comb};
  assign p1_add_152989_comb = {{1{p1_sel_152127_comb[15]}}, p1_sel_152127_comb} + {{1{p1_sel_152128_comb[15]}}, p1_sel_152128_comb};
  assign p1_add_152990_comb = {{1{p1_sel_152129_comb[15]}}, p1_sel_152129_comb} + {{1{p1_sel_152130_comb[15]}}, p1_sel_152130_comb};
  assign p1_add_152991_comb = {{1{p1_sel_152131_comb[15]}}, p1_sel_152131_comb} + {{1{p1_sel_152132_comb[15]}}, p1_sel_152132_comb};
  assign p1_add_152992_comb = {{1{p1_sel_152133_comb[15]}}, p1_sel_152133_comb} + {{1{p1_sel_152134_comb[15]}}, p1_sel_152134_comb};
  assign p1_add_152993_comb = {{1{p1_sel_152135_comb[15]}}, p1_sel_152135_comb} + {{1{p1_sel_152136_comb[15]}}, p1_sel_152136_comb};
  assign p1_add_152994_comb = {{1{p1_sel_152137_comb[15]}}, p1_sel_152137_comb} + {{1{p1_sel_152138_comb[15]}}, p1_sel_152138_comb};
  assign p1_add_152995_comb = {{1{p1_sel_152139_comb[15]}}, p1_sel_152139_comb} + {{1{p1_sel_152140_comb[15]}}, p1_sel_152140_comb};
  assign p1_add_152996_comb = {{1{p1_sel_152141_comb[15]}}, p1_sel_152141_comb} + {{1{p1_sel_152142_comb[15]}}, p1_sel_152142_comb};
  assign p1_add_152997_comb = {{1{p1_sel_152143_comb[15]}}, p1_sel_152143_comb} + {{1{p1_sel_152144_comb[15]}}, p1_sel_152144_comb};
  assign p1_add_152998_comb = {{1{p1_sel_152145_comb[15]}}, p1_sel_152145_comb} + {{1{p1_sel_152146_comb[15]}}, p1_sel_152146_comb};
  assign p1_add_152999_comb = {{1{p1_sel_152147_comb[15]}}, p1_sel_152147_comb} + {{1{p1_sel_152148_comb[15]}}, p1_sel_152148_comb};
  assign p1_add_153000_comb = {{1{p1_sel_152149_comb[15]}}, p1_sel_152149_comb} + {{1{p1_sel_152150_comb[15]}}, p1_sel_152150_comb};
  assign p1_add_153001_comb = {{1{p1_sel_152151_comb[15]}}, p1_sel_152151_comb} + {{1{p1_sel_152152_comb[15]}}, p1_sel_152152_comb};
  assign p1_add_153002_comb = {{1{p1_sel_152153_comb[15]}}, p1_sel_152153_comb} + {{1{p1_sel_152154_comb[15]}}, p1_sel_152154_comb};
  assign p1_add_153003_comb = {{1{p1_sel_152155_comb[15]}}, p1_sel_152155_comb} + {{1{p1_sel_152156_comb[15]}}, p1_sel_152156_comb};
  assign p1_add_153004_comb = {{1{p1_sel_152157_comb[15]}}, p1_sel_152157_comb} + {{1{p1_sel_152158_comb[15]}}, p1_sel_152158_comb};
  assign p1_add_153005_comb = {{1{p1_sel_152159_comb[15]}}, p1_sel_152159_comb} + {{1{p1_sel_152160_comb[15]}}, p1_sel_152160_comb};
  assign p1_add_153006_comb = {{1{p1_sel_152161_comb[15]}}, p1_sel_152161_comb} + {{1{p1_sel_152162_comb[15]}}, p1_sel_152162_comb};
  assign p1_add_153007_comb = {{1{p1_sel_152163_comb[15]}}, p1_sel_152163_comb} + {{1{p1_sel_152164_comb[15]}}, p1_sel_152164_comb};
  assign p1_add_153008_comb = {{1{p1_sel_152165_comb[15]}}, p1_sel_152165_comb} + {{1{p1_sel_152166_comb[15]}}, p1_sel_152166_comb};
  assign p1_add_153009_comb = {{1{p1_sel_152167_comb[15]}}, p1_sel_152167_comb} + {{1{p1_sel_152168_comb[15]}}, p1_sel_152168_comb};
  assign p1_add_153010_comb = {{1{p1_sel_152169_comb[15]}}, p1_sel_152169_comb} + {{1{p1_sel_152170_comb[15]}}, p1_sel_152170_comb};
  assign p1_add_153011_comb = {{1{p1_sel_152171_comb[15]}}, p1_sel_152171_comb} + {{1{p1_sel_152172_comb[15]}}, p1_sel_152172_comb};
  assign p1_add_153012_comb = {{1{p1_sel_152173_comb[15]}}, p1_sel_152173_comb} + {{1{p1_sel_152174_comb[15]}}, p1_sel_152174_comb};
  assign p1_add_153013_comb = {{1{p1_sel_152175_comb[15]}}, p1_sel_152175_comb} + {{1{p1_sel_152176_comb[15]}}, p1_sel_152176_comb};
  assign p1_add_153014_comb = {{1{p1_sel_152177_comb[15]}}, p1_sel_152177_comb} + {{1{p1_sel_152178_comb[15]}}, p1_sel_152178_comb};
  assign p1_add_153015_comb = {{1{p1_sel_152179_comb[15]}}, p1_sel_152179_comb} + {{1{p1_sel_152180_comb[15]}}, p1_sel_152180_comb};
  assign p1_add_153016_comb = {{1{p1_sel_152181_comb[15]}}, p1_sel_152181_comb} + {{1{p1_sel_152182_comb[15]}}, p1_sel_152182_comb};
  assign p1_add_153017_comb = {{1{p1_sel_152183_comb[15]}}, p1_sel_152183_comb} + {{1{p1_sel_152184_comb[15]}}, p1_sel_152184_comb};
  assign p1_add_153018_comb = {{1{p1_sel_152185_comb[15]}}, p1_sel_152185_comb} + {{1{p1_sel_152186_comb[15]}}, p1_sel_152186_comb};
  assign p1_add_153019_comb = {{1{p1_sel_152187_comb[15]}}, p1_sel_152187_comb} + {{1{p1_sel_152188_comb[15]}}, p1_sel_152188_comb};
  assign p1_add_153020_comb = {{1{p1_sel_152189_comb[15]}}, p1_sel_152189_comb} + {{1{p1_sel_152190_comb[15]}}, p1_sel_152190_comb};
  assign p1_add_153021_comb = {{1{p1_sel_152191_comb[15]}}, p1_sel_152191_comb} + {{1{p1_sel_152192_comb[15]}}, p1_sel_152192_comb};
  assign p1_add_153022_comb = {{1{p1_sel_152193_comb[15]}}, p1_sel_152193_comb} + {{1{p1_sel_152194_comb[15]}}, p1_sel_152194_comb};
  assign p1_add_153023_comb = {{1{p1_sel_152195_comb[15]}}, p1_sel_152195_comb} + {{1{p1_sel_152196_comb[15]}}, p1_sel_152196_comb};
  assign p1_add_153024_comb = {{1{p1_sel_152197_comb[15]}}, p1_sel_152197_comb} + {{1{p1_sel_152198_comb[15]}}, p1_sel_152198_comb};
  assign p1_add_153025_comb = {{1{p1_sel_152199_comb[15]}}, p1_sel_152199_comb} + {{1{p1_sel_152200_comb[15]}}, p1_sel_152200_comb};
  assign p1_add_153026_comb = {{1{p1_sel_152201_comb[15]}}, p1_sel_152201_comb} + {{1{p1_sel_152202_comb[15]}}, p1_sel_152202_comb};
  assign p1_add_153027_comb = {{1{p1_sel_152203_comb[15]}}, p1_sel_152203_comb} + {{1{p1_sel_152204_comb[15]}}, p1_sel_152204_comb};
  assign p1_add_153028_comb = {{1{p1_sel_152205_comb[15]}}, p1_sel_152205_comb} + {{1{p1_sel_152206_comb[15]}}, p1_sel_152206_comb};
  assign p1_add_153029_comb = {{1{p1_sel_152207_comb[15]}}, p1_sel_152207_comb} + {{1{p1_sel_152208_comb[15]}}, p1_sel_152208_comb};
  assign p1_add_153030_comb = {{1{p1_sel_152209_comb[15]}}, p1_sel_152209_comb} + {{1{p1_sel_152210_comb[15]}}, p1_sel_152210_comb};
  assign p1_add_153031_comb = {{1{p1_sel_152211_comb[15]}}, p1_sel_152211_comb} + {{1{p1_sel_152212_comb[15]}}, p1_sel_152212_comb};
  assign p1_add_153032_comb = {{1{p1_sel_152213_comb[15]}}, p1_sel_152213_comb} + {{1{p1_sel_152214_comb[15]}}, p1_sel_152214_comb};
  assign p1_add_153033_comb = {{1{p1_sel_152215_comb[15]}}, p1_sel_152215_comb} + {{1{p1_sel_152216_comb[15]}}, p1_sel_152216_comb};
  assign p1_add_153034_comb = {{1{p1_sel_152217_comb[15]}}, p1_sel_152217_comb} + {{1{p1_sel_152218_comb[15]}}, p1_sel_152218_comb};
  assign p1_add_153035_comb = {{1{p1_sel_152219_comb[15]}}, p1_sel_152219_comb} + {{1{p1_sel_152220_comb[15]}}, p1_sel_152220_comb};
  assign p1_add_153036_comb = {{1{p1_sel_152221_comb[15]}}, p1_sel_152221_comb} + {{1{p1_sel_152222_comb[15]}}, p1_sel_152222_comb};
  assign p1_add_153037_comb = {{1{p1_sel_152223_comb[15]}}, p1_sel_152223_comb} + {{1{p1_sel_152224_comb[15]}}, p1_sel_152224_comb};
  assign p1_add_153038_comb = {{1{p1_sel_152225_comb[15]}}, p1_sel_152225_comb} + {{1{p1_sel_152226_comb[15]}}, p1_sel_152226_comb};
  assign p1_add_153039_comb = {{1{p1_sel_152227_comb[15]}}, p1_sel_152227_comb} + {{1{p1_sel_152228_comb[15]}}, p1_sel_152228_comb};
  assign p1_add_153040_comb = {{1{p1_sel_152229_comb[15]}}, p1_sel_152229_comb} + {{1{p1_sel_152230_comb[15]}}, p1_sel_152230_comb};
  assign p1_add_153041_comb = {{1{p1_sel_152231_comb[15]}}, p1_sel_152231_comb} + {{1{p1_sel_152232_comb[15]}}, p1_sel_152232_comb};
  assign p1_add_153042_comb = {{1{p1_sel_152233_comb[15]}}, p1_sel_152233_comb} + {{1{p1_sel_152234_comb[15]}}, p1_sel_152234_comb};
  assign p1_add_153043_comb = {{1{p1_sel_152235_comb[15]}}, p1_sel_152235_comb} + {{1{p1_sel_152236_comb[15]}}, p1_sel_152236_comb};
  assign p1_add_153044_comb = {{1{p1_sel_152237_comb[15]}}, p1_sel_152237_comb} + {{1{p1_sel_152238_comb[15]}}, p1_sel_152238_comb};
  assign p1_add_153045_comb = {{1{p1_sel_152239_comb[15]}}, p1_sel_152239_comb} + {{1{p1_sel_152240_comb[15]}}, p1_sel_152240_comb};
  assign p1_add_153046_comb = {{1{p1_sel_152241_comb[15]}}, p1_sel_152241_comb} + {{1{p1_sel_152242_comb[15]}}, p1_sel_152242_comb};
  assign p1_add_153047_comb = {{1{p1_sel_152243_comb[15]}}, p1_sel_152243_comb} + {{1{p1_sel_152244_comb[15]}}, p1_sel_152244_comb};
  assign p1_add_153048_comb = {{1{p1_sel_152245_comb[15]}}, p1_sel_152245_comb} + {{1{p1_sel_152246_comb[15]}}, p1_sel_152246_comb};
  assign p1_add_153049_comb = {{1{p1_sel_152247_comb[15]}}, p1_sel_152247_comb} + {{1{p1_sel_152248_comb[15]}}, p1_sel_152248_comb};
  assign p1_add_153050_comb = {{1{p1_sel_152249_comb[15]}}, p1_sel_152249_comb} + {{1{p1_sel_152250_comb[15]}}, p1_sel_152250_comb};
  assign p1_add_153051_comb = {{1{p1_sel_152251_comb[15]}}, p1_sel_152251_comb} + {{1{p1_sel_152252_comb[15]}}, p1_sel_152252_comb};
  assign p1_add_153052_comb = {{1{p1_sel_152253_comb[15]}}, p1_sel_152253_comb} + {{1{p1_sel_152254_comb[15]}}, p1_sel_152254_comb};
  assign p1_add_153053_comb = {{1{p1_sel_152255_comb[15]}}, p1_sel_152255_comb} + {{1{p1_sel_152256_comb[15]}}, p1_sel_152256_comb};
  assign p1_add_153054_comb = {{1{p1_sel_152257_comb[15]}}, p1_sel_152257_comb} + {{1{p1_sel_152258_comb[15]}}, p1_sel_152258_comb};
  assign p1_add_153055_comb = {{1{p1_sel_152259_comb[15]}}, p1_sel_152259_comb} + {{1{p1_sel_152260_comb[15]}}, p1_sel_152260_comb};
  assign p1_add_153056_comb = {{1{p1_sel_152261_comb[15]}}, p1_sel_152261_comb} + {{1{p1_sel_152262_comb[15]}}, p1_sel_152262_comb};
  assign p1_add_153057_comb = {{1{p1_sel_152263_comb[15]}}, p1_sel_152263_comb} + {{1{p1_sel_152264_comb[15]}}, p1_sel_152264_comb};
  assign p1_add_153058_comb = {{1{p1_sel_152265_comb[15]}}, p1_sel_152265_comb} + {{1{p1_sel_152266_comb[15]}}, p1_sel_152266_comb};
  assign p1_add_153059_comb = {{1{p1_sel_152267_comb[15]}}, p1_sel_152267_comb} + {{1{p1_sel_152268_comb[15]}}, p1_sel_152268_comb};
  assign p1_add_153060_comb = {{1{p1_sel_152269_comb[15]}}, p1_sel_152269_comb} + {{1{p1_sel_152270_comb[15]}}, p1_sel_152270_comb};
  assign p1_add_153061_comb = {{1{p1_sel_152271_comb[15]}}, p1_sel_152271_comb} + {{1{p1_sel_152272_comb[15]}}, p1_sel_152272_comb};
  assign p1_add_153062_comb = {{1{p1_sel_152273_comb[15]}}, p1_sel_152273_comb} + {{1{p1_sel_152274_comb[15]}}, p1_sel_152274_comb};
  assign p1_add_153063_comb = {{1{p1_sel_152275_comb[15]}}, p1_sel_152275_comb} + {{1{p1_sel_152276_comb[15]}}, p1_sel_152276_comb};
  assign p1_add_153064_comb = {{1{p1_sel_152277_comb[15]}}, p1_sel_152277_comb} + {{1{p1_sel_152278_comb[15]}}, p1_sel_152278_comb};
  assign p1_add_153065_comb = {{1{p1_sel_152279_comb[15]}}, p1_sel_152279_comb} + {{1{p1_sel_152280_comb[15]}}, p1_sel_152280_comb};
  assign p1_add_153066_comb = {{1{p1_sel_152281_comb[15]}}, p1_sel_152281_comb} + {{1{p1_sel_152282_comb[15]}}, p1_sel_152282_comb};
  assign p1_add_153067_comb = {{1{p1_sel_152283_comb[15]}}, p1_sel_152283_comb} + {{1{p1_sel_152284_comb[15]}}, p1_sel_152284_comb};
  assign p1_add_153068_comb = {{1{p1_sel_152285_comb[15]}}, p1_sel_152285_comb} + {{1{p1_sel_152286_comb[15]}}, p1_sel_152286_comb};
  assign p1_add_153069_comb = {{1{p1_sel_152287_comb[15]}}, p1_sel_152287_comb} + {{1{p1_sel_152288_comb[15]}}, p1_sel_152288_comb};
  assign p1_add_153070_comb = {{1{p1_sel_152289_comb[15]}}, p1_sel_152289_comb} + {{1{p1_sel_152290_comb[15]}}, p1_sel_152290_comb};
  assign p1_add_153071_comb = {{1{p1_sel_152291_comb[15]}}, p1_sel_152291_comb} + {{1{p1_sel_152292_comb[15]}}, p1_sel_152292_comb};
  assign p1_add_153072_comb = {{1{p1_sel_152293_comb[15]}}, p1_sel_152293_comb} + {{1{p1_sel_152294_comb[15]}}, p1_sel_152294_comb};
  assign p1_add_153073_comb = {{1{p1_sel_152295_comb[15]}}, p1_sel_152295_comb} + {{1{p1_sel_152296_comb[15]}}, p1_sel_152296_comb};
  assign p1_add_153074_comb = {{1{p1_sel_152297_comb[15]}}, p1_sel_152297_comb} + {{1{p1_sel_152298_comb[15]}}, p1_sel_152298_comb};
  assign p1_add_153075_comb = {{1{p1_sel_152299_comb[15]}}, p1_sel_152299_comb} + {{1{p1_sel_152300_comb[15]}}, p1_sel_152300_comb};
  assign p1_add_153076_comb = {{1{p1_sel_152301_comb[15]}}, p1_sel_152301_comb} + {{1{p1_sel_152302_comb[15]}}, p1_sel_152302_comb};
  assign p1_add_153077_comb = {{1{p1_sel_152303_comb[15]}}, p1_sel_152303_comb} + {{1{p1_sel_152304_comb[15]}}, p1_sel_152304_comb};
  assign p1_add_153078_comb = {{1{p1_sel_152305_comb[15]}}, p1_sel_152305_comb} + {{1{p1_sel_152306_comb[15]}}, p1_sel_152306_comb};
  assign p1_add_153079_comb = {{1{p1_sel_152307_comb[15]}}, p1_sel_152307_comb} + {{1{p1_sel_152308_comb[15]}}, p1_sel_152308_comb};
  assign p1_add_153080_comb = {{1{p1_sel_152309_comb[15]}}, p1_sel_152309_comb} + {{1{p1_sel_152310_comb[15]}}, p1_sel_152310_comb};
  assign p1_add_153081_comb = {{1{p1_sel_152311_comb[15]}}, p1_sel_152311_comb} + {{1{p1_sel_152312_comb[15]}}, p1_sel_152312_comb};
  assign p1_add_153082_comb = {{1{p1_sel_152313_comb[15]}}, p1_sel_152313_comb} + {{1{p1_sel_152314_comb[15]}}, p1_sel_152314_comb};
  assign p1_add_153083_comb = {{1{p1_sel_152315_comb[15]}}, p1_sel_152315_comb} + {{1{p1_sel_152316_comb[15]}}, p1_sel_152316_comb};
  assign p1_add_153084_comb = {{1{p1_sel_152317_comb[15]}}, p1_sel_152317_comb} + {{1{p1_sel_152318_comb[15]}}, p1_sel_152318_comb};
  assign p1_add_153085_comb = {{1{p1_sel_152319_comb[15]}}, p1_sel_152319_comb} + {{1{p1_sel_152320_comb[15]}}, p1_sel_152320_comb};
  assign p1_add_153086_comb = {{1{p1_sel_152321_comb[15]}}, p1_sel_152321_comb} + {{1{p1_sel_152322_comb[15]}}, p1_sel_152322_comb};
  assign p1_add_153087_comb = {{1{p1_sel_152323_comb[15]}}, p1_sel_152323_comb} + {{1{p1_sel_152324_comb[15]}}, p1_sel_152324_comb};
  assign p1_add_153088_comb = {{1{p1_sel_152325_comb[15]}}, p1_sel_152325_comb} + {{1{p1_sel_152326_comb[15]}}, p1_sel_152326_comb};
  assign p1_add_153089_comb = {{1{p1_sel_152327_comb[15]}}, p1_sel_152327_comb} + {{1{p1_sel_152328_comb[15]}}, p1_sel_152328_comb};
  assign p1_add_153090_comb = {{1{p1_sel_152329_comb[15]}}, p1_sel_152329_comb} + {{1{p1_sel_152330_comb[15]}}, p1_sel_152330_comb};
  assign p1_add_153091_comb = {{1{p1_sel_152331_comb[15]}}, p1_sel_152331_comb} + {{1{p1_sel_152332_comb[15]}}, p1_sel_152332_comb};
  assign p1_add_153092_comb = {{1{p1_sel_152333_comb[15]}}, p1_sel_152333_comb} + {{1{p1_sel_152334_comb[15]}}, p1_sel_152334_comb};
  assign p1_add_153093_comb = {{1{p1_sel_152335_comb[15]}}, p1_sel_152335_comb} + {{1{p1_sel_152336_comb[15]}}, p1_sel_152336_comb};
  assign p1_add_153094_comb = {{1{p1_sel_152337_comb[15]}}, p1_sel_152337_comb} + {{1{p1_sel_152338_comb[15]}}, p1_sel_152338_comb};
  assign p1_add_153095_comb = {{1{p1_sel_152339_comb[15]}}, p1_sel_152339_comb} + {{1{p1_sel_152340_comb[15]}}, p1_sel_152340_comb};
  assign p1_add_153096_comb = {{1{p1_sel_152341_comb[15]}}, p1_sel_152341_comb} + {{1{p1_sel_152342_comb[15]}}, p1_sel_152342_comb};
  assign p1_add_153097_comb = {{1{p1_sel_152343_comb[15]}}, p1_sel_152343_comb} + {{1{p1_sel_152344_comb[15]}}, p1_sel_152344_comb};
  assign p1_add_153098_comb = {{1{p1_sel_152345_comb[15]}}, p1_sel_152345_comb} + {{1{p1_sel_152346_comb[15]}}, p1_sel_152346_comb};
  assign p1_add_153099_comb = {{1{p1_sel_152347_comb[15]}}, p1_sel_152347_comb} + {{1{p1_sel_152348_comb[15]}}, p1_sel_152348_comb};
  assign p1_add_153100_comb = {{1{p1_sel_152349_comb[15]}}, p1_sel_152349_comb} + {{1{p1_sel_152350_comb[15]}}, p1_sel_152350_comb};
  assign p1_add_153101_comb = {{1{p1_sel_152351_comb[15]}}, p1_sel_152351_comb} + {{1{p1_sel_152352_comb[15]}}, p1_sel_152352_comb};
  assign p1_add_153102_comb = {{1{p1_sel_152353_comb[15]}}, p1_sel_152353_comb} + {{1{p1_sel_152354_comb[15]}}, p1_sel_152354_comb};
  assign p1_add_153103_comb = {{1{p1_sel_152355_comb[15]}}, p1_sel_152355_comb} + {{1{p1_sel_152356_comb[15]}}, p1_sel_152356_comb};
  assign p1_add_153104_comb = {{1{p1_sel_152357_comb[15]}}, p1_sel_152357_comb} + {{1{p1_sel_152358_comb[15]}}, p1_sel_152358_comb};
  assign p1_add_153105_comb = {{1{p1_sel_152359_comb[15]}}, p1_sel_152359_comb} + {{1{p1_sel_152360_comb[15]}}, p1_sel_152360_comb};
  assign p1_add_153106_comb = {{1{p1_sel_152361_comb[15]}}, p1_sel_152361_comb} + {{1{p1_sel_152362_comb[15]}}, p1_sel_152362_comb};
  assign p1_add_153107_comb = {{1{p1_sel_152363_comb[15]}}, p1_sel_152363_comb} + {{1{p1_sel_152364_comb[15]}}, p1_sel_152364_comb};
  assign p1_add_153108_comb = {{1{p1_sel_152365_comb[15]}}, p1_sel_152365_comb} + {{1{p1_sel_152366_comb[15]}}, p1_sel_152366_comb};
  assign p1_add_153109_comb = {{1{p1_sel_152367_comb[15]}}, p1_sel_152367_comb} + {{1{p1_sel_152368_comb[15]}}, p1_sel_152368_comb};
  assign p1_add_153110_comb = {{1{p1_sel_152369_comb[15]}}, p1_sel_152369_comb} + {{1{p1_sel_152370_comb[15]}}, p1_sel_152370_comb};
  assign p1_add_153111_comb = {{1{p1_sel_152371_comb[15]}}, p1_sel_152371_comb} + {{1{p1_sel_152372_comb[15]}}, p1_sel_152372_comb};
  assign p1_add_153112_comb = {{1{p1_sel_152373_comb[15]}}, p1_sel_152373_comb} + {{1{p1_sel_152374_comb[15]}}, p1_sel_152374_comb};
  assign p1_add_153113_comb = {{1{p1_sel_152375_comb[15]}}, p1_sel_152375_comb} + {{1{p1_sel_152376_comb[15]}}, p1_sel_152376_comb};
  assign p1_add_153114_comb = {{1{p1_sel_152377_comb[15]}}, p1_sel_152377_comb} + {{1{p1_sel_152378_comb[15]}}, p1_sel_152378_comb};
  assign p1_add_153115_comb = {{1{p1_sel_152379_comb[15]}}, p1_sel_152379_comb} + {{1{p1_sel_152380_comb[15]}}, p1_sel_152380_comb};
  assign p1_add_153116_comb = {{1{p1_sel_152381_comb[15]}}, p1_sel_152381_comb} + {{1{p1_sel_152382_comb[15]}}, p1_sel_152382_comb};
  assign p1_add_153117_comb = {{1{p1_sel_152383_comb[15]}}, p1_sel_152383_comb} + {{1{p1_sel_152384_comb[15]}}, p1_sel_152384_comb};
  assign p1_add_153118_comb = {{1{p1_sel_152385_comb[15]}}, p1_sel_152385_comb} + {{1{p1_sel_152386_comb[15]}}, p1_sel_152386_comb};
  assign p1_add_153119_comb = {{1{p1_sel_152387_comb[15]}}, p1_sel_152387_comb} + {{1{p1_sel_152388_comb[15]}}, p1_sel_152388_comb};
  assign p1_add_153120_comb = {{1{p1_sel_152389_comb[15]}}, p1_sel_152389_comb} + {{1{p1_sel_152390_comb[15]}}, p1_sel_152390_comb};
  assign p1_add_153121_comb = {{1{p1_sel_152391_comb[15]}}, p1_sel_152391_comb} + {{1{p1_sel_152392_comb[15]}}, p1_sel_152392_comb};
  assign p1_add_153122_comb = {{1{p1_sel_152393_comb[15]}}, p1_sel_152393_comb} + {{1{p1_sel_152394_comb[15]}}, p1_sel_152394_comb};
  assign p1_add_153123_comb = {{1{p1_sel_152395_comb[15]}}, p1_sel_152395_comb} + {{1{p1_sel_152396_comb[15]}}, p1_sel_152396_comb};
  assign p1_add_153124_comb = {{1{p1_sel_152397_comb[15]}}, p1_sel_152397_comb} + {{1{p1_sel_152398_comb[15]}}, p1_sel_152398_comb};
  assign p1_add_153125_comb = {{1{p1_sel_152399_comb[15]}}, p1_sel_152399_comb} + {{1{p1_sel_152400_comb[15]}}, p1_sel_152400_comb};
  assign p1_add_153126_comb = {{1{p1_sel_152401_comb[15]}}, p1_sel_152401_comb} + {{1{p1_sel_152402_comb[15]}}, p1_sel_152402_comb};
  assign p1_add_153127_comb = {{1{p1_sel_152403_comb[15]}}, p1_sel_152403_comb} + {{1{p1_sel_152404_comb[15]}}, p1_sel_152404_comb};
  assign p1_add_153128_comb = {{1{p1_sel_152405_comb[15]}}, p1_sel_152405_comb} + {{1{p1_sel_152406_comb[15]}}, p1_sel_152406_comb};
  assign p1_add_153129_comb = {{1{p1_sel_152407_comb[15]}}, p1_sel_152407_comb} + {{1{p1_sel_152408_comb[15]}}, p1_sel_152408_comb};
  assign p1_add_153130_comb = {{1{p1_sel_152409_comb[15]}}, p1_sel_152409_comb} + {{1{p1_sel_152410_comb[15]}}, p1_sel_152410_comb};
  assign p1_sum__526_comb = p1_sum__524_comb + p1_sum__525_comb;
  assign p1_sum__470_comb = p1_sum__468_comb + p1_sum__469_comb;
  assign p1_sum__414_comb = p1_sum__412_comb + p1_sum__413_comb;
  assign p1_sum__358_comb = p1_sum__356_comb + p1_sum__357_comb;
  assign p1_sum__302_comb = p1_sum__300_comb + p1_sum__301_comb;
  assign p1_sum__246_comb = p1_sum__244_comb + p1_sum__245_comb;
  assign p1_sum__190_comb = p1_sum__188_comb + p1_sum__189_comb;
  assign p1_sum__134_comb = p1_sum__132_comb + p1_sum__133_comb;
  assign p1_sum__1580_comb = {{8{p1_add_152907_comb[16]}}, p1_add_152907_comb};
  assign p1_sum__1581_comb = {{8{p1_add_152908_comb[16]}}, p1_add_152908_comb};
  assign p1_sum__1582_comb = {{8{p1_add_152909_comb[16]}}, p1_add_152909_comb};
  assign p1_sum__1583_comb = {{8{p1_add_152910_comb[16]}}, p1_add_152910_comb};
  assign p1_sum__1552_comb = {{8{p1_add_152911_comb[16]}}, p1_add_152911_comb};
  assign p1_sum__1553_comb = {{8{p1_add_152912_comb[16]}}, p1_add_152912_comb};
  assign p1_sum__1554_comb = {{8{p1_add_152913_comb[16]}}, p1_add_152913_comb};
  assign p1_sum__1555_comb = {{8{p1_add_152914_comb[16]}}, p1_add_152914_comb};
  assign p1_sum__1524_comb = {{8{p1_add_152915_comb[16]}}, p1_add_152915_comb};
  assign p1_sum__1525_comb = {{8{p1_add_152916_comb[16]}}, p1_add_152916_comb};
  assign p1_sum__1526_comb = {{8{p1_add_152917_comb[16]}}, p1_add_152917_comb};
  assign p1_sum__1527_comb = {{8{p1_add_152918_comb[16]}}, p1_add_152918_comb};
  assign p1_sum__1496_comb = {{8{p1_add_152919_comb[16]}}, p1_add_152919_comb};
  assign p1_sum__1497_comb = {{8{p1_add_152920_comb[16]}}, p1_add_152920_comb};
  assign p1_sum__1498_comb = {{8{p1_add_152921_comb[16]}}, p1_add_152921_comb};
  assign p1_sum__1499_comb = {{8{p1_add_152922_comb[16]}}, p1_add_152922_comb};
  assign p1_sum__1468_comb = {{8{p1_add_152923_comb[16]}}, p1_add_152923_comb};
  assign p1_sum__1469_comb = {{8{p1_add_152924_comb[16]}}, p1_add_152924_comb};
  assign p1_sum__1470_comb = {{8{p1_add_152925_comb[16]}}, p1_add_152925_comb};
  assign p1_sum__1471_comb = {{8{p1_add_152926_comb[16]}}, p1_add_152926_comb};
  assign p1_sum__1440_comb = {{8{p1_add_152927_comb[16]}}, p1_add_152927_comb};
  assign p1_sum__1441_comb = {{8{p1_add_152928_comb[16]}}, p1_add_152928_comb};
  assign p1_sum__1442_comb = {{8{p1_add_152929_comb[16]}}, p1_add_152929_comb};
  assign p1_sum__1443_comb = {{8{p1_add_152930_comb[16]}}, p1_add_152930_comb};
  assign p1_sum__1412_comb = {{8{p1_add_152931_comb[16]}}, p1_add_152931_comb};
  assign p1_sum__1413_comb = {{8{p1_add_152932_comb[16]}}, p1_add_152932_comb};
  assign p1_sum__1414_comb = {{8{p1_add_152933_comb[16]}}, p1_add_152933_comb};
  assign p1_sum__1415_comb = {{8{p1_add_152934_comb[16]}}, p1_add_152934_comb};
  assign p1_sum__1384_comb = {{8{p1_add_152935_comb[16]}}, p1_add_152935_comb};
  assign p1_sum__1385_comb = {{8{p1_add_152936_comb[16]}}, p1_add_152936_comb};
  assign p1_sum__1386_comb = {{8{p1_add_152937_comb[16]}}, p1_add_152937_comb};
  assign p1_sum__1387_comb = {{8{p1_add_152938_comb[16]}}, p1_add_152938_comb};
  assign p1_sum__1576_comb = {{8{p1_add_152939_comb[16]}}, p1_add_152939_comb};
  assign p1_sum__1577_comb = {{8{p1_add_152940_comb[16]}}, p1_add_152940_comb};
  assign p1_sum__1578_comb = {{8{p1_add_152941_comb[16]}}, p1_add_152941_comb};
  assign p1_sum__1579_comb = {{8{p1_add_152942_comb[16]}}, p1_add_152942_comb};
  assign p1_sum__1548_comb = {{8{p1_add_152943_comb[16]}}, p1_add_152943_comb};
  assign p1_sum__1549_comb = {{8{p1_add_152944_comb[16]}}, p1_add_152944_comb};
  assign p1_sum__1550_comb = {{8{p1_add_152945_comb[16]}}, p1_add_152945_comb};
  assign p1_sum__1551_comb = {{8{p1_add_152946_comb[16]}}, p1_add_152946_comb};
  assign p1_sum__1520_comb = {{8{p1_add_152947_comb[16]}}, p1_add_152947_comb};
  assign p1_sum__1521_comb = {{8{p1_add_152948_comb[16]}}, p1_add_152948_comb};
  assign p1_sum__1522_comb = {{8{p1_add_152949_comb[16]}}, p1_add_152949_comb};
  assign p1_sum__1523_comb = {{8{p1_add_152950_comb[16]}}, p1_add_152950_comb};
  assign p1_sum__1492_comb = {{8{p1_add_152951_comb[16]}}, p1_add_152951_comb};
  assign p1_sum__1493_comb = {{8{p1_add_152952_comb[16]}}, p1_add_152952_comb};
  assign p1_sum__1494_comb = {{8{p1_add_152953_comb[16]}}, p1_add_152953_comb};
  assign p1_sum__1495_comb = {{8{p1_add_152954_comb[16]}}, p1_add_152954_comb};
  assign p1_sum__1464_comb = {{8{p1_add_152955_comb[16]}}, p1_add_152955_comb};
  assign p1_sum__1465_comb = {{8{p1_add_152956_comb[16]}}, p1_add_152956_comb};
  assign p1_sum__1466_comb = {{8{p1_add_152957_comb[16]}}, p1_add_152957_comb};
  assign p1_sum__1467_comb = {{8{p1_add_152958_comb[16]}}, p1_add_152958_comb};
  assign p1_sum__1436_comb = {{8{p1_add_152959_comb[16]}}, p1_add_152959_comb};
  assign p1_sum__1437_comb = {{8{p1_add_152960_comb[16]}}, p1_add_152960_comb};
  assign p1_sum__1438_comb = {{8{p1_add_152961_comb[16]}}, p1_add_152961_comb};
  assign p1_sum__1439_comb = {{8{p1_add_152962_comb[16]}}, p1_add_152962_comb};
  assign p1_sum__1408_comb = {{8{p1_add_152963_comb[16]}}, p1_add_152963_comb};
  assign p1_sum__1409_comb = {{8{p1_add_152964_comb[16]}}, p1_add_152964_comb};
  assign p1_sum__1410_comb = {{8{p1_add_152965_comb[16]}}, p1_add_152965_comb};
  assign p1_sum__1411_comb = {{8{p1_add_152966_comb[16]}}, p1_add_152966_comb};
  assign p1_sum__1380_comb = {{8{p1_add_152967_comb[16]}}, p1_add_152967_comb};
  assign p1_sum__1381_comb = {{8{p1_add_152968_comb[16]}}, p1_add_152968_comb};
  assign p1_sum__1382_comb = {{8{p1_add_152969_comb[16]}}, p1_add_152969_comb};
  assign p1_sum__1383_comb = {{8{p1_add_152970_comb[16]}}, p1_add_152970_comb};
  assign p1_sum__1572_comb = {{8{p1_add_152971_comb[16]}}, p1_add_152971_comb};
  assign p1_sum__1573_comb = {{8{p1_add_152972_comb[16]}}, p1_add_152972_comb};
  assign p1_sum__1574_comb = {{8{p1_add_152973_comb[16]}}, p1_add_152973_comb};
  assign p1_sum__1575_comb = {{8{p1_add_152974_comb[16]}}, p1_add_152974_comb};
  assign p1_sum__1544_comb = {{8{p1_add_152975_comb[16]}}, p1_add_152975_comb};
  assign p1_sum__1545_comb = {{8{p1_add_152976_comb[16]}}, p1_add_152976_comb};
  assign p1_sum__1546_comb = {{8{p1_add_152977_comb[16]}}, p1_add_152977_comb};
  assign p1_sum__1547_comb = {{8{p1_add_152978_comb[16]}}, p1_add_152978_comb};
  assign p1_sum__1516_comb = {{8{p1_add_152979_comb[16]}}, p1_add_152979_comb};
  assign p1_sum__1517_comb = {{8{p1_add_152980_comb[16]}}, p1_add_152980_comb};
  assign p1_sum__1518_comb = {{8{p1_add_152981_comb[16]}}, p1_add_152981_comb};
  assign p1_sum__1519_comb = {{8{p1_add_152982_comb[16]}}, p1_add_152982_comb};
  assign p1_sum__1488_comb = {{8{p1_add_152983_comb[16]}}, p1_add_152983_comb};
  assign p1_sum__1489_comb = {{8{p1_add_152984_comb[16]}}, p1_add_152984_comb};
  assign p1_sum__1490_comb = {{8{p1_add_152985_comb[16]}}, p1_add_152985_comb};
  assign p1_sum__1491_comb = {{8{p1_add_152986_comb[16]}}, p1_add_152986_comb};
  assign p1_sum__1460_comb = {{8{p1_add_152987_comb[16]}}, p1_add_152987_comb};
  assign p1_sum__1461_comb = {{8{p1_add_152988_comb[16]}}, p1_add_152988_comb};
  assign p1_sum__1462_comb = {{8{p1_add_152989_comb[16]}}, p1_add_152989_comb};
  assign p1_sum__1463_comb = {{8{p1_add_152990_comb[16]}}, p1_add_152990_comb};
  assign p1_sum__1432_comb = {{8{p1_add_152991_comb[16]}}, p1_add_152991_comb};
  assign p1_sum__1433_comb = {{8{p1_add_152992_comb[16]}}, p1_add_152992_comb};
  assign p1_sum__1434_comb = {{8{p1_add_152993_comb[16]}}, p1_add_152993_comb};
  assign p1_sum__1435_comb = {{8{p1_add_152994_comb[16]}}, p1_add_152994_comb};
  assign p1_sum__1404_comb = {{8{p1_add_152995_comb[16]}}, p1_add_152995_comb};
  assign p1_sum__1405_comb = {{8{p1_add_152996_comb[16]}}, p1_add_152996_comb};
  assign p1_sum__1406_comb = {{8{p1_add_152997_comb[16]}}, p1_add_152997_comb};
  assign p1_sum__1407_comb = {{8{p1_add_152998_comb[16]}}, p1_add_152998_comb};
  assign p1_sum__1376_comb = {{8{p1_add_152999_comb[16]}}, p1_add_152999_comb};
  assign p1_sum__1377_comb = {{8{p1_add_153000_comb[16]}}, p1_add_153000_comb};
  assign p1_sum__1378_comb = {{8{p1_add_153001_comb[16]}}, p1_add_153001_comb};
  assign p1_sum__1379_comb = {{8{p1_add_153002_comb[16]}}, p1_add_153002_comb};
  assign p1_sum__1568_comb = {{8{p1_add_153003_comb[16]}}, p1_add_153003_comb};
  assign p1_sum__1569_comb = {{8{p1_add_153004_comb[16]}}, p1_add_153004_comb};
  assign p1_sum__1570_comb = {{8{p1_add_153005_comb[16]}}, p1_add_153005_comb};
  assign p1_sum__1571_comb = {{8{p1_add_153006_comb[16]}}, p1_add_153006_comb};
  assign p1_sum__1540_comb = {{8{p1_add_153007_comb[16]}}, p1_add_153007_comb};
  assign p1_sum__1541_comb = {{8{p1_add_153008_comb[16]}}, p1_add_153008_comb};
  assign p1_sum__1542_comb = {{8{p1_add_153009_comb[16]}}, p1_add_153009_comb};
  assign p1_sum__1543_comb = {{8{p1_add_153010_comb[16]}}, p1_add_153010_comb};
  assign p1_sum__1512_comb = {{8{p1_add_153011_comb[16]}}, p1_add_153011_comb};
  assign p1_sum__1513_comb = {{8{p1_add_153012_comb[16]}}, p1_add_153012_comb};
  assign p1_sum__1514_comb = {{8{p1_add_153013_comb[16]}}, p1_add_153013_comb};
  assign p1_sum__1515_comb = {{8{p1_add_153014_comb[16]}}, p1_add_153014_comb};
  assign p1_sum__1484_comb = {{8{p1_add_153015_comb[16]}}, p1_add_153015_comb};
  assign p1_sum__1485_comb = {{8{p1_add_153016_comb[16]}}, p1_add_153016_comb};
  assign p1_sum__1486_comb = {{8{p1_add_153017_comb[16]}}, p1_add_153017_comb};
  assign p1_sum__1487_comb = {{8{p1_add_153018_comb[16]}}, p1_add_153018_comb};
  assign p1_sum__1456_comb = {{8{p1_add_153019_comb[16]}}, p1_add_153019_comb};
  assign p1_sum__1457_comb = {{8{p1_add_153020_comb[16]}}, p1_add_153020_comb};
  assign p1_sum__1458_comb = {{8{p1_add_153021_comb[16]}}, p1_add_153021_comb};
  assign p1_sum__1459_comb = {{8{p1_add_153022_comb[16]}}, p1_add_153022_comb};
  assign p1_sum__1428_comb = {{8{p1_add_153023_comb[16]}}, p1_add_153023_comb};
  assign p1_sum__1429_comb = {{8{p1_add_153024_comb[16]}}, p1_add_153024_comb};
  assign p1_sum__1430_comb = {{8{p1_add_153025_comb[16]}}, p1_add_153025_comb};
  assign p1_sum__1431_comb = {{8{p1_add_153026_comb[16]}}, p1_add_153026_comb};
  assign p1_sum__1400_comb = {{8{p1_add_153027_comb[16]}}, p1_add_153027_comb};
  assign p1_sum__1401_comb = {{8{p1_add_153028_comb[16]}}, p1_add_153028_comb};
  assign p1_sum__1402_comb = {{8{p1_add_153029_comb[16]}}, p1_add_153029_comb};
  assign p1_sum__1403_comb = {{8{p1_add_153030_comb[16]}}, p1_add_153030_comb};
  assign p1_sum__1372_comb = {{8{p1_add_153031_comb[16]}}, p1_add_153031_comb};
  assign p1_sum__1373_comb = {{8{p1_add_153032_comb[16]}}, p1_add_153032_comb};
  assign p1_sum__1374_comb = {{8{p1_add_153033_comb[16]}}, p1_add_153033_comb};
  assign p1_sum__1375_comb = {{8{p1_add_153034_comb[16]}}, p1_add_153034_comb};
  assign p1_sum__1564_comb = {{8{p1_add_153035_comb[16]}}, p1_add_153035_comb};
  assign p1_sum__1565_comb = {{8{p1_add_153036_comb[16]}}, p1_add_153036_comb};
  assign p1_sum__1566_comb = {{8{p1_add_153037_comb[16]}}, p1_add_153037_comb};
  assign p1_sum__1567_comb = {{8{p1_add_153038_comb[16]}}, p1_add_153038_comb};
  assign p1_sum__1536_comb = {{8{p1_add_153039_comb[16]}}, p1_add_153039_comb};
  assign p1_sum__1537_comb = {{8{p1_add_153040_comb[16]}}, p1_add_153040_comb};
  assign p1_sum__1538_comb = {{8{p1_add_153041_comb[16]}}, p1_add_153041_comb};
  assign p1_sum__1539_comb = {{8{p1_add_153042_comb[16]}}, p1_add_153042_comb};
  assign p1_sum__1508_comb = {{8{p1_add_153043_comb[16]}}, p1_add_153043_comb};
  assign p1_sum__1509_comb = {{8{p1_add_153044_comb[16]}}, p1_add_153044_comb};
  assign p1_sum__1510_comb = {{8{p1_add_153045_comb[16]}}, p1_add_153045_comb};
  assign p1_sum__1511_comb = {{8{p1_add_153046_comb[16]}}, p1_add_153046_comb};
  assign p1_sum__1480_comb = {{8{p1_add_153047_comb[16]}}, p1_add_153047_comb};
  assign p1_sum__1481_comb = {{8{p1_add_153048_comb[16]}}, p1_add_153048_comb};
  assign p1_sum__1482_comb = {{8{p1_add_153049_comb[16]}}, p1_add_153049_comb};
  assign p1_sum__1483_comb = {{8{p1_add_153050_comb[16]}}, p1_add_153050_comb};
  assign p1_sum__1452_comb = {{8{p1_add_153051_comb[16]}}, p1_add_153051_comb};
  assign p1_sum__1453_comb = {{8{p1_add_153052_comb[16]}}, p1_add_153052_comb};
  assign p1_sum__1454_comb = {{8{p1_add_153053_comb[16]}}, p1_add_153053_comb};
  assign p1_sum__1455_comb = {{8{p1_add_153054_comb[16]}}, p1_add_153054_comb};
  assign p1_sum__1424_comb = {{8{p1_add_153055_comb[16]}}, p1_add_153055_comb};
  assign p1_sum__1425_comb = {{8{p1_add_153056_comb[16]}}, p1_add_153056_comb};
  assign p1_sum__1426_comb = {{8{p1_add_153057_comb[16]}}, p1_add_153057_comb};
  assign p1_sum__1427_comb = {{8{p1_add_153058_comb[16]}}, p1_add_153058_comb};
  assign p1_sum__1396_comb = {{8{p1_add_153059_comb[16]}}, p1_add_153059_comb};
  assign p1_sum__1397_comb = {{8{p1_add_153060_comb[16]}}, p1_add_153060_comb};
  assign p1_sum__1398_comb = {{8{p1_add_153061_comb[16]}}, p1_add_153061_comb};
  assign p1_sum__1399_comb = {{8{p1_add_153062_comb[16]}}, p1_add_153062_comb};
  assign p1_sum__1368_comb = {{8{p1_add_153063_comb[16]}}, p1_add_153063_comb};
  assign p1_sum__1369_comb = {{8{p1_add_153064_comb[16]}}, p1_add_153064_comb};
  assign p1_sum__1370_comb = {{8{p1_add_153065_comb[16]}}, p1_add_153065_comb};
  assign p1_sum__1371_comb = {{8{p1_add_153066_comb[16]}}, p1_add_153066_comb};
  assign p1_sum__1560_comb = {{8{p1_add_153067_comb[16]}}, p1_add_153067_comb};
  assign p1_sum__1561_comb = {{8{p1_add_153068_comb[16]}}, p1_add_153068_comb};
  assign p1_sum__1562_comb = {{8{p1_add_153069_comb[16]}}, p1_add_153069_comb};
  assign p1_sum__1563_comb = {{8{p1_add_153070_comb[16]}}, p1_add_153070_comb};
  assign p1_sum__1532_comb = {{8{p1_add_153071_comb[16]}}, p1_add_153071_comb};
  assign p1_sum__1533_comb = {{8{p1_add_153072_comb[16]}}, p1_add_153072_comb};
  assign p1_sum__1534_comb = {{8{p1_add_153073_comb[16]}}, p1_add_153073_comb};
  assign p1_sum__1535_comb = {{8{p1_add_153074_comb[16]}}, p1_add_153074_comb};
  assign p1_sum__1504_comb = {{8{p1_add_153075_comb[16]}}, p1_add_153075_comb};
  assign p1_sum__1505_comb = {{8{p1_add_153076_comb[16]}}, p1_add_153076_comb};
  assign p1_sum__1506_comb = {{8{p1_add_153077_comb[16]}}, p1_add_153077_comb};
  assign p1_sum__1507_comb = {{8{p1_add_153078_comb[16]}}, p1_add_153078_comb};
  assign p1_sum__1476_comb = {{8{p1_add_153079_comb[16]}}, p1_add_153079_comb};
  assign p1_sum__1477_comb = {{8{p1_add_153080_comb[16]}}, p1_add_153080_comb};
  assign p1_sum__1478_comb = {{8{p1_add_153081_comb[16]}}, p1_add_153081_comb};
  assign p1_sum__1479_comb = {{8{p1_add_153082_comb[16]}}, p1_add_153082_comb};
  assign p1_sum__1448_comb = {{8{p1_add_153083_comb[16]}}, p1_add_153083_comb};
  assign p1_sum__1449_comb = {{8{p1_add_153084_comb[16]}}, p1_add_153084_comb};
  assign p1_sum__1450_comb = {{8{p1_add_153085_comb[16]}}, p1_add_153085_comb};
  assign p1_sum__1451_comb = {{8{p1_add_153086_comb[16]}}, p1_add_153086_comb};
  assign p1_sum__1420_comb = {{8{p1_add_153087_comb[16]}}, p1_add_153087_comb};
  assign p1_sum__1421_comb = {{8{p1_add_153088_comb[16]}}, p1_add_153088_comb};
  assign p1_sum__1422_comb = {{8{p1_add_153089_comb[16]}}, p1_add_153089_comb};
  assign p1_sum__1423_comb = {{8{p1_add_153090_comb[16]}}, p1_add_153090_comb};
  assign p1_sum__1392_comb = {{8{p1_add_153091_comb[16]}}, p1_add_153091_comb};
  assign p1_sum__1393_comb = {{8{p1_add_153092_comb[16]}}, p1_add_153092_comb};
  assign p1_sum__1394_comb = {{8{p1_add_153093_comb[16]}}, p1_add_153093_comb};
  assign p1_sum__1395_comb = {{8{p1_add_153094_comb[16]}}, p1_add_153094_comb};
  assign p1_sum__1364_comb = {{8{p1_add_153095_comb[16]}}, p1_add_153095_comb};
  assign p1_sum__1365_comb = {{8{p1_add_153096_comb[16]}}, p1_add_153096_comb};
  assign p1_sum__1366_comb = {{8{p1_add_153097_comb[16]}}, p1_add_153097_comb};
  assign p1_sum__1367_comb = {{8{p1_add_153098_comb[16]}}, p1_add_153098_comb};
  assign p1_sum__1556_comb = {{8{p1_add_153099_comb[16]}}, p1_add_153099_comb};
  assign p1_sum__1557_comb = {{8{p1_add_153100_comb[16]}}, p1_add_153100_comb};
  assign p1_sum__1558_comb = {{8{p1_add_153101_comb[16]}}, p1_add_153101_comb};
  assign p1_sum__1559_comb = {{8{p1_add_153102_comb[16]}}, p1_add_153102_comb};
  assign p1_sum__1528_comb = {{8{p1_add_153103_comb[16]}}, p1_add_153103_comb};
  assign p1_sum__1529_comb = {{8{p1_add_153104_comb[16]}}, p1_add_153104_comb};
  assign p1_sum__1530_comb = {{8{p1_add_153105_comb[16]}}, p1_add_153105_comb};
  assign p1_sum__1531_comb = {{8{p1_add_153106_comb[16]}}, p1_add_153106_comb};
  assign p1_sum__1500_comb = {{8{p1_add_153107_comb[16]}}, p1_add_153107_comb};
  assign p1_sum__1501_comb = {{8{p1_add_153108_comb[16]}}, p1_add_153108_comb};
  assign p1_sum__1502_comb = {{8{p1_add_153109_comb[16]}}, p1_add_153109_comb};
  assign p1_sum__1503_comb = {{8{p1_add_153110_comb[16]}}, p1_add_153110_comb};
  assign p1_sum__1472_comb = {{8{p1_add_153111_comb[16]}}, p1_add_153111_comb};
  assign p1_sum__1473_comb = {{8{p1_add_153112_comb[16]}}, p1_add_153112_comb};
  assign p1_sum__1474_comb = {{8{p1_add_153113_comb[16]}}, p1_add_153113_comb};
  assign p1_sum__1475_comb = {{8{p1_add_153114_comb[16]}}, p1_add_153114_comb};
  assign p1_sum__1444_comb = {{8{p1_add_153115_comb[16]}}, p1_add_153115_comb};
  assign p1_sum__1445_comb = {{8{p1_add_153116_comb[16]}}, p1_add_153116_comb};
  assign p1_sum__1446_comb = {{8{p1_add_153117_comb[16]}}, p1_add_153117_comb};
  assign p1_sum__1447_comb = {{8{p1_add_153118_comb[16]}}, p1_add_153118_comb};
  assign p1_sum__1416_comb = {{8{p1_add_153119_comb[16]}}, p1_add_153119_comb};
  assign p1_sum__1417_comb = {{8{p1_add_153120_comb[16]}}, p1_add_153120_comb};
  assign p1_sum__1418_comb = {{8{p1_add_153121_comb[16]}}, p1_add_153121_comb};
  assign p1_sum__1419_comb = {{8{p1_add_153122_comb[16]}}, p1_add_153122_comb};
  assign p1_sum__1388_comb = {{8{p1_add_153123_comb[16]}}, p1_add_153123_comb};
  assign p1_sum__1389_comb = {{8{p1_add_153124_comb[16]}}, p1_add_153124_comb};
  assign p1_sum__1390_comb = {{8{p1_add_153125_comb[16]}}, p1_add_153125_comb};
  assign p1_sum__1391_comb = {{8{p1_add_153126_comb[16]}}, p1_add_153126_comb};
  assign p1_sum__1360_comb = {{8{p1_add_153127_comb[16]}}, p1_add_153127_comb};
  assign p1_sum__1361_comb = {{8{p1_add_153128_comb[16]}}, p1_add_153128_comb};
  assign p1_sum__1362_comb = {{8{p1_add_153129_comb[16]}}, p1_add_153129_comb};
  assign p1_sum__1363_comb = {{8{p1_add_153130_comb[16]}}, p1_add_153130_comb};
  assign p1_umul_153371_comb = umul32b_32b_x_7b(p1_sum__526_comb, 7'h5b);
  assign p1_umul_153372_comb = umul32b_32b_x_7b(p1_sum__470_comb, 7'h5b);
  assign p1_umul_153373_comb = umul32b_32b_x_7b(p1_sum__414_comb, 7'h5b);
  assign p1_umul_153374_comb = umul32b_32b_x_7b(p1_sum__358_comb, 7'h5b);
  assign p1_umul_153375_comb = umul32b_32b_x_7b(p1_sum__302_comb, 7'h5b);
  assign p1_umul_153376_comb = umul32b_32b_x_7b(p1_sum__246_comb, 7'h5b);
  assign p1_umul_153377_comb = umul32b_32b_x_7b(p1_sum__190_comb, 7'h5b);
  assign p1_umul_153378_comb = umul32b_32b_x_7b(p1_sum__134_comb, 7'h5b);
  assign p1_sum__1246_comb = p1_sum__1580_comb + p1_sum__1581_comb;
  assign p1_sum__1247_comb = p1_sum__1582_comb + p1_sum__1583_comb;
  assign p1_sum__1232_comb = p1_sum__1552_comb + p1_sum__1553_comb;
  assign p1_sum__1233_comb = p1_sum__1554_comb + p1_sum__1555_comb;
  assign p1_sum__1218_comb = p1_sum__1524_comb + p1_sum__1525_comb;
  assign p1_sum__1219_comb = p1_sum__1526_comb + p1_sum__1527_comb;
  assign p1_sum__1204_comb = p1_sum__1496_comb + p1_sum__1497_comb;
  assign p1_sum__1205_comb = p1_sum__1498_comb + p1_sum__1499_comb;
  assign p1_sum__1190_comb = p1_sum__1468_comb + p1_sum__1469_comb;
  assign p1_sum__1191_comb = p1_sum__1470_comb + p1_sum__1471_comb;
  assign p1_sum__1176_comb = p1_sum__1440_comb + p1_sum__1441_comb;
  assign p1_sum__1177_comb = p1_sum__1442_comb + p1_sum__1443_comb;
  assign p1_sum__1162_comb = p1_sum__1412_comb + p1_sum__1413_comb;
  assign p1_sum__1163_comb = p1_sum__1414_comb + p1_sum__1415_comb;
  assign p1_sum__1148_comb = p1_sum__1384_comb + p1_sum__1385_comb;
  assign p1_sum__1149_comb = p1_sum__1386_comb + p1_sum__1387_comb;
  assign p1_sum__1244_comb = p1_sum__1576_comb + p1_sum__1577_comb;
  assign p1_sum__1245_comb = p1_sum__1578_comb + p1_sum__1579_comb;
  assign p1_sum__1230_comb = p1_sum__1548_comb + p1_sum__1549_comb;
  assign p1_sum__1231_comb = p1_sum__1550_comb + p1_sum__1551_comb;
  assign p1_sum__1216_comb = p1_sum__1520_comb + p1_sum__1521_comb;
  assign p1_sum__1217_comb = p1_sum__1522_comb + p1_sum__1523_comb;
  assign p1_sum__1202_comb = p1_sum__1492_comb + p1_sum__1493_comb;
  assign p1_sum__1203_comb = p1_sum__1494_comb + p1_sum__1495_comb;
  assign p1_sum__1188_comb = p1_sum__1464_comb + p1_sum__1465_comb;
  assign p1_sum__1189_comb = p1_sum__1466_comb + p1_sum__1467_comb;
  assign p1_sum__1174_comb = p1_sum__1436_comb + p1_sum__1437_comb;
  assign p1_sum__1175_comb = p1_sum__1438_comb + p1_sum__1439_comb;
  assign p1_sum__1160_comb = p1_sum__1408_comb + p1_sum__1409_comb;
  assign p1_sum__1161_comb = p1_sum__1410_comb + p1_sum__1411_comb;
  assign p1_sum__1146_comb = p1_sum__1380_comb + p1_sum__1381_comb;
  assign p1_sum__1147_comb = p1_sum__1382_comb + p1_sum__1383_comb;
  assign p1_sum__1242_comb = p1_sum__1572_comb + p1_sum__1573_comb;
  assign p1_sum__1243_comb = p1_sum__1574_comb + p1_sum__1575_comb;
  assign p1_sum__1228_comb = p1_sum__1544_comb + p1_sum__1545_comb;
  assign p1_sum__1229_comb = p1_sum__1546_comb + p1_sum__1547_comb;
  assign p1_sum__1214_comb = p1_sum__1516_comb + p1_sum__1517_comb;
  assign p1_sum__1215_comb = p1_sum__1518_comb + p1_sum__1519_comb;
  assign p1_sum__1200_comb = p1_sum__1488_comb + p1_sum__1489_comb;
  assign p1_sum__1201_comb = p1_sum__1490_comb + p1_sum__1491_comb;
  assign p1_sum__1186_comb = p1_sum__1460_comb + p1_sum__1461_comb;
  assign p1_sum__1187_comb = p1_sum__1462_comb + p1_sum__1463_comb;
  assign p1_sum__1172_comb = p1_sum__1432_comb + p1_sum__1433_comb;
  assign p1_sum__1173_comb = p1_sum__1434_comb + p1_sum__1435_comb;
  assign p1_sum__1158_comb = p1_sum__1404_comb + p1_sum__1405_comb;
  assign p1_sum__1159_comb = p1_sum__1406_comb + p1_sum__1407_comb;
  assign p1_sum__1144_comb = p1_sum__1376_comb + p1_sum__1377_comb;
  assign p1_sum__1145_comb = p1_sum__1378_comb + p1_sum__1379_comb;
  assign p1_sum__1240_comb = p1_sum__1568_comb + p1_sum__1569_comb;
  assign p1_sum__1241_comb = p1_sum__1570_comb + p1_sum__1571_comb;
  assign p1_sum__1226_comb = p1_sum__1540_comb + p1_sum__1541_comb;
  assign p1_sum__1227_comb = p1_sum__1542_comb + p1_sum__1543_comb;
  assign p1_sum__1212_comb = p1_sum__1512_comb + p1_sum__1513_comb;
  assign p1_sum__1213_comb = p1_sum__1514_comb + p1_sum__1515_comb;
  assign p1_sum__1198_comb = p1_sum__1484_comb + p1_sum__1485_comb;
  assign p1_sum__1199_comb = p1_sum__1486_comb + p1_sum__1487_comb;
  assign p1_sum__1184_comb = p1_sum__1456_comb + p1_sum__1457_comb;
  assign p1_sum__1185_comb = p1_sum__1458_comb + p1_sum__1459_comb;
  assign p1_sum__1170_comb = p1_sum__1428_comb + p1_sum__1429_comb;
  assign p1_sum__1171_comb = p1_sum__1430_comb + p1_sum__1431_comb;
  assign p1_sum__1156_comb = p1_sum__1400_comb + p1_sum__1401_comb;
  assign p1_sum__1157_comb = p1_sum__1402_comb + p1_sum__1403_comb;
  assign p1_sum__1142_comb = p1_sum__1372_comb + p1_sum__1373_comb;
  assign p1_sum__1143_comb = p1_sum__1374_comb + p1_sum__1375_comb;
  assign p1_sum__1238_comb = p1_sum__1564_comb + p1_sum__1565_comb;
  assign p1_sum__1239_comb = p1_sum__1566_comb + p1_sum__1567_comb;
  assign p1_sum__1224_comb = p1_sum__1536_comb + p1_sum__1537_comb;
  assign p1_sum__1225_comb = p1_sum__1538_comb + p1_sum__1539_comb;
  assign p1_sum__1210_comb = p1_sum__1508_comb + p1_sum__1509_comb;
  assign p1_sum__1211_comb = p1_sum__1510_comb + p1_sum__1511_comb;
  assign p1_sum__1196_comb = p1_sum__1480_comb + p1_sum__1481_comb;
  assign p1_sum__1197_comb = p1_sum__1482_comb + p1_sum__1483_comb;
  assign p1_sum__1182_comb = p1_sum__1452_comb + p1_sum__1453_comb;
  assign p1_sum__1183_comb = p1_sum__1454_comb + p1_sum__1455_comb;
  assign p1_sum__1168_comb = p1_sum__1424_comb + p1_sum__1425_comb;
  assign p1_sum__1169_comb = p1_sum__1426_comb + p1_sum__1427_comb;
  assign p1_sum__1154_comb = p1_sum__1396_comb + p1_sum__1397_comb;
  assign p1_sum__1155_comb = p1_sum__1398_comb + p1_sum__1399_comb;
  assign p1_sum__1140_comb = p1_sum__1368_comb + p1_sum__1369_comb;
  assign p1_sum__1141_comb = p1_sum__1370_comb + p1_sum__1371_comb;
  assign p1_sum__1236_comb = p1_sum__1560_comb + p1_sum__1561_comb;
  assign p1_sum__1237_comb = p1_sum__1562_comb + p1_sum__1563_comb;
  assign p1_sum__1222_comb = p1_sum__1532_comb + p1_sum__1533_comb;
  assign p1_sum__1223_comb = p1_sum__1534_comb + p1_sum__1535_comb;
  assign p1_sum__1208_comb = p1_sum__1504_comb + p1_sum__1505_comb;
  assign p1_sum__1209_comb = p1_sum__1506_comb + p1_sum__1507_comb;
  assign p1_sum__1194_comb = p1_sum__1476_comb + p1_sum__1477_comb;
  assign p1_sum__1195_comb = p1_sum__1478_comb + p1_sum__1479_comb;
  assign p1_sum__1180_comb = p1_sum__1448_comb + p1_sum__1449_comb;
  assign p1_sum__1181_comb = p1_sum__1450_comb + p1_sum__1451_comb;
  assign p1_sum__1166_comb = p1_sum__1420_comb + p1_sum__1421_comb;
  assign p1_sum__1167_comb = p1_sum__1422_comb + p1_sum__1423_comb;
  assign p1_sum__1152_comb = p1_sum__1392_comb + p1_sum__1393_comb;
  assign p1_sum__1153_comb = p1_sum__1394_comb + p1_sum__1395_comb;
  assign p1_sum__1138_comb = p1_sum__1364_comb + p1_sum__1365_comb;
  assign p1_sum__1139_comb = p1_sum__1366_comb + p1_sum__1367_comb;
  assign p1_sum__1234_comb = p1_sum__1556_comb + p1_sum__1557_comb;
  assign p1_sum__1235_comb = p1_sum__1558_comb + p1_sum__1559_comb;
  assign p1_sum__1220_comb = p1_sum__1528_comb + p1_sum__1529_comb;
  assign p1_sum__1221_comb = p1_sum__1530_comb + p1_sum__1531_comb;
  assign p1_sum__1206_comb = p1_sum__1500_comb + p1_sum__1501_comb;
  assign p1_sum__1207_comb = p1_sum__1502_comb + p1_sum__1503_comb;
  assign p1_sum__1192_comb = p1_sum__1472_comb + p1_sum__1473_comb;
  assign p1_sum__1193_comb = p1_sum__1474_comb + p1_sum__1475_comb;
  assign p1_sum__1178_comb = p1_sum__1444_comb + p1_sum__1445_comb;
  assign p1_sum__1179_comb = p1_sum__1446_comb + p1_sum__1447_comb;
  assign p1_sum__1164_comb = p1_sum__1416_comb + p1_sum__1417_comb;
  assign p1_sum__1165_comb = p1_sum__1418_comb + p1_sum__1419_comb;
  assign p1_sum__1150_comb = p1_sum__1388_comb + p1_sum__1389_comb;
  assign p1_sum__1151_comb = p1_sum__1390_comb + p1_sum__1391_comb;
  assign p1_sum__1136_comb = p1_sum__1360_comb + p1_sum__1361_comb;
  assign p1_sum__1137_comb = p1_sum__1362_comb + p1_sum__1363_comb;
  assign p1_sum__1079_comb = p1_sum__1246_comb + p1_sum__1247_comb;
  assign p1_sum__1072_comb = p1_sum__1232_comb + p1_sum__1233_comb;
  assign p1_sum__1065_comb = p1_sum__1218_comb + p1_sum__1219_comb;
  assign p1_sum__1058_comb = p1_sum__1204_comb + p1_sum__1205_comb;
  assign p1_sum__1051_comb = p1_sum__1190_comb + p1_sum__1191_comb;
  assign p1_sum__1044_comb = p1_sum__1176_comb + p1_sum__1177_comb;
  assign p1_sum__1037_comb = p1_sum__1162_comb + p1_sum__1163_comb;
  assign p1_sum__1030_comb = p1_sum__1148_comb + p1_sum__1149_comb;
  assign p1_sum__1078_comb = p1_sum__1244_comb + p1_sum__1245_comb;
  assign p1_sum__1071_comb = p1_sum__1230_comb + p1_sum__1231_comb;
  assign p1_sum__1064_comb = p1_sum__1216_comb + p1_sum__1217_comb;
  assign p1_sum__1057_comb = p1_sum__1202_comb + p1_sum__1203_comb;
  assign p1_sum__1050_comb = p1_sum__1188_comb + p1_sum__1189_comb;
  assign p1_sum__1043_comb = p1_sum__1174_comb + p1_sum__1175_comb;
  assign p1_sum__1036_comb = p1_sum__1160_comb + p1_sum__1161_comb;
  assign p1_sum__1029_comb = p1_sum__1146_comb + p1_sum__1147_comb;
  assign p1_sum__1077_comb = p1_sum__1242_comb + p1_sum__1243_comb;
  assign p1_sum__1070_comb = p1_sum__1228_comb + p1_sum__1229_comb;
  assign p1_sum__1063_comb = p1_sum__1214_comb + p1_sum__1215_comb;
  assign p1_sum__1056_comb = p1_sum__1200_comb + p1_sum__1201_comb;
  assign p1_sum__1049_comb = p1_sum__1186_comb + p1_sum__1187_comb;
  assign p1_sum__1042_comb = p1_sum__1172_comb + p1_sum__1173_comb;
  assign p1_sum__1035_comb = p1_sum__1158_comb + p1_sum__1159_comb;
  assign p1_sum__1028_comb = p1_sum__1144_comb + p1_sum__1145_comb;
  assign p1_sum__1076_comb = p1_sum__1240_comb + p1_sum__1241_comb;
  assign p1_sum__1069_comb = p1_sum__1226_comb + p1_sum__1227_comb;
  assign p1_sum__1062_comb = p1_sum__1212_comb + p1_sum__1213_comb;
  assign p1_sum__1055_comb = p1_sum__1198_comb + p1_sum__1199_comb;
  assign p1_sum__1048_comb = p1_sum__1184_comb + p1_sum__1185_comb;
  assign p1_sum__1041_comb = p1_sum__1170_comb + p1_sum__1171_comb;
  assign p1_sum__1034_comb = p1_sum__1156_comb + p1_sum__1157_comb;
  assign p1_sum__1027_comb = p1_sum__1142_comb + p1_sum__1143_comb;
  assign p1_sum__1075_comb = p1_sum__1238_comb + p1_sum__1239_comb;
  assign p1_sum__1068_comb = p1_sum__1224_comb + p1_sum__1225_comb;
  assign p1_sum__1061_comb = p1_sum__1210_comb + p1_sum__1211_comb;
  assign p1_sum__1054_comb = p1_sum__1196_comb + p1_sum__1197_comb;
  assign p1_sum__1047_comb = p1_sum__1182_comb + p1_sum__1183_comb;
  assign p1_sum__1040_comb = p1_sum__1168_comb + p1_sum__1169_comb;
  assign p1_sum__1033_comb = p1_sum__1154_comb + p1_sum__1155_comb;
  assign p1_sum__1026_comb = p1_sum__1140_comb + p1_sum__1141_comb;
  assign p1_sum__1074_comb = p1_sum__1236_comb + p1_sum__1237_comb;
  assign p1_sum__1067_comb = p1_sum__1222_comb + p1_sum__1223_comb;
  assign p1_sum__1060_comb = p1_sum__1208_comb + p1_sum__1209_comb;
  assign p1_sum__1053_comb = p1_sum__1194_comb + p1_sum__1195_comb;
  assign p1_sum__1046_comb = p1_sum__1180_comb + p1_sum__1181_comb;
  assign p1_sum__1039_comb = p1_sum__1166_comb + p1_sum__1167_comb;
  assign p1_sum__1032_comb = p1_sum__1152_comb + p1_sum__1153_comb;
  assign p1_sum__1025_comb = p1_sum__1138_comb + p1_sum__1139_comb;
  assign p1_sum__1073_comb = p1_sum__1234_comb + p1_sum__1235_comb;
  assign p1_sum__1066_comb = p1_sum__1220_comb + p1_sum__1221_comb;
  assign p1_sum__1059_comb = p1_sum__1206_comb + p1_sum__1207_comb;
  assign p1_sum__1052_comb = p1_sum__1192_comb + p1_sum__1193_comb;
  assign p1_sum__1045_comb = p1_sum__1178_comb + p1_sum__1179_comb;
  assign p1_sum__1038_comb = p1_sum__1164_comb + p1_sum__1165_comb;
  assign p1_sum__1031_comb = p1_sum__1150_comb + p1_sum__1151_comb;
  assign p1_sum__1024_comb = p1_sum__1136_comb + p1_sum__1137_comb;
  assign p1_add_153619_comb = p1_umul_153371_comb[31:7] + 25'h000_0001;
  assign p1_add_153620_comb = p1_umul_153372_comb[31:7] + 25'h000_0001;
  assign p1_add_153621_comb = p1_umul_153373_comb[31:7] + 25'h000_0001;
  assign p1_add_153622_comb = p1_umul_153374_comb[31:7] + 25'h000_0001;
  assign p1_add_153623_comb = p1_umul_153375_comb[31:7] + 25'h000_0001;
  assign p1_add_153624_comb = p1_umul_153376_comb[31:7] + 25'h000_0001;
  assign p1_add_153625_comb = p1_umul_153377_comb[31:7] + 25'h000_0001;
  assign p1_add_153626_comb = p1_umul_153378_comb[31:7] + 25'h000_0001;
  assign p1_add_153627_comb = p1_sum__1079_comb + 25'h000_0001;
  assign p1_add_153628_comb = p1_sum__1072_comb + 25'h000_0001;
  assign p1_add_153629_comb = p1_sum__1065_comb + 25'h000_0001;
  assign p1_add_153630_comb = p1_sum__1058_comb + 25'h000_0001;
  assign p1_add_153631_comb = p1_sum__1051_comb + 25'h000_0001;
  assign p1_add_153632_comb = p1_sum__1044_comb + 25'h000_0001;
  assign p1_add_153633_comb = p1_sum__1037_comb + 25'h000_0001;
  assign p1_add_153634_comb = p1_sum__1030_comb + 25'h000_0001;
  assign p1_add_153635_comb = p1_sum__1078_comb + 25'h000_0001;
  assign p1_add_153636_comb = p1_sum__1071_comb + 25'h000_0001;
  assign p1_add_153637_comb = p1_sum__1064_comb + 25'h000_0001;
  assign p1_add_153638_comb = p1_sum__1057_comb + 25'h000_0001;
  assign p1_add_153639_comb = p1_sum__1050_comb + 25'h000_0001;
  assign p1_add_153640_comb = p1_sum__1043_comb + 25'h000_0001;
  assign p1_add_153641_comb = p1_sum__1036_comb + 25'h000_0001;
  assign p1_add_153642_comb = p1_sum__1029_comb + 25'h000_0001;
  assign p1_add_153643_comb = p1_sum__1077_comb + 25'h000_0001;
  assign p1_add_153644_comb = p1_sum__1070_comb + 25'h000_0001;
  assign p1_add_153645_comb = p1_sum__1063_comb + 25'h000_0001;
  assign p1_add_153646_comb = p1_sum__1056_comb + 25'h000_0001;
  assign p1_add_153647_comb = p1_sum__1049_comb + 25'h000_0001;
  assign p1_add_153648_comb = p1_sum__1042_comb + 25'h000_0001;
  assign p1_add_153649_comb = p1_sum__1035_comb + 25'h000_0001;
  assign p1_add_153650_comb = p1_sum__1028_comb + 25'h000_0001;
  assign p1_add_153651_comb = p1_sum__1076_comb + 25'h000_0001;
  assign p1_add_153652_comb = p1_sum__1069_comb + 25'h000_0001;
  assign p1_add_153653_comb = p1_sum__1062_comb + 25'h000_0001;
  assign p1_add_153654_comb = p1_sum__1055_comb + 25'h000_0001;
  assign p1_add_153655_comb = p1_sum__1048_comb + 25'h000_0001;
  assign p1_add_153656_comb = p1_sum__1041_comb + 25'h000_0001;
  assign p1_add_153657_comb = p1_sum__1034_comb + 25'h000_0001;
  assign p1_add_153658_comb = p1_sum__1027_comb + 25'h000_0001;
  assign p1_add_153659_comb = p1_sum__1075_comb + 25'h000_0001;
  assign p1_add_153660_comb = p1_sum__1068_comb + 25'h000_0001;
  assign p1_add_153661_comb = p1_sum__1061_comb + 25'h000_0001;
  assign p1_add_153662_comb = p1_sum__1054_comb + 25'h000_0001;
  assign p1_add_153663_comb = p1_sum__1047_comb + 25'h000_0001;
  assign p1_add_153664_comb = p1_sum__1040_comb + 25'h000_0001;
  assign p1_add_153665_comb = p1_sum__1033_comb + 25'h000_0001;
  assign p1_add_153666_comb = p1_sum__1026_comb + 25'h000_0001;
  assign p1_add_153667_comb = p1_sum__1074_comb + 25'h000_0001;
  assign p1_add_153668_comb = p1_sum__1067_comb + 25'h000_0001;
  assign p1_add_153669_comb = p1_sum__1060_comb + 25'h000_0001;
  assign p1_add_153670_comb = p1_sum__1053_comb + 25'h000_0001;
  assign p1_add_153671_comb = p1_sum__1046_comb + 25'h000_0001;
  assign p1_add_153672_comb = p1_sum__1039_comb + 25'h000_0001;
  assign p1_add_153673_comb = p1_sum__1032_comb + 25'h000_0001;
  assign p1_add_153674_comb = p1_sum__1025_comb + 25'h000_0001;
  assign p1_add_153675_comb = p1_sum__1073_comb + 25'h000_0001;
  assign p1_add_153676_comb = p1_sum__1066_comb + 25'h000_0001;
  assign p1_add_153677_comb = p1_sum__1059_comb + 25'h000_0001;
  assign p1_add_153678_comb = p1_sum__1052_comb + 25'h000_0001;
  assign p1_add_153679_comb = p1_sum__1045_comb + 25'h000_0001;
  assign p1_add_153680_comb = p1_sum__1038_comb + 25'h000_0001;
  assign p1_add_153681_comb = p1_sum__1031_comb + 25'h000_0001;
  assign p1_add_153682_comb = p1_sum__1024_comb + 25'h000_0001;
  assign p1_clipped__320_comb = $signed(p1_add_153619_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153619_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153619_comb[16:8]);
  assign p1_clipped__321_comb = $signed(p1_add_153620_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153620_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153620_comb[16:8]);
  assign p1_clipped__322_comb = $signed(p1_add_153621_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153621_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153621_comb[16:8]);
  assign p1_clipped__323_comb = $signed(p1_add_153622_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153622_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153622_comb[16:8]);
  assign p1_clipped__324_comb = $signed(p1_add_153623_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153623_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153623_comb[16:8]);
  assign p1_clipped__325_comb = $signed(p1_add_153624_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153624_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153624_comb[16:8]);
  assign p1_clipped__326_comb = $signed(p1_add_153625_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153625_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153625_comb[16:8]);
  assign p1_clipped__327_comb = $signed(p1_add_153626_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153626_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153626_comb[16:8]);
  assign p1_clipped__328_comb = $signed(p1_add_153627_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153627_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153627_comb[16:8]);
  assign p1_clipped__329_comb = $signed(p1_add_153628_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153628_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153628_comb[16:8]);
  assign p1_clipped__330_comb = $signed(p1_add_153629_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153629_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153629_comb[16:8]);
  assign p1_clipped__331_comb = $signed(p1_add_153630_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153630_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153630_comb[16:8]);
  assign p1_clipped__332_comb = $signed(p1_add_153631_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153631_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153631_comb[16:8]);
  assign p1_clipped__333_comb = $signed(p1_add_153632_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153632_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153632_comb[16:8]);
  assign p1_clipped__334_comb = $signed(p1_add_153633_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153633_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153633_comb[16:8]);
  assign p1_clipped__335_comb = $signed(p1_add_153634_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153634_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153634_comb[16:8]);
  assign p1_clipped__336_comb = $signed(p1_add_153635_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153635_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153635_comb[16:8]);
  assign p1_clipped__337_comb = $signed(p1_add_153636_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153636_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153636_comb[16:8]);
  assign p1_clipped__338_comb = $signed(p1_add_153637_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153637_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153637_comb[16:8]);
  assign p1_clipped__339_comb = $signed(p1_add_153638_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153638_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153638_comb[16:8]);
  assign p1_clipped__340_comb = $signed(p1_add_153639_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153639_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153639_comb[16:8]);
  assign p1_clipped__341_comb = $signed(p1_add_153640_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153640_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153640_comb[16:8]);
  assign p1_clipped__342_comb = $signed(p1_add_153641_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153641_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153641_comb[16:8]);
  assign p1_clipped__343_comb = $signed(p1_add_153642_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153642_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153642_comb[16:8]);
  assign p1_clipped__344_comb = $signed(p1_add_153643_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153643_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153643_comb[16:8]);
  assign p1_clipped__345_comb = $signed(p1_add_153644_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153644_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153644_comb[16:8]);
  assign p1_clipped__346_comb = $signed(p1_add_153645_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153645_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153645_comb[16:8]);
  assign p1_clipped__347_comb = $signed(p1_add_153646_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153646_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153646_comb[16:8]);
  assign p1_clipped__348_comb = $signed(p1_add_153647_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153647_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153647_comb[16:8]);
  assign p1_clipped__349_comb = $signed(p1_add_153648_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153648_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153648_comb[16:8]);
  assign p1_clipped__350_comb = $signed(p1_add_153649_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153649_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153649_comb[16:8]);
  assign p1_clipped__351_comb = $signed(p1_add_153650_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153650_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153650_comb[16:8]);
  assign p1_clipped__352_comb = $signed(p1_add_153651_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153651_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153651_comb[16:8]);
  assign p1_clipped__353_comb = $signed(p1_add_153652_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153652_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153652_comb[16:8]);
  assign p1_clipped__354_comb = $signed(p1_add_153653_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153653_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153653_comb[16:8]);
  assign p1_clipped__355_comb = $signed(p1_add_153654_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153654_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153654_comb[16:8]);
  assign p1_clipped__356_comb = $signed(p1_add_153655_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153655_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153655_comb[16:8]);
  assign p1_clipped__357_comb = $signed(p1_add_153656_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153656_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153656_comb[16:8]);
  assign p1_clipped__358_comb = $signed(p1_add_153657_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153657_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153657_comb[16:8]);
  assign p1_clipped__359_comb = $signed(p1_add_153658_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153658_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153658_comb[16:8]);
  assign p1_clipped__360_comb = $signed(p1_add_153659_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153659_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153659_comb[16:8]);
  assign p1_clipped__361_comb = $signed(p1_add_153660_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153660_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153660_comb[16:8]);
  assign p1_clipped__362_comb = $signed(p1_add_153661_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153661_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153661_comb[16:8]);
  assign p1_clipped__363_comb = $signed(p1_add_153662_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153662_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153662_comb[16:8]);
  assign p1_clipped__364_comb = $signed(p1_add_153663_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153663_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153663_comb[16:8]);
  assign p1_clipped__365_comb = $signed(p1_add_153664_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153664_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153664_comb[16:8]);
  assign p1_clipped__366_comb = $signed(p1_add_153665_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153665_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153665_comb[16:8]);
  assign p1_clipped__367_comb = $signed(p1_add_153666_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153666_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153666_comb[16:8]);
  assign p1_clipped__368_comb = $signed(p1_add_153667_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153667_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153667_comb[16:8]);
  assign p1_clipped__369_comb = $signed(p1_add_153668_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153668_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153668_comb[16:8]);
  assign p1_clipped__370_comb = $signed(p1_add_153669_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153669_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153669_comb[16:8]);
  assign p1_clipped__371_comb = $signed(p1_add_153670_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153670_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153670_comb[16:8]);
  assign p1_clipped__372_comb = $signed(p1_add_153671_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153671_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153671_comb[16:8]);
  assign p1_clipped__373_comb = $signed(p1_add_153672_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153672_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153672_comb[16:8]);
  assign p1_clipped__374_comb = $signed(p1_add_153673_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153673_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153673_comb[16:8]);
  assign p1_clipped__375_comb = $signed(p1_add_153674_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153674_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153674_comb[16:8]);
  assign p1_clipped__376_comb = $signed(p1_add_153675_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153675_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153675_comb[16:8]);
  assign p1_clipped__377_comb = $signed(p1_add_153676_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153676_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153676_comb[16:8]);
  assign p1_clipped__378_comb = $signed(p1_add_153677_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153677_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153677_comb[16:8]);
  assign p1_clipped__379_comb = $signed(p1_add_153678_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153678_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153678_comb[16:8]);
  assign p1_clipped__380_comb = $signed(p1_add_153679_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153679_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153679_comb[16:8]);
  assign p1_clipped__381_comb = $signed(p1_add_153680_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153680_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153680_comb[16:8]);
  assign p1_clipped__382_comb = $signed(p1_add_153681_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153681_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153681_comb[16:8]);
  assign p1_clipped__383_comb = $signed(p1_add_153682_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p1_add_153682_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p1_add_153682_comb[16:8]);
  assign p1_add_154451_comb = {{1{p1_clipped__320_comb[8]}}, p1_clipped__320_comb} + 10'h001;
  assign p1_add_154452_comb = {{1{p1_clipped__321_comb[8]}}, p1_clipped__321_comb} + 10'h001;
  assign p1_add_154453_comb = {{1{p1_clipped__322_comb[8]}}, p1_clipped__322_comb} + 10'h001;
  assign p1_add_154454_comb = {{1{p1_clipped__323_comb[8]}}, p1_clipped__323_comb} + 10'h001;
  assign p1_add_154455_comb = {{1{p1_clipped__324_comb[8]}}, p1_clipped__324_comb} + 10'h001;
  assign p1_add_154456_comb = {{1{p1_clipped__325_comb[8]}}, p1_clipped__325_comb} + 10'h001;
  assign p1_add_154457_comb = {{1{p1_clipped__326_comb[8]}}, p1_clipped__326_comb} + 10'h001;
  assign p1_add_154458_comb = {{1{p1_clipped__327_comb[8]}}, p1_clipped__327_comb} + 10'h001;
  assign p1_add_154459_comb = {{1{p1_clipped__328_comb[8]}}, p1_clipped__328_comb} + 10'h001;
  assign p1_add_154460_comb = {{1{p1_clipped__329_comb[8]}}, p1_clipped__329_comb} + 10'h001;
  assign p1_add_154461_comb = {{1{p1_clipped__330_comb[8]}}, p1_clipped__330_comb} + 10'h001;
  assign p1_add_154462_comb = {{1{p1_clipped__331_comb[8]}}, p1_clipped__331_comb} + 10'h001;
  assign p1_add_154463_comb = {{1{p1_clipped__332_comb[8]}}, p1_clipped__332_comb} + 10'h001;
  assign p1_add_154464_comb = {{1{p1_clipped__333_comb[8]}}, p1_clipped__333_comb} + 10'h001;
  assign p1_add_154465_comb = {{1{p1_clipped__334_comb[8]}}, p1_clipped__334_comb} + 10'h001;
  assign p1_add_154466_comb = {{1{p1_clipped__335_comb[8]}}, p1_clipped__335_comb} + 10'h001;
  assign p1_add_154467_comb = {{1{p1_clipped__336_comb[8]}}, p1_clipped__336_comb} + 10'h001;
  assign p1_add_154468_comb = {{1{p1_clipped__337_comb[8]}}, p1_clipped__337_comb} + 10'h001;
  assign p1_add_154469_comb = {{1{p1_clipped__338_comb[8]}}, p1_clipped__338_comb} + 10'h001;
  assign p1_add_154470_comb = {{1{p1_clipped__339_comb[8]}}, p1_clipped__339_comb} + 10'h001;
  assign p1_add_154471_comb = {{1{p1_clipped__340_comb[8]}}, p1_clipped__340_comb} + 10'h001;
  assign p1_add_154472_comb = {{1{p1_clipped__341_comb[8]}}, p1_clipped__341_comb} + 10'h001;
  assign p1_add_154473_comb = {{1{p1_clipped__342_comb[8]}}, p1_clipped__342_comb} + 10'h001;
  assign p1_add_154474_comb = {{1{p1_clipped__343_comb[8]}}, p1_clipped__343_comb} + 10'h001;
  assign p1_add_154475_comb = {{1{p1_clipped__344_comb[8]}}, p1_clipped__344_comb} + 10'h001;
  assign p1_add_154476_comb = {{1{p1_clipped__345_comb[8]}}, p1_clipped__345_comb} + 10'h001;
  assign p1_add_154477_comb = {{1{p1_clipped__346_comb[8]}}, p1_clipped__346_comb} + 10'h001;
  assign p1_add_154478_comb = {{1{p1_clipped__347_comb[8]}}, p1_clipped__347_comb} + 10'h001;
  assign p1_add_154479_comb = {{1{p1_clipped__348_comb[8]}}, p1_clipped__348_comb} + 10'h001;
  assign p1_add_154480_comb = {{1{p1_clipped__349_comb[8]}}, p1_clipped__349_comb} + 10'h001;
  assign p1_add_154481_comb = {{1{p1_clipped__350_comb[8]}}, p1_clipped__350_comb} + 10'h001;
  assign p1_add_154482_comb = {{1{p1_clipped__351_comb[8]}}, p1_clipped__351_comb} + 10'h001;
  assign p1_add_154483_comb = {{1{p1_clipped__352_comb[8]}}, p1_clipped__352_comb} + 10'h001;
  assign p1_add_154484_comb = {{1{p1_clipped__353_comb[8]}}, p1_clipped__353_comb} + 10'h001;
  assign p1_add_154485_comb = {{1{p1_clipped__354_comb[8]}}, p1_clipped__354_comb} + 10'h001;
  assign p1_add_154486_comb = {{1{p1_clipped__355_comb[8]}}, p1_clipped__355_comb} + 10'h001;
  assign p1_add_154487_comb = {{1{p1_clipped__356_comb[8]}}, p1_clipped__356_comb} + 10'h001;
  assign p1_add_154488_comb = {{1{p1_clipped__357_comb[8]}}, p1_clipped__357_comb} + 10'h001;
  assign p1_add_154489_comb = {{1{p1_clipped__358_comb[8]}}, p1_clipped__358_comb} + 10'h001;
  assign p1_add_154490_comb = {{1{p1_clipped__359_comb[8]}}, p1_clipped__359_comb} + 10'h001;
  assign p1_add_154491_comb = {{1{p1_clipped__360_comb[8]}}, p1_clipped__360_comb} + 10'h001;
  assign p1_add_154492_comb = {{1{p1_clipped__361_comb[8]}}, p1_clipped__361_comb} + 10'h001;
  assign p1_add_154493_comb = {{1{p1_clipped__362_comb[8]}}, p1_clipped__362_comb} + 10'h001;
  assign p1_add_154494_comb = {{1{p1_clipped__363_comb[8]}}, p1_clipped__363_comb} + 10'h001;
  assign p1_add_154495_comb = {{1{p1_clipped__364_comb[8]}}, p1_clipped__364_comb} + 10'h001;
  assign p1_add_154496_comb = {{1{p1_clipped__365_comb[8]}}, p1_clipped__365_comb} + 10'h001;
  assign p1_add_154497_comb = {{1{p1_clipped__366_comb[8]}}, p1_clipped__366_comb} + 10'h001;
  assign p1_add_154498_comb = {{1{p1_clipped__367_comb[8]}}, p1_clipped__367_comb} + 10'h001;
  assign p1_add_154499_comb = {{1{p1_clipped__368_comb[8]}}, p1_clipped__368_comb} + 10'h001;
  assign p1_add_154500_comb = {{1{p1_clipped__369_comb[8]}}, p1_clipped__369_comb} + 10'h001;
  assign p1_add_154501_comb = {{1{p1_clipped__370_comb[8]}}, p1_clipped__370_comb} + 10'h001;
  assign p1_add_154502_comb = {{1{p1_clipped__371_comb[8]}}, p1_clipped__371_comb} + 10'h001;
  assign p1_add_154503_comb = {{1{p1_clipped__372_comb[8]}}, p1_clipped__372_comb} + 10'h001;
  assign p1_add_154504_comb = {{1{p1_clipped__373_comb[8]}}, p1_clipped__373_comb} + 10'h001;
  assign p1_add_154505_comb = {{1{p1_clipped__374_comb[8]}}, p1_clipped__374_comb} + 10'h001;
  assign p1_add_154506_comb = {{1{p1_clipped__375_comb[8]}}, p1_clipped__375_comb} + 10'h001;
  assign p1_add_154507_comb = {{1{p1_clipped__376_comb[8]}}, p1_clipped__376_comb} + 10'h001;
  assign p1_add_154508_comb = {{1{p1_clipped__377_comb[8]}}, p1_clipped__377_comb} + 10'h001;
  assign p1_add_154509_comb = {{1{p1_clipped__378_comb[8]}}, p1_clipped__378_comb} + 10'h001;
  assign p1_add_154510_comb = {{1{p1_clipped__379_comb[8]}}, p1_clipped__379_comb} + 10'h001;
  assign p1_add_154511_comb = {{1{p1_clipped__380_comb[8]}}, p1_clipped__380_comb} + 10'h001;
  assign p1_add_154512_comb = {{1{p1_clipped__381_comb[8]}}, p1_clipped__381_comb} + 10'h001;
  assign p1_add_154513_comb = {{1{p1_clipped__382_comb[8]}}, p1_clipped__382_comb} + 10'h001;
  assign p1_add_154514_comb = {{1{p1_clipped__383_comb[8]}}, p1_clipped__383_comb} + 10'h001;
  assign p1_bit_slice_154515_comb = p1_add_154451_comb[9:8];
  assign p1_bit_slice_154516_comb = p1_add_154452_comb[9:8];
  assign p1_bit_slice_154517_comb = p1_add_154453_comb[9:8];
  assign p1_bit_slice_154518_comb = p1_add_154454_comb[9:8];
  assign p1_bit_slice_154519_comb = p1_add_154455_comb[9:8];
  assign p1_bit_slice_154520_comb = p1_add_154456_comb[9:8];
  assign p1_bit_slice_154521_comb = p1_add_154457_comb[9:8];
  assign p1_bit_slice_154522_comb = p1_add_154458_comb[9:8];
  assign p1_bit_slice_154523_comb = p1_add_154459_comb[9:8];
  assign p1_bit_slice_154524_comb = p1_add_154460_comb[9:8];
  assign p1_bit_slice_154525_comb = p1_add_154461_comb[9:8];
  assign p1_bit_slice_154526_comb = p1_add_154462_comb[9:8];
  assign p1_bit_slice_154527_comb = p1_add_154463_comb[9:8];
  assign p1_bit_slice_154528_comb = p1_add_154464_comb[9:8];
  assign p1_bit_slice_154529_comb = p1_add_154465_comb[9:8];
  assign p1_bit_slice_154530_comb = p1_add_154466_comb[9:8];
  assign p1_bit_slice_154531_comb = p1_add_154467_comb[9:8];
  assign p1_bit_slice_154532_comb = p1_add_154468_comb[9:8];
  assign p1_bit_slice_154533_comb = p1_add_154469_comb[9:8];
  assign p1_bit_slice_154534_comb = p1_add_154470_comb[9:8];
  assign p1_bit_slice_154535_comb = p1_add_154471_comb[9:8];
  assign p1_bit_slice_154536_comb = p1_add_154472_comb[9:8];
  assign p1_bit_slice_154537_comb = p1_add_154473_comb[9:8];
  assign p1_bit_slice_154538_comb = p1_add_154474_comb[9:8];
  assign p1_bit_slice_154539_comb = p1_add_154475_comb[9:8];
  assign p1_bit_slice_154540_comb = p1_add_154476_comb[9:8];
  assign p1_bit_slice_154541_comb = p1_add_154477_comb[9:8];
  assign p1_bit_slice_154542_comb = p1_add_154478_comb[9:8];
  assign p1_bit_slice_154543_comb = p1_add_154479_comb[9:8];
  assign p1_bit_slice_154544_comb = p1_add_154480_comb[9:8];
  assign p1_bit_slice_154545_comb = p1_add_154481_comb[9:8];
  assign p1_bit_slice_154546_comb = p1_add_154482_comb[9:8];
  assign p1_bit_slice_154547_comb = p1_add_154483_comb[9:8];
  assign p1_bit_slice_154548_comb = p1_add_154484_comb[9:8];
  assign p1_bit_slice_154549_comb = p1_add_154485_comb[9:8];
  assign p1_bit_slice_154550_comb = p1_add_154486_comb[9:8];
  assign p1_bit_slice_154551_comb = p1_add_154487_comb[9:8];
  assign p1_bit_slice_154552_comb = p1_add_154488_comb[9:8];
  assign p1_bit_slice_154553_comb = p1_add_154489_comb[9:8];
  assign p1_bit_slice_154554_comb = p1_add_154490_comb[9:8];
  assign p1_bit_slice_154555_comb = p1_add_154491_comb[9:8];
  assign p1_bit_slice_154556_comb = p1_add_154492_comb[9:8];
  assign p1_bit_slice_154557_comb = p1_add_154493_comb[9:8];
  assign p1_bit_slice_154558_comb = p1_add_154494_comb[9:8];
  assign p1_bit_slice_154559_comb = p1_add_154495_comb[9:8];
  assign p1_bit_slice_154560_comb = p1_add_154496_comb[9:8];
  assign p1_bit_slice_154561_comb = p1_add_154497_comb[9:8];
  assign p1_bit_slice_154562_comb = p1_add_154498_comb[9:8];
  assign p1_bit_slice_154563_comb = p1_add_154499_comb[9:8];
  assign p1_bit_slice_154564_comb = p1_add_154500_comb[9:8];
  assign p1_bit_slice_154565_comb = p1_add_154501_comb[9:8];
  assign p1_bit_slice_154566_comb = p1_add_154502_comb[9:8];
  assign p1_bit_slice_154567_comb = p1_add_154503_comb[9:8];
  assign p1_bit_slice_154568_comb = p1_add_154504_comb[9:8];
  assign p1_bit_slice_154569_comb = p1_add_154505_comb[9:8];
  assign p1_bit_slice_154570_comb = p1_add_154506_comb[9:8];
  assign p1_bit_slice_154571_comb = p1_add_154507_comb[9:8];
  assign p1_bit_slice_154572_comb = p1_add_154508_comb[9:8];
  assign p1_bit_slice_154573_comb = p1_add_154509_comb[9:8];
  assign p1_bit_slice_154574_comb = p1_add_154510_comb[9:8];
  assign p1_bit_slice_154575_comb = p1_add_154511_comb[9:8];
  assign p1_bit_slice_154576_comb = p1_add_154512_comb[9:8];
  assign p1_bit_slice_154577_comb = p1_add_154513_comb[9:8];
  assign p1_bit_slice_154578_comb = p1_add_154514_comb[9:8];
  assign p1_add_154707_comb = {{1{p1_bit_slice_154515_comb[1]}}, p1_bit_slice_154515_comb} + 3'h1;
  assign p1_add_154708_comb = {{1{p1_bit_slice_154516_comb[1]}}, p1_bit_slice_154516_comb} + 3'h1;
  assign p1_add_154709_comb = {{1{p1_bit_slice_154517_comb[1]}}, p1_bit_slice_154517_comb} + 3'h1;
  assign p1_add_154710_comb = {{1{p1_bit_slice_154518_comb[1]}}, p1_bit_slice_154518_comb} + 3'h1;
  assign p1_add_154711_comb = {{1{p1_bit_slice_154519_comb[1]}}, p1_bit_slice_154519_comb} + 3'h1;
  assign p1_add_154712_comb = {{1{p1_bit_slice_154520_comb[1]}}, p1_bit_slice_154520_comb} + 3'h1;
  assign p1_add_154713_comb = {{1{p1_bit_slice_154521_comb[1]}}, p1_bit_slice_154521_comb} + 3'h1;
  assign p1_add_154714_comb = {{1{p1_bit_slice_154522_comb[1]}}, p1_bit_slice_154522_comb} + 3'h1;
  assign p1_add_154715_comb = {{1{p1_bit_slice_154523_comb[1]}}, p1_bit_slice_154523_comb} + 3'h1;
  assign p1_add_154716_comb = {{1{p1_bit_slice_154524_comb[1]}}, p1_bit_slice_154524_comb} + 3'h1;
  assign p1_add_154717_comb = {{1{p1_bit_slice_154525_comb[1]}}, p1_bit_slice_154525_comb} + 3'h1;
  assign p1_add_154718_comb = {{1{p1_bit_slice_154526_comb[1]}}, p1_bit_slice_154526_comb} + 3'h1;
  assign p1_add_154719_comb = {{1{p1_bit_slice_154527_comb[1]}}, p1_bit_slice_154527_comb} + 3'h1;
  assign p1_add_154720_comb = {{1{p1_bit_slice_154528_comb[1]}}, p1_bit_slice_154528_comb} + 3'h1;
  assign p1_add_154721_comb = {{1{p1_bit_slice_154529_comb[1]}}, p1_bit_slice_154529_comb} + 3'h1;
  assign p1_add_154722_comb = {{1{p1_bit_slice_154530_comb[1]}}, p1_bit_slice_154530_comb} + 3'h1;
  assign p1_add_154723_comb = {{1{p1_bit_slice_154531_comb[1]}}, p1_bit_slice_154531_comb} + 3'h1;
  assign p1_add_154724_comb = {{1{p1_bit_slice_154532_comb[1]}}, p1_bit_slice_154532_comb} + 3'h1;
  assign p1_add_154725_comb = {{1{p1_bit_slice_154533_comb[1]}}, p1_bit_slice_154533_comb} + 3'h1;
  assign p1_add_154726_comb = {{1{p1_bit_slice_154534_comb[1]}}, p1_bit_slice_154534_comb} + 3'h1;
  assign p1_add_154727_comb = {{1{p1_bit_slice_154535_comb[1]}}, p1_bit_slice_154535_comb} + 3'h1;
  assign p1_add_154728_comb = {{1{p1_bit_slice_154536_comb[1]}}, p1_bit_slice_154536_comb} + 3'h1;
  assign p1_add_154729_comb = {{1{p1_bit_slice_154537_comb[1]}}, p1_bit_slice_154537_comb} + 3'h1;
  assign p1_add_154730_comb = {{1{p1_bit_slice_154538_comb[1]}}, p1_bit_slice_154538_comb} + 3'h1;
  assign p1_add_154731_comb = {{1{p1_bit_slice_154539_comb[1]}}, p1_bit_slice_154539_comb} + 3'h1;
  assign p1_add_154732_comb = {{1{p1_bit_slice_154540_comb[1]}}, p1_bit_slice_154540_comb} + 3'h1;
  assign p1_add_154733_comb = {{1{p1_bit_slice_154541_comb[1]}}, p1_bit_slice_154541_comb} + 3'h1;
  assign p1_add_154734_comb = {{1{p1_bit_slice_154542_comb[1]}}, p1_bit_slice_154542_comb} + 3'h1;
  assign p1_add_154735_comb = {{1{p1_bit_slice_154543_comb[1]}}, p1_bit_slice_154543_comb} + 3'h1;
  assign p1_add_154736_comb = {{1{p1_bit_slice_154544_comb[1]}}, p1_bit_slice_154544_comb} + 3'h1;
  assign p1_add_154737_comb = {{1{p1_bit_slice_154545_comb[1]}}, p1_bit_slice_154545_comb} + 3'h1;
  assign p1_add_154738_comb = {{1{p1_bit_slice_154546_comb[1]}}, p1_bit_slice_154546_comb} + 3'h1;
  assign p1_add_154739_comb = {{1{p1_bit_slice_154547_comb[1]}}, p1_bit_slice_154547_comb} + 3'h1;
  assign p1_add_154740_comb = {{1{p1_bit_slice_154548_comb[1]}}, p1_bit_slice_154548_comb} + 3'h1;
  assign p1_add_154741_comb = {{1{p1_bit_slice_154549_comb[1]}}, p1_bit_slice_154549_comb} + 3'h1;
  assign p1_add_154742_comb = {{1{p1_bit_slice_154550_comb[1]}}, p1_bit_slice_154550_comb} + 3'h1;
  assign p1_add_154743_comb = {{1{p1_bit_slice_154551_comb[1]}}, p1_bit_slice_154551_comb} + 3'h1;
  assign p1_add_154744_comb = {{1{p1_bit_slice_154552_comb[1]}}, p1_bit_slice_154552_comb} + 3'h1;
  assign p1_add_154745_comb = {{1{p1_bit_slice_154553_comb[1]}}, p1_bit_slice_154553_comb} + 3'h1;
  assign p1_add_154746_comb = {{1{p1_bit_slice_154554_comb[1]}}, p1_bit_slice_154554_comb} + 3'h1;
  assign p1_add_154747_comb = {{1{p1_bit_slice_154555_comb[1]}}, p1_bit_slice_154555_comb} + 3'h1;
  assign p1_add_154748_comb = {{1{p1_bit_slice_154556_comb[1]}}, p1_bit_slice_154556_comb} + 3'h1;
  assign p1_add_154749_comb = {{1{p1_bit_slice_154557_comb[1]}}, p1_bit_slice_154557_comb} + 3'h1;
  assign p1_add_154750_comb = {{1{p1_bit_slice_154558_comb[1]}}, p1_bit_slice_154558_comb} + 3'h1;
  assign p1_add_154751_comb = {{1{p1_bit_slice_154559_comb[1]}}, p1_bit_slice_154559_comb} + 3'h1;
  assign p1_add_154752_comb = {{1{p1_bit_slice_154560_comb[1]}}, p1_bit_slice_154560_comb} + 3'h1;
  assign p1_add_154753_comb = {{1{p1_bit_slice_154561_comb[1]}}, p1_bit_slice_154561_comb} + 3'h1;
  assign p1_add_154754_comb = {{1{p1_bit_slice_154562_comb[1]}}, p1_bit_slice_154562_comb} + 3'h1;
  assign p1_add_154755_comb = {{1{p1_bit_slice_154563_comb[1]}}, p1_bit_slice_154563_comb} + 3'h1;
  assign p1_add_154756_comb = {{1{p1_bit_slice_154564_comb[1]}}, p1_bit_slice_154564_comb} + 3'h1;
  assign p1_add_154757_comb = {{1{p1_bit_slice_154565_comb[1]}}, p1_bit_slice_154565_comb} + 3'h1;
  assign p1_add_154758_comb = {{1{p1_bit_slice_154566_comb[1]}}, p1_bit_slice_154566_comb} + 3'h1;
  assign p1_add_154759_comb = {{1{p1_bit_slice_154567_comb[1]}}, p1_bit_slice_154567_comb} + 3'h1;
  assign p1_add_154760_comb = {{1{p1_bit_slice_154568_comb[1]}}, p1_bit_slice_154568_comb} + 3'h1;
  assign p1_add_154761_comb = {{1{p1_bit_slice_154569_comb[1]}}, p1_bit_slice_154569_comb} + 3'h1;
  assign p1_add_154762_comb = {{1{p1_bit_slice_154570_comb[1]}}, p1_bit_slice_154570_comb} + 3'h1;
  assign p1_add_154763_comb = {{1{p1_bit_slice_154571_comb[1]}}, p1_bit_slice_154571_comb} + 3'h1;
  assign p1_add_154764_comb = {{1{p1_bit_slice_154572_comb[1]}}, p1_bit_slice_154572_comb} + 3'h1;
  assign p1_add_154765_comb = {{1{p1_bit_slice_154573_comb[1]}}, p1_bit_slice_154573_comb} + 3'h1;
  assign p1_add_154766_comb = {{1{p1_bit_slice_154574_comb[1]}}, p1_bit_slice_154574_comb} + 3'h1;
  assign p1_add_154767_comb = {{1{p1_bit_slice_154575_comb[1]}}, p1_bit_slice_154575_comb} + 3'h1;
  assign p1_add_154768_comb = {{1{p1_bit_slice_154576_comb[1]}}, p1_bit_slice_154576_comb} + 3'h1;
  assign p1_add_154769_comb = {{1{p1_bit_slice_154577_comb[1]}}, p1_bit_slice_154577_comb} + 3'h1;
  assign p1_add_154770_comb = {{1{p1_bit_slice_154578_comb[1]}}, p1_bit_slice_154578_comb} + 3'h1;
  assign p1_clipped__136_comb = p1_add_154707_comb[1] ? 8'hff : {p1_add_154707_comb[0], p1_add_154451_comb[7:1]};
  assign p1_clipped__152_comb = p1_add_154708_comb[1] ? 8'hff : {p1_add_154708_comb[0], p1_add_154452_comb[7:1]};
  assign p1_clipped__168_comb = p1_add_154709_comb[1] ? 8'hff : {p1_add_154709_comb[0], p1_add_154453_comb[7:1]};
  assign p1_clipped__184_comb = p1_add_154710_comb[1] ? 8'hff : {p1_add_154710_comb[0], p1_add_154454_comb[7:1]};
  assign p1_clipped__200_comb = p1_add_154711_comb[1] ? 8'hff : {p1_add_154711_comb[0], p1_add_154455_comb[7:1]};
  assign p1_clipped__216_comb = p1_add_154712_comb[1] ? 8'hff : {p1_add_154712_comb[0], p1_add_154456_comb[7:1]};
  assign p1_clipped__232_comb = p1_add_154713_comb[1] ? 8'hff : {p1_add_154713_comb[0], p1_add_154457_comb[7:1]};
  assign p1_clipped__248_comb = p1_add_154714_comb[1] ? 8'hff : {p1_add_154714_comb[0], p1_add_154458_comb[7:1]};
  assign p1_clipped__137_comb = p1_add_154715_comb[1] ? 8'hff : {p1_add_154715_comb[0], p1_add_154459_comb[7:1]};
  assign p1_clipped__153_comb = p1_add_154716_comb[1] ? 8'hff : {p1_add_154716_comb[0], p1_add_154460_comb[7:1]};
  assign p1_clipped__169_comb = p1_add_154717_comb[1] ? 8'hff : {p1_add_154717_comb[0], p1_add_154461_comb[7:1]};
  assign p1_clipped__185_comb = p1_add_154718_comb[1] ? 8'hff : {p1_add_154718_comb[0], p1_add_154462_comb[7:1]};
  assign p1_clipped__201_comb = p1_add_154719_comb[1] ? 8'hff : {p1_add_154719_comb[0], p1_add_154463_comb[7:1]};
  assign p1_clipped__217_comb = p1_add_154720_comb[1] ? 8'hff : {p1_add_154720_comb[0], p1_add_154464_comb[7:1]};
  assign p1_clipped__233_comb = p1_add_154721_comb[1] ? 8'hff : {p1_add_154721_comb[0], p1_add_154465_comb[7:1]};
  assign p1_clipped__249_comb = p1_add_154722_comb[1] ? 8'hff : {p1_add_154722_comb[0], p1_add_154466_comb[7:1]};
  assign p1_clipped__138_comb = p1_add_154723_comb[1] ? 8'hff : {p1_add_154723_comb[0], p1_add_154467_comb[7:1]};
  assign p1_clipped__154_comb = p1_add_154724_comb[1] ? 8'hff : {p1_add_154724_comb[0], p1_add_154468_comb[7:1]};
  assign p1_clipped__170_comb = p1_add_154725_comb[1] ? 8'hff : {p1_add_154725_comb[0], p1_add_154469_comb[7:1]};
  assign p1_clipped__186_comb = p1_add_154726_comb[1] ? 8'hff : {p1_add_154726_comb[0], p1_add_154470_comb[7:1]};
  assign p1_clipped__202_comb = p1_add_154727_comb[1] ? 8'hff : {p1_add_154727_comb[0], p1_add_154471_comb[7:1]};
  assign p1_clipped__218_comb = p1_add_154728_comb[1] ? 8'hff : {p1_add_154728_comb[0], p1_add_154472_comb[7:1]};
  assign p1_clipped__234_comb = p1_add_154729_comb[1] ? 8'hff : {p1_add_154729_comb[0], p1_add_154473_comb[7:1]};
  assign p1_clipped__250_comb = p1_add_154730_comb[1] ? 8'hff : {p1_add_154730_comb[0], p1_add_154474_comb[7:1]};
  assign p1_clipped__139_comb = p1_add_154731_comb[1] ? 8'hff : {p1_add_154731_comb[0], p1_add_154475_comb[7:1]};
  assign p1_clipped__155_comb = p1_add_154732_comb[1] ? 8'hff : {p1_add_154732_comb[0], p1_add_154476_comb[7:1]};
  assign p1_clipped__171_comb = p1_add_154733_comb[1] ? 8'hff : {p1_add_154733_comb[0], p1_add_154477_comb[7:1]};
  assign p1_clipped__187_comb = p1_add_154734_comb[1] ? 8'hff : {p1_add_154734_comb[0], p1_add_154478_comb[7:1]};
  assign p1_clipped__203_comb = p1_add_154735_comb[1] ? 8'hff : {p1_add_154735_comb[0], p1_add_154479_comb[7:1]};
  assign p1_clipped__219_comb = p1_add_154736_comb[1] ? 8'hff : {p1_add_154736_comb[0], p1_add_154480_comb[7:1]};
  assign p1_clipped__235_comb = p1_add_154737_comb[1] ? 8'hff : {p1_add_154737_comb[0], p1_add_154481_comb[7:1]};
  assign p1_clipped__251_comb = p1_add_154738_comb[1] ? 8'hff : {p1_add_154738_comb[0], p1_add_154482_comb[7:1]};
  assign p1_clipped__140_comb = p1_add_154739_comb[1] ? 8'hff : {p1_add_154739_comb[0], p1_add_154483_comb[7:1]};
  assign p1_clipped__156_comb = p1_add_154740_comb[1] ? 8'hff : {p1_add_154740_comb[0], p1_add_154484_comb[7:1]};
  assign p1_clipped__172_comb = p1_add_154741_comb[1] ? 8'hff : {p1_add_154741_comb[0], p1_add_154485_comb[7:1]};
  assign p1_clipped__188_comb = p1_add_154742_comb[1] ? 8'hff : {p1_add_154742_comb[0], p1_add_154486_comb[7:1]};
  assign p1_clipped__204_comb = p1_add_154743_comb[1] ? 8'hff : {p1_add_154743_comb[0], p1_add_154487_comb[7:1]};
  assign p1_clipped__220_comb = p1_add_154744_comb[1] ? 8'hff : {p1_add_154744_comb[0], p1_add_154488_comb[7:1]};
  assign p1_clipped__236_comb = p1_add_154745_comb[1] ? 8'hff : {p1_add_154745_comb[0], p1_add_154489_comb[7:1]};
  assign p1_clipped__252_comb = p1_add_154746_comb[1] ? 8'hff : {p1_add_154746_comb[0], p1_add_154490_comb[7:1]};
  assign p1_clipped__141_comb = p1_add_154747_comb[1] ? 8'hff : {p1_add_154747_comb[0], p1_add_154491_comb[7:1]};
  assign p1_clipped__157_comb = p1_add_154748_comb[1] ? 8'hff : {p1_add_154748_comb[0], p1_add_154492_comb[7:1]};
  assign p1_clipped__173_comb = p1_add_154749_comb[1] ? 8'hff : {p1_add_154749_comb[0], p1_add_154493_comb[7:1]};
  assign p1_clipped__189_comb = p1_add_154750_comb[1] ? 8'hff : {p1_add_154750_comb[0], p1_add_154494_comb[7:1]};
  assign p1_clipped__205_comb = p1_add_154751_comb[1] ? 8'hff : {p1_add_154751_comb[0], p1_add_154495_comb[7:1]};
  assign p1_clipped__221_comb = p1_add_154752_comb[1] ? 8'hff : {p1_add_154752_comb[0], p1_add_154496_comb[7:1]};
  assign p1_clipped__237_comb = p1_add_154753_comb[1] ? 8'hff : {p1_add_154753_comb[0], p1_add_154497_comb[7:1]};
  assign p1_clipped__253_comb = p1_add_154754_comb[1] ? 8'hff : {p1_add_154754_comb[0], p1_add_154498_comb[7:1]};
  assign p1_clipped__142_comb = p1_add_154755_comb[1] ? 8'hff : {p1_add_154755_comb[0], p1_add_154499_comb[7:1]};
  assign p1_clipped__158_comb = p1_add_154756_comb[1] ? 8'hff : {p1_add_154756_comb[0], p1_add_154500_comb[7:1]};
  assign p1_clipped__174_comb = p1_add_154757_comb[1] ? 8'hff : {p1_add_154757_comb[0], p1_add_154501_comb[7:1]};
  assign p1_clipped__190_comb = p1_add_154758_comb[1] ? 8'hff : {p1_add_154758_comb[0], p1_add_154502_comb[7:1]};
  assign p1_clipped__206_comb = p1_add_154759_comb[1] ? 8'hff : {p1_add_154759_comb[0], p1_add_154503_comb[7:1]};
  assign p1_clipped__222_comb = p1_add_154760_comb[1] ? 8'hff : {p1_add_154760_comb[0], p1_add_154504_comb[7:1]};
  assign p1_clipped__238_comb = p1_add_154761_comb[1] ? 8'hff : {p1_add_154761_comb[0], p1_add_154505_comb[7:1]};
  assign p1_clipped__254_comb = p1_add_154762_comb[1] ? 8'hff : {p1_add_154762_comb[0], p1_add_154506_comb[7:1]};
  assign p1_clipped__143_comb = p1_add_154763_comb[1] ? 8'hff : {p1_add_154763_comb[0], p1_add_154507_comb[7:1]};
  assign p1_clipped__159_comb = p1_add_154764_comb[1] ? 8'hff : {p1_add_154764_comb[0], p1_add_154508_comb[7:1]};
  assign p1_clipped__175_comb = p1_add_154765_comb[1] ? 8'hff : {p1_add_154765_comb[0], p1_add_154509_comb[7:1]};
  assign p1_clipped__191_comb = p1_add_154766_comb[1] ? 8'hff : {p1_add_154766_comb[0], p1_add_154510_comb[7:1]};
  assign p1_clipped__207_comb = p1_add_154767_comb[1] ? 8'hff : {p1_add_154767_comb[0], p1_add_154511_comb[7:1]};
  assign p1_clipped__223_comb = p1_add_154768_comb[1] ? 8'hff : {p1_add_154768_comb[0], p1_add_154512_comb[7:1]};
  assign p1_clipped__239_comb = p1_add_154769_comb[1] ? 8'hff : {p1_add_154769_comb[0], p1_add_154513_comb[7:1]};
  assign p1_clipped__255_comb = p1_add_154770_comb[1] ? 8'hff : {p1_add_154770_comb[0], p1_add_154514_comb[7:1]};
  assign p1_array_155155_comb[0] = p1_clipped__136_comb;
  assign p1_array_155155_comb[1] = p1_clipped__152_comb;
  assign p1_array_155155_comb[2] = p1_clipped__168_comb;
  assign p1_array_155155_comb[3] = p1_clipped__184_comb;
  assign p1_array_155155_comb[4] = p1_clipped__200_comb;
  assign p1_array_155155_comb[5] = p1_clipped__216_comb;
  assign p1_array_155155_comb[6] = p1_clipped__232_comb;
  assign p1_array_155155_comb[7] = p1_clipped__248_comb;
  assign p1_array_155156_comb[0] = p1_clipped__137_comb;
  assign p1_array_155156_comb[1] = p1_clipped__153_comb;
  assign p1_array_155156_comb[2] = p1_clipped__169_comb;
  assign p1_array_155156_comb[3] = p1_clipped__185_comb;
  assign p1_array_155156_comb[4] = p1_clipped__201_comb;
  assign p1_array_155156_comb[5] = p1_clipped__217_comb;
  assign p1_array_155156_comb[6] = p1_clipped__233_comb;
  assign p1_array_155156_comb[7] = p1_clipped__249_comb;
  assign p1_array_155157_comb[0] = p1_clipped__138_comb;
  assign p1_array_155157_comb[1] = p1_clipped__154_comb;
  assign p1_array_155157_comb[2] = p1_clipped__170_comb;
  assign p1_array_155157_comb[3] = p1_clipped__186_comb;
  assign p1_array_155157_comb[4] = p1_clipped__202_comb;
  assign p1_array_155157_comb[5] = p1_clipped__218_comb;
  assign p1_array_155157_comb[6] = p1_clipped__234_comb;
  assign p1_array_155157_comb[7] = p1_clipped__250_comb;
  assign p1_array_155158_comb[0] = p1_clipped__139_comb;
  assign p1_array_155158_comb[1] = p1_clipped__155_comb;
  assign p1_array_155158_comb[2] = p1_clipped__171_comb;
  assign p1_array_155158_comb[3] = p1_clipped__187_comb;
  assign p1_array_155158_comb[4] = p1_clipped__203_comb;
  assign p1_array_155158_comb[5] = p1_clipped__219_comb;
  assign p1_array_155158_comb[6] = p1_clipped__235_comb;
  assign p1_array_155158_comb[7] = p1_clipped__251_comb;
  assign p1_array_155159_comb[0] = p1_clipped__140_comb;
  assign p1_array_155159_comb[1] = p1_clipped__156_comb;
  assign p1_array_155159_comb[2] = p1_clipped__172_comb;
  assign p1_array_155159_comb[3] = p1_clipped__188_comb;
  assign p1_array_155159_comb[4] = p1_clipped__204_comb;
  assign p1_array_155159_comb[5] = p1_clipped__220_comb;
  assign p1_array_155159_comb[6] = p1_clipped__236_comb;
  assign p1_array_155159_comb[7] = p1_clipped__252_comb;
  assign p1_array_155160_comb[0] = p1_clipped__141_comb;
  assign p1_array_155160_comb[1] = p1_clipped__157_comb;
  assign p1_array_155160_comb[2] = p1_clipped__173_comb;
  assign p1_array_155160_comb[3] = p1_clipped__189_comb;
  assign p1_array_155160_comb[4] = p1_clipped__205_comb;
  assign p1_array_155160_comb[5] = p1_clipped__221_comb;
  assign p1_array_155160_comb[6] = p1_clipped__237_comb;
  assign p1_array_155160_comb[7] = p1_clipped__253_comb;
  assign p1_array_155161_comb[0] = p1_clipped__142_comb;
  assign p1_array_155161_comb[1] = p1_clipped__158_comb;
  assign p1_array_155161_comb[2] = p1_clipped__174_comb;
  assign p1_array_155161_comb[3] = p1_clipped__190_comb;
  assign p1_array_155161_comb[4] = p1_clipped__206_comb;
  assign p1_array_155161_comb[5] = p1_clipped__222_comb;
  assign p1_array_155161_comb[6] = p1_clipped__238_comb;
  assign p1_array_155161_comb[7] = p1_clipped__254_comb;
  assign p1_array_155162_comb[0] = p1_clipped__143_comb;
  assign p1_array_155162_comb[1] = p1_clipped__159_comb;
  assign p1_array_155162_comb[2] = p1_clipped__175_comb;
  assign p1_array_155162_comb[3] = p1_clipped__191_comb;
  assign p1_array_155162_comb[4] = p1_clipped__207_comb;
  assign p1_array_155162_comb[5] = p1_clipped__223_comb;
  assign p1_array_155162_comb[6] = p1_clipped__239_comb;
  assign p1_array_155162_comb[7] = p1_clipped__255_comb;
  assign p1_col_transformed_comb[0][0] = p1_array_155155_comb[0];
  assign p1_col_transformed_comb[0][1] = p1_array_155155_comb[1];
  assign p1_col_transformed_comb[0][2] = p1_array_155155_comb[2];
  assign p1_col_transformed_comb[0][3] = p1_array_155155_comb[3];
  assign p1_col_transformed_comb[0][4] = p1_array_155155_comb[4];
  assign p1_col_transformed_comb[0][5] = p1_array_155155_comb[5];
  assign p1_col_transformed_comb[0][6] = p1_array_155155_comb[6];
  assign p1_col_transformed_comb[0][7] = p1_array_155155_comb[7];
  assign p1_col_transformed_comb[1][0] = p1_array_155156_comb[0];
  assign p1_col_transformed_comb[1][1] = p1_array_155156_comb[1];
  assign p1_col_transformed_comb[1][2] = p1_array_155156_comb[2];
  assign p1_col_transformed_comb[1][3] = p1_array_155156_comb[3];
  assign p1_col_transformed_comb[1][4] = p1_array_155156_comb[4];
  assign p1_col_transformed_comb[1][5] = p1_array_155156_comb[5];
  assign p1_col_transformed_comb[1][6] = p1_array_155156_comb[6];
  assign p1_col_transformed_comb[1][7] = p1_array_155156_comb[7];
  assign p1_col_transformed_comb[2][0] = p1_array_155157_comb[0];
  assign p1_col_transformed_comb[2][1] = p1_array_155157_comb[1];
  assign p1_col_transformed_comb[2][2] = p1_array_155157_comb[2];
  assign p1_col_transformed_comb[2][3] = p1_array_155157_comb[3];
  assign p1_col_transformed_comb[2][4] = p1_array_155157_comb[4];
  assign p1_col_transformed_comb[2][5] = p1_array_155157_comb[5];
  assign p1_col_transformed_comb[2][6] = p1_array_155157_comb[6];
  assign p1_col_transformed_comb[2][7] = p1_array_155157_comb[7];
  assign p1_col_transformed_comb[3][0] = p1_array_155158_comb[0];
  assign p1_col_transformed_comb[3][1] = p1_array_155158_comb[1];
  assign p1_col_transformed_comb[3][2] = p1_array_155158_comb[2];
  assign p1_col_transformed_comb[3][3] = p1_array_155158_comb[3];
  assign p1_col_transformed_comb[3][4] = p1_array_155158_comb[4];
  assign p1_col_transformed_comb[3][5] = p1_array_155158_comb[5];
  assign p1_col_transformed_comb[3][6] = p1_array_155158_comb[6];
  assign p1_col_transformed_comb[3][7] = p1_array_155158_comb[7];
  assign p1_col_transformed_comb[4][0] = p1_array_155159_comb[0];
  assign p1_col_transformed_comb[4][1] = p1_array_155159_comb[1];
  assign p1_col_transformed_comb[4][2] = p1_array_155159_comb[2];
  assign p1_col_transformed_comb[4][3] = p1_array_155159_comb[3];
  assign p1_col_transformed_comb[4][4] = p1_array_155159_comb[4];
  assign p1_col_transformed_comb[4][5] = p1_array_155159_comb[5];
  assign p1_col_transformed_comb[4][6] = p1_array_155159_comb[6];
  assign p1_col_transformed_comb[4][7] = p1_array_155159_comb[7];
  assign p1_col_transformed_comb[5][0] = p1_array_155160_comb[0];
  assign p1_col_transformed_comb[5][1] = p1_array_155160_comb[1];
  assign p1_col_transformed_comb[5][2] = p1_array_155160_comb[2];
  assign p1_col_transformed_comb[5][3] = p1_array_155160_comb[3];
  assign p1_col_transformed_comb[5][4] = p1_array_155160_comb[4];
  assign p1_col_transformed_comb[5][5] = p1_array_155160_comb[5];
  assign p1_col_transformed_comb[5][6] = p1_array_155160_comb[6];
  assign p1_col_transformed_comb[5][7] = p1_array_155160_comb[7];
  assign p1_col_transformed_comb[6][0] = p1_array_155161_comb[0];
  assign p1_col_transformed_comb[6][1] = p1_array_155161_comb[1];
  assign p1_col_transformed_comb[6][2] = p1_array_155161_comb[2];
  assign p1_col_transformed_comb[6][3] = p1_array_155161_comb[3];
  assign p1_col_transformed_comb[6][4] = p1_array_155161_comb[4];
  assign p1_col_transformed_comb[6][5] = p1_array_155161_comb[5];
  assign p1_col_transformed_comb[6][6] = p1_array_155161_comb[6];
  assign p1_col_transformed_comb[6][7] = p1_array_155161_comb[7];
  assign p1_col_transformed_comb[7][0] = p1_array_155162_comb[0];
  assign p1_col_transformed_comb[7][1] = p1_array_155162_comb[1];
  assign p1_col_transformed_comb[7][2] = p1_array_155162_comb[2];
  assign p1_col_transformed_comb[7][3] = p1_array_155162_comb[3];
  assign p1_col_transformed_comb[7][4] = p1_array_155162_comb[4];
  assign p1_col_transformed_comb[7][5] = p1_array_155162_comb[5];
  assign p1_col_transformed_comb[7][6] = p1_array_155162_comb[6];
  assign p1_col_transformed_comb[7][7] = p1_array_155162_comb[7];

  // Registers for pipe stage 1:
  reg [7:0] p1_col_transformed[0:7][0:7];
  always @ (posedge clk) begin
    p1_col_transformed[0][0] <= p1_col_transformed_comb[0][0];
    p1_col_transformed[0][1] <= p1_col_transformed_comb[0][1];
    p1_col_transformed[0][2] <= p1_col_transformed_comb[0][2];
    p1_col_transformed[0][3] <= p1_col_transformed_comb[0][3];
    p1_col_transformed[0][4] <= p1_col_transformed_comb[0][4];
    p1_col_transformed[0][5] <= p1_col_transformed_comb[0][5];
    p1_col_transformed[0][6] <= p1_col_transformed_comb[0][6];
    p1_col_transformed[0][7] <= p1_col_transformed_comb[0][7];
    p1_col_transformed[1][0] <= p1_col_transformed_comb[1][0];
    p1_col_transformed[1][1] <= p1_col_transformed_comb[1][1];
    p1_col_transformed[1][2] <= p1_col_transformed_comb[1][2];
    p1_col_transformed[1][3] <= p1_col_transformed_comb[1][3];
    p1_col_transformed[1][4] <= p1_col_transformed_comb[1][4];
    p1_col_transformed[1][5] <= p1_col_transformed_comb[1][5];
    p1_col_transformed[1][6] <= p1_col_transformed_comb[1][6];
    p1_col_transformed[1][7] <= p1_col_transformed_comb[1][7];
    p1_col_transformed[2][0] <= p1_col_transformed_comb[2][0];
    p1_col_transformed[2][1] <= p1_col_transformed_comb[2][1];
    p1_col_transformed[2][2] <= p1_col_transformed_comb[2][2];
    p1_col_transformed[2][3] <= p1_col_transformed_comb[2][3];
    p1_col_transformed[2][4] <= p1_col_transformed_comb[2][4];
    p1_col_transformed[2][5] <= p1_col_transformed_comb[2][5];
    p1_col_transformed[2][6] <= p1_col_transformed_comb[2][6];
    p1_col_transformed[2][7] <= p1_col_transformed_comb[2][7];
    p1_col_transformed[3][0] <= p1_col_transformed_comb[3][0];
    p1_col_transformed[3][1] <= p1_col_transformed_comb[3][1];
    p1_col_transformed[3][2] <= p1_col_transformed_comb[3][2];
    p1_col_transformed[3][3] <= p1_col_transformed_comb[3][3];
    p1_col_transformed[3][4] <= p1_col_transformed_comb[3][4];
    p1_col_transformed[3][5] <= p1_col_transformed_comb[3][5];
    p1_col_transformed[3][6] <= p1_col_transformed_comb[3][6];
    p1_col_transformed[3][7] <= p1_col_transformed_comb[3][7];
    p1_col_transformed[4][0] <= p1_col_transformed_comb[4][0];
    p1_col_transformed[4][1] <= p1_col_transformed_comb[4][1];
    p1_col_transformed[4][2] <= p1_col_transformed_comb[4][2];
    p1_col_transformed[4][3] <= p1_col_transformed_comb[4][3];
    p1_col_transformed[4][4] <= p1_col_transformed_comb[4][4];
    p1_col_transformed[4][5] <= p1_col_transformed_comb[4][5];
    p1_col_transformed[4][6] <= p1_col_transformed_comb[4][6];
    p1_col_transformed[4][7] <= p1_col_transformed_comb[4][7];
    p1_col_transformed[5][0] <= p1_col_transformed_comb[5][0];
    p1_col_transformed[5][1] <= p1_col_transformed_comb[5][1];
    p1_col_transformed[5][2] <= p1_col_transformed_comb[5][2];
    p1_col_transformed[5][3] <= p1_col_transformed_comb[5][3];
    p1_col_transformed[5][4] <= p1_col_transformed_comb[5][4];
    p1_col_transformed[5][5] <= p1_col_transformed_comb[5][5];
    p1_col_transformed[5][6] <= p1_col_transformed_comb[5][6];
    p1_col_transformed[5][7] <= p1_col_transformed_comb[5][7];
    p1_col_transformed[6][0] <= p1_col_transformed_comb[6][0];
    p1_col_transformed[6][1] <= p1_col_transformed_comb[6][1];
    p1_col_transformed[6][2] <= p1_col_transformed_comb[6][2];
    p1_col_transformed[6][3] <= p1_col_transformed_comb[6][3];
    p1_col_transformed[6][4] <= p1_col_transformed_comb[6][4];
    p1_col_transformed[6][5] <= p1_col_transformed_comb[6][5];
    p1_col_transformed[6][6] <= p1_col_transformed_comb[6][6];
    p1_col_transformed[6][7] <= p1_col_transformed_comb[6][7];
    p1_col_transformed[7][0] <= p1_col_transformed_comb[7][0];
    p1_col_transformed[7][1] <= p1_col_transformed_comb[7][1];
    p1_col_transformed[7][2] <= p1_col_transformed_comb[7][2];
    p1_col_transformed[7][3] <= p1_col_transformed_comb[7][3];
    p1_col_transformed[7][4] <= p1_col_transformed_comb[7][4];
    p1_col_transformed[7][5] <= p1_col_transformed_comb[7][5];
    p1_col_transformed[7][6] <= p1_col_transformed_comb[7][6];
    p1_col_transformed[7][7] <= p1_col_transformed_comb[7][7];
  end
  assign out = {{p1_col_transformed[7][7], p1_col_transformed[7][6], p1_col_transformed[7][5], p1_col_transformed[7][4], p1_col_transformed[7][3], p1_col_transformed[7][2], p1_col_transformed[7][1], p1_col_transformed[7][0]}, {p1_col_transformed[6][7], p1_col_transformed[6][6], p1_col_transformed[6][5], p1_col_transformed[6][4], p1_col_transformed[6][3], p1_col_transformed[6][2], p1_col_transformed[6][1], p1_col_transformed[6][0]}, {p1_col_transformed[5][7], p1_col_transformed[5][6], p1_col_transformed[5][5], p1_col_transformed[5][4], p1_col_transformed[5][3], p1_col_transformed[5][2], p1_col_transformed[5][1], p1_col_transformed[5][0]}, {p1_col_transformed[4][7], p1_col_transformed[4][6], p1_col_transformed[4][5], p1_col_transformed[4][4], p1_col_transformed[4][3], p1_col_transformed[4][2], p1_col_transformed[4][1], p1_col_transformed[4][0]}, {p1_col_transformed[3][7], p1_col_transformed[3][6], p1_col_transformed[3][5], p1_col_transformed[3][4], p1_col_transformed[3][3], p1_col_transformed[3][2], p1_col_transformed[3][1], p1_col_transformed[3][0]}, {p1_col_transformed[2][7], p1_col_transformed[2][6], p1_col_transformed[2][5], p1_col_transformed[2][4], p1_col_transformed[2][3], p1_col_transformed[2][2], p1_col_transformed[2][1], p1_col_transformed[2][0]}, {p1_col_transformed[1][7], p1_col_transformed[1][6], p1_col_transformed[1][5], p1_col_transformed[1][4], p1_col_transformed[1][3], p1_col_transformed[1][2], p1_col_transformed[1][1], p1_col_transformed[1][0]}, {p1_col_transformed[0][7], p1_col_transformed[0][6], p1_col_transformed[0][5], p1_col_transformed[0][4], p1_col_transformed[0][3], p1_col_transformed[0][2], p1_col_transformed[0][1], p1_col_transformed[0][0]}};
endmodule
