module Zigzag_reorder(
  input wire clk,
  input wire [639:0] matrix,
  input wire is_enable,
  output wire [639:0] out
);
  wire [9:0] ZERO64[0:63];
  assign ZERO64[0] = 10'h000;
  assign ZERO64[1] = 10'h000;
  assign ZERO64[2] = 10'h000;
  assign ZERO64[3] = 10'h000;
  assign ZERO64[4] = 10'h000;
  assign ZERO64[5] = 10'h000;
  assign ZERO64[6] = 10'h000;
  assign ZERO64[7] = 10'h000;
  assign ZERO64[8] = 10'h000;
  assign ZERO64[9] = 10'h000;
  assign ZERO64[10] = 10'h000;
  assign ZERO64[11] = 10'h000;
  assign ZERO64[12] = 10'h000;
  assign ZERO64[13] = 10'h000;
  assign ZERO64[14] = 10'h000;
  assign ZERO64[15] = 10'h000;
  assign ZERO64[16] = 10'h000;
  assign ZERO64[17] = 10'h000;
  assign ZERO64[18] = 10'h000;
  assign ZERO64[19] = 10'h000;
  assign ZERO64[20] = 10'h000;
  assign ZERO64[21] = 10'h000;
  assign ZERO64[22] = 10'h000;
  assign ZERO64[23] = 10'h000;
  assign ZERO64[24] = 10'h000;
  assign ZERO64[25] = 10'h000;
  assign ZERO64[26] = 10'h000;
  assign ZERO64[27] = 10'h000;
  assign ZERO64[28] = 10'h000;
  assign ZERO64[29] = 10'h000;
  assign ZERO64[30] = 10'h000;
  assign ZERO64[31] = 10'h000;
  assign ZERO64[32] = 10'h000;
  assign ZERO64[33] = 10'h000;
  assign ZERO64[34] = 10'h000;
  assign ZERO64[35] = 10'h000;
  assign ZERO64[36] = 10'h000;
  assign ZERO64[37] = 10'h000;
  assign ZERO64[38] = 10'h000;
  assign ZERO64[39] = 10'h000;
  assign ZERO64[40] = 10'h000;
  assign ZERO64[41] = 10'h000;
  assign ZERO64[42] = 10'h000;
  assign ZERO64[43] = 10'h000;
  assign ZERO64[44] = 10'h000;
  assign ZERO64[45] = 10'h000;
  assign ZERO64[46] = 10'h000;
  assign ZERO64[47] = 10'h000;
  assign ZERO64[48] = 10'h000;
  assign ZERO64[49] = 10'h000;
  assign ZERO64[50] = 10'h000;
  assign ZERO64[51] = 10'h000;
  assign ZERO64[52] = 10'h000;
  assign ZERO64[53] = 10'h000;
  assign ZERO64[54] = 10'h000;
  assign ZERO64[55] = 10'h000;
  assign ZERO64[56] = 10'h000;
  assign ZERO64[57] = 10'h000;
  assign ZERO64[58] = 10'h000;
  assign ZERO64[59] = 10'h000;
  assign ZERO64[60] = 10'h000;
  assign ZERO64[61] = 10'h000;
  assign ZERO64[62] = 10'h000;
  assign ZERO64[63] = 10'h000;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg p0_is_enable;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_is_enable <= is_enable;
  end

  // ===== Pipe stage 1:
  wire [9:0] p1_array_1507_comb[0:63];
  wire [9:0] p1_sel_1508_comb[0:63];
  assign p1_array_1507_comb[0] = p0_matrix[3'h7][3'h7];
  assign p1_array_1507_comb[1] = p0_matrix[3'h7][3'h6];
  assign p1_array_1507_comb[2] = p0_matrix[3'h6][3'h7];
  assign p1_array_1507_comb[3] = p0_matrix[3'h5][3'h7];
  assign p1_array_1507_comb[4] = p0_matrix[3'h6][3'h6];
  assign p1_array_1507_comb[5] = p0_matrix[3'h7][3'h5];
  assign p1_array_1507_comb[6] = p0_matrix[3'h7][3'h4];
  assign p1_array_1507_comb[7] = p0_matrix[3'h6][3'h5];
  assign p1_array_1507_comb[8] = p0_matrix[3'h5][3'h6];
  assign p1_array_1507_comb[9] = p0_matrix[3'h4][3'h7];
  assign p1_array_1507_comb[10] = p0_matrix[3'h3][3'h7];
  assign p1_array_1507_comb[11] = p0_matrix[3'h4][3'h6];
  assign p1_array_1507_comb[12] = p0_matrix[3'h5][3'h5];
  assign p1_array_1507_comb[13] = p0_matrix[3'h6][3'h4];
  assign p1_array_1507_comb[14] = p0_matrix[3'h7][3'h3];
  assign p1_array_1507_comb[15] = p0_matrix[3'h7][3'h2];
  assign p1_array_1507_comb[16] = p0_matrix[3'h6][3'h3];
  assign p1_array_1507_comb[17] = p0_matrix[3'h5][3'h4];
  assign p1_array_1507_comb[18] = p0_matrix[3'h4][3'h5];
  assign p1_array_1507_comb[19] = p0_matrix[3'h3][3'h6];
  assign p1_array_1507_comb[20] = p0_matrix[3'h2][3'h7];
  assign p1_array_1507_comb[21] = p0_matrix[3'h1][3'h7];
  assign p1_array_1507_comb[22] = p0_matrix[3'h2][3'h6];
  assign p1_array_1507_comb[23] = p0_matrix[3'h3][3'h5];
  assign p1_array_1507_comb[24] = p0_matrix[3'h4][3'h4];
  assign p1_array_1507_comb[25] = p0_matrix[3'h5][3'h3];
  assign p1_array_1507_comb[26] = p0_matrix[3'h6][3'h2];
  assign p1_array_1507_comb[27] = p0_matrix[3'h7][3'h1];
  assign p1_array_1507_comb[28] = p0_matrix[3'h7][3'h0];
  assign p1_array_1507_comb[29] = p0_matrix[3'h6][3'h1];
  assign p1_array_1507_comb[30] = p0_matrix[3'h5][3'h2];
  assign p1_array_1507_comb[31] = p0_matrix[3'h4][3'h3];
  assign p1_array_1507_comb[32] = p0_matrix[3'h3][3'h4];
  assign p1_array_1507_comb[33] = p0_matrix[3'h2][3'h5];
  assign p1_array_1507_comb[34] = p0_matrix[3'h1][3'h6];
  assign p1_array_1507_comb[35] = p0_matrix[3'h0][3'h7];
  assign p1_array_1507_comb[36] = p0_matrix[3'h0][3'h6];
  assign p1_array_1507_comb[37] = p0_matrix[3'h1][3'h5];
  assign p1_array_1507_comb[38] = p0_matrix[3'h2][3'h4];
  assign p1_array_1507_comb[39] = p0_matrix[3'h3][3'h3];
  assign p1_array_1507_comb[40] = p0_matrix[3'h4][3'h2];
  assign p1_array_1507_comb[41] = p0_matrix[3'h5][3'h1];
  assign p1_array_1507_comb[42] = p0_matrix[3'h6][3'h0];
  assign p1_array_1507_comb[43] = p0_matrix[3'h5][3'h0];
  assign p1_array_1507_comb[44] = p0_matrix[3'h4][3'h1];
  assign p1_array_1507_comb[45] = p0_matrix[3'h3][3'h2];
  assign p1_array_1507_comb[46] = p0_matrix[3'h2][3'h3];
  assign p1_array_1507_comb[47] = p0_matrix[3'h1][3'h4];
  assign p1_array_1507_comb[48] = p0_matrix[3'h0][3'h5];
  assign p1_array_1507_comb[49] = p0_matrix[3'h0][3'h4];
  assign p1_array_1507_comb[50] = p0_matrix[3'h1][3'h3];
  assign p1_array_1507_comb[51] = p0_matrix[3'h2][3'h2];
  assign p1_array_1507_comb[52] = p0_matrix[3'h3][3'h1];
  assign p1_array_1507_comb[53] = p0_matrix[3'h4][3'h0];
  assign p1_array_1507_comb[54] = p0_matrix[3'h3][3'h0];
  assign p1_array_1507_comb[55] = p0_matrix[3'h2][3'h1];
  assign p1_array_1507_comb[56] = p0_matrix[3'h1][3'h2];
  assign p1_array_1507_comb[57] = p0_matrix[3'h0][3'h3];
  assign p1_array_1507_comb[58] = p0_matrix[3'h0][3'h2];
  assign p1_array_1507_comb[59] = p0_matrix[3'h1][3'h1];
  assign p1_array_1507_comb[60] = p0_matrix[3'h2][3'h0];
  assign p1_array_1507_comb[61] = p0_matrix[3'h1][3'h0];
  assign p1_array_1507_comb[62] = p0_matrix[3'h0][3'h1];
  assign p1_array_1507_comb[63] = p0_matrix[3'h0][3'h0];
  assign p1_sel_1508_comb[0] = p0_is_enable == 1'h0 ? ZERO64[0] : p1_array_1507_comb[0];
  assign p1_sel_1508_comb[1] = p0_is_enable == 1'h0 ? ZERO64[1] : p1_array_1507_comb[1];
  assign p1_sel_1508_comb[2] = p0_is_enable == 1'h0 ? ZERO64[2] : p1_array_1507_comb[2];
  assign p1_sel_1508_comb[3] = p0_is_enable == 1'h0 ? ZERO64[3] : p1_array_1507_comb[3];
  assign p1_sel_1508_comb[4] = p0_is_enable == 1'h0 ? ZERO64[4] : p1_array_1507_comb[4];
  assign p1_sel_1508_comb[5] = p0_is_enable == 1'h0 ? ZERO64[5] : p1_array_1507_comb[5];
  assign p1_sel_1508_comb[6] = p0_is_enable == 1'h0 ? ZERO64[6] : p1_array_1507_comb[6];
  assign p1_sel_1508_comb[7] = p0_is_enable == 1'h0 ? ZERO64[7] : p1_array_1507_comb[7];
  assign p1_sel_1508_comb[8] = p0_is_enable == 1'h0 ? ZERO64[8] : p1_array_1507_comb[8];
  assign p1_sel_1508_comb[9] = p0_is_enable == 1'h0 ? ZERO64[9] : p1_array_1507_comb[9];
  assign p1_sel_1508_comb[10] = p0_is_enable == 1'h0 ? ZERO64[10] : p1_array_1507_comb[10];
  assign p1_sel_1508_comb[11] = p0_is_enable == 1'h0 ? ZERO64[11] : p1_array_1507_comb[11];
  assign p1_sel_1508_comb[12] = p0_is_enable == 1'h0 ? ZERO64[12] : p1_array_1507_comb[12];
  assign p1_sel_1508_comb[13] = p0_is_enable == 1'h0 ? ZERO64[13] : p1_array_1507_comb[13];
  assign p1_sel_1508_comb[14] = p0_is_enable == 1'h0 ? ZERO64[14] : p1_array_1507_comb[14];
  assign p1_sel_1508_comb[15] = p0_is_enable == 1'h0 ? ZERO64[15] : p1_array_1507_comb[15];
  assign p1_sel_1508_comb[16] = p0_is_enable == 1'h0 ? ZERO64[16] : p1_array_1507_comb[16];
  assign p1_sel_1508_comb[17] = p0_is_enable == 1'h0 ? ZERO64[17] : p1_array_1507_comb[17];
  assign p1_sel_1508_comb[18] = p0_is_enable == 1'h0 ? ZERO64[18] : p1_array_1507_comb[18];
  assign p1_sel_1508_comb[19] = p0_is_enable == 1'h0 ? ZERO64[19] : p1_array_1507_comb[19];
  assign p1_sel_1508_comb[20] = p0_is_enable == 1'h0 ? ZERO64[20] : p1_array_1507_comb[20];
  assign p1_sel_1508_comb[21] = p0_is_enable == 1'h0 ? ZERO64[21] : p1_array_1507_comb[21];
  assign p1_sel_1508_comb[22] = p0_is_enable == 1'h0 ? ZERO64[22] : p1_array_1507_comb[22];
  assign p1_sel_1508_comb[23] = p0_is_enable == 1'h0 ? ZERO64[23] : p1_array_1507_comb[23];
  assign p1_sel_1508_comb[24] = p0_is_enable == 1'h0 ? ZERO64[24] : p1_array_1507_comb[24];
  assign p1_sel_1508_comb[25] = p0_is_enable == 1'h0 ? ZERO64[25] : p1_array_1507_comb[25];
  assign p1_sel_1508_comb[26] = p0_is_enable == 1'h0 ? ZERO64[26] : p1_array_1507_comb[26];
  assign p1_sel_1508_comb[27] = p0_is_enable == 1'h0 ? ZERO64[27] : p1_array_1507_comb[27];
  assign p1_sel_1508_comb[28] = p0_is_enable == 1'h0 ? ZERO64[28] : p1_array_1507_comb[28];
  assign p1_sel_1508_comb[29] = p0_is_enable == 1'h0 ? ZERO64[29] : p1_array_1507_comb[29];
  assign p1_sel_1508_comb[30] = p0_is_enable == 1'h0 ? ZERO64[30] : p1_array_1507_comb[30];
  assign p1_sel_1508_comb[31] = p0_is_enable == 1'h0 ? ZERO64[31] : p1_array_1507_comb[31];
  assign p1_sel_1508_comb[32] = p0_is_enable == 1'h0 ? ZERO64[32] : p1_array_1507_comb[32];
  assign p1_sel_1508_comb[33] = p0_is_enable == 1'h0 ? ZERO64[33] : p1_array_1507_comb[33];
  assign p1_sel_1508_comb[34] = p0_is_enable == 1'h0 ? ZERO64[34] : p1_array_1507_comb[34];
  assign p1_sel_1508_comb[35] = p0_is_enable == 1'h0 ? ZERO64[35] : p1_array_1507_comb[35];
  assign p1_sel_1508_comb[36] = p0_is_enable == 1'h0 ? ZERO64[36] : p1_array_1507_comb[36];
  assign p1_sel_1508_comb[37] = p0_is_enable == 1'h0 ? ZERO64[37] : p1_array_1507_comb[37];
  assign p1_sel_1508_comb[38] = p0_is_enable == 1'h0 ? ZERO64[38] : p1_array_1507_comb[38];
  assign p1_sel_1508_comb[39] = p0_is_enable == 1'h0 ? ZERO64[39] : p1_array_1507_comb[39];
  assign p1_sel_1508_comb[40] = p0_is_enable == 1'h0 ? ZERO64[40] : p1_array_1507_comb[40];
  assign p1_sel_1508_comb[41] = p0_is_enable == 1'h0 ? ZERO64[41] : p1_array_1507_comb[41];
  assign p1_sel_1508_comb[42] = p0_is_enable == 1'h0 ? ZERO64[42] : p1_array_1507_comb[42];
  assign p1_sel_1508_comb[43] = p0_is_enable == 1'h0 ? ZERO64[43] : p1_array_1507_comb[43];
  assign p1_sel_1508_comb[44] = p0_is_enable == 1'h0 ? ZERO64[44] : p1_array_1507_comb[44];
  assign p1_sel_1508_comb[45] = p0_is_enable == 1'h0 ? ZERO64[45] : p1_array_1507_comb[45];
  assign p1_sel_1508_comb[46] = p0_is_enable == 1'h0 ? ZERO64[46] : p1_array_1507_comb[46];
  assign p1_sel_1508_comb[47] = p0_is_enable == 1'h0 ? ZERO64[47] : p1_array_1507_comb[47];
  assign p1_sel_1508_comb[48] = p0_is_enable == 1'h0 ? ZERO64[48] : p1_array_1507_comb[48];
  assign p1_sel_1508_comb[49] = p0_is_enable == 1'h0 ? ZERO64[49] : p1_array_1507_comb[49];
  assign p1_sel_1508_comb[50] = p0_is_enable == 1'h0 ? ZERO64[50] : p1_array_1507_comb[50];
  assign p1_sel_1508_comb[51] = p0_is_enable == 1'h0 ? ZERO64[51] : p1_array_1507_comb[51];
  assign p1_sel_1508_comb[52] = p0_is_enable == 1'h0 ? ZERO64[52] : p1_array_1507_comb[52];
  assign p1_sel_1508_comb[53] = p0_is_enable == 1'h0 ? ZERO64[53] : p1_array_1507_comb[53];
  assign p1_sel_1508_comb[54] = p0_is_enable == 1'h0 ? ZERO64[54] : p1_array_1507_comb[54];
  assign p1_sel_1508_comb[55] = p0_is_enable == 1'h0 ? ZERO64[55] : p1_array_1507_comb[55];
  assign p1_sel_1508_comb[56] = p0_is_enable == 1'h0 ? ZERO64[56] : p1_array_1507_comb[56];
  assign p1_sel_1508_comb[57] = p0_is_enable == 1'h0 ? ZERO64[57] : p1_array_1507_comb[57];
  assign p1_sel_1508_comb[58] = p0_is_enable == 1'h0 ? ZERO64[58] : p1_array_1507_comb[58];
  assign p1_sel_1508_comb[59] = p0_is_enable == 1'h0 ? ZERO64[59] : p1_array_1507_comb[59];
  assign p1_sel_1508_comb[60] = p0_is_enable == 1'h0 ? ZERO64[60] : p1_array_1507_comb[60];
  assign p1_sel_1508_comb[61] = p0_is_enable == 1'h0 ? ZERO64[61] : p1_array_1507_comb[61];
  assign p1_sel_1508_comb[62] = p0_is_enable == 1'h0 ? ZERO64[62] : p1_array_1507_comb[62];
  assign p1_sel_1508_comb[63] = p0_is_enable == 1'h0 ? ZERO64[63] : p1_array_1507_comb[63];

  // Registers for pipe stage 1:
  reg [9:0] p1_sel_1508[0:63];
  always @ (posedge clk) begin
    p1_sel_1508[0] <= p1_sel_1508_comb[0];
    p1_sel_1508[1] <= p1_sel_1508_comb[1];
    p1_sel_1508[2] <= p1_sel_1508_comb[2];
    p1_sel_1508[3] <= p1_sel_1508_comb[3];
    p1_sel_1508[4] <= p1_sel_1508_comb[4];
    p1_sel_1508[5] <= p1_sel_1508_comb[5];
    p1_sel_1508[6] <= p1_sel_1508_comb[6];
    p1_sel_1508[7] <= p1_sel_1508_comb[7];
    p1_sel_1508[8] <= p1_sel_1508_comb[8];
    p1_sel_1508[9] <= p1_sel_1508_comb[9];
    p1_sel_1508[10] <= p1_sel_1508_comb[10];
    p1_sel_1508[11] <= p1_sel_1508_comb[11];
    p1_sel_1508[12] <= p1_sel_1508_comb[12];
    p1_sel_1508[13] <= p1_sel_1508_comb[13];
    p1_sel_1508[14] <= p1_sel_1508_comb[14];
    p1_sel_1508[15] <= p1_sel_1508_comb[15];
    p1_sel_1508[16] <= p1_sel_1508_comb[16];
    p1_sel_1508[17] <= p1_sel_1508_comb[17];
    p1_sel_1508[18] <= p1_sel_1508_comb[18];
    p1_sel_1508[19] <= p1_sel_1508_comb[19];
    p1_sel_1508[20] <= p1_sel_1508_comb[20];
    p1_sel_1508[21] <= p1_sel_1508_comb[21];
    p1_sel_1508[22] <= p1_sel_1508_comb[22];
    p1_sel_1508[23] <= p1_sel_1508_comb[23];
    p1_sel_1508[24] <= p1_sel_1508_comb[24];
    p1_sel_1508[25] <= p1_sel_1508_comb[25];
    p1_sel_1508[26] <= p1_sel_1508_comb[26];
    p1_sel_1508[27] <= p1_sel_1508_comb[27];
    p1_sel_1508[28] <= p1_sel_1508_comb[28];
    p1_sel_1508[29] <= p1_sel_1508_comb[29];
    p1_sel_1508[30] <= p1_sel_1508_comb[30];
    p1_sel_1508[31] <= p1_sel_1508_comb[31];
    p1_sel_1508[32] <= p1_sel_1508_comb[32];
    p1_sel_1508[33] <= p1_sel_1508_comb[33];
    p1_sel_1508[34] <= p1_sel_1508_comb[34];
    p1_sel_1508[35] <= p1_sel_1508_comb[35];
    p1_sel_1508[36] <= p1_sel_1508_comb[36];
    p1_sel_1508[37] <= p1_sel_1508_comb[37];
    p1_sel_1508[38] <= p1_sel_1508_comb[38];
    p1_sel_1508[39] <= p1_sel_1508_comb[39];
    p1_sel_1508[40] <= p1_sel_1508_comb[40];
    p1_sel_1508[41] <= p1_sel_1508_comb[41];
    p1_sel_1508[42] <= p1_sel_1508_comb[42];
    p1_sel_1508[43] <= p1_sel_1508_comb[43];
    p1_sel_1508[44] <= p1_sel_1508_comb[44];
    p1_sel_1508[45] <= p1_sel_1508_comb[45];
    p1_sel_1508[46] <= p1_sel_1508_comb[46];
    p1_sel_1508[47] <= p1_sel_1508_comb[47];
    p1_sel_1508[48] <= p1_sel_1508_comb[48];
    p1_sel_1508[49] <= p1_sel_1508_comb[49];
    p1_sel_1508[50] <= p1_sel_1508_comb[50];
    p1_sel_1508[51] <= p1_sel_1508_comb[51];
    p1_sel_1508[52] <= p1_sel_1508_comb[52];
    p1_sel_1508[53] <= p1_sel_1508_comb[53];
    p1_sel_1508[54] <= p1_sel_1508_comb[54];
    p1_sel_1508[55] <= p1_sel_1508_comb[55];
    p1_sel_1508[56] <= p1_sel_1508_comb[56];
    p1_sel_1508[57] <= p1_sel_1508_comb[57];
    p1_sel_1508[58] <= p1_sel_1508_comb[58];
    p1_sel_1508[59] <= p1_sel_1508_comb[59];
    p1_sel_1508[60] <= p1_sel_1508_comb[60];
    p1_sel_1508[61] <= p1_sel_1508_comb[61];
    p1_sel_1508[62] <= p1_sel_1508_comb[62];
    p1_sel_1508[63] <= p1_sel_1508_comb[63];
  end
  assign out = {p1_sel_1508[63], p1_sel_1508[62], p1_sel_1508[61], p1_sel_1508[60], p1_sel_1508[59], p1_sel_1508[58], p1_sel_1508[57], p1_sel_1508[56], p1_sel_1508[55], p1_sel_1508[54], p1_sel_1508[53], p1_sel_1508[52], p1_sel_1508[51], p1_sel_1508[50], p1_sel_1508[49], p1_sel_1508[48], p1_sel_1508[47], p1_sel_1508[46], p1_sel_1508[45], p1_sel_1508[44], p1_sel_1508[43], p1_sel_1508[42], p1_sel_1508[41], p1_sel_1508[40], p1_sel_1508[39], p1_sel_1508[38], p1_sel_1508[37], p1_sel_1508[36], p1_sel_1508[35], p1_sel_1508[34], p1_sel_1508[33], p1_sel_1508[32], p1_sel_1508[31], p1_sel_1508[30], p1_sel_1508[29], p1_sel_1508[28], p1_sel_1508[27], p1_sel_1508[26], p1_sel_1508[25], p1_sel_1508[24], p1_sel_1508[23], p1_sel_1508[22], p1_sel_1508[21], p1_sel_1508[20], p1_sel_1508[19], p1_sel_1508[18], p1_sel_1508[17], p1_sel_1508[16], p1_sel_1508[15], p1_sel_1508[14], p1_sel_1508[13], p1_sel_1508[12], p1_sel_1508[11], p1_sel_1508[10], p1_sel_1508[9], p1_sel_1508[8], p1_sel_1508[7], p1_sel_1508[6], p1_sel_1508[5], p1_sel_1508[4], p1_sel_1508[3], p1_sel_1508[2], p1_sel_1508[1], p1_sel_1508[0]};
endmodule
