module dct_1d_s10(
  input wire clk,
  input wire [79:0] x,
  output wire [79:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [15:0] smul16b_8b_x_9b (input reg [7:0] lhs, input reg [8:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [15:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul16b_8b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_8b (input reg [7:0] lhs, input reg [7:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_6b (input reg [7:0] lhs, input reg [5:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [23:0] umul24b_24b_x_7b (input reg [23:0] lhs, input reg [6:0] rhs);
    begin
      umul24b_24b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [9:0] x_unflattened[0:7];
  assign x_unflattened[0] = x[9:0];
  assign x_unflattened[1] = x[19:10];
  assign x_unflattened[2] = x[29:20];
  assign x_unflattened[3] = x[39:30];
  assign x_unflattened[4] = x[49:40];
  assign x_unflattened[5] = x[59:50];
  assign x_unflattened[6] = x[69:60];
  assign x_unflattened[7] = x[79:70];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_x[0:7];
  always @ (posedge clk) begin
    p0_x[0] <= x_unflattened[0];
    p0_x[1] <= x_unflattened[1];
    p0_x[2] <= x_unflattened[2];
    p0_x[3] <= x_unflattened[3];
    p0_x[4] <= x_unflattened[4];
    p0_x[5] <= x_unflattened[5];
    p0_x[6] <= x_unflattened[6];
    p0_x[7] <= x_unflattened[7];
  end

  // ===== Pipe stage 1:
  wire [9:0] p1_array_index_5797_comb;
  wire [9:0] p1_array_index_5798_comb;
  wire [9:0] p1_array_index_5799_comb;
  wire [9:0] p1_array_index_5800_comb;
  wire [9:0] p1_array_index_5801_comb;
  wire [9:0] p1_array_index_5802_comb;
  wire [9:0] p1_array_index_5803_comb;
  wire [9:0] p1_array_index_5804_comb;
  wire [7:0] p1_concat_5829_comb;
  wire [7:0] p1_concat_5831_comb;
  wire [7:0] p1_concat_5833_comb;
  wire [7:0] p1_concat_5835_comb;
  wire [7:0] p1_concat_5838_comb;
  wire [7:0] p1_concat_5840_comb;
  wire [7:0] p1_concat_5844_comb;
  wire [7:0] p1_concat_5846_comb;
  wire [15:0] p1_smul_3154_NarrowedMult__comb;
  wire [15:0] p1_smul_3153_NarrowedMult__comb;
  wire [15:0] p1_smul_3148_NarrowedMult__comb;
  wire [15:0] p1_smul_3147_NarrowedMult__comb;
  wire [15:0] p1_smul_3146_NarrowedMult__comb;
  wire [15:0] p1_smul_3144_NarrowedMult__comb;
  wire [15:0] p1_smul_3141_NarrowedMult__comb;
  wire [15:0] p1_smul_3139_NarrowedMult__comb;
  wire [15:0] p1_smul_3129_NarrowedMult__comb;
  wire [15:0] p1_smul_3127_NarrowedMult__comb;
  wire [15:0] p1_smul_3126_NarrowedMult__comb;
  wire [15:0] p1_smul_3124_NarrowedMult__comb;
  wire [15:0] p1_smul_3120_NarrowedMult__comb;
  wire [15:0] p1_smul_3119_NarrowedMult__comb;
  wire [15:0] p1_smul_3118_NarrowedMult__comb;
  wire [15:0] p1_smul_3117_NarrowedMult__comb;
  wire [14:0] p1_smul_3113_NarrowedMult__comb;
  wire [14:0] p1_smul_3112_NarrowedMult__comb;
  wire [14:0] p1_smul_3109_NarrowedMult__comb;
  wire [14:0] p1_smul_3108_NarrowedMult__comb;
  wire [14:0] p1_smul_3106_NarrowedMult__comb;
  wire [14:0] p1_smul_3104_NarrowedMult__comb;
  wire [14:0] p1_smul_3101_NarrowedMult__comb;
  wire [14:0] p1_smul_3099_NarrowedMult__comb;
  wire [14:0] p1_smul_3152_NarrowedMult__comb;
  wire [13:0] p1_smul_3168_NarrowedMult__comb;
  wire [13:0] p1_smul_3170_NarrowedMult__comb;
  wire [14:0] p1_smul_3149_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_5909_comb;
  wire [13:0] p1_smul_3189_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_5911_comb;
  wire [14:0] p1_smul_3143_NarrowedMult__comb;
  wire [14:0] p1_smul_3142_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_5914_comb;
  wire [13:0] p1_smul_3209_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_5916_comb;
  wire [14:0] p1_smul_3130_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_5926_comb;
  wire [13:0] p1_smul_3256_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_5928_comb;
  wire [14:0] p1_bit_slice_5929_comb;
  wire [13:0] p1_smul_3266_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_5931_comb;
  wire [14:0] p1_smul_3123_NarrowedMult__comb;
  wire [13:0] p1_smul_3277_NarrowedMult__comb;
  wire [14:0] p1_smul_3121_NarrowedMult__comb;
  wire [14:0] p1_smul_3116_NarrowedMult__comb;
  wire [13:0] p1_smul_3305_NarrowedMult__comb;
  wire [13:0] p1_smul_3114_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_5956_comb;
  wire [13:0] p1_bit_slice_5957_comb;
  wire [13:0] p1_smul_3111_NarrowedMult__comb;
  wire [13:0] p1_smul_3110_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_5960_comb;
  wire [13:0] p1_bit_slice_5961_comb;
  wire [13:0] p1_smul_3107_NarrowedMult__comb;
  wire [15:0] p1_smul_3138_NarrowedMult__comb;
  wire [15:0] p1_smul_3137_NarrowedMult__comb;
  wire [15:0] p1_smul_3136_NarrowedMult__comb;
  wire [15:0] p1_smul_3135_NarrowedMult__comb;
  wire [15:0] p1_smul_3134_NarrowedMult__comb;
  wire [15:0] p1_smul_3133_NarrowedMult__comb;
  wire [15:0] p1_smul_3132_NarrowedMult__comb;
  wire [15:0] p1_smul_3131_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_5987_comb;
  wire [13:0] p1_smul_3105_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_5989_comb;
  wire [13:0] p1_smul_3103_NarrowedMult__comb;
  wire [13:0] p1_smul_3102_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_5992_comb;
  wire [13:0] p1_smul_3100_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_5994_comb;
  wire [16:0] p1_add_5949_comb;
  wire [16:0] p1_add_5954_comb;
  wire [16:0] p1_add_5997_comb;
  wire [16:0] p1_add_5998_comb;
  wire [15:0] p1_bit_slice_6009_comb;
  wire [15:0] p1_add_6010_comb;
  wire [15:0] p1_add_6011_comb;
  wire [15:0] p1_bit_slice_6012_comb;
  wire [15:0] p1_add_6021_comb;
  wire p1_bit_slice_6022_comb;
  wire [15:0] p1_add_6023_comb;
  wire p1_bit_slice_6024_comb;
  wire [15:0] p1_add_6025_comb;
  wire p1_bit_slice_6026_comb;
  wire [15:0] p1_add_6027_comb;
  wire p1_bit_slice_6028_comb;
  wire [15:0] p1_add_6037_comb;
  wire p1_bit_slice_6038_comb;
  wire [15:0] p1_add_6039_comb;
  wire p1_bit_slice_6040_comb;
  wire [15:0] p1_add_6041_comb;
  wire p1_bit_slice_6042_comb;
  wire [15:0] p1_add_6043_comb;
  wire p1_bit_slice_6044_comb;
  wire [15:0] p1_add_6053_comb;
  wire [15:0] p1_bit_slice_6054_comb;
  wire [15:0] p1_bit_slice_6055_comb;
  wire [15:0] p1_add_6056_comb;
  wire [8:0] p1_add_6057_comb;
  wire [8:0] p1_add_6058_comb;
  wire [8:0] p1_add_6059_comb;
  wire [8:0] p1_add_6060_comb;
  wire [14:0] p1_add_6061_comb;
  wire p1_bit_slice_6062_comb;
  wire [14:0] p1_add_6063_comb;
  wire p1_bit_slice_6064_comb;
  wire [14:0] p1_add_6065_comb;
  wire p1_bit_slice_6066_comb;
  wire [14:0] p1_add_6067_comb;
  wire p1_bit_slice_6068_comb;
  wire [16:0] p1_add_6069_comb;
  wire [16:0] p1_add_6070_comb;
  wire [16:0] p1_add_6071_comb;
  wire [16:0] p1_add_6072_comb;
  wire [14:0] p1_add_6073_comb;
  wire p1_bit_slice_6074_comb;
  wire [14:0] p1_add_6075_comb;
  wire p1_bit_slice_6076_comb;
  wire [14:0] p1_add_6077_comb;
  wire p1_bit_slice_6078_comb;
  wire [14:0] p1_add_6079_comb;
  wire p1_bit_slice_6080_comb;
  wire p1_bit_slice_6081_comb;
  wire p1_bit_slice_6082_comb;
  wire p1_bit_slice_6083_comb;
  wire p1_bit_slice_6084_comb;
  assign p1_array_index_5797_comb = p0_x[3'h0];
  assign p1_array_index_5798_comb = p0_x[3'h1];
  assign p1_array_index_5799_comb = p0_x[3'h6];
  assign p1_array_index_5800_comb = p0_x[3'h7];
  assign p1_array_index_5801_comb = p0_x[3'h2];
  assign p1_array_index_5802_comb = p0_x[3'h5];
  assign p1_array_index_5803_comb = p0_x[3'h3];
  assign p1_array_index_5804_comb = p0_x[3'h4];
  assign p1_concat_5829_comb = {~p1_array_index_5797_comb[7], p1_array_index_5797_comb[6:0]};
  assign p1_concat_5831_comb = {~p1_array_index_5798_comb[7], p1_array_index_5798_comb[6:0]};
  assign p1_concat_5833_comb = {~p1_array_index_5799_comb[7], p1_array_index_5799_comb[6:0]};
  assign p1_concat_5835_comb = {~p1_array_index_5800_comb[7], p1_array_index_5800_comb[6:0]};
  assign p1_concat_5838_comb = {~p1_array_index_5801_comb[7], p1_array_index_5801_comb[6:0]};
  assign p1_concat_5840_comb = {~p1_array_index_5802_comb[7], p1_array_index_5802_comb[6:0]};
  assign p1_concat_5844_comb = {~p1_array_index_5803_comb[7], p1_array_index_5803_comb[6:0]};
  assign p1_concat_5846_comb = {~p1_array_index_5804_comb[7], p1_array_index_5804_comb[6:0]};
  assign p1_smul_3154_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5829_comb, 9'h0fb);
  assign p1_smul_3153_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5831_comb, 9'h0d5);
  assign p1_smul_3148_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5833_comb, 9'h12b);
  assign p1_smul_3147_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5835_comb, 9'h105);
  assign p1_smul_3146_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5829_comb, 9'h0d5);
  assign p1_smul_3144_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5838_comb, 9'h105);
  assign p1_smul_3141_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5840_comb, 9'h0fb);
  assign p1_smul_3139_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5835_comb, 9'h12b);
  assign p1_smul_3129_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5831_comb, 9'h105);
  assign p1_smul_3127_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5844_comb, 9'h0d5);
  assign p1_smul_3126_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5846_comb, 9'h0d5);
  assign p1_smul_3124_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5833_comb, 9'h105);
  assign p1_smul_3120_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5838_comb, 9'h0d5);
  assign p1_smul_3119_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5844_comb, 9'h105);
  assign p1_smul_3118_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5846_comb, 9'h105);
  assign p1_smul_3117_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5840_comb, 9'h0d5);
  assign p1_smul_3113_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5831_comb, 7'h31);
  assign p1_smul_3112_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5838_comb, 7'h4f);
  assign p1_smul_3109_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5840_comb, 7'h4f);
  assign p1_smul_3108_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5833_comb, 7'h31);
  assign p1_smul_3106_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5829_comb, 7'h31);
  assign p1_smul_3104_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5838_comb, 7'h31);
  assign p1_smul_3101_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5840_comb, 7'h31);
  assign p1_smul_3099_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5835_comb, 7'h31);
  assign p1_smul_3152_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5838_comb, 8'h47);
  assign p1_smul_3168_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5844_comb, 6'h19);
  assign p1_smul_3170_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5846_comb, 6'h27);
  assign p1_smul_3149_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5840_comb, 8'hb9);
  assign p1_bit_slice_5909_comb = p1_smul_3146_NarrowedMult__comb[15:1];
  assign p1_smul_3189_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5831_comb, 6'h27);
  assign p1_bit_slice_5911_comb = p1_smul_3144_NarrowedMult__comb[15:1];
  assign p1_smul_3143_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5844_comb, 8'hb9);
  assign p1_smul_3142_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5846_comb, 8'h47);
  assign p1_bit_slice_5914_comb = p1_smul_3141_NarrowedMult__comb[15:1];
  assign p1_smul_3209_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5833_comb, 6'h19);
  assign p1_bit_slice_5916_comb = p1_smul_3139_NarrowedMult__comb[15:1];
  assign p1_smul_3130_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5829_comb, 8'h47);
  assign p1_bit_slice_5926_comb = p1_smul_3129_NarrowedMult__comb[15:1];
  assign p1_smul_3256_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5838_comb, 6'h27);
  assign p1_bit_slice_5928_comb = p1_smul_3127_NarrowedMult__comb[15:1];
  assign p1_bit_slice_5929_comb = p1_smul_3126_NarrowedMult__comb[15:1];
  assign p1_smul_3266_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5840_comb, 6'h27);
  assign p1_bit_slice_5931_comb = p1_smul_3124_NarrowedMult__comb[15:1];
  assign p1_smul_3123_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5835_comb, 8'h47);
  assign p1_smul_3277_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5829_comb, 6'h19);
  assign p1_smul_3121_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5831_comb, 8'hb9);
  assign p1_smul_3116_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5833_comb, 8'hb9);
  assign p1_smul_3305_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5835_comb, 6'h19);
  assign p1_smul_3114_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5829_comb, 7'h3b);
  assign p1_bit_slice_5956_comb = p1_smul_3113_NarrowedMult__comb[14:1];
  assign p1_bit_slice_5957_comb = p1_smul_3112_NarrowedMult__comb[14:1];
  assign p1_smul_3111_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5844_comb, 7'h45);
  assign p1_smul_3110_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5846_comb, 7'h45);
  assign p1_bit_slice_5960_comb = p1_smul_3109_NarrowedMult__comb[14:1];
  assign p1_bit_slice_5961_comb = p1_smul_3108_NarrowedMult__comb[14:1];
  assign p1_smul_3107_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5835_comb, 7'h3b);
  assign p1_smul_3138_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5829_comb, 9'h0b5);
  assign p1_smul_3137_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5831_comb, 9'h14b);
  assign p1_smul_3136_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5838_comb, 9'h14b);
  assign p1_smul_3135_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5844_comb, 9'h0b5);
  assign p1_smul_3134_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5846_comb, 9'h0b5);
  assign p1_smul_3133_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5840_comb, 9'h14b);
  assign p1_smul_3132_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5833_comb, 9'h14b);
  assign p1_smul_3131_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5835_comb, 9'h0b5);
  assign p1_bit_slice_5987_comb = p1_smul_3106_NarrowedMult__comb[14:1];
  assign p1_smul_3105_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5831_comb, 7'h45);
  assign p1_bit_slice_5989_comb = p1_smul_3104_NarrowedMult__comb[14:1];
  assign p1_smul_3103_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5844_comb, 7'h3b);
  assign p1_smul_3102_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5846_comb, 7'h3b);
  assign p1_bit_slice_5992_comb = p1_smul_3101_NarrowedMult__comb[14:1];
  assign p1_smul_3100_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5833_comb, 7'h45);
  assign p1_bit_slice_5994_comb = p1_smul_3099_NarrowedMult__comb[14:1];
  assign p1_add_5949_comb = {{1{p1_smul_3154_NarrowedMult__comb[15]}}, p1_smul_3154_NarrowedMult__comb} + {{1{p1_smul_3153_NarrowedMult__comb[15]}}, p1_smul_3153_NarrowedMult__comb};
  assign p1_add_5954_comb = {{1{p1_smul_3148_NarrowedMult__comb[15]}}, p1_smul_3148_NarrowedMult__comb} + {{1{p1_smul_3147_NarrowedMult__comb[15]}}, p1_smul_3147_NarrowedMult__comb};
  assign p1_add_5997_comb = {{1{p1_smul_3120_NarrowedMult__comb[15]}}, p1_smul_3120_NarrowedMult__comb} + {{1{p1_smul_3119_NarrowedMult__comb[15]}}, p1_smul_3119_NarrowedMult__comb};
  assign p1_add_5998_comb = {{1{p1_smul_3118_NarrowedMult__comb[15]}}, p1_smul_3118_NarrowedMult__comb} + {{1{p1_smul_3117_NarrowedMult__comb[15]}}, p1_smul_3117_NarrowedMult__comb};
  assign p1_bit_slice_6009_comb = p1_add_5949_comb[16:1];
  assign p1_add_6010_comb = {{1{p1_smul_3152_NarrowedMult__comb[14]}}, p1_smul_3152_NarrowedMult__comb} + {{2{p1_smul_3168_NarrowedMult__comb[13]}}, p1_smul_3168_NarrowedMult__comb};
  assign p1_add_6011_comb = {{2{p1_smul_3170_NarrowedMult__comb[13]}}, p1_smul_3170_NarrowedMult__comb} + {{1{p1_smul_3149_NarrowedMult__comb[14]}}, p1_smul_3149_NarrowedMult__comb};
  assign p1_bit_slice_6012_comb = p1_add_5954_comb[16:1];
  assign p1_add_6021_comb = {{1{p1_bit_slice_5909_comb[14]}}, p1_bit_slice_5909_comb} + {{2{p1_smul_3189_NarrowedMult__comb[13]}}, p1_smul_3189_NarrowedMult__comb};
  assign p1_bit_slice_6022_comb = p1_smul_3146_NarrowedMult__comb[0];
  assign p1_add_6023_comb = {{1{p1_bit_slice_5911_comb[14]}}, p1_bit_slice_5911_comb} + {{1{p1_smul_3143_NarrowedMult__comb[14]}}, p1_smul_3143_NarrowedMult__comb};
  assign p1_bit_slice_6024_comb = p1_smul_3144_NarrowedMult__comb[0];
  assign p1_add_6025_comb = {{1{p1_smul_3142_NarrowedMult__comb[14]}}, p1_smul_3142_NarrowedMult__comb} + {{1{p1_bit_slice_5914_comb[14]}}, p1_bit_slice_5914_comb};
  assign p1_bit_slice_6026_comb = p1_smul_3141_NarrowedMult__comb[0];
  assign p1_add_6027_comb = {{2{p1_smul_3209_NarrowedMult__comb[13]}}, p1_smul_3209_NarrowedMult__comb} + {{1{p1_bit_slice_5916_comb[14]}}, p1_bit_slice_5916_comb};
  assign p1_bit_slice_6028_comb = p1_smul_3139_NarrowedMult__comb[0];
  assign p1_add_6037_comb = {{1{p1_smul_3130_NarrowedMult__comb[14]}}, p1_smul_3130_NarrowedMult__comb} + {{1{p1_bit_slice_5926_comb[14]}}, p1_bit_slice_5926_comb};
  assign p1_bit_slice_6038_comb = p1_smul_3129_NarrowedMult__comb[0];
  assign p1_add_6039_comb = {{2{p1_smul_3256_NarrowedMult__comb[13]}}, p1_smul_3256_NarrowedMult__comb} + {{1{p1_bit_slice_5928_comb[14]}}, p1_bit_slice_5928_comb};
  assign p1_bit_slice_6040_comb = p1_smul_3127_NarrowedMult__comb[0];
  assign p1_add_6041_comb = {{1{p1_bit_slice_5929_comb[14]}}, p1_bit_slice_5929_comb} + {{2{p1_smul_3266_NarrowedMult__comb[13]}}, p1_smul_3266_NarrowedMult__comb};
  assign p1_bit_slice_6042_comb = p1_smul_3126_NarrowedMult__comb[0];
  assign p1_add_6043_comb = {{1{p1_bit_slice_5931_comb[14]}}, p1_bit_slice_5931_comb} + {{1{p1_smul_3123_NarrowedMult__comb[14]}}, p1_smul_3123_NarrowedMult__comb};
  assign p1_bit_slice_6044_comb = p1_smul_3124_NarrowedMult__comb[0];
  assign p1_add_6053_comb = {{2{p1_smul_3277_NarrowedMult__comb[13]}}, p1_smul_3277_NarrowedMult__comb} + {{1{p1_smul_3121_NarrowedMult__comb[14]}}, p1_smul_3121_NarrowedMult__comb};
  assign p1_bit_slice_6054_comb = p1_add_5997_comb[16:1];
  assign p1_bit_slice_6055_comb = p1_add_5998_comb[16:1];
  assign p1_add_6056_comb = {{1{p1_smul_3116_NarrowedMult__comb[14]}}, p1_smul_3116_NarrowedMult__comb} + {{2{p1_smul_3305_NarrowedMult__comb[13]}}, p1_smul_3305_NarrowedMult__comb};
  assign p1_add_6057_comb = {{1{p1_concat_5829_comb[7]}}, p1_concat_5829_comb} + {{1{p1_concat_5831_comb[7]}}, p1_concat_5831_comb};
  assign p1_add_6058_comb = {{1{p1_concat_5838_comb[7]}}, p1_concat_5838_comb} + {{1{p1_concat_5844_comb[7]}}, p1_concat_5844_comb};
  assign p1_add_6059_comb = {{1{p1_concat_5846_comb[7]}}, p1_concat_5846_comb} + {{1{p1_concat_5840_comb[7]}}, p1_concat_5840_comb};
  assign p1_add_6060_comb = {{1{p1_concat_5833_comb[7]}}, p1_concat_5833_comb} + {{1{p1_concat_5835_comb[7]}}, p1_concat_5835_comb};
  assign p1_add_6061_comb = {{1{p1_smul_3114_NarrowedMult__comb[13]}}, p1_smul_3114_NarrowedMult__comb} + {{1{p1_bit_slice_5956_comb[13]}}, p1_bit_slice_5956_comb};
  assign p1_bit_slice_6062_comb = p1_smul_3113_NarrowedMult__comb[0];
  assign p1_add_6063_comb = {{1{p1_bit_slice_5957_comb[13]}}, p1_bit_slice_5957_comb} + {{1{p1_smul_3111_NarrowedMult__comb[13]}}, p1_smul_3111_NarrowedMult__comb};
  assign p1_bit_slice_6064_comb = p1_smul_3112_NarrowedMult__comb[0];
  assign p1_add_6065_comb = {{1{p1_smul_3110_NarrowedMult__comb[13]}}, p1_smul_3110_NarrowedMult__comb} + {{1{p1_bit_slice_5960_comb[13]}}, p1_bit_slice_5960_comb};
  assign p1_bit_slice_6066_comb = p1_smul_3109_NarrowedMult__comb[0];
  assign p1_add_6067_comb = {{1{p1_bit_slice_5961_comb[13]}}, p1_bit_slice_5961_comb} + {{1{p1_smul_3107_NarrowedMult__comb[13]}}, p1_smul_3107_NarrowedMult__comb};
  assign p1_bit_slice_6068_comb = p1_smul_3108_NarrowedMult__comb[0];
  assign p1_add_6069_comb = {{1{p1_smul_3138_NarrowedMult__comb[15]}}, p1_smul_3138_NarrowedMult__comb} + {{1{p1_smul_3137_NarrowedMult__comb[15]}}, p1_smul_3137_NarrowedMult__comb};
  assign p1_add_6070_comb = {{1{p1_smul_3136_NarrowedMult__comb[15]}}, p1_smul_3136_NarrowedMult__comb} + {{1{p1_smul_3135_NarrowedMult__comb[15]}}, p1_smul_3135_NarrowedMult__comb};
  assign p1_add_6071_comb = {{1{p1_smul_3134_NarrowedMult__comb[15]}}, p1_smul_3134_NarrowedMult__comb} + {{1{p1_smul_3133_NarrowedMult__comb[15]}}, p1_smul_3133_NarrowedMult__comb};
  assign p1_add_6072_comb = {{1{p1_smul_3132_NarrowedMult__comb[15]}}, p1_smul_3132_NarrowedMult__comb} + {{1{p1_smul_3131_NarrowedMult__comb[15]}}, p1_smul_3131_NarrowedMult__comb};
  assign p1_add_6073_comb = {{1{p1_bit_slice_5987_comb[13]}}, p1_bit_slice_5987_comb} + {{1{p1_smul_3105_NarrowedMult__comb[13]}}, p1_smul_3105_NarrowedMult__comb};
  assign p1_bit_slice_6074_comb = p1_smul_3106_NarrowedMult__comb[0];
  assign p1_add_6075_comb = {{1{p1_bit_slice_5989_comb[13]}}, p1_bit_slice_5989_comb} + {{1{p1_smul_3103_NarrowedMult__comb[13]}}, p1_smul_3103_NarrowedMult__comb};
  assign p1_bit_slice_6076_comb = p1_smul_3104_NarrowedMult__comb[0];
  assign p1_add_6077_comb = {{1{p1_smul_3102_NarrowedMult__comb[13]}}, p1_smul_3102_NarrowedMult__comb} + {{1{p1_bit_slice_5992_comb[13]}}, p1_bit_slice_5992_comb};
  assign p1_bit_slice_6078_comb = p1_smul_3101_NarrowedMult__comb[0];
  assign p1_add_6079_comb = {{1{p1_smul_3100_NarrowedMult__comb[13]}}, p1_smul_3100_NarrowedMult__comb} + {{1{p1_bit_slice_5994_comb[13]}}, p1_bit_slice_5994_comb};
  assign p1_bit_slice_6080_comb = p1_smul_3099_NarrowedMult__comb[0];
  assign p1_bit_slice_6081_comb = p1_add_5949_comb[0];
  assign p1_bit_slice_6082_comb = p1_add_5954_comb[0];
  assign p1_bit_slice_6083_comb = p1_add_5997_comb[0];
  assign p1_bit_slice_6084_comb = p1_add_5998_comb[0];

  // Registers for pipe stage 1:
  reg [15:0] p1_bit_slice_6009;
  reg [15:0] p1_add_6010;
  reg [15:0] p1_add_6011;
  reg [15:0] p1_bit_slice_6012;
  reg [15:0] p1_add_6021;
  reg p1_bit_slice_6022;
  reg [15:0] p1_add_6023;
  reg p1_bit_slice_6024;
  reg [15:0] p1_add_6025;
  reg p1_bit_slice_6026;
  reg [15:0] p1_add_6027;
  reg p1_bit_slice_6028;
  reg [15:0] p1_add_6037;
  reg p1_bit_slice_6038;
  reg [15:0] p1_add_6039;
  reg p1_bit_slice_6040;
  reg [15:0] p1_add_6041;
  reg p1_bit_slice_6042;
  reg [15:0] p1_add_6043;
  reg p1_bit_slice_6044;
  reg [15:0] p1_add_6053;
  reg [15:0] p1_bit_slice_6054;
  reg [15:0] p1_bit_slice_6055;
  reg [15:0] p1_add_6056;
  reg [8:0] p1_add_6057;
  reg [8:0] p1_add_6058;
  reg [8:0] p1_add_6059;
  reg [8:0] p1_add_6060;
  reg [14:0] p1_add_6061;
  reg p1_bit_slice_6062;
  reg [14:0] p1_add_6063;
  reg p1_bit_slice_6064;
  reg [14:0] p1_add_6065;
  reg p1_bit_slice_6066;
  reg [14:0] p1_add_6067;
  reg p1_bit_slice_6068;
  reg [16:0] p1_add_6069;
  reg [16:0] p1_add_6070;
  reg [16:0] p1_add_6071;
  reg [16:0] p1_add_6072;
  reg [14:0] p1_add_6073;
  reg p1_bit_slice_6074;
  reg [14:0] p1_add_6075;
  reg p1_bit_slice_6076;
  reg [14:0] p1_add_6077;
  reg p1_bit_slice_6078;
  reg [14:0] p1_add_6079;
  reg p1_bit_slice_6080;
  reg p1_bit_slice_6081;
  reg p1_bit_slice_6082;
  reg p1_bit_slice_6083;
  reg p1_bit_slice_6084;
  always @ (posedge clk) begin
    p1_bit_slice_6009 <= p1_bit_slice_6009_comb;
    p1_add_6010 <= p1_add_6010_comb;
    p1_add_6011 <= p1_add_6011_comb;
    p1_bit_slice_6012 <= p1_bit_slice_6012_comb;
    p1_add_6021 <= p1_add_6021_comb;
    p1_bit_slice_6022 <= p1_bit_slice_6022_comb;
    p1_add_6023 <= p1_add_6023_comb;
    p1_bit_slice_6024 <= p1_bit_slice_6024_comb;
    p1_add_6025 <= p1_add_6025_comb;
    p1_bit_slice_6026 <= p1_bit_slice_6026_comb;
    p1_add_6027 <= p1_add_6027_comb;
    p1_bit_slice_6028 <= p1_bit_slice_6028_comb;
    p1_add_6037 <= p1_add_6037_comb;
    p1_bit_slice_6038 <= p1_bit_slice_6038_comb;
    p1_add_6039 <= p1_add_6039_comb;
    p1_bit_slice_6040 <= p1_bit_slice_6040_comb;
    p1_add_6041 <= p1_add_6041_comb;
    p1_bit_slice_6042 <= p1_bit_slice_6042_comb;
    p1_add_6043 <= p1_add_6043_comb;
    p1_bit_slice_6044 <= p1_bit_slice_6044_comb;
    p1_add_6053 <= p1_add_6053_comb;
    p1_bit_slice_6054 <= p1_bit_slice_6054_comb;
    p1_bit_slice_6055 <= p1_bit_slice_6055_comb;
    p1_add_6056 <= p1_add_6056_comb;
    p1_add_6057 <= p1_add_6057_comb;
    p1_add_6058 <= p1_add_6058_comb;
    p1_add_6059 <= p1_add_6059_comb;
    p1_add_6060 <= p1_add_6060_comb;
    p1_add_6061 <= p1_add_6061_comb;
    p1_bit_slice_6062 <= p1_bit_slice_6062_comb;
    p1_add_6063 <= p1_add_6063_comb;
    p1_bit_slice_6064 <= p1_bit_slice_6064_comb;
    p1_add_6065 <= p1_add_6065_comb;
    p1_bit_slice_6066 <= p1_bit_slice_6066_comb;
    p1_add_6067 <= p1_add_6067_comb;
    p1_bit_slice_6068 <= p1_bit_slice_6068_comb;
    p1_add_6069 <= p1_add_6069_comb;
    p1_add_6070 <= p1_add_6070_comb;
    p1_add_6071 <= p1_add_6071_comb;
    p1_add_6072 <= p1_add_6072_comb;
    p1_add_6073 <= p1_add_6073_comb;
    p1_bit_slice_6074 <= p1_bit_slice_6074_comb;
    p1_add_6075 <= p1_add_6075_comb;
    p1_bit_slice_6076 <= p1_bit_slice_6076_comb;
    p1_add_6077 <= p1_add_6077_comb;
    p1_bit_slice_6078 <= p1_bit_slice_6078_comb;
    p1_add_6079 <= p1_add_6079_comb;
    p1_bit_slice_6080 <= p1_bit_slice_6080_comb;
    p1_bit_slice_6081 <= p1_bit_slice_6081_comb;
    p1_bit_slice_6082 <= p1_bit_slice_6082_comb;
    p1_bit_slice_6083 <= p1_bit_slice_6083_comb;
    p1_bit_slice_6084 <= p1_bit_slice_6084_comb;
  end

  // ===== Pipe stage 2:
  wire [16:0] p2_concat_6193_comb;
  wire [16:0] p2_concat_6194_comb;
  wire [16:0] p2_concat_6195_comb;
  wire [16:0] p2_concat_6196_comb;
  wire [16:0] p2_concat_6197_comb;
  wire [16:0] p2_concat_6198_comb;
  wire [16:0] p2_concat_6199_comb;
  wire [16:0] p2_concat_6200_comb;
  wire [15:0] p2_concat_6211_comb;
  wire [15:0] p2_concat_6212_comb;
  wire [15:0] p2_concat_6213_comb;
  wire [15:0] p2_concat_6214_comb;
  wire [24:0] p2_sum__97_comb;
  wire [24:0] p2_sum__98_comb;
  wire [24:0] p2_sum__99_comb;
  wire [24:0] p2_sum__100_comb;
  wire [15:0] p2_concat_6227_comb;
  wire [15:0] p2_concat_6228_comb;
  wire [15:0] p2_concat_6229_comb;
  wire [15:0] p2_concat_6230_comb;
  wire [23:0] p2_add_6209_comb;
  wire [23:0] p2_add_6210_comb;
  wire [24:0] p2_sum__101_comb;
  wire [24:0] p2_sum__102_comb;
  wire [24:0] p2_sum__103_comb;
  wire [24:0] p2_sum__104_comb;
  wire [24:0] p2_sum__93_comb;
  wire [24:0] p2_sum__94_comb;
  wire [24:0] p2_sum__95_comb;
  wire [24:0] p2_sum__96_comb;
  wire [23:0] p2_add_6231_comb;
  wire [23:0] p2_add_6232_comb;
  wire [23:0] p2_add_6233_comb;
  wire [23:0] p2_add_6234_comb;
  wire [24:0] p2_sum__77_comb;
  wire [24:0] p2_sum__78_comb;
  wire [24:0] p2_sum__83_comb;
  wire [24:0] p2_sum__84_comb;
  wire [24:0] p2_sum__79_comb;
  wire [24:0] p2_sum__80_comb;
  wire [24:0] p2_sum__75_comb;
  wire [24:0] p2_sum__76_comb;
  wire [24:0] p2_sum__71_comb;
  wire [24:0] p2_sum__72_comb;
  wire [23:0] p2_add_6253_comb;
  wire [23:0] p2_add_6257_comb;
  wire [23:0] p2_add_6258_comb;
  wire [24:0] p2_sum__67_comb;
  wire [23:0] p2_add_6265_comb;
  wire [23:0] p2_add_6266_comb;
  wire [24:0] p2_sum__70_comb;
  wire [24:0] p2_sum__68_comb;
  wire [24:0] p2_sum__66_comb;
  wire [24:0] p2_sum__64_comb;
  wire [23:0] p2_umul_2636_NarrowedMult__comb;
  wire [23:0] p2_add_6271_comb;
  wire [24:0] p2_add_6273_comb;
  wire [23:0] p2_add_6275_comb;
  wire [24:0] p2_add_6270_comb;
  wire [24:0] p2_add_6272_comb;
  wire [24:0] p2_add_6274_comb;
  wire [24:0] p2_add_6276_comb;
  wire [16:0] p2_bit_slice_6277_comb;
  wire [16:0] p2_bit_slice_6279_comb;
  wire [16:0] p2_bit_slice_6281_comb;
  wire [16:0] p2_bit_slice_6283_comb;
  wire [16:0] p2_bit_slice_6278_comb;
  wire [16:0] p2_bit_slice_6280_comb;
  wire [16:0] p2_bit_slice_6282_comb;
  wire [16:0] p2_bit_slice_6284_comb;
  wire [17:0] p2_add_6301_comb;
  wire [17:0] p2_add_6303_comb;
  wire [17:0] p2_add_6305_comb;
  wire [17:0] p2_add_6307_comb;
  wire [17:0] p2_add_6302_comb;
  wire [17:0] p2_add_6304_comb;
  wire [17:0] p2_add_6306_comb;
  wire [17:0] p2_add_6308_comb;
  wire [9:0] p2_bit_slice_6309_comb;
  wire [9:0] p2_bit_slice_6310_comb;
  wire [9:0] p2_bit_slice_6311_comb;
  wire [9:0] p2_bit_slice_6312_comb;
  wire [6:0] p2_bit_slice_6313_comb;
  wire [6:0] p2_bit_slice_6314_comb;
  wire [6:0] p2_bit_slice_6315_comb;
  wire [6:0] p2_bit_slice_6316_comb;
  assign p2_concat_6193_comb = {p1_add_6021, p1_bit_slice_6022};
  assign p2_concat_6194_comb = {p1_add_6023, p1_bit_slice_6024};
  assign p2_concat_6195_comb = {p1_add_6025, p1_bit_slice_6026};
  assign p2_concat_6196_comb = {p1_add_6027, p1_bit_slice_6028};
  assign p2_concat_6197_comb = {p1_add_6037, p1_bit_slice_6038};
  assign p2_concat_6198_comb = {p1_add_6039, p1_bit_slice_6040};
  assign p2_concat_6199_comb = {p1_add_6041, p1_bit_slice_6042};
  assign p2_concat_6200_comb = {p1_add_6043, p1_bit_slice_6044};
  assign p2_concat_6211_comb = {p1_add_6061, p1_bit_slice_6062};
  assign p2_concat_6212_comb = {p1_add_6063, p1_bit_slice_6064};
  assign p2_concat_6213_comb = {p1_add_6065, p1_bit_slice_6066};
  assign p2_concat_6214_comb = {p1_add_6067, p1_bit_slice_6068};
  assign p2_sum__97_comb = {{8{p1_add_6069[16]}}, p1_add_6069};
  assign p2_sum__98_comb = {{8{p1_add_6070[16]}}, p1_add_6070};
  assign p2_sum__99_comb = {{8{p1_add_6071[16]}}, p1_add_6071};
  assign p2_sum__100_comb = {{8{p1_add_6072[16]}}, p1_add_6072};
  assign p2_concat_6227_comb = {p1_add_6073, p1_bit_slice_6074};
  assign p2_concat_6228_comb = {p1_add_6075, p1_bit_slice_6076};
  assign p2_concat_6229_comb = {p1_add_6077, p1_bit_slice_6078};
  assign p2_concat_6230_comb = {p1_add_6079, p1_bit_slice_6080};
  assign p2_add_6209_comb = {{8{p1_bit_slice_6009[15]}}, p1_bit_slice_6009} + {{8{p1_add_6010[15]}}, p1_add_6010};
  assign p2_add_6210_comb = {{8{p1_add_6011[15]}}, p1_add_6011} + {{8{p1_bit_slice_6012[15]}}, p1_bit_slice_6012};
  assign p2_sum__101_comb = {{8{p2_concat_6193_comb[16]}}, p2_concat_6193_comb};
  assign p2_sum__102_comb = {{8{p2_concat_6194_comb[16]}}, p2_concat_6194_comb};
  assign p2_sum__103_comb = {{8{p2_concat_6195_comb[16]}}, p2_concat_6195_comb};
  assign p2_sum__104_comb = {{8{p2_concat_6196_comb[16]}}, p2_concat_6196_comb};
  assign p2_sum__93_comb = {{8{p2_concat_6197_comb[16]}}, p2_concat_6197_comb};
  assign p2_sum__94_comb = {{8{p2_concat_6198_comb[16]}}, p2_concat_6198_comb};
  assign p2_sum__95_comb = {{8{p2_concat_6199_comb[16]}}, p2_concat_6199_comb};
  assign p2_sum__96_comb = {{8{p2_concat_6200_comb[16]}}, p2_concat_6200_comb};
  assign p2_add_6231_comb = {{8{p1_add_6053[15]}}, p1_add_6053} + {{8{p1_bit_slice_6054[15]}}, p1_bit_slice_6054};
  assign p2_add_6232_comb = {{8{p1_bit_slice_6055[15]}}, p1_bit_slice_6055} + {{8{p1_add_6056[15]}}, p1_add_6056};
  assign p2_add_6233_comb = {{15{p1_add_6057[8]}}, p1_add_6057} + {{15{p1_add_6058[8]}}, p1_add_6058};
  assign p2_add_6234_comb = {{15{p1_add_6059[8]}}, p1_add_6059} + {{15{p1_add_6060[8]}}, p1_add_6060};
  assign p2_sum__77_comb = p2_sum__97_comb + p2_sum__98_comb;
  assign p2_sum__78_comb = p2_sum__99_comb + p2_sum__100_comb;
  assign p2_sum__83_comb = {p2_add_6209_comb, p1_bit_slice_6081};
  assign p2_sum__84_comb = {p2_add_6210_comb, p1_bit_slice_6082};
  assign p2_sum__79_comb = p2_sum__101_comb + p2_sum__102_comb;
  assign p2_sum__80_comb = p2_sum__103_comb + p2_sum__104_comb;
  assign p2_sum__75_comb = p2_sum__93_comb + p2_sum__94_comb;
  assign p2_sum__76_comb = p2_sum__95_comb + p2_sum__96_comb;
  assign p2_sum__71_comb = {p2_add_6231_comb, p1_bit_slice_6083};
  assign p2_sum__72_comb = {p2_add_6232_comb, p1_bit_slice_6084};
  assign p2_add_6253_comb = p2_add_6233_comb + p2_add_6234_comb;
  assign p2_add_6257_comb = {{8{p2_concat_6211_comb[15]}}, p2_concat_6211_comb} + {{8{p2_concat_6212_comb[15]}}, p2_concat_6212_comb};
  assign p2_add_6258_comb = {{8{p2_concat_6213_comb[15]}}, p2_concat_6213_comb} + {{8{p2_concat_6214_comb[15]}}, p2_concat_6214_comb};
  assign p2_sum__67_comb = p2_sum__77_comb + p2_sum__78_comb;
  assign p2_add_6265_comb = {{8{p2_concat_6227_comb[15]}}, p2_concat_6227_comb} + {{8{p2_concat_6228_comb[15]}}, p2_concat_6228_comb};
  assign p2_add_6266_comb = {{8{p2_concat_6229_comb[15]}}, p2_concat_6229_comb} + {{8{p2_concat_6230_comb[15]}}, p2_concat_6230_comb};
  assign p2_sum__70_comb = p2_sum__83_comb + p2_sum__84_comb;
  assign p2_sum__68_comb = p2_sum__79_comb + p2_sum__80_comb;
  assign p2_sum__66_comb = p2_sum__75_comb + p2_sum__76_comb;
  assign p2_sum__64_comb = p2_sum__71_comb + p2_sum__72_comb;
  assign p2_umul_2636_NarrowedMult__comb = umul24b_24b_x_7b(p2_add_6253_comb, 7'h5b);
  assign p2_add_6271_comb = p2_add_6257_comb + p2_add_6258_comb;
  assign p2_add_6273_comb = p2_sum__67_comb + 25'h000_0001;
  assign p2_add_6275_comb = p2_add_6265_comb + p2_add_6266_comb;
  assign p2_add_6270_comb = p2_sum__70_comb + 25'h000_0001;
  assign p2_add_6272_comb = p2_sum__68_comb + 25'h000_0001;
  assign p2_add_6274_comb = p2_sum__66_comb + 25'h000_0001;
  assign p2_add_6276_comb = p2_sum__64_comb + 25'h000_0001;
  assign p2_bit_slice_6277_comb = p2_umul_2636_NarrowedMult__comb[23:7];
  assign p2_bit_slice_6279_comb = p2_add_6271_comb[23:7];
  assign p2_bit_slice_6281_comb = p2_add_6273_comb[24:8];
  assign p2_bit_slice_6283_comb = p2_add_6275_comb[23:7];
  assign p2_bit_slice_6278_comb = p2_add_6270_comb[24:8];
  assign p2_bit_slice_6280_comb = p2_add_6272_comb[24:8];
  assign p2_bit_slice_6282_comb = p2_add_6274_comb[24:8];
  assign p2_bit_slice_6284_comb = p2_add_6276_comb[24:8];
  assign p2_add_6301_comb = {{1{p2_bit_slice_6277_comb[16]}}, p2_bit_slice_6277_comb} + 18'h0_0001;
  assign p2_add_6303_comb = {{1{p2_bit_slice_6279_comb[16]}}, p2_bit_slice_6279_comb} + 18'h0_0001;
  assign p2_add_6305_comb = {{1{p2_bit_slice_6281_comb[16]}}, p2_bit_slice_6281_comb} + 18'h0_0001;
  assign p2_add_6307_comb = {{1{p2_bit_slice_6283_comb[16]}}, p2_bit_slice_6283_comb} + 18'h0_0001;
  assign p2_add_6302_comb = {{1{p2_bit_slice_6278_comb[16]}}, p2_bit_slice_6278_comb} + 18'h0_0001;
  assign p2_add_6304_comb = {{1{p2_bit_slice_6280_comb[16]}}, p2_bit_slice_6280_comb} + 18'h0_0001;
  assign p2_add_6306_comb = {{1{p2_bit_slice_6282_comb[16]}}, p2_bit_slice_6282_comb} + 18'h0_0001;
  assign p2_add_6308_comb = {{1{p2_bit_slice_6284_comb[16]}}, p2_bit_slice_6284_comb} + 18'h0_0001;
  assign p2_bit_slice_6309_comb = p2_add_6301_comb[17:8];
  assign p2_bit_slice_6310_comb = p2_add_6303_comb[17:8];
  assign p2_bit_slice_6311_comb = p2_add_6305_comb[17:8];
  assign p2_bit_slice_6312_comb = p2_add_6307_comb[17:8];
  assign p2_bit_slice_6313_comb = p2_add_6301_comb[7:1];
  assign p2_bit_slice_6314_comb = p2_add_6303_comb[7:1];
  assign p2_bit_slice_6315_comb = p2_add_6305_comb[7:1];
  assign p2_bit_slice_6316_comb = p2_add_6307_comb[7:1];

  // Registers for pipe stage 2:
  reg [17:0] p2_add_6302;
  reg [17:0] p2_add_6304;
  reg [17:0] p2_add_6306;
  reg [17:0] p2_add_6308;
  reg [9:0] p2_bit_slice_6309;
  reg [9:0] p2_bit_slice_6310;
  reg [9:0] p2_bit_slice_6311;
  reg [9:0] p2_bit_slice_6312;
  reg [6:0] p2_bit_slice_6313;
  reg [6:0] p2_bit_slice_6314;
  reg [6:0] p2_bit_slice_6315;
  reg [6:0] p2_bit_slice_6316;
  always @ (posedge clk) begin
    p2_add_6302 <= p2_add_6302_comb;
    p2_add_6304 <= p2_add_6304_comb;
    p2_add_6306 <= p2_add_6306_comb;
    p2_add_6308 <= p2_add_6308_comb;
    p2_bit_slice_6309 <= p2_bit_slice_6309_comb;
    p2_bit_slice_6310 <= p2_bit_slice_6310_comb;
    p2_bit_slice_6311 <= p2_bit_slice_6311_comb;
    p2_bit_slice_6312 <= p2_bit_slice_6312_comb;
    p2_bit_slice_6313 <= p2_bit_slice_6313_comb;
    p2_bit_slice_6314 <= p2_bit_slice_6314_comb;
    p2_bit_slice_6315 <= p2_bit_slice_6315_comb;
    p2_bit_slice_6316 <= p2_bit_slice_6316_comb;
  end

  // ===== Pipe stage 3:
  wire [9:0] p3_bit_slice_6341_comb;
  wire [9:0] p3_bit_slice_6342_comb;
  wire [9:0] p3_bit_slice_6343_comb;
  wire [9:0] p3_bit_slice_6344_comb;
  wire [10:0] p3_add_6361_comb;
  wire [10:0] p3_add_6362_comb;
  wire [10:0] p3_add_6364_comb;
  wire [10:0] p3_add_6365_comb;
  wire [10:0] p3_add_6367_comb;
  wire [10:0] p3_add_6368_comb;
  wire [10:0] p3_add_6370_comb;
  wire [10:0] p3_add_6371_comb;
  wire [17:0] p3_concat_6373_comb;
  wire [17:0] p3_concat_6376_comb;
  wire [17:0] p3_concat_6379_comb;
  wire [17:0] p3_concat_6382_comb;
  wire [17:0] p3_concat_6385_comb;
  wire [17:0] p3_concat_6388_comb;
  wire [17:0] p3_concat_6391_comb;
  wire [17:0] p3_concat_6394_comb;
  wire [9:0] p3_clipped__8_comb;
  wire [9:0] p3_clipped__9_comb;
  wire [9:0] p3_clipped__10_comb;
  wire [9:0] p3_clipped__11_comb;
  wire [9:0] p3_clipped__12_comb;
  wire [9:0] p3_clipped__13_comb;
  wire [9:0] p3_clipped__14_comb;
  wire [9:0] p3_clipped__15_comb;
  wire [9:0] p3_result_comb[0:7];
  assign p3_bit_slice_6341_comb = p2_add_6302[17:8];
  assign p3_bit_slice_6342_comb = p2_add_6304[17:8];
  assign p3_bit_slice_6343_comb = p2_add_6306[17:8];
  assign p3_bit_slice_6344_comb = p2_add_6308[17:8];
  assign p3_add_6361_comb = {{1{p2_bit_slice_6309[9]}}, p2_bit_slice_6309} + 11'h001;
  assign p3_add_6362_comb = {{1{p3_bit_slice_6341_comb[9]}}, p3_bit_slice_6341_comb} + 11'h001;
  assign p3_add_6364_comb = {{1{p2_bit_slice_6310[9]}}, p2_bit_slice_6310} + 11'h001;
  assign p3_add_6365_comb = {{1{p3_bit_slice_6342_comb[9]}}, p3_bit_slice_6342_comb} + 11'h001;
  assign p3_add_6367_comb = {{1{p2_bit_slice_6311[9]}}, p2_bit_slice_6311} + 11'h001;
  assign p3_add_6368_comb = {{1{p3_bit_slice_6343_comb[9]}}, p3_bit_slice_6343_comb} + 11'h001;
  assign p3_add_6370_comb = {{1{p2_bit_slice_6312[9]}}, p2_bit_slice_6312} + 11'h001;
  assign p3_add_6371_comb = {{1{p3_bit_slice_6344_comb[9]}}, p3_bit_slice_6344_comb} + 11'h001;
  assign p3_concat_6373_comb = {p3_add_6361_comb, p2_bit_slice_6313};
  assign p3_concat_6376_comb = {p3_add_6362_comb, p2_add_6302[7:1]};
  assign p3_concat_6379_comb = {p3_add_6364_comb, p2_bit_slice_6314};
  assign p3_concat_6382_comb = {p3_add_6365_comb, p2_add_6304[7:1]};
  assign p3_concat_6385_comb = {p3_add_6367_comb, p2_bit_slice_6315};
  assign p3_concat_6388_comb = {p3_add_6368_comb, p2_add_6306[7:1]};
  assign p3_concat_6391_comb = {p3_add_6370_comb, p2_bit_slice_6316};
  assign p3_concat_6394_comb = {p3_add_6371_comb, p2_add_6308[7:1]};
  assign p3_clipped__8_comb = $signed(p3_concat_6373_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_6373_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_6361_comb[2:0], p2_bit_slice_6313});
  assign p3_clipped__9_comb = $signed(p3_concat_6376_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_6376_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_6362_comb[2:0], p2_add_6302[7:1]});
  assign p3_clipped__10_comb = $signed(p3_concat_6379_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_6379_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_6364_comb[2:0], p2_bit_slice_6314});
  assign p3_clipped__11_comb = $signed(p3_concat_6382_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_6382_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_6365_comb[2:0], p2_add_6304[7:1]});
  assign p3_clipped__12_comb = $signed(p3_concat_6385_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_6385_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_6367_comb[2:0], p2_bit_slice_6315});
  assign p3_clipped__13_comb = $signed(p3_concat_6388_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_6388_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_6368_comb[2:0], p2_add_6306[7:1]});
  assign p3_clipped__14_comb = $signed(p3_concat_6391_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_6391_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_6370_comb[2:0], p2_bit_slice_6316});
  assign p3_clipped__15_comb = $signed(p3_concat_6394_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_6394_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_6371_comb[2:0], p2_add_6308[7:1]});
  assign p3_result_comb[0] = p3_clipped__8_comb;
  assign p3_result_comb[1] = p3_clipped__9_comb;
  assign p3_result_comb[2] = p3_clipped__10_comb;
  assign p3_result_comb[3] = p3_clipped__11_comb;
  assign p3_result_comb[4] = p3_clipped__12_comb;
  assign p3_result_comb[5] = p3_clipped__13_comb;
  assign p3_result_comb[6] = p3_clipped__14_comb;
  assign p3_result_comb[7] = p3_clipped__15_comb;

  // Registers for pipe stage 3:
  reg [9:0] p3_result[0:7];
  always @ (posedge clk) begin
    p3_result[0] <= p3_result_comb[0];
    p3_result[1] <= p3_result_comb[1];
    p3_result[2] <= p3_result_comb[2];
    p3_result[3] <= p3_result_comb[3];
    p3_result[4] <= p3_result_comb[4];
    p3_result[5] <= p3_result_comb[5];
    p3_result[6] <= p3_result_comb[6];
    p3_result[7] <= p3_result_comb[7];
  end
  assign out = {p3_result[7], p3_result[6], p3_result[5], p3_result[4], p3_result[3], p3_result[2], p3_result[1], p3_result[0]};
endmodule
