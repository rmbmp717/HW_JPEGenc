module Huffman_DCenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire is_luminance,
  output wire [32:0] out
);
  wire [7:0] literal_807[0:12];
  assign literal_807[0] = 8'h01;
  assign literal_807[1] = 8'h00;
  assign literal_807[2] = 8'h04;
  assign literal_807[3] = 8'h05;
  assign literal_807[4] = 8'h0c;
  assign literal_807[5] = 8'h0d;
  assign literal_807[6] = 8'h0e;
  assign literal_807[7] = 8'h1e;
  assign literal_807[8] = 8'h3e;
  assign literal_807[9] = 8'h7e;
  assign literal_807[10] = 8'hfe;
  assign literal_807[11] = 8'hfe;
  assign literal_807[12] = 8'h00;
  wire [7:0] literal_809[0:12];
  assign literal_809[0] = 8'h06;
  assign literal_809[1] = 8'h05;
  assign literal_809[2] = 8'h03;
  assign literal_809[3] = 8'h02;
  assign literal_809[4] = 8'h00;
  assign literal_809[5] = 8'h01;
  assign literal_809[6] = 8'h04;
  assign literal_809[7] = 8'h0e;
  assign literal_809[8] = 8'h1e;
  assign literal_809[9] = 8'h3e;
  assign literal_809[10] = 8'h7e;
  assign literal_809[11] = 8'hfe;
  assign literal_809[12] = 8'h00;
  wire [3:0] literal_810[0:12];
  assign literal_810[0] = 4'h2;
  assign literal_810[1] = 4'h2;
  assign literal_810[2] = 4'h3;
  assign literal_810[3] = 4'h3;
  assign literal_810[4] = 4'h4;
  assign literal_810[5] = 4'h4;
  assign literal_810[6] = 4'h4;
  assign literal_810[7] = 4'h5;
  assign literal_810[8] = 4'h6;
  assign literal_810[9] = 4'h7;
  assign literal_810[10] = 4'h8;
  assign literal_810[11] = 4'h9;
  assign literal_810[12] = 4'h0;
  wire [3:0] literal_811[0:12];
  assign literal_811[0] = 4'h3;
  assign literal_811[1] = 4'h3;
  assign literal_811[2] = 4'h3;
  assign literal_811[3] = 4'h3;
  assign literal_811[4] = 4'h3;
  assign literal_811[5] = 4'h3;
  assign literal_811[6] = 4'h3;
  assign literal_811[7] = 4'h4;
  assign literal_811[8] = 4'h5;
  assign literal_811[9] = 4'h6;
  assign literal_811[10] = 4'h7;
  assign literal_811[11] = 4'h8;
  assign literal_811[12] = 4'h0;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [9:0] p1_dc_comb;
  wire [7:0] p1_bin_value__1_comb;
  wire [7:0] p1_bin_value_comb;
  wire [7:0] p1_dc_abs_comb;
  wire p1_BoolList_squeezed_const_msb_bits_comb;
  wire [2:0] p1_sel_786_comb;
  wire p1_BoolList_squeezed_const_msb_bits__1_comb;
  wire [3:0] p1_concat_798_comb;
  wire [3:0] p1_Length_squeezed_const_msb_bits_comb;
  wire [7:0] p1_Code_size_comb;
  wire [3:0] p1_bit_slice_808_comb;
  wire [5:0] p1_BoolList_squeezed_squeezed_comb;
  wire [2:0] p1_Length_squeezed_squeezed_comb;
  wire [7:0] p1_flipped_comb;
  wire [8:0] p1_BoolList_comb;
  wire [7:0] p1_Length_comb;
  wire [7:0] p1_Code_list_comb;
  wire [32:0] p1_tuple_830_comb;
  assign p1_dc_comb = p0_matrix[3'h0][3'h0];
  assign p1_bin_value__1_comb = p1_dc_comb[7:0];
  assign p1_bin_value_comb = -p1_bin_value__1_comb;
  assign p1_dc_abs_comb = p1_dc_comb[9] ? p1_bin_value_comb : p1_bin_value__1_comb;
  assign p1_BoolList_squeezed_const_msb_bits_comb = 1'h0;
  assign p1_sel_786_comb = |p1_dc_abs_comb[7:3] ? 3'h4 : {p1_BoolList_squeezed_const_msb_bits_comb, |p1_dc_abs_comb[7:2] ? 2'h3 : (|p1_dc_abs_comb[7:1] ? 2'h2 : 2'h1)};
  assign p1_BoolList_squeezed_const_msb_bits__1_comb = 1'h0;
  assign p1_concat_798_comb = {p1_BoolList_squeezed_const_msb_bits__1_comb, |p1_dc_abs_comb[7:6] ? 3'h7 : (|p1_dc_abs_comb[7:5] ? 3'h6 : (|p1_dc_abs_comb[7:4] ? 3'h5 : p1_sel_786_comb))};
  assign p1_Length_squeezed_const_msb_bits_comb = 4'h0;
  assign p1_Code_size_comb = {p1_Length_squeezed_const_msb_bits_comb, p1_dc_abs_comb[7] ? 4'h8 : p1_concat_798_comb} & {8{p1_dc_abs_comb != 8'h00}};
  assign p1_bit_slice_808_comb = p1_Code_size_comb[3:0];
  assign p1_BoolList_squeezed_squeezed_comb = p0_is_luminance ? literal_809[p1_bit_slice_808_comb > 4'hc ? 4'hc : p1_bit_slice_808_comb][5:0] : literal_807[p1_bit_slice_808_comb > 4'hc ? 4'hc : p1_bit_slice_808_comb][5:0];
  assign p1_Length_squeezed_squeezed_comb = p0_is_luminance ? literal_811[p1_bit_slice_808_comb > 4'hc ? 4'hc : p1_bit_slice_808_comb][2:0] : literal_810[p1_bit_slice_808_comb > 4'hc ? 4'hc : p1_bit_slice_808_comb][2:0];
  assign p1_flipped_comb = ~p1_bin_value_comb;
  assign p1_BoolList_comb = {3'h0, p1_BoolList_squeezed_squeezed_comb};
  assign p1_Length_comb = {5'h00, p1_Length_squeezed_squeezed_comb};
  assign p1_Code_list_comb = $signed(p1_dc_comb) <= $signed(10'h000) ? p1_flipped_comb : p1_bin_value__1_comb;
  assign p1_tuple_830_comb = {p1_BoolList_comb, p1_Length_comb, p1_Code_list_comb, p1_Code_size_comb};

  // Registers for pipe stage 1:
  reg [32:0] p1_tuple_830;
  always @ (posedge clk) begin
    p1_tuple_830 <= p1_tuple_830_comb;
  end
  assign out = p1_tuple_830;
endmodule
