module dct_1d_s12(
  input wire clk,
  input wire [95:0] x,
  output wire [95:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [20:0] smul21b_12b_x_9b (input reg [11:0] lhs, input reg [8:0] rhs);
    reg signed [11:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [20:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul21b_12b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [19:0] smul20b_12b_x_8b (input reg [11:0] lhs, input reg [7:0] rhs);
    reg signed [11:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [19:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul20b_12b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [17:0] smul18b_12b_x_6b (input reg [11:0] lhs, input reg [5:0] rhs);
    reg signed [11:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [17:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul18b_12b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [18:0] smul19b_12b_x_7b (input reg [11:0] lhs, input reg [6:0] rhs);
    reg signed [11:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [18:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul19b_12b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_7b (input reg [31:0] lhs, input reg [6:0] rhs);
    begin
      umul32b_32b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [11:0] x_unflattened[0:7];
  assign x_unflattened[0] = x[11:0];
  assign x_unflattened[1] = x[23:12];
  assign x_unflattened[2] = x[35:24];
  assign x_unflattened[3] = x[47:36];
  assign x_unflattened[4] = x[59:48];
  assign x_unflattened[5] = x[71:60];
  assign x_unflattened[6] = x[83:72];
  assign x_unflattened[7] = x[95:84];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [11:0] p0_x[0:7];
  always @ (posedge clk) begin
    p0_x[0] <= x_unflattened[0];
    p0_x[1] <= x_unflattened[1];
    p0_x[2] <= x_unflattened[2];
    p0_x[3] <= x_unflattened[3];
    p0_x[4] <= x_unflattened[4];
    p0_x[5] <= x_unflattened[5];
    p0_x[6] <= x_unflattened[6];
    p0_x[7] <= x_unflattened[7];
  end

  // ===== Pipe stage 1:
  wire [11:0] p1_array_index_5005_comb;
  wire [11:0] p1_array_index_4993_comb;
  wire [11:0] p1_array_index_4999_comb;
  wire [11:0] p1_array_index_5009_comb;
  wire [11:0] p1_array_index_4995_comb;
  wire [11:0] p1_array_index_4989_comb;
  wire [11:0] p1_array_index_4991_comb;
  wire [11:0] p1_array_index_4997_comb;
  wire [20:0] p1_smul_5069_comb;
  wire [20:0] p1_smul_5070_comb;
  wire [20:0] p1_smul_5077_comb;
  wire [20:0] p1_smul_5078_comb;
  wire [20:0] p1_smul_5094_comb;
  wire [19:0] p1_smul_2602_NarrowedMult__comb;
  wire [19:0] p1_smul_2604_NarrowedMult__comb;
  wire [20:0] p1_smul_5097_comb;
  wire [20:0] p1_smul_5101_comb;
  wire [20:0] p1_smul_5102_comb;
  wire [20:0] p1_smul_5103_comb;
  wire [20:0] p1_smul_5104_comb;
  wire [20:0] p1_smul_5105_comb;
  wire [20:0] p1_smul_5106_comb;
  wire [20:0] p1_smul_5107_comb;
  wire [20:0] p1_smul_5108_comb;
  wire [19:0] p1_smul_2628_NarrowedMult__comb;
  wire [20:0] p1_smul_5110_comb;
  wire [20:0] p1_smul_5117_comb;
  wire [19:0] p1_smul_2642_NarrowedMult__comb;
  wire [20:0] p1_smul_5134_comb;
  wire [20:0] p1_smul_5135_comb;
  wire [20:0] p1_smul_5136_comb;
  wire [20:0] p1_smul_5137_comb;
  wire [17:0] p1_smul_2570_NarrowedMult__comb;
  wire [17:0] p1_smul_2572_NarrowedMult__comb;
  wire [18:0] p1_smul_2582_NarrowedMult__comb;
  wire [18:0] p1_smul_2584_NarrowedMult__comb;
  wire [18:0] p1_smul_2590_NarrowedMult__comb;
  wire [18:0] p1_smul_2592_NarrowedMult__comb;
  wire [17:0] p1_smul_2598_NarrowedMult__comb;
  wire [17:0] p1_smul_2608_NarrowedMult__comb;
  wire [17:0] p1_smul_2632_NarrowedMult__comb;
  wire [17:0] p1_smul_2638_NarrowedMult__comb;
  wire [18:0] p1_smul_2644_NarrowedMult__comb;
  wire [18:0] p1_smul_2648_NarrowedMult__comb;
  wire [18:0] p1_smul_2654_NarrowedMult__comb;
  wire [18:0] p1_smul_2658_NarrowedMult__comb;
  wire [17:0] p1_smul_2660_NarrowedMult__comb;
  wire [17:0] p1_smul_2674_NarrowedMult__comb;
  wire [19:0] p1_smul_2568_NarrowedMult__comb;
  wire [19:0] p1_smul_2574_NarrowedMult__comb;
  wire [18:0] p1_smul_2580_NarrowedMult__comb;
  wire [18:0] p1_smul_2586_NarrowedMult__comb;
  wire [18:0] p1_smul_2588_NarrowedMult__comb;
  wire [18:0] p1_smul_2594_NarrowedMult__comb;
  wire [20:0] p1_smul_5091_comb;
  wire [20:0] p1_smul_5100_comb;
  wire [20:0] p1_smul_5113_comb;
  wire [20:0] p1_smul_5114_comb;
  wire [18:0] p1_smul_2646_NarrowedMult__comb;
  wire [18:0] p1_smul_2650_NarrowedMult__comb;
  wire [18:0] p1_smul_2652_NarrowedMult__comb;
  wire [18:0] p1_smul_2656_NarrowedMult__comb;
  wire [19:0] p1_smul_2662_NarrowedMult__comb;
  wire [19:0] p1_smul_2672_NarrowedMult__comb;
  wire [12:0] p1_add_5245_comb;
  wire [12:0] p1_add_5246_comb;
  wire [12:0] p1_add_5247_comb;
  wire [12:0] p1_add_5248_comb;
  wire [13:0] p1_add_5249_comb;
  wire [13:0] p1_add_5250_comb;
  wire [13:0] p1_add_5255_comb;
  wire [13:0] p1_add_5256_comb;
  wire [13:0] p1_add_5267_comb;
  wire [13:0] p1_add_5268_comb;
  wire [13:0] p1_add_5269_comb;
  wire [13:0] p1_add_5270_comb;
  wire [13:0] p1_add_5273_comb;
  wire [13:0] p1_add_5274_comb;
  wire [13:0] p1_add_5275_comb;
  wire [13:0] p1_add_5276_comb;
  wire [13:0] p1_add_5277_comb;
  wire [13:0] p1_add_5278_comb;
  wire [13:0] p1_add_5279_comb;
  wire [13:0] p1_add_5280_comb;
  wire [13:0] p1_add_5281_comb;
  wire [13:0] p1_add_5282_comb;
  wire [13:0] p1_add_5287_comb;
  wire [13:0] p1_add_5288_comb;
  wire [13:0] p1_add_5299_comb;
  wire [13:0] p1_add_5300_comb;
  wire [13:0] p1_add_5301_comb;
  wire [13:0] p1_add_5302_comb;
  wire [31:0] p1_sum__8_comb;
  wire [31:0] p1_sum__9_comb;
  wire [31:0] p1_sum__10_comb;
  wire [31:0] p1_sum__11_comb;
  wire [11:0] p1_add_5155_comb;
  wire [11:0] p1_add_5156_comb;
  wire [12:0] p1_add_5165_comb;
  wire [12:0] p1_add_5166_comb;
  wire [12:0] p1_add_5171_comb;
  wire [12:0] p1_add_5172_comb;
  wire [11:0] p1_add_5177_comb;
  wire [11:0] p1_add_5186_comb;
  wire [11:0] p1_add_5209_comb;
  wire [11:0] p1_add_5214_comb;
  wire [12:0] p1_add_5219_comb;
  wire [12:0] p1_add_5222_comb;
  wire [12:0] p1_add_5227_comb;
  wire [12:0] p1_add_5230_comb;
  wire [11:0] p1_add_5231_comb;
  wire [11:0] p1_add_5244_comb;
  wire [13:0] p1_add_5251_comb;
  wire [13:0] p1_add_5254_comb;
  wire [13:0] p1_add_5257_comb;
  wire [13:0] p1_add_5260_comb;
  wire [13:0] p1_add_5261_comb;
  wire [13:0] p1_add_5264_comb;
  wire [13:0] p1_add_5265_comb;
  wire [13:0] p1_add_5272_comb;
  wire [13:0] p1_add_5284_comb;
  wire [13:0] p1_add_5285_comb;
  wire [13:0] p1_add_5290_comb;
  wire [13:0] p1_add_5292_comb;
  wire [13:0] p1_add_5293_comb;
  wire [13:0] p1_add_5295_comb;
  wire [13:0] p1_add_5298_comb;
  wire [13:0] p1_add_5303_comb;
  wire [31:0] p1_sum__12_comb;
  wire [31:0] p1_sum__13_comb;
  wire [10:0] p1_bit_slice_5252_comb;
  wire [10:0] p1_bit_slice_5253_comb;
  wire [11:0] p1_bit_slice_5258_comb;
  wire [11:0] p1_bit_slice_5259_comb;
  wire [11:0] p1_bit_slice_5262_comb;
  wire [11:0] p1_bit_slice_5263_comb;
  wire [10:0] p1_bit_slice_5266_comb;
  wire [10:0] p1_bit_slice_5271_comb;
  wire [10:0] p1_bit_slice_5283_comb;
  wire [10:0] p1_bit_slice_5286_comb;
  wire [11:0] p1_bit_slice_5289_comb;
  wire [11:0] p1_bit_slice_5291_comb;
  wire [11:0] p1_bit_slice_5294_comb;
  wire [11:0] p1_bit_slice_5296_comb;
  wire [10:0] p1_bit_slice_5297_comb;
  wire [10:0] p1_bit_slice_5304_comb;
  wire [12:0] p1_bit_slice_5311_comb;
  wire [12:0] p1_bit_slice_5312_comb;
  wire [12:0] p1_bit_slice_5315_comb;
  wire [12:0] p1_bit_slice_5316_comb;
  wire [12:0] p1_bit_slice_5317_comb;
  wire [12:0] p1_bit_slice_5318_comb;
  wire [12:0] p1_bit_slice_5319_comb;
  wire [12:0] p1_bit_slice_5324_comb;
  wire [12:0] p1_bit_slice_5335_comb;
  wire [12:0] p1_bit_slice_5336_comb;
  wire [12:0] p1_bit_slice_5339_comb;
  wire [12:0] p1_bit_slice_5340_comb;
  wire [12:0] p1_bit_slice_5341_comb;
  wire [12:0] p1_bit_slice_5342_comb;
  wire [12:0] p1_bit_slice_5343_comb;
  wire [12:0] p1_bit_slice_5348_comb;
  wire [12:0] p1_add_5351_comb;
  wire [12:0] p1_add_5352_comb;
  wire [12:0] p1_add_5353_comb;
  wire [12:0] p1_add_5354_comb;
  wire [12:0] p1_add_5355_comb;
  wire [12:0] p1_add_5356_comb;
  wire [12:0] p1_add_5357_comb;
  wire [12:0] p1_add_5358_comb;
  wire [12:0] p1_add_5359_comb;
  wire [12:0] p1_add_5360_comb;
  wire [12:0] p1_add_5361_comb;
  wire [12:0] p1_add_5362_comb;
  wire [31:0] p1_sum__14_comb;
  assign p1_array_index_5005_comb = p0_x[3'h0];
  assign p1_array_index_4993_comb = p0_x[3'h1];
  assign p1_array_index_4999_comb = p0_x[3'h6];
  assign p1_array_index_5009_comb = p0_x[3'h7];
  assign p1_array_index_4995_comb = p0_x[3'h2];
  assign p1_array_index_4989_comb = p0_x[3'h3];
  assign p1_array_index_4991_comb = p0_x[3'h4];
  assign p1_array_index_4997_comb = p0_x[3'h5];
  assign p1_smul_5069_comb = smul21b_12b_x_9b(p1_array_index_5005_comb, 9'h0fb);
  assign p1_smul_5070_comb = smul21b_12b_x_9b(p1_array_index_4993_comb, 9'h0d5);
  assign p1_smul_5077_comb = smul21b_12b_x_9b(p1_array_index_4999_comb, 9'h12b);
  assign p1_smul_5078_comb = smul21b_12b_x_9b(p1_array_index_5009_comb, 9'h105);
  assign p1_smul_5094_comb = smul21b_12b_x_9b(p1_array_index_4995_comb, 9'h105);
  assign p1_smul_2602_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_4989_comb, 8'hb9);
  assign p1_smul_2604_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_4991_comb, 8'h47);
  assign p1_smul_5097_comb = smul21b_12b_x_9b(p1_array_index_4997_comb, 9'h0fb);
  assign p1_smul_5101_comb = smul21b_12b_x_9b(p1_array_index_5005_comb, 9'h0b5);
  assign p1_smul_5102_comb = smul21b_12b_x_9b(p1_array_index_4993_comb, 9'h14b);
  assign p1_smul_5103_comb = smul21b_12b_x_9b(p1_array_index_4995_comb, 9'h14b);
  assign p1_smul_5104_comb = smul21b_12b_x_9b(p1_array_index_4989_comb, 9'h0b5);
  assign p1_smul_5105_comb = smul21b_12b_x_9b(p1_array_index_4991_comb, 9'h0b5);
  assign p1_smul_5106_comb = smul21b_12b_x_9b(p1_array_index_4997_comb, 9'h14b);
  assign p1_smul_5107_comb = smul21b_12b_x_9b(p1_array_index_4999_comb, 9'h14b);
  assign p1_smul_5108_comb = smul21b_12b_x_9b(p1_array_index_5009_comb, 9'h0b5);
  assign p1_smul_2628_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_5005_comb, 8'h47);
  assign p1_smul_5110_comb = smul21b_12b_x_9b(p1_array_index_4993_comb, 9'h105);
  assign p1_smul_5117_comb = smul21b_12b_x_9b(p1_array_index_4999_comb, 9'h105);
  assign p1_smul_2642_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_5009_comb, 8'h47);
  assign p1_smul_5134_comb = smul21b_12b_x_9b(p1_array_index_4995_comb, 9'h0d5);
  assign p1_smul_5135_comb = smul21b_12b_x_9b(p1_array_index_4989_comb, 9'h105);
  assign p1_smul_5136_comb = smul21b_12b_x_9b(p1_array_index_4991_comb, 9'h105);
  assign p1_smul_5137_comb = smul21b_12b_x_9b(p1_array_index_4997_comb, 9'h0d5);
  assign p1_smul_2570_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_4989_comb, 6'h19);
  assign p1_smul_2572_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_4991_comb, 6'h27);
  assign p1_smul_2582_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4993_comb, 7'h31);
  assign p1_smul_2584_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4995_comb, 7'h4f);
  assign p1_smul_2590_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4997_comb, 7'h4f);
  assign p1_smul_2592_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4999_comb, 7'h31);
  assign p1_smul_2598_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_4993_comb, 6'h27);
  assign p1_smul_2608_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_4999_comb, 6'h19);
  assign p1_smul_2632_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_4995_comb, 6'h27);
  assign p1_smul_2638_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_4997_comb, 6'h27);
  assign p1_smul_2644_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_5005_comb, 7'h31);
  assign p1_smul_2648_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4995_comb, 7'h31);
  assign p1_smul_2654_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4997_comb, 7'h31);
  assign p1_smul_2658_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_5009_comb, 7'h31);
  assign p1_smul_2660_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_5005_comb, 6'h19);
  assign p1_smul_2674_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_5009_comb, 6'h19);
  assign p1_smul_2568_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_4995_comb, 8'h47);
  assign p1_smul_2574_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_4997_comb, 8'hb9);
  assign p1_smul_2580_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_5005_comb, 7'h3b);
  assign p1_smul_2586_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4989_comb, 7'h45);
  assign p1_smul_2588_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4991_comb, 7'h45);
  assign p1_smul_2594_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_5009_comb, 7'h3b);
  assign p1_smul_5091_comb = smul21b_12b_x_9b(p1_array_index_5005_comb, 9'h0d5);
  assign p1_smul_5100_comb = smul21b_12b_x_9b(p1_array_index_5009_comb, 9'h12b);
  assign p1_smul_5113_comb = smul21b_12b_x_9b(p1_array_index_4989_comb, 9'h0d5);
  assign p1_smul_5114_comb = smul21b_12b_x_9b(p1_array_index_4991_comb, 9'h0d5);
  assign p1_smul_2646_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4993_comb, 7'h45);
  assign p1_smul_2650_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4989_comb, 7'h3b);
  assign p1_smul_2652_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4991_comb, 7'h3b);
  assign p1_smul_2656_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_4999_comb, 7'h45);
  assign p1_smul_2662_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_4993_comb, 8'hb9);
  assign p1_smul_2672_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_4999_comb, 8'hb9);
  assign p1_add_5245_comb = {{1{p1_array_index_5005_comb[11]}}, p1_array_index_5005_comb} + {{1{p1_array_index_4993_comb[11]}}, p1_array_index_4993_comb};
  assign p1_add_5246_comb = {{1{p1_array_index_4995_comb[11]}}, p1_array_index_4995_comb} + {{1{p1_array_index_4989_comb[11]}}, p1_array_index_4989_comb};
  assign p1_add_5247_comb = {{1{p1_array_index_4991_comb[11]}}, p1_array_index_4991_comb} + {{1{p1_array_index_4997_comb[11]}}, p1_array_index_4997_comb};
  assign p1_add_5248_comb = {{1{p1_array_index_4999_comb[11]}}, p1_array_index_4999_comb} + {{1{p1_array_index_5009_comb[11]}}, p1_array_index_5009_comb};
  assign p1_add_5249_comb = p1_smul_5069_comb[20:7] + 14'h0001;
  assign p1_add_5250_comb = p1_smul_5070_comb[20:7] + 14'h0001;
  assign p1_add_5255_comb = p1_smul_5077_comb[20:7] + 14'h0001;
  assign p1_add_5256_comb = p1_smul_5078_comb[20:7] + 14'h0001;
  assign p1_add_5267_comb = p1_smul_5094_comb[20:7] + 14'h0001;
  assign p1_add_5268_comb = p1_smul_2602_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_5269_comb = p1_smul_2604_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_5270_comb = p1_smul_5097_comb[20:7] + 14'h0001;
  assign p1_add_5273_comb = p1_smul_5101_comb[20:7] + 14'h0001;
  assign p1_add_5274_comb = p1_smul_5102_comb[20:7] + 14'h0001;
  assign p1_add_5275_comb = p1_smul_5103_comb[20:7] + 14'h0001;
  assign p1_add_5276_comb = p1_smul_5104_comb[20:7] + 14'h0001;
  assign p1_add_5277_comb = p1_smul_5105_comb[20:7] + 14'h0001;
  assign p1_add_5278_comb = p1_smul_5106_comb[20:7] + 14'h0001;
  assign p1_add_5279_comb = p1_smul_5107_comb[20:7] + 14'h0001;
  assign p1_add_5280_comb = p1_smul_5108_comb[20:7] + 14'h0001;
  assign p1_add_5281_comb = p1_smul_2628_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_5282_comb = p1_smul_5110_comb[20:7] + 14'h0001;
  assign p1_add_5287_comb = p1_smul_5117_comb[20:7] + 14'h0001;
  assign p1_add_5288_comb = p1_smul_2642_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_5299_comb = p1_smul_5134_comb[20:7] + 14'h0001;
  assign p1_add_5300_comb = p1_smul_5135_comb[20:7] + 14'h0001;
  assign p1_add_5301_comb = p1_smul_5136_comb[20:7] + 14'h0001;
  assign p1_add_5302_comb = p1_smul_5137_comb[20:7] + 14'h0001;
  assign p1_sum__8_comb = {{19{p1_add_5245_comb[12]}}, p1_add_5245_comb};
  assign p1_sum__9_comb = {{19{p1_add_5246_comb[12]}}, p1_add_5246_comb};
  assign p1_sum__10_comb = {{19{p1_add_5247_comb[12]}}, p1_add_5247_comb};
  assign p1_sum__11_comb = {{19{p1_add_5248_comb[12]}}, p1_add_5248_comb};
  assign p1_add_5155_comb = p1_smul_2570_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_5156_comb = p1_smul_2572_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_5165_comb = p1_smul_2582_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_5166_comb = p1_smul_2584_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_5171_comb = p1_smul_2590_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_5172_comb = p1_smul_2592_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_5177_comb = p1_smul_2598_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_5186_comb = p1_smul_2608_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_5209_comb = p1_smul_2632_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_5214_comb = p1_smul_2638_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_5219_comb = p1_smul_2644_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_5222_comb = p1_smul_2648_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_5227_comb = p1_smul_2654_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_5230_comb = p1_smul_2658_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_5231_comb = p1_smul_2660_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_5244_comb = p1_smul_2674_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_5251_comb = p1_smul_2568_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_5254_comb = p1_smul_2574_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_5257_comb = p1_smul_2580_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_5260_comb = p1_smul_2586_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_5261_comb = p1_smul_2588_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_5264_comb = p1_smul_2594_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_5265_comb = p1_smul_5091_comb[20:7] + 14'h0001;
  assign p1_add_5272_comb = p1_smul_5100_comb[20:7] + 14'h0001;
  assign p1_add_5284_comb = p1_smul_5113_comb[20:7] + 14'h0001;
  assign p1_add_5285_comb = p1_smul_5114_comb[20:7] + 14'h0001;
  assign p1_add_5290_comb = p1_smul_2646_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_5292_comb = p1_smul_2650_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_5293_comb = p1_smul_2652_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_5295_comb = p1_smul_2656_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_5298_comb = p1_smul_2662_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_5303_comb = p1_smul_2672_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_sum__12_comb = p1_sum__8_comb + p1_sum__9_comb;
  assign p1_sum__13_comb = p1_sum__10_comb + p1_sum__11_comb;
  assign p1_bit_slice_5252_comb = p1_add_5155_comb[11:1];
  assign p1_bit_slice_5253_comb = p1_add_5156_comb[11:1];
  assign p1_bit_slice_5258_comb = p1_add_5165_comb[12:1];
  assign p1_bit_slice_5259_comb = p1_add_5166_comb[12:1];
  assign p1_bit_slice_5262_comb = p1_add_5171_comb[12:1];
  assign p1_bit_slice_5263_comb = p1_add_5172_comb[12:1];
  assign p1_bit_slice_5266_comb = p1_add_5177_comb[11:1];
  assign p1_bit_slice_5271_comb = p1_add_5186_comb[11:1];
  assign p1_bit_slice_5283_comb = p1_add_5209_comb[11:1];
  assign p1_bit_slice_5286_comb = p1_add_5214_comb[11:1];
  assign p1_bit_slice_5289_comb = p1_add_5219_comb[12:1];
  assign p1_bit_slice_5291_comb = p1_add_5222_comb[12:1];
  assign p1_bit_slice_5294_comb = p1_add_5227_comb[12:1];
  assign p1_bit_slice_5296_comb = p1_add_5230_comb[12:1];
  assign p1_bit_slice_5297_comb = p1_add_5231_comb[11:1];
  assign p1_bit_slice_5304_comb = p1_add_5244_comb[11:1];
  assign p1_bit_slice_5311_comb = p1_add_5251_comb[13:1];
  assign p1_bit_slice_5312_comb = p1_add_5254_comb[13:1];
  assign p1_bit_slice_5315_comb = p1_add_5257_comb[13:1];
  assign p1_bit_slice_5316_comb = p1_add_5260_comb[13:1];
  assign p1_bit_slice_5317_comb = p1_add_5261_comb[13:1];
  assign p1_bit_slice_5318_comb = p1_add_5264_comb[13:1];
  assign p1_bit_slice_5319_comb = p1_add_5265_comb[13:1];
  assign p1_bit_slice_5324_comb = p1_add_5272_comb[13:1];
  assign p1_bit_slice_5335_comb = p1_add_5284_comb[13:1];
  assign p1_bit_slice_5336_comb = p1_add_5285_comb[13:1];
  assign p1_bit_slice_5339_comb = p1_add_5290_comb[13:1];
  assign p1_bit_slice_5340_comb = p1_add_5292_comb[13:1];
  assign p1_bit_slice_5341_comb = p1_add_5293_comb[13:1];
  assign p1_bit_slice_5342_comb = p1_add_5295_comb[13:1];
  assign p1_bit_slice_5343_comb = p1_add_5298_comb[13:1];
  assign p1_bit_slice_5348_comb = p1_add_5303_comb[13:1];
  assign p1_add_5351_comb = p1_add_5249_comb[13:1] + p1_add_5250_comb[13:1];
  assign p1_add_5352_comb = p1_add_5255_comb[13:1] + p1_add_5256_comb[13:1];
  assign p1_add_5353_comb = p1_add_5267_comb[13:1] + p1_add_5268_comb[13:1];
  assign p1_add_5354_comb = p1_add_5269_comb[13:1] + p1_add_5270_comb[13:1];
  assign p1_add_5355_comb = p1_add_5273_comb[13:1] + p1_add_5274_comb[13:1];
  assign p1_add_5356_comb = p1_add_5275_comb[13:1] + p1_add_5276_comb[13:1];
  assign p1_add_5357_comb = p1_add_5277_comb[13:1] + p1_add_5278_comb[13:1];
  assign p1_add_5358_comb = p1_add_5279_comb[13:1] + p1_add_5280_comb[13:1];
  assign p1_add_5359_comb = p1_add_5281_comb[13:1] + p1_add_5282_comb[13:1];
  assign p1_add_5360_comb = p1_add_5287_comb[13:1] + p1_add_5288_comb[13:1];
  assign p1_add_5361_comb = p1_add_5299_comb[13:1] + p1_add_5300_comb[13:1];
  assign p1_add_5362_comb = p1_add_5301_comb[13:1] + p1_add_5302_comb[13:1];
  assign p1_sum__14_comb = p1_sum__12_comb + p1_sum__13_comb;

  // Registers for pipe stage 1:
  reg [10:0] p1_bit_slice_5252;
  reg [10:0] p1_bit_slice_5253;
  reg [11:0] p1_bit_slice_5258;
  reg [11:0] p1_bit_slice_5259;
  reg [11:0] p1_bit_slice_5262;
  reg [11:0] p1_bit_slice_5263;
  reg [10:0] p1_bit_slice_5266;
  reg [10:0] p1_bit_slice_5271;
  reg [10:0] p1_bit_slice_5283;
  reg [10:0] p1_bit_slice_5286;
  reg [11:0] p1_bit_slice_5289;
  reg [11:0] p1_bit_slice_5291;
  reg [11:0] p1_bit_slice_5294;
  reg [11:0] p1_bit_slice_5296;
  reg [10:0] p1_bit_slice_5297;
  reg [10:0] p1_bit_slice_5304;
  reg [12:0] p1_bit_slice_5311;
  reg [12:0] p1_bit_slice_5312;
  reg [12:0] p1_bit_slice_5315;
  reg [12:0] p1_bit_slice_5316;
  reg [12:0] p1_bit_slice_5317;
  reg [12:0] p1_bit_slice_5318;
  reg [12:0] p1_bit_slice_5319;
  reg [12:0] p1_bit_slice_5324;
  reg [12:0] p1_bit_slice_5335;
  reg [12:0] p1_bit_slice_5336;
  reg [12:0] p1_bit_slice_5339;
  reg [12:0] p1_bit_slice_5340;
  reg [12:0] p1_bit_slice_5341;
  reg [12:0] p1_bit_slice_5342;
  reg [12:0] p1_bit_slice_5343;
  reg [12:0] p1_bit_slice_5348;
  reg [12:0] p1_add_5351;
  reg [12:0] p1_add_5352;
  reg [12:0] p1_add_5353;
  reg [12:0] p1_add_5354;
  reg [12:0] p1_add_5355;
  reg [12:0] p1_add_5356;
  reg [12:0] p1_add_5357;
  reg [12:0] p1_add_5358;
  reg [12:0] p1_add_5359;
  reg [12:0] p1_add_5360;
  reg [12:0] p1_add_5361;
  reg [12:0] p1_add_5362;
  reg [31:0] p1_sum__14;
  always @ (posedge clk) begin
    p1_bit_slice_5252 <= p1_bit_slice_5252_comb;
    p1_bit_slice_5253 <= p1_bit_slice_5253_comb;
    p1_bit_slice_5258 <= p1_bit_slice_5258_comb;
    p1_bit_slice_5259 <= p1_bit_slice_5259_comb;
    p1_bit_slice_5262 <= p1_bit_slice_5262_comb;
    p1_bit_slice_5263 <= p1_bit_slice_5263_comb;
    p1_bit_slice_5266 <= p1_bit_slice_5266_comb;
    p1_bit_slice_5271 <= p1_bit_slice_5271_comb;
    p1_bit_slice_5283 <= p1_bit_slice_5283_comb;
    p1_bit_slice_5286 <= p1_bit_slice_5286_comb;
    p1_bit_slice_5289 <= p1_bit_slice_5289_comb;
    p1_bit_slice_5291 <= p1_bit_slice_5291_comb;
    p1_bit_slice_5294 <= p1_bit_slice_5294_comb;
    p1_bit_slice_5296 <= p1_bit_slice_5296_comb;
    p1_bit_slice_5297 <= p1_bit_slice_5297_comb;
    p1_bit_slice_5304 <= p1_bit_slice_5304_comb;
    p1_bit_slice_5311 <= p1_bit_slice_5311_comb;
    p1_bit_slice_5312 <= p1_bit_slice_5312_comb;
    p1_bit_slice_5315 <= p1_bit_slice_5315_comb;
    p1_bit_slice_5316 <= p1_bit_slice_5316_comb;
    p1_bit_slice_5317 <= p1_bit_slice_5317_comb;
    p1_bit_slice_5318 <= p1_bit_slice_5318_comb;
    p1_bit_slice_5319 <= p1_bit_slice_5319_comb;
    p1_bit_slice_5324 <= p1_bit_slice_5324_comb;
    p1_bit_slice_5335 <= p1_bit_slice_5335_comb;
    p1_bit_slice_5336 <= p1_bit_slice_5336_comb;
    p1_bit_slice_5339 <= p1_bit_slice_5339_comb;
    p1_bit_slice_5340 <= p1_bit_slice_5340_comb;
    p1_bit_slice_5341 <= p1_bit_slice_5341_comb;
    p1_bit_slice_5342 <= p1_bit_slice_5342_comb;
    p1_bit_slice_5343 <= p1_bit_slice_5343_comb;
    p1_bit_slice_5348 <= p1_bit_slice_5348_comb;
    p1_add_5351 <= p1_add_5351_comb;
    p1_add_5352 <= p1_add_5352_comb;
    p1_add_5353 <= p1_add_5353_comb;
    p1_add_5354 <= p1_add_5354_comb;
    p1_add_5355 <= p1_add_5355_comb;
    p1_add_5356 <= p1_add_5356_comb;
    p1_add_5357 <= p1_add_5357_comb;
    p1_add_5358 <= p1_add_5358_comb;
    p1_add_5359 <= p1_add_5359_comb;
    p1_add_5360 <= p1_add_5360_comb;
    p1_add_5361 <= p1_add_5361_comb;
    p1_add_5362 <= p1_add_5362_comb;
    p1_sum__14 <= p1_sum__14_comb;
  end

  // ===== Pipe stage 2:
  wire [24:0] p2_sum__97_comb;
  wire [24:0] p2_sum__98_comb;
  wire [24:0] p2_sum__99_comb;
  wire [24:0] p2_sum__100_comb;
  wire [31:0] p2_umul_5515_comb;
  wire [12:0] p2_add_5470_comb;
  wire [12:0] p2_add_5471_comb;
  wire [12:0] p2_add_5472_comb;
  wire [12:0] p2_add_5473_comb;
  wire [12:0] p2_add_5474_comb;
  wire [12:0] p2_add_5475_comb;
  wire [12:0] p2_add_5476_comb;
  wire [12:0] p2_add_5477_comb;
  wire [12:0] p2_add_5478_comb;
  wire [12:0] p2_add_5479_comb;
  wire [12:0] p2_add_5480_comb;
  wire [12:0] p2_add_5481_comb;
  wire [12:0] p2_add_5482_comb;
  wire [12:0] p2_add_5483_comb;
  wire [12:0] p2_add_5484_comb;
  wire [12:0] p2_add_5485_comb;
  wire [24:0] p2_sum__77_comb;
  wire [24:0] p2_sum__78_comb;
  wire [24:0] p2_sum__109_comb;
  wire [24:0] p2_sum__110_comb;
  wire [24:0] p2_sum__111_comb;
  wire [24:0] p2_sum__112_comb;
  wire [24:0] p2_sum__105_comb;
  wire [24:0] p2_sum__106_comb;
  wire [24:0] p2_sum__107_comb;
  wire [24:0] p2_sum__108_comb;
  wire [24:0] p2_sum__101_comb;
  wire [24:0] p2_sum__102_comb;
  wire [24:0] p2_sum__103_comb;
  wire [24:0] p2_sum__104_comb;
  wire [24:0] p2_sum__93_comb;
  wire [24:0] p2_sum__94_comb;
  wire [24:0] p2_sum__95_comb;
  wire [24:0] p2_sum__96_comb;
  wire [24:0] p2_sum__89_comb;
  wire [24:0] p2_sum__90_comb;
  wire [24:0] p2_sum__91_comb;
  wire [24:0] p2_sum__92_comb;
  wire [24:0] p2_sum__85_comb;
  wire [24:0] p2_sum__86_comb;
  wire [24:0] p2_sum__87_comb;
  wire [24:0] p2_sum__88_comb;
  wire [24:0] p2_sum__67_comb;
  wire [24:0] p2_add_5546_comb;
  wire [24:0] p2_sum__83_comb;
  wire [24:0] p2_sum__84_comb;
  wire [24:0] p2_sum__81_comb;
  wire [24:0] p2_sum__82_comb;
  wire [24:0] p2_sum__79_comb;
  wire [24:0] p2_sum__80_comb;
  wire [24:0] p2_sum__75_comb;
  wire [24:0] p2_sum__76_comb;
  wire [24:0] p2_sum__73_comb;
  wire [24:0] p2_sum__74_comb;
  wire [24:0] p2_sum__71_comb;
  wire [24:0] p2_sum__72_comb;
  wire [24:0] p2_add_5550_comb;
  wire [24:0] p2_sum__70_comb;
  wire [24:0] p2_sum__69_comb;
  wire [24:0] p2_sum__68_comb;
  wire [24:0] p2_sum__66_comb;
  wire [24:0] p2_sum__65_comb;
  wire [24:0] p2_sum__64_comb;
  wire [24:0] p2_add_5547_comb;
  wire [24:0] p2_add_5548_comb;
  wire [24:0] p2_add_5549_comb;
  wire [24:0] p2_add_5551_comb;
  wire [24:0] p2_add_5552_comb;
  wire [24:0] p2_add_5553_comb;
  wire p2_sgt_5563_comb;
  wire [11:0] p2_bit_slice_5564_comb;
  wire p2_slt_5565_comb;
  wire [11:0] p2_sel_5566_comb;
  wire p2_slt_5567_comb;
  assign p2_sum__97_comb = {{12{p1_add_5355[12]}}, p1_add_5355};
  assign p2_sum__98_comb = {{12{p1_add_5356[12]}}, p1_add_5356};
  assign p2_sum__99_comb = {{12{p1_add_5357[12]}}, p1_add_5357};
  assign p2_sum__100_comb = {{12{p1_add_5358[12]}}, p1_add_5358};
  assign p2_umul_5515_comb = umul32b_32b_x_7b(p1_sum__14, 7'h5b);
  assign p2_add_5470_comb = p1_bit_slice_5311 + {{2{p1_bit_slice_5252[10]}}, p1_bit_slice_5252};
  assign p2_add_5471_comb = {{2{p1_bit_slice_5253[10]}}, p1_bit_slice_5253} + p1_bit_slice_5312;
  assign p2_add_5472_comb = p1_bit_slice_5315 + {{1{p1_bit_slice_5258[11]}}, p1_bit_slice_5258};
  assign p2_add_5473_comb = {{1{p1_bit_slice_5259[11]}}, p1_bit_slice_5259} + p1_bit_slice_5316;
  assign p2_add_5474_comb = p1_bit_slice_5317 + {{1{p1_bit_slice_5262[11]}}, p1_bit_slice_5262};
  assign p2_add_5475_comb = {{1{p1_bit_slice_5263[11]}}, p1_bit_slice_5263} + p1_bit_slice_5318;
  assign p2_add_5476_comb = p1_bit_slice_5319 + {{2{p1_bit_slice_5266[10]}}, p1_bit_slice_5266};
  assign p2_add_5477_comb = {{2{p1_bit_slice_5271[10]}}, p1_bit_slice_5271} + p1_bit_slice_5324;
  assign p2_add_5478_comb = {{2{p1_bit_slice_5283[10]}}, p1_bit_slice_5283} + p1_bit_slice_5335;
  assign p2_add_5479_comb = p1_bit_slice_5336 + {{2{p1_bit_slice_5286[10]}}, p1_bit_slice_5286};
  assign p2_add_5480_comb = {{1{p1_bit_slice_5289[11]}}, p1_bit_slice_5289} + p1_bit_slice_5339;
  assign p2_add_5481_comb = {{1{p1_bit_slice_5291[11]}}, p1_bit_slice_5291} + p1_bit_slice_5340;
  assign p2_add_5482_comb = p1_bit_slice_5341 + {{1{p1_bit_slice_5294[11]}}, p1_bit_slice_5294};
  assign p2_add_5483_comb = p1_bit_slice_5342 + {{1{p1_bit_slice_5296[11]}}, p1_bit_slice_5296};
  assign p2_add_5484_comb = {{2{p1_bit_slice_5297[10]}}, p1_bit_slice_5297} + p1_bit_slice_5343;
  assign p2_add_5485_comb = p1_bit_slice_5348 + {{2{p1_bit_slice_5304[10]}}, p1_bit_slice_5304};
  assign p2_sum__77_comb = p2_sum__97_comb + p2_sum__98_comb;
  assign p2_sum__78_comb = p2_sum__99_comb + p2_sum__100_comb;
  assign p2_sum__109_comb = {{12{p1_add_5351[12]}}, p1_add_5351};
  assign p2_sum__110_comb = {{12{p2_add_5470_comb[12]}}, p2_add_5470_comb};
  assign p2_sum__111_comb = {{12{p2_add_5471_comb[12]}}, p2_add_5471_comb};
  assign p2_sum__112_comb = {{12{p1_add_5352[12]}}, p1_add_5352};
  assign p2_sum__105_comb = {{12{p2_add_5472_comb[12]}}, p2_add_5472_comb};
  assign p2_sum__106_comb = {{12{p2_add_5473_comb[12]}}, p2_add_5473_comb};
  assign p2_sum__107_comb = {{12{p2_add_5474_comb[12]}}, p2_add_5474_comb};
  assign p2_sum__108_comb = {{12{p2_add_5475_comb[12]}}, p2_add_5475_comb};
  assign p2_sum__101_comb = {{12{p2_add_5476_comb[12]}}, p2_add_5476_comb};
  assign p2_sum__102_comb = {{12{p1_add_5353[12]}}, p1_add_5353};
  assign p2_sum__103_comb = {{12{p1_add_5354[12]}}, p1_add_5354};
  assign p2_sum__104_comb = {{12{p2_add_5477_comb[12]}}, p2_add_5477_comb};
  assign p2_sum__93_comb = {{12{p1_add_5359[12]}}, p1_add_5359};
  assign p2_sum__94_comb = {{12{p2_add_5478_comb[12]}}, p2_add_5478_comb};
  assign p2_sum__95_comb = {{12{p2_add_5479_comb[12]}}, p2_add_5479_comb};
  assign p2_sum__96_comb = {{12{p1_add_5360[12]}}, p1_add_5360};
  assign p2_sum__89_comb = {{12{p2_add_5480_comb[12]}}, p2_add_5480_comb};
  assign p2_sum__90_comb = {{12{p2_add_5481_comb[12]}}, p2_add_5481_comb};
  assign p2_sum__91_comb = {{12{p2_add_5482_comb[12]}}, p2_add_5482_comb};
  assign p2_sum__92_comb = {{12{p2_add_5483_comb[12]}}, p2_add_5483_comb};
  assign p2_sum__85_comb = {{12{p2_add_5484_comb[12]}}, p2_add_5484_comb};
  assign p2_sum__86_comb = {{12{p1_add_5361[12]}}, p1_add_5361};
  assign p2_sum__87_comb = {{12{p1_add_5362[12]}}, p1_add_5362};
  assign p2_sum__88_comb = {{12{p2_add_5485_comb[12]}}, p2_add_5485_comb};
  assign p2_sum__67_comb = p2_sum__77_comb + p2_sum__78_comb;
  assign p2_add_5546_comb = p2_umul_5515_comb[31:7] + 25'h000_0001;
  assign p2_sum__83_comb = p2_sum__109_comb + p2_sum__110_comb;
  assign p2_sum__84_comb = p2_sum__111_comb + p2_sum__112_comb;
  assign p2_sum__81_comb = p2_sum__105_comb + p2_sum__106_comb;
  assign p2_sum__82_comb = p2_sum__107_comb + p2_sum__108_comb;
  assign p2_sum__79_comb = p2_sum__101_comb + p2_sum__102_comb;
  assign p2_sum__80_comb = p2_sum__103_comb + p2_sum__104_comb;
  assign p2_sum__75_comb = p2_sum__93_comb + p2_sum__94_comb;
  assign p2_sum__76_comb = p2_sum__95_comb + p2_sum__96_comb;
  assign p2_sum__73_comb = p2_sum__89_comb + p2_sum__90_comb;
  assign p2_sum__74_comb = p2_sum__91_comb + p2_sum__92_comb;
  assign p2_sum__71_comb = p2_sum__85_comb + p2_sum__86_comb;
  assign p2_sum__72_comb = p2_sum__87_comb + p2_sum__88_comb;
  assign p2_add_5550_comb = p2_sum__67_comb + 25'h000_0001;
  assign p2_sum__70_comb = p2_sum__83_comb + p2_sum__84_comb;
  assign p2_sum__69_comb = p2_sum__81_comb + p2_sum__82_comb;
  assign p2_sum__68_comb = p2_sum__79_comb + p2_sum__80_comb;
  assign p2_sum__66_comb = p2_sum__75_comb + p2_sum__76_comb;
  assign p2_sum__65_comb = p2_sum__73_comb + p2_sum__74_comb;
  assign p2_sum__64_comb = p2_sum__71_comb + p2_sum__72_comb;
  assign p2_add_5547_comb = p2_sum__70_comb + 25'h000_0001;
  assign p2_add_5548_comb = p2_sum__69_comb + 25'h000_0001;
  assign p2_add_5549_comb = p2_sum__68_comb + 25'h000_0001;
  assign p2_add_5551_comb = p2_sum__66_comb + 25'h000_0001;
  assign p2_add_5552_comb = p2_sum__65_comb + 25'h000_0001;
  assign p2_add_5553_comb = p2_sum__64_comb + 25'h000_0001;
  assign p2_sgt_5563_comb = $signed(p2_add_5550_comb[24:1]) > $signed(24'h00_07ff);
  assign p2_bit_slice_5564_comb = p2_add_5550_comb[12:1];
  assign p2_slt_5565_comb = $signed(p2_add_5546_comb[24:1]) < $signed(24'hff_f800);
  assign p2_sel_5566_comb = $signed(p2_add_5546_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p2_add_5546_comb[12:1];
  assign p2_slt_5567_comb = $signed(p2_add_5550_comb[24:1]) < $signed(24'hff_f800);

  // Registers for pipe stage 2:
  reg [24:0] p2_add_5547;
  reg [24:0] p2_add_5548;
  reg [24:0] p2_add_5549;
  reg [24:0] p2_add_5551;
  reg [24:0] p2_add_5552;
  reg [24:0] p2_add_5553;
  reg p2_sgt_5563;
  reg [11:0] p2_bit_slice_5564;
  reg p2_slt_5565;
  reg [11:0] p2_sel_5566;
  reg p2_slt_5567;
  always @ (posedge clk) begin
    p2_add_5547 <= p2_add_5547_comb;
    p2_add_5548 <= p2_add_5548_comb;
    p2_add_5549 <= p2_add_5549_comb;
    p2_add_5551 <= p2_add_5551_comb;
    p2_add_5552 <= p2_add_5552_comb;
    p2_add_5553 <= p2_add_5553_comb;
    p2_sgt_5563 <= p2_sgt_5563_comb;
    p2_bit_slice_5564 <= p2_bit_slice_5564_comb;
    p2_slt_5565 <= p2_slt_5565_comb;
    p2_sel_5566 <= p2_sel_5566_comb;
    p2_slt_5567 <= p2_slt_5567_comb;
  end

  // ===== Pipe stage 3:
  wire [11:0] p3_clipped__8_comb;
  wire [11:0] p3_clipped__9_comb;
  wire [11:0] p3_clipped__10_comb;
  wire [11:0] p3_clipped__11_comb;
  wire [11:0] p3_clipped__12_comb;
  wire [11:0] p3_clipped__13_comb;
  wire [11:0] p3_clipped__14_comb;
  wire [11:0] p3_clipped__15_comb;
  wire [11:0] p3_result_comb[0:7];
  assign p3_clipped__8_comb = p2_slt_5565 ? 12'h800 : p2_sel_5566;
  assign p3_clipped__9_comb = $signed(p2_add_5547[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p2_add_5547[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p2_add_5547[12:1]);
  assign p3_clipped__10_comb = $signed(p2_add_5548[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p2_add_5548[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p2_add_5548[12:1]);
  assign p3_clipped__11_comb = $signed(p2_add_5549[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p2_add_5549[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p2_add_5549[12:1]);
  assign p3_clipped__12_comb = p2_slt_5567 ? 12'h800 : (p2_sgt_5563 ? 12'h7ff : p2_bit_slice_5564);
  assign p3_clipped__13_comb = $signed(p2_add_5551[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p2_add_5551[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p2_add_5551[12:1]);
  assign p3_clipped__14_comb = $signed(p2_add_5552[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p2_add_5552[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p2_add_5552[12:1]);
  assign p3_clipped__15_comb = $signed(p2_add_5553[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p2_add_5553[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p2_add_5553[12:1]);
  assign p3_result_comb[0] = p3_clipped__8_comb;
  assign p3_result_comb[1] = p3_clipped__9_comb;
  assign p3_result_comb[2] = p3_clipped__10_comb;
  assign p3_result_comb[3] = p3_clipped__11_comb;
  assign p3_result_comb[4] = p3_clipped__12_comb;
  assign p3_result_comb[5] = p3_clipped__13_comb;
  assign p3_result_comb[6] = p3_clipped__14_comb;
  assign p3_result_comb[7] = p3_clipped__15_comb;

  // Registers for pipe stage 3:
  reg [11:0] p3_result[0:7];
  always @ (posedge clk) begin
    p3_result[0] <= p3_result_comb[0];
    p3_result[1] <= p3_result_comb[1];
    p3_result[2] <= p3_result_comb[2];
    p3_result[3] <= p3_result_comb[3];
    p3_result[4] <= p3_result_comb[4];
    p3_result[5] <= p3_result_comb[5];
    p3_result[6] <= p3_result_comb[6];
    p3_result[7] <= p3_result_comb[7];
  end
  assign out = {p3_result[7], p3_result[6], p3_result[5], p3_result[4], p3_result[3], p3_result[2], p3_result[1], p3_result[0]};
endmodule
