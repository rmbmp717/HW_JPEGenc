module Huffman_ACenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [35:0] out
);
  wire [4:0] literal_9079[0:251];
  assign literal_9079[0] = 5'h02;
  assign literal_9079[1] = 5'h02;
  assign literal_9079[2] = 5'h03;
  assign literal_9079[3] = 5'h04;
  assign literal_9079[4] = 5'h05;
  assign literal_9079[5] = 5'h07;
  assign literal_9079[6] = 5'h08;
  assign literal_9079[7] = 5'h0e;
  assign literal_9079[8] = 5'h10;
  assign literal_9079[9] = 5'h10;
  assign literal_9079[10] = 5'h10;
  assign literal_9079[11] = 5'h00;
  assign literal_9079[12] = 5'h00;
  assign literal_9079[13] = 5'h00;
  assign literal_9079[14] = 5'h00;
  assign literal_9079[15] = 5'h00;
  assign literal_9079[16] = 5'h00;
  assign literal_9079[17] = 5'h03;
  assign literal_9079[18] = 5'h06;
  assign literal_9079[19] = 5'h07;
  assign literal_9079[20] = 5'h09;
  assign literal_9079[21] = 5'h0b;
  assign literal_9079[22] = 5'h0d;
  assign literal_9079[23] = 5'h10;
  assign literal_9079[24] = 5'h10;
  assign literal_9079[25] = 5'h10;
  assign literal_9079[26] = 5'h10;
  assign literal_9079[27] = 5'h00;
  assign literal_9079[28] = 5'h00;
  assign literal_9079[29] = 5'h00;
  assign literal_9079[30] = 5'h00;
  assign literal_9079[31] = 5'h00;
  assign literal_9079[32] = 5'h00;
  assign literal_9079[33] = 5'h05;
  assign literal_9079[34] = 5'h07;
  assign literal_9079[35] = 5'h0a;
  assign literal_9079[36] = 5'h0c;
  assign literal_9079[37] = 5'h0d;
  assign literal_9079[38] = 5'h10;
  assign literal_9079[39] = 5'h10;
  assign literal_9079[40] = 5'h10;
  assign literal_9079[41] = 5'h10;
  assign literal_9079[42] = 5'h10;
  assign literal_9079[43] = 5'h00;
  assign literal_9079[44] = 5'h00;
  assign literal_9079[45] = 5'h00;
  assign literal_9079[46] = 5'h00;
  assign literal_9079[47] = 5'h00;
  assign literal_9079[48] = 5'h00;
  assign literal_9079[49] = 5'h06;
  assign literal_9079[50] = 5'h08;
  assign literal_9079[51] = 5'h0b;
  assign literal_9079[52] = 5'h0c;
  assign literal_9079[53] = 5'h0f;
  assign literal_9079[54] = 5'h10;
  assign literal_9079[55] = 5'h10;
  assign literal_9079[56] = 5'h10;
  assign literal_9079[57] = 5'h10;
  assign literal_9079[58] = 5'h10;
  assign literal_9079[59] = 5'h00;
  assign literal_9079[60] = 5'h00;
  assign literal_9079[61] = 5'h00;
  assign literal_9079[62] = 5'h00;
  assign literal_9079[63] = 5'h00;
  assign literal_9079[64] = 5'h00;
  assign literal_9079[65] = 5'h06;
  assign literal_9079[66] = 5'h0a;
  assign literal_9079[67] = 5'h0c;
  assign literal_9079[68] = 5'h0f;
  assign literal_9079[69] = 5'h10;
  assign literal_9079[70] = 5'h10;
  assign literal_9079[71] = 5'h10;
  assign literal_9079[72] = 5'h10;
  assign literal_9079[73] = 5'h10;
  assign literal_9079[74] = 5'h10;
  assign literal_9079[75] = 5'h00;
  assign literal_9079[76] = 5'h00;
  assign literal_9079[77] = 5'h00;
  assign literal_9079[78] = 5'h00;
  assign literal_9079[79] = 5'h00;
  assign literal_9079[80] = 5'h00;
  assign literal_9079[81] = 5'h07;
  assign literal_9079[82] = 5'h0b;
  assign literal_9079[83] = 5'h0d;
  assign literal_9079[84] = 5'h10;
  assign literal_9079[85] = 5'h10;
  assign literal_9079[86] = 5'h10;
  assign literal_9079[87] = 5'h10;
  assign literal_9079[88] = 5'h10;
  assign literal_9079[89] = 5'h10;
  assign literal_9079[90] = 5'h10;
  assign literal_9079[91] = 5'h00;
  assign literal_9079[92] = 5'h00;
  assign literal_9079[93] = 5'h00;
  assign literal_9079[94] = 5'h00;
  assign literal_9079[95] = 5'h00;
  assign literal_9079[96] = 5'h00;
  assign literal_9079[97] = 5'h07;
  assign literal_9079[98] = 5'h0b;
  assign literal_9079[99] = 5'h0d;
  assign literal_9079[100] = 5'h10;
  assign literal_9079[101] = 5'h10;
  assign literal_9079[102] = 5'h10;
  assign literal_9079[103] = 5'h10;
  assign literal_9079[104] = 5'h10;
  assign literal_9079[105] = 5'h10;
  assign literal_9079[106] = 5'h10;
  assign literal_9079[107] = 5'h00;
  assign literal_9079[108] = 5'h00;
  assign literal_9079[109] = 5'h00;
  assign literal_9079[110] = 5'h00;
  assign literal_9079[111] = 5'h00;
  assign literal_9079[112] = 5'h00;
  assign literal_9079[113] = 5'h08;
  assign literal_9079[114] = 5'h0b;
  assign literal_9079[115] = 5'h0e;
  assign literal_9079[116] = 5'h10;
  assign literal_9079[117] = 5'h10;
  assign literal_9079[118] = 5'h10;
  assign literal_9079[119] = 5'h10;
  assign literal_9079[120] = 5'h10;
  assign literal_9079[121] = 5'h10;
  assign literal_9079[122] = 5'h10;
  assign literal_9079[123] = 5'h00;
  assign literal_9079[124] = 5'h00;
  assign literal_9079[125] = 5'h00;
  assign literal_9079[126] = 5'h00;
  assign literal_9079[127] = 5'h00;
  assign literal_9079[128] = 5'h00;
  assign literal_9079[129] = 5'h08;
  assign literal_9079[130] = 5'h0c;
  assign literal_9079[131] = 5'h10;
  assign literal_9079[132] = 5'h10;
  assign literal_9079[133] = 5'h10;
  assign literal_9079[134] = 5'h10;
  assign literal_9079[135] = 5'h10;
  assign literal_9079[136] = 5'h10;
  assign literal_9079[137] = 5'h10;
  assign literal_9079[138] = 5'h10;
  assign literal_9079[139] = 5'h00;
  assign literal_9079[140] = 5'h00;
  assign literal_9079[141] = 5'h00;
  assign literal_9079[142] = 5'h00;
  assign literal_9079[143] = 5'h00;
  assign literal_9079[144] = 5'h00;
  assign literal_9079[145] = 5'h08;
  assign literal_9079[146] = 5'h0d;
  assign literal_9079[147] = 5'h10;
  assign literal_9079[148] = 5'h10;
  assign literal_9079[149] = 5'h10;
  assign literal_9079[150] = 5'h10;
  assign literal_9079[151] = 5'h10;
  assign literal_9079[152] = 5'h10;
  assign literal_9079[153] = 5'h10;
  assign literal_9079[154] = 5'h10;
  assign literal_9079[155] = 5'h00;
  assign literal_9079[156] = 5'h00;
  assign literal_9079[157] = 5'h00;
  assign literal_9079[158] = 5'h00;
  assign literal_9079[159] = 5'h00;
  assign literal_9079[160] = 5'h00;
  assign literal_9079[161] = 5'h09;
  assign literal_9079[162] = 5'h0d;
  assign literal_9079[163] = 5'h10;
  assign literal_9079[164] = 5'h10;
  assign literal_9079[165] = 5'h10;
  assign literal_9079[166] = 5'h10;
  assign literal_9079[167] = 5'h10;
  assign literal_9079[168] = 5'h10;
  assign literal_9079[169] = 5'h10;
  assign literal_9079[170] = 5'h10;
  assign literal_9079[171] = 5'h00;
  assign literal_9079[172] = 5'h00;
  assign literal_9079[173] = 5'h00;
  assign literal_9079[174] = 5'h00;
  assign literal_9079[175] = 5'h00;
  assign literal_9079[176] = 5'h00;
  assign literal_9079[177] = 5'h09;
  assign literal_9079[178] = 5'h0d;
  assign literal_9079[179] = 5'h10;
  assign literal_9079[180] = 5'h10;
  assign literal_9079[181] = 5'h10;
  assign literal_9079[182] = 5'h10;
  assign literal_9079[183] = 5'h10;
  assign literal_9079[184] = 5'h10;
  assign literal_9079[185] = 5'h10;
  assign literal_9079[186] = 5'h10;
  assign literal_9079[187] = 5'h00;
  assign literal_9079[188] = 5'h00;
  assign literal_9079[189] = 5'h00;
  assign literal_9079[190] = 5'h00;
  assign literal_9079[191] = 5'h00;
  assign literal_9079[192] = 5'h00;
  assign literal_9079[193] = 5'h0a;
  assign literal_9079[194] = 5'h0d;
  assign literal_9079[195] = 5'h10;
  assign literal_9079[196] = 5'h10;
  assign literal_9079[197] = 5'h10;
  assign literal_9079[198] = 5'h10;
  assign literal_9079[199] = 5'h10;
  assign literal_9079[200] = 5'h10;
  assign literal_9079[201] = 5'h10;
  assign literal_9079[202] = 5'h10;
  assign literal_9079[203] = 5'h00;
  assign literal_9079[204] = 5'h00;
  assign literal_9079[205] = 5'h00;
  assign literal_9079[206] = 5'h00;
  assign literal_9079[207] = 5'h00;
  assign literal_9079[208] = 5'h00;
  assign literal_9079[209] = 5'h0a;
  assign literal_9079[210] = 5'h0e;
  assign literal_9079[211] = 5'h10;
  assign literal_9079[212] = 5'h10;
  assign literal_9079[213] = 5'h10;
  assign literal_9079[214] = 5'h10;
  assign literal_9079[215] = 5'h10;
  assign literal_9079[216] = 5'h10;
  assign literal_9079[217] = 5'h10;
  assign literal_9079[218] = 5'h10;
  assign literal_9079[219] = 5'h00;
  assign literal_9079[220] = 5'h00;
  assign literal_9079[221] = 5'h00;
  assign literal_9079[222] = 5'h00;
  assign literal_9079[223] = 5'h00;
  assign literal_9079[224] = 5'h00;
  assign literal_9079[225] = 5'h0a;
  assign literal_9079[226] = 5'h0f;
  assign literal_9079[227] = 5'h10;
  assign literal_9079[228] = 5'h10;
  assign literal_9079[229] = 5'h10;
  assign literal_9079[230] = 5'h10;
  assign literal_9079[231] = 5'h10;
  assign literal_9079[232] = 5'h10;
  assign literal_9079[233] = 5'h10;
  assign literal_9079[234] = 5'h10;
  assign literal_9079[235] = 5'h00;
  assign literal_9079[236] = 5'h00;
  assign literal_9079[237] = 5'h00;
  assign literal_9079[238] = 5'h00;
  assign literal_9079[239] = 5'h00;
  assign literal_9079[240] = 5'h09;
  assign literal_9079[241] = 5'h0b;
  assign literal_9079[242] = 5'h10;
  assign literal_9079[243] = 5'h10;
  assign literal_9079[244] = 5'h10;
  assign literal_9079[245] = 5'h10;
  assign literal_9079[246] = 5'h10;
  assign literal_9079[247] = 5'h10;
  assign literal_9079[248] = 5'h10;
  assign literal_9079[249] = 5'h10;
  assign literal_9079[250] = 5'h10;
  assign literal_9079[251] = 5'h00;
  wire [4:0] literal_9081[0:251];
  assign literal_9081[0] = 5'h04;
  assign literal_9081[1] = 5'h02;
  assign literal_9081[2] = 5'h02;
  assign literal_9081[3] = 5'h03;
  assign literal_9081[4] = 5'h04;
  assign literal_9081[5] = 5'h05;
  assign literal_9081[6] = 5'h07;
  assign literal_9081[7] = 5'h09;
  assign literal_9081[8] = 5'h10;
  assign literal_9081[9] = 5'h10;
  assign literal_9081[10] = 5'h10;
  assign literal_9081[11] = 5'h00;
  assign literal_9081[12] = 5'h00;
  assign literal_9081[13] = 5'h00;
  assign literal_9081[14] = 5'h00;
  assign literal_9081[15] = 5'h00;
  assign literal_9081[16] = 5'h00;
  assign literal_9081[17] = 5'h04;
  assign literal_9081[18] = 5'h05;
  assign literal_9081[19] = 5'h07;
  assign literal_9081[20] = 5'h09;
  assign literal_9081[21] = 5'h0a;
  assign literal_9081[22] = 5'h0b;
  assign literal_9081[23] = 5'h10;
  assign literal_9081[24] = 5'h10;
  assign literal_9081[25] = 5'h10;
  assign literal_9081[26] = 5'h10;
  assign literal_9081[27] = 5'h00;
  assign literal_9081[28] = 5'h00;
  assign literal_9081[29] = 5'h00;
  assign literal_9081[30] = 5'h00;
  assign literal_9081[31] = 5'h00;
  assign literal_9081[32] = 5'h00;
  assign literal_9081[33] = 5'h05;
  assign literal_9081[34] = 5'h08;
  assign literal_9081[35] = 5'h0a;
  assign literal_9081[36] = 5'h0c;
  assign literal_9081[37] = 5'h0e;
  assign literal_9081[38] = 5'h10;
  assign literal_9081[39] = 5'h10;
  assign literal_9081[40] = 5'h10;
  assign literal_9081[41] = 5'h10;
  assign literal_9081[42] = 5'h10;
  assign literal_9081[43] = 5'h00;
  assign literal_9081[44] = 5'h00;
  assign literal_9081[45] = 5'h00;
  assign literal_9081[46] = 5'h00;
  assign literal_9081[47] = 5'h00;
  assign literal_9081[48] = 5'h00;
  assign literal_9081[49] = 5'h06;
  assign literal_9081[50] = 5'h09;
  assign literal_9081[51] = 5'h0b;
  assign literal_9081[52] = 5'h0e;
  assign literal_9081[53] = 5'h10;
  assign literal_9081[54] = 5'h10;
  assign literal_9081[55] = 5'h10;
  assign literal_9081[56] = 5'h10;
  assign literal_9081[57] = 5'h10;
  assign literal_9081[58] = 5'h10;
  assign literal_9081[59] = 5'h00;
  assign literal_9081[60] = 5'h00;
  assign literal_9081[61] = 5'h00;
  assign literal_9081[62] = 5'h00;
  assign literal_9081[63] = 5'h00;
  assign literal_9081[64] = 5'h00;
  assign literal_9081[65] = 5'h06;
  assign literal_9081[66] = 5'h0a;
  assign literal_9081[67] = 5'h0e;
  assign literal_9081[68] = 5'h10;
  assign literal_9081[69] = 5'h10;
  assign literal_9081[70] = 5'h10;
  assign literal_9081[71] = 5'h10;
  assign literal_9081[72] = 5'h10;
  assign literal_9081[73] = 5'h10;
  assign literal_9081[74] = 5'h10;
  assign literal_9081[75] = 5'h00;
  assign literal_9081[76] = 5'h00;
  assign literal_9081[77] = 5'h00;
  assign literal_9081[78] = 5'h00;
  assign literal_9081[79] = 5'h00;
  assign literal_9081[80] = 5'h00;
  assign literal_9081[81] = 5'h07;
  assign literal_9081[82] = 5'h0a;
  assign literal_9081[83] = 5'h0e;
  assign literal_9081[84] = 5'h10;
  assign literal_9081[85] = 5'h10;
  assign literal_9081[86] = 5'h10;
  assign literal_9081[87] = 5'h10;
  assign literal_9081[88] = 5'h10;
  assign literal_9081[89] = 5'h10;
  assign literal_9081[90] = 5'h10;
  assign literal_9081[91] = 5'h00;
  assign literal_9081[92] = 5'h00;
  assign literal_9081[93] = 5'h00;
  assign literal_9081[94] = 5'h00;
  assign literal_9081[95] = 5'h00;
  assign literal_9081[96] = 5'h00;
  assign literal_9081[97] = 5'h07;
  assign literal_9081[98] = 5'h0c;
  assign literal_9081[99] = 5'h0f;
  assign literal_9081[100] = 5'h10;
  assign literal_9081[101] = 5'h10;
  assign literal_9081[102] = 5'h10;
  assign literal_9081[103] = 5'h10;
  assign literal_9081[104] = 5'h10;
  assign literal_9081[105] = 5'h10;
  assign literal_9081[106] = 5'h10;
  assign literal_9081[107] = 5'h00;
  assign literal_9081[108] = 5'h00;
  assign literal_9081[109] = 5'h00;
  assign literal_9081[110] = 5'h00;
  assign literal_9081[111] = 5'h00;
  assign literal_9081[112] = 5'h00;
  assign literal_9081[113] = 5'h08;
  assign literal_9081[114] = 5'h0c;
  assign literal_9081[115] = 5'h10;
  assign literal_9081[116] = 5'h10;
  assign literal_9081[117] = 5'h10;
  assign literal_9081[118] = 5'h10;
  assign literal_9081[119] = 5'h10;
  assign literal_9081[120] = 5'h10;
  assign literal_9081[121] = 5'h10;
  assign literal_9081[122] = 5'h10;
  assign literal_9081[123] = 5'h00;
  assign literal_9081[124] = 5'h00;
  assign literal_9081[125] = 5'h00;
  assign literal_9081[126] = 5'h00;
  assign literal_9081[127] = 5'h00;
  assign literal_9081[128] = 5'h00;
  assign literal_9081[129] = 5'h09;
  assign literal_9081[130] = 5'h0d;
  assign literal_9081[131] = 5'h10;
  assign literal_9081[132] = 5'h10;
  assign literal_9081[133] = 5'h10;
  assign literal_9081[134] = 5'h10;
  assign literal_9081[135] = 5'h10;
  assign literal_9081[136] = 5'h10;
  assign literal_9081[137] = 5'h10;
  assign literal_9081[138] = 5'h10;
  assign literal_9081[139] = 5'h00;
  assign literal_9081[140] = 5'h00;
  assign literal_9081[141] = 5'h00;
  assign literal_9081[142] = 5'h00;
  assign literal_9081[143] = 5'h00;
  assign literal_9081[144] = 5'h00;
  assign literal_9081[145] = 5'h09;
  assign literal_9081[146] = 5'h0e;
  assign literal_9081[147] = 5'h10;
  assign literal_9081[148] = 5'h10;
  assign literal_9081[149] = 5'h10;
  assign literal_9081[150] = 5'h10;
  assign literal_9081[151] = 5'h10;
  assign literal_9081[152] = 5'h10;
  assign literal_9081[153] = 5'h10;
  assign literal_9081[154] = 5'h10;
  assign literal_9081[155] = 5'h00;
  assign literal_9081[156] = 5'h00;
  assign literal_9081[157] = 5'h00;
  assign literal_9081[158] = 5'h00;
  assign literal_9081[159] = 5'h00;
  assign literal_9081[160] = 5'h00;
  assign literal_9081[161] = 5'h09;
  assign literal_9081[162] = 5'h0e;
  assign literal_9081[163] = 5'h10;
  assign literal_9081[164] = 5'h10;
  assign literal_9081[165] = 5'h10;
  assign literal_9081[166] = 5'h10;
  assign literal_9081[167] = 5'h10;
  assign literal_9081[168] = 5'h10;
  assign literal_9081[169] = 5'h10;
  assign literal_9081[170] = 5'h10;
  assign literal_9081[171] = 5'h00;
  assign literal_9081[172] = 5'h00;
  assign literal_9081[173] = 5'h00;
  assign literal_9081[174] = 5'h00;
  assign literal_9081[175] = 5'h00;
  assign literal_9081[176] = 5'h00;
  assign literal_9081[177] = 5'h0a;
  assign literal_9081[178] = 5'h0f;
  assign literal_9081[179] = 5'h10;
  assign literal_9081[180] = 5'h10;
  assign literal_9081[181] = 5'h10;
  assign literal_9081[182] = 5'h10;
  assign literal_9081[183] = 5'h10;
  assign literal_9081[184] = 5'h10;
  assign literal_9081[185] = 5'h10;
  assign literal_9081[186] = 5'h10;
  assign literal_9081[187] = 5'h00;
  assign literal_9081[188] = 5'h00;
  assign literal_9081[189] = 5'h00;
  assign literal_9081[190] = 5'h00;
  assign literal_9081[191] = 5'h00;
  assign literal_9081[192] = 5'h00;
  assign literal_9081[193] = 5'h0a;
  assign literal_9081[194] = 5'h10;
  assign literal_9081[195] = 5'h10;
  assign literal_9081[196] = 5'h10;
  assign literal_9081[197] = 5'h10;
  assign literal_9081[198] = 5'h10;
  assign literal_9081[199] = 5'h10;
  assign literal_9081[200] = 5'h10;
  assign literal_9081[201] = 5'h10;
  assign literal_9081[202] = 5'h10;
  assign literal_9081[203] = 5'h00;
  assign literal_9081[204] = 5'h00;
  assign literal_9081[205] = 5'h00;
  assign literal_9081[206] = 5'h00;
  assign literal_9081[207] = 5'h00;
  assign literal_9081[208] = 5'h00;
  assign literal_9081[209] = 5'h0a;
  assign literal_9081[210] = 5'h10;
  assign literal_9081[211] = 5'h10;
  assign literal_9081[212] = 5'h10;
  assign literal_9081[213] = 5'h10;
  assign literal_9081[214] = 5'h10;
  assign literal_9081[215] = 5'h10;
  assign literal_9081[216] = 5'h10;
  assign literal_9081[217] = 5'h10;
  assign literal_9081[218] = 5'h10;
  assign literal_9081[219] = 5'h00;
  assign literal_9081[220] = 5'h00;
  assign literal_9081[221] = 5'h00;
  assign literal_9081[222] = 5'h00;
  assign literal_9081[223] = 5'h00;
  assign literal_9081[224] = 5'h00;
  assign literal_9081[225] = 5'h0b;
  assign literal_9081[226] = 5'h10;
  assign literal_9081[227] = 5'h10;
  assign literal_9081[228] = 5'h10;
  assign literal_9081[229] = 5'h10;
  assign literal_9081[230] = 5'h10;
  assign literal_9081[231] = 5'h10;
  assign literal_9081[232] = 5'h10;
  assign literal_9081[233] = 5'h10;
  assign literal_9081[234] = 5'h10;
  assign literal_9081[235] = 5'h00;
  assign literal_9081[236] = 5'h00;
  assign literal_9081[237] = 5'h00;
  assign literal_9081[238] = 5'h00;
  assign literal_9081[239] = 5'h00;
  assign literal_9081[240] = 5'h0c;
  assign literal_9081[241] = 5'h0d;
  assign literal_9081[242] = 5'h10;
  assign literal_9081[243] = 5'h10;
  assign literal_9081[244] = 5'h10;
  assign literal_9081[245] = 5'h10;
  assign literal_9081[246] = 5'h10;
  assign literal_9081[247] = 5'h10;
  assign literal_9081[248] = 5'h10;
  assign literal_9081[249] = 5'h10;
  assign literal_9081[250] = 5'h10;
  assign literal_9081[251] = 5'h00;
  wire [15:0] literal_9082[0:251];
  assign literal_9082[0] = 16'h0001;
  assign literal_9082[1] = 16'h0000;
  assign literal_9082[2] = 16'h0004;
  assign literal_9082[3] = 16'h000c;
  assign literal_9082[4] = 16'h001a;
  assign literal_9082[5] = 16'h0076;
  assign literal_9082[6] = 16'h00f6;
  assign literal_9082[7] = 16'h3fe0;
  assign literal_9082[8] = 16'hff96;
  assign literal_9082[9] = 16'hff97;
  assign literal_9082[10] = 16'hff98;
  assign literal_9082[11] = 16'h0000;
  assign literal_9082[12] = 16'h0000;
  assign literal_9082[13] = 16'h0000;
  assign literal_9082[14] = 16'h0000;
  assign literal_9082[15] = 16'h0000;
  assign literal_9082[16] = 16'h0000;
  assign literal_9082[17] = 16'h0005;
  assign literal_9082[18] = 16'h0038;
  assign literal_9082[19] = 16'h0078;
  assign literal_9082[20] = 16'h01f9;
  assign literal_9082[21] = 16'h07f2;
  assign literal_9082[22] = 16'h1fe8;
  assign literal_9082[23] = 16'hff93;
  assign literal_9082[24] = 16'hff99;
  assign literal_9082[25] = 16'hff9a;
  assign literal_9082[26] = 16'hff9e;
  assign literal_9082[27] = 16'h0000;
  assign literal_9082[28] = 16'h0000;
  assign literal_9082[29] = 16'h0000;
  assign literal_9082[30] = 16'h0000;
  assign literal_9082[31] = 16'h0000;
  assign literal_9082[32] = 16'h0000;
  assign literal_9082[33] = 16'h001b;
  assign literal_9082[34] = 16'h007a;
  assign literal_9082[35] = 16'h03f7;
  assign literal_9082[36] = 16'h0ff0;
  assign literal_9082[37] = 16'h1feb;
  assign literal_9082[38] = 16'hff9b;
  assign literal_9082[39] = 16'hff9f;
  assign literal_9082[40] = 16'hffa8;
  assign literal_9082[41] = 16'hffa9;
  assign literal_9082[42] = 16'hfff1;
  assign literal_9082[43] = 16'h0000;
  assign literal_9082[44] = 16'h0000;
  assign literal_9082[45] = 16'h0000;
  assign literal_9082[46] = 16'h0000;
  assign literal_9082[47] = 16'h0000;
  assign literal_9082[48] = 16'h0000;
  assign literal_9082[49] = 16'h0039;
  assign literal_9082[50] = 16'h00fa;
  assign literal_9082[51] = 16'h07f7;
  assign literal_9082[52] = 16'h0ff1;
  assign literal_9082[53] = 16'h7fc6;
  assign literal_9082[54] = 16'hff9c;
  assign literal_9082[55] = 16'hffa3;
  assign literal_9082[56] = 16'hffd7;
  assign literal_9082[57] = 16'hffe4;
  assign literal_9082[58] = 16'hfff2;
  assign literal_9082[59] = 16'h0000;
  assign literal_9082[60] = 16'h0000;
  assign literal_9082[61] = 16'h0000;
  assign literal_9082[62] = 16'h0000;
  assign literal_9082[63] = 16'h0000;
  assign literal_9082[64] = 16'h0000;
  assign literal_9082[65] = 16'h003a;
  assign literal_9082[66] = 16'h03f8;
  assign literal_9082[67] = 16'h0ff2;
  assign literal_9082[68] = 16'h7fc8;
  assign literal_9082[69] = 16'hff9d;
  assign literal_9082[70] = 16'hffbf;
  assign literal_9082[71] = 16'hffcb;
  assign literal_9082[72] = 16'hffd8;
  assign literal_9082[73] = 16'hffe5;
  assign literal_9082[74] = 16'hfff3;
  assign literal_9082[75] = 16'h0000;
  assign literal_9082[76] = 16'h0000;
  assign literal_9082[77] = 16'h0000;
  assign literal_9082[78] = 16'h0000;
  assign literal_9082[79] = 16'h0000;
  assign literal_9082[80] = 16'h0000;
  assign literal_9082[81] = 16'h0077;
  assign literal_9082[82] = 16'h07f3;
  assign literal_9082[83] = 16'h1fea;
  assign literal_9082[84] = 16'hff94;
  assign literal_9082[85] = 16'hffa2;
  assign literal_9082[86] = 16'hffc0;
  assign literal_9082[87] = 16'hffcc;
  assign literal_9082[88] = 16'hffd9;
  assign literal_9082[89] = 16'hffe6;
  assign literal_9082[90] = 16'hfff4;
  assign literal_9082[91] = 16'h0000;
  assign literal_9082[92] = 16'h0000;
  assign literal_9082[93] = 16'h0000;
  assign literal_9082[94] = 16'h0000;
  assign literal_9082[95] = 16'h0000;
  assign literal_9082[96] = 16'h0000;
  assign literal_9082[97] = 16'h0079;
  assign literal_9082[98] = 16'h07f4;
  assign literal_9082[99] = 16'h1fed;
  assign literal_9082[100] = 16'hffa0;
  assign literal_9082[101] = 16'hffb5;
  assign literal_9082[102] = 16'hffc1;
  assign literal_9082[103] = 16'hffcd;
  assign literal_9082[104] = 16'hffda;
  assign literal_9082[105] = 16'hffe7;
  assign literal_9082[106] = 16'hfff5;
  assign literal_9082[107] = 16'h0000;
  assign literal_9082[108] = 16'h0000;
  assign literal_9082[109] = 16'h0000;
  assign literal_9082[110] = 16'h0000;
  assign literal_9082[111] = 16'h0000;
  assign literal_9082[112] = 16'h0000;
  assign literal_9082[113] = 16'h00f7;
  assign literal_9082[114] = 16'h07f5;
  assign literal_9082[115] = 16'h3fe1;
  assign literal_9082[116] = 16'hffa1;
  assign literal_9082[117] = 16'hffb6;
  assign literal_9082[118] = 16'hffc2;
  assign literal_9082[119] = 16'hffce;
  assign literal_9082[120] = 16'hffdb;
  assign literal_9082[121] = 16'hffe8;
  assign literal_9082[122] = 16'hfff6;
  assign literal_9082[123] = 16'h0000;
  assign literal_9082[124] = 16'h0000;
  assign literal_9082[125] = 16'h0000;
  assign literal_9082[126] = 16'h0000;
  assign literal_9082[127] = 16'h0000;
  assign literal_9082[128] = 16'h0000;
  assign literal_9082[129] = 16'h00f8;
  assign literal_9082[130] = 16'h0ff3;
  assign literal_9082[131] = 16'hff92;
  assign literal_9082[132] = 16'hffad;
  assign literal_9082[133] = 16'hffb7;
  assign literal_9082[134] = 16'hffc3;
  assign literal_9082[135] = 16'hffcf;
  assign literal_9082[136] = 16'hffdc;
  assign literal_9082[137] = 16'hffe9;
  assign literal_9082[138] = 16'hfff7;
  assign literal_9082[139] = 16'h0000;
  assign literal_9082[140] = 16'h0000;
  assign literal_9082[141] = 16'h0000;
  assign literal_9082[142] = 16'h0000;
  assign literal_9082[143] = 16'h0000;
  assign literal_9082[144] = 16'h0000;
  assign literal_9082[145] = 16'h00f9;
  assign literal_9082[146] = 16'h1fe9;
  assign literal_9082[147] = 16'hff95;
  assign literal_9082[148] = 16'hffae;
  assign literal_9082[149] = 16'hffb8;
  assign literal_9082[150] = 16'hffc4;
  assign literal_9082[151] = 16'hffd0;
  assign literal_9082[152] = 16'hffdd;
  assign literal_9082[153] = 16'hffea;
  assign literal_9082[154] = 16'hfff8;
  assign literal_9082[155] = 16'h0000;
  assign literal_9082[156] = 16'h0000;
  assign literal_9082[157] = 16'h0000;
  assign literal_9082[158] = 16'h0000;
  assign literal_9082[159] = 16'h0000;
  assign literal_9082[160] = 16'h0000;
  assign literal_9082[161] = 16'h01f6;
  assign literal_9082[162] = 16'h1fec;
  assign literal_9082[163] = 16'hffa5;
  assign literal_9082[164] = 16'hffaf;
  assign literal_9082[165] = 16'hffb9;
  assign literal_9082[166] = 16'hffc5;
  assign literal_9082[167] = 16'hffd1;
  assign literal_9082[168] = 16'hffde;
  assign literal_9082[169] = 16'hffeb;
  assign literal_9082[170] = 16'hfff9;
  assign literal_9082[171] = 16'h0000;
  assign literal_9082[172] = 16'h0000;
  assign literal_9082[173] = 16'h0000;
  assign literal_9082[174] = 16'h0000;
  assign literal_9082[175] = 16'h0000;
  assign literal_9082[176] = 16'h0000;
  assign literal_9082[177] = 16'h01f7;
  assign literal_9082[178] = 16'h1fee;
  assign literal_9082[179] = 16'hffa6;
  assign literal_9082[180] = 16'hffb0;
  assign literal_9082[181] = 16'hffba;
  assign literal_9082[182] = 16'hffc6;
  assign literal_9082[183] = 16'hffd2;
  assign literal_9082[184] = 16'hffdf;
  assign literal_9082[185] = 16'hffec;
  assign literal_9082[186] = 16'hfffa;
  assign literal_9082[187] = 16'h0000;
  assign literal_9082[188] = 16'h0000;
  assign literal_9082[189] = 16'h0000;
  assign literal_9082[190] = 16'h0000;
  assign literal_9082[191] = 16'h0000;
  assign literal_9082[192] = 16'h0000;
  assign literal_9082[193] = 16'h03f4;
  assign literal_9082[194] = 16'h1fef;
  assign literal_9082[195] = 16'hffa7;
  assign literal_9082[196] = 16'hffb1;
  assign literal_9082[197] = 16'hffbb;
  assign literal_9082[198] = 16'hffc7;
  assign literal_9082[199] = 16'hffd3;
  assign literal_9082[200] = 16'hffe0;
  assign literal_9082[201] = 16'hffed;
  assign literal_9082[202] = 16'hfffb;
  assign literal_9082[203] = 16'h0000;
  assign literal_9082[204] = 16'h0000;
  assign literal_9082[205] = 16'h0000;
  assign literal_9082[206] = 16'h0000;
  assign literal_9082[207] = 16'h0000;
  assign literal_9082[208] = 16'h0000;
  assign literal_9082[209] = 16'h03f5;
  assign literal_9082[210] = 16'h3fe2;
  assign literal_9082[211] = 16'hffaa;
  assign literal_9082[212] = 16'hffb2;
  assign literal_9082[213] = 16'hffbc;
  assign literal_9082[214] = 16'hffc8;
  assign literal_9082[215] = 16'hffd4;
  assign literal_9082[216] = 16'hffe1;
  assign literal_9082[217] = 16'hffee;
  assign literal_9082[218] = 16'hfffc;
  assign literal_9082[219] = 16'h0000;
  assign literal_9082[220] = 16'h0000;
  assign literal_9082[221] = 16'h0000;
  assign literal_9082[222] = 16'h0000;
  assign literal_9082[223] = 16'h0000;
  assign literal_9082[224] = 16'h0000;
  assign literal_9082[225] = 16'h03f6;
  assign literal_9082[226] = 16'h7fc7;
  assign literal_9082[227] = 16'hffab;
  assign literal_9082[228] = 16'hffb3;
  assign literal_9082[229] = 16'hffbd;
  assign literal_9082[230] = 16'hffc9;
  assign literal_9082[231] = 16'hffd5;
  assign literal_9082[232] = 16'hffe2;
  assign literal_9082[233] = 16'hffef;
  assign literal_9082[234] = 16'hfffd;
  assign literal_9082[235] = 16'h0000;
  assign literal_9082[236] = 16'h0000;
  assign literal_9082[237] = 16'h0000;
  assign literal_9082[238] = 16'h0000;
  assign literal_9082[239] = 16'h0000;
  assign literal_9082[240] = 16'h01f8;
  assign literal_9082[241] = 16'h07f6;
  assign literal_9082[242] = 16'hffa4;
  assign literal_9082[243] = 16'hffac;
  assign literal_9082[244] = 16'hffb4;
  assign literal_9082[245] = 16'hffbe;
  assign literal_9082[246] = 16'hffca;
  assign literal_9082[247] = 16'hffd6;
  assign literal_9082[248] = 16'hffe3;
  assign literal_9082[249] = 16'hfff0;
  assign literal_9082[250] = 16'hfffe;
  assign literal_9082[251] = 16'h0000;
  wire [15:0] literal_9083[0:251];
  assign literal_9083[0] = 16'h000c;
  assign literal_9083[1] = 16'h0000;
  assign literal_9083[2] = 16'h0001;
  assign literal_9083[3] = 16'h0004;
  assign literal_9083[4] = 16'h000b;
  assign literal_9083[5] = 16'h001a;
  assign literal_9083[6] = 16'h0079;
  assign literal_9083[7] = 16'h01f9;
  assign literal_9083[8] = 16'hff9c;
  assign literal_9083[9] = 16'hff9f;
  assign literal_9083[10] = 16'hffa0;
  assign literal_9083[11] = 16'h0000;
  assign literal_9083[12] = 16'h0000;
  assign literal_9083[13] = 16'h0000;
  assign literal_9083[14] = 16'h0000;
  assign literal_9083[15] = 16'h0000;
  assign literal_9083[16] = 16'h0000;
  assign literal_9083[17] = 16'h000a;
  assign literal_9083[18] = 16'h001c;
  assign literal_9083[19] = 16'h007a;
  assign literal_9083[20] = 16'h01f5;
  assign literal_9083[21] = 16'h03f4;
  assign literal_9083[22] = 16'h07f8;
  assign literal_9083[23] = 16'hff95;
  assign literal_9083[24] = 16'hffa1;
  assign literal_9083[25] = 16'hffa2;
  assign literal_9083[26] = 16'hffad;
  assign literal_9083[27] = 16'h0000;
  assign literal_9083[28] = 16'h0000;
  assign literal_9083[29] = 16'h0000;
  assign literal_9083[30] = 16'h0000;
  assign literal_9083[31] = 16'h0000;
  assign literal_9083[32] = 16'h0000;
  assign literal_9083[33] = 16'h001b;
  assign literal_9083[34] = 16'h00f8;
  assign literal_9083[35] = 16'h03f7;
  assign literal_9083[36] = 16'h0ff4;
  assign literal_9083[37] = 16'h3fdc;
  assign literal_9083[38] = 16'hff9d;
  assign literal_9083[39] = 16'hff90;
  assign literal_9083[40] = 16'hffac;
  assign literal_9083[41] = 16'hffe3;
  assign literal_9083[42] = 16'hfff1;
  assign literal_9083[43] = 16'h0000;
  assign literal_9083[44] = 16'h0000;
  assign literal_9083[45] = 16'h0000;
  assign literal_9083[46] = 16'h0000;
  assign literal_9083[47] = 16'h0000;
  assign literal_9083[48] = 16'h0000;
  assign literal_9083[49] = 16'h003a;
  assign literal_9083[50] = 16'h01f6;
  assign literal_9083[51] = 16'h07f7;
  assign literal_9083[52] = 16'h3fde;
  assign literal_9083[53] = 16'hff8e;
  assign literal_9083[54] = 16'hff94;
  assign literal_9083[55] = 16'hffc9;
  assign literal_9083[56] = 16'hffd6;
  assign literal_9083[57] = 16'hffe4;
  assign literal_9083[58] = 16'hfff2;
  assign literal_9083[59] = 16'h0000;
  assign literal_9083[60] = 16'h0000;
  assign literal_9083[61] = 16'h0000;
  assign literal_9083[62] = 16'h0000;
  assign literal_9083[63] = 16'h0000;
  assign literal_9083[64] = 16'h0000;
  assign literal_9083[65] = 16'h003b;
  assign literal_9083[66] = 16'h03f6;
  assign literal_9083[67] = 16'h3fdd;
  assign literal_9083[68] = 16'hff8f;
  assign literal_9083[69] = 16'hffa5;
  assign literal_9083[70] = 16'hffa6;
  assign literal_9083[71] = 16'hffca;
  assign literal_9083[72] = 16'hffd7;
  assign literal_9083[73] = 16'hffe5;
  assign literal_9083[74] = 16'hfff3;
  assign literal_9083[75] = 16'h0000;
  assign literal_9083[76] = 16'h0000;
  assign literal_9083[77] = 16'h0000;
  assign literal_9083[78] = 16'h0000;
  assign literal_9083[79] = 16'h0000;
  assign literal_9083[80] = 16'h0000;
  assign literal_9083[81] = 16'h0078;
  assign literal_9083[82] = 16'h03f9;
  assign literal_9083[83] = 16'h3fdf;
  assign literal_9083[84] = 16'hff96;
  assign literal_9083[85] = 16'hffab;
  assign literal_9083[86] = 16'hffa9;
  assign literal_9083[87] = 16'hffcb;
  assign literal_9083[88] = 16'hffd8;
  assign literal_9083[89] = 16'hffe6;
  assign literal_9083[90] = 16'hfff4;
  assign literal_9083[91] = 16'h0000;
  assign literal_9083[92] = 16'h0000;
  assign literal_9083[93] = 16'h0000;
  assign literal_9083[94] = 16'h0000;
  assign literal_9083[95] = 16'h0000;
  assign literal_9083[96] = 16'h0000;
  assign literal_9083[97] = 16'h007b;
  assign literal_9083[98] = 16'h0ff2;
  assign literal_9083[99] = 16'h7fc5;
  assign literal_9083[100] = 16'hff97;
  assign literal_9083[101] = 16'hffb5;
  assign literal_9083[102] = 16'hffbf;
  assign literal_9083[103] = 16'hffcc;
  assign literal_9083[104] = 16'hffd9;
  assign literal_9083[105] = 16'hffe7;
  assign literal_9083[106] = 16'hfff5;
  assign literal_9083[107] = 16'h0000;
  assign literal_9083[108] = 16'h0000;
  assign literal_9083[109] = 16'h0000;
  assign literal_9083[110] = 16'h0000;
  assign literal_9083[111] = 16'h0000;
  assign literal_9083[112] = 16'h0000;
  assign literal_9083[113] = 16'h00f9;
  assign literal_9083[114] = 16'h0ff5;
  assign literal_9083[115] = 16'hff8c;
  assign literal_9083[116] = 16'hff98;
  assign literal_9083[117] = 16'hffb6;
  assign literal_9083[118] = 16'hffc0;
  assign literal_9083[119] = 16'hffcd;
  assign literal_9083[120] = 16'hffda;
  assign literal_9083[121] = 16'hffe8;
  assign literal_9083[122] = 16'hfff6;
  assign literal_9083[123] = 16'h0000;
  assign literal_9083[124] = 16'h0000;
  assign literal_9083[125] = 16'h0000;
  assign literal_9083[126] = 16'h0000;
  assign literal_9083[127] = 16'h0000;
  assign literal_9083[128] = 16'h0000;
  assign literal_9083[129] = 16'h01f4;
  assign literal_9083[130] = 16'h1fec;
  assign literal_9083[131] = 16'hff9e;
  assign literal_9083[132] = 16'hffa3;
  assign literal_9083[133] = 16'hffb7;
  assign literal_9083[134] = 16'hffc1;
  assign literal_9083[135] = 16'hffce;
  assign literal_9083[136] = 16'hffdb;
  assign literal_9083[137] = 16'hffe9;
  assign literal_9083[138] = 16'hfff7;
  assign literal_9083[139] = 16'h0000;
  assign literal_9083[140] = 16'h0000;
  assign literal_9083[141] = 16'h0000;
  assign literal_9083[142] = 16'h0000;
  assign literal_9083[143] = 16'h0000;
  assign literal_9083[144] = 16'h0000;
  assign literal_9083[145] = 16'h01f7;
  assign literal_9083[146] = 16'h3fe0;
  assign literal_9083[147] = 16'hff91;
  assign literal_9083[148] = 16'hffa4;
  assign literal_9083[149] = 16'hffb8;
  assign literal_9083[150] = 16'hffc2;
  assign literal_9083[151] = 16'hffcf;
  assign literal_9083[152] = 16'hffdc;
  assign literal_9083[153] = 16'hffea;
  assign literal_9083[154] = 16'hfff8;
  assign literal_9083[155] = 16'h0000;
  assign literal_9083[156] = 16'h0000;
  assign literal_9083[157] = 16'h0000;
  assign literal_9083[158] = 16'h0000;
  assign literal_9083[159] = 16'h0000;
  assign literal_9083[160] = 16'h0000;
  assign literal_9083[161] = 16'h01f8;
  assign literal_9083[162] = 16'h3fe1;
  assign literal_9083[163] = 16'hff92;
  assign literal_9083[164] = 16'hffa7;
  assign literal_9083[165] = 16'hffb9;
  assign literal_9083[166] = 16'hffc3;
  assign literal_9083[167] = 16'hffd0;
  assign literal_9083[168] = 16'hffdd;
  assign literal_9083[169] = 16'hffeb;
  assign literal_9083[170] = 16'hfff9;
  assign literal_9083[171] = 16'h0000;
  assign literal_9083[172] = 16'h0000;
  assign literal_9083[173] = 16'h0000;
  assign literal_9083[174] = 16'h0000;
  assign literal_9083[175] = 16'h0000;
  assign literal_9083[176] = 16'h0000;
  assign literal_9083[177] = 16'h03f5;
  assign literal_9083[178] = 16'h7fc4;
  assign literal_9083[179] = 16'hff93;
  assign literal_9083[180] = 16'hffa8;
  assign literal_9083[181] = 16'hffba;
  assign literal_9083[182] = 16'hffc4;
  assign literal_9083[183] = 16'hffd1;
  assign literal_9083[184] = 16'hffde;
  assign literal_9083[185] = 16'hffec;
  assign literal_9083[186] = 16'hfffa;
  assign literal_9083[187] = 16'h0000;
  assign literal_9083[188] = 16'h0000;
  assign literal_9083[189] = 16'h0000;
  assign literal_9083[190] = 16'h0000;
  assign literal_9083[191] = 16'h0000;
  assign literal_9083[192] = 16'h0000;
  assign literal_9083[193] = 16'h03f8;
  assign literal_9083[194] = 16'hff8d;
  assign literal_9083[195] = 16'hff99;
  assign literal_9083[196] = 16'hffb1;
  assign literal_9083[197] = 16'hffbb;
  assign literal_9083[198] = 16'hffc5;
  assign literal_9083[199] = 16'hffd2;
  assign literal_9083[200] = 16'hffdf;
  assign literal_9083[201] = 16'hffed;
  assign literal_9083[202] = 16'hfffb;
  assign literal_9083[203] = 16'h0000;
  assign literal_9083[204] = 16'h0000;
  assign literal_9083[205] = 16'h0000;
  assign literal_9083[206] = 16'h0000;
  assign literal_9083[207] = 16'h0000;
  assign literal_9083[208] = 16'h0000;
  assign literal_9083[209] = 16'h03fa;
  assign literal_9083[210] = 16'hff9a;
  assign literal_9083[211] = 16'hffaa;
  assign literal_9083[212] = 16'hffb2;
  assign literal_9083[213] = 16'hffbc;
  assign literal_9083[214] = 16'hffc6;
  assign literal_9083[215] = 16'hffd3;
  assign literal_9083[216] = 16'hffe0;
  assign literal_9083[217] = 16'hffee;
  assign literal_9083[218] = 16'hfffc;
  assign literal_9083[219] = 16'h0000;
  assign literal_9083[220] = 16'h0000;
  assign literal_9083[221] = 16'h0000;
  assign literal_9083[222] = 16'h0000;
  assign literal_9083[223] = 16'h0000;
  assign literal_9083[224] = 16'h0000;
  assign literal_9083[225] = 16'h07f6;
  assign literal_9083[226] = 16'hff9b;
  assign literal_9083[227] = 16'hffaf;
  assign literal_9083[228] = 16'hffb3;
  assign literal_9083[229] = 16'hffbd;
  assign literal_9083[230] = 16'hffc7;
  assign literal_9083[231] = 16'hffd4;
  assign literal_9083[232] = 16'hffe1;
  assign literal_9083[233] = 16'hffef;
  assign literal_9083[234] = 16'hfffd;
  assign literal_9083[235] = 16'h0000;
  assign literal_9083[236] = 16'h0000;
  assign literal_9083[237] = 16'h0000;
  assign literal_9083[238] = 16'h0000;
  assign literal_9083[239] = 16'h0000;
  assign literal_9083[240] = 16'h0ff3;
  assign literal_9083[241] = 16'h1fed;
  assign literal_9083[242] = 16'hffae;
  assign literal_9083[243] = 16'hffb0;
  assign literal_9083[244] = 16'hffb4;
  assign literal_9083[245] = 16'hffbe;
  assign literal_9083[246] = 16'hffc8;
  assign literal_9083[247] = 16'hffd5;
  assign literal_9083[248] = 16'hffe2;
  assign literal_9083[249] = 16'hfff0;
  assign literal_9083[250] = 16'hfffe;
  assign literal_9083[251] = 16'h0000;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [9:0] p1_row0_comb[0:7];
  wire [9:0] p1_row1_comb[0:7];
  wire [9:0] p1_array_concat_8141_comb[0:15];
  wire [9:0] p1_row2_comb[0:7];
  wire [9:0] p1_array_concat_8144_comb[0:23];
  wire [9:0] p1_row3_comb[0:7];
  wire [2:0] p1_idx_u8__4_squeezed_comb;
  wire [9:0] p1_array_concat_8147_comb[0:31];
  wire [9:0] p1_row4_comb[0:7];
  wire [2:0] p1_idx_u8__5_squeezed_comb;
  wire [9:0] p1_array_concat_8150_comb[0:39];
  wire [9:0] p1_row5_comb[0:7];
  wire [2:0] p1_idx_u8__6_squeezed_comb;
  wire [7:0] p1_idx_u8__1_comb;
  wire [7:0] p1_idx_u8__3_comb;
  wire [7:0] p1_idx_u8__5_comb;
  wire [7:0] p1_idx_u8__7_comb;
  wire [7:0] p1_idx_u8__9_comb;
  wire [7:0] p1_idx_u8__11_comb;
  wire [7:0] p1_idx_u8__13_comb;
  wire [9:0] p1_array_concat_8156_comb[0:47];
  wire [9:0] p1_row6_comb[0:7];
  wire [2:0] p1_idx_u8__7_squeezed_comb;
  wire [6:0] p1_add_8159_comb;
  wire [7:0] p1_actual_index__1_comb;
  wire [6:0] p1_add_8274_comb;
  wire [7:0] p1_actual_index__3_comb;
  wire [5:0] p1_add_8257_comb;
  wire [7:0] p1_actual_index__5_comb;
  wire [6:0] p1_add_8241_comb;
  wire [7:0] p1_actual_index__7_comb;
  wire [7:0] p1_actual_index__9_comb;
  wire [6:0] p1_add_8192_comb;
  wire [7:0] p1_actual_index__11_comb;
  wire [7:0] p1_actual_index__13_comb;
  wire [7:0] p1_idx_u8__15_comb;
  wire [7:0] p1_idx_u8__17_comb;
  wire [7:0] p1_idx_u8__19_comb;
  wire [7:0] p1_idx_u8__21_comb;
  wire [7:0] p1_idx_u8__23_comb;
  wire [7:0] p1_idx_u8__25_comb;
  wire [7:0] p1_idx_u8__27_comb;
  wire [7:0] p1_idx_u8__29_comb;
  wire [7:0] p1_idx_u8__31_comb;
  wire [7:0] p1_idx_u8__33_comb;
  wire [7:0] p1_idx_u8__35_comb;
  wire [7:0] p1_idx_u8__37_comb;
  wire [7:0] p1_idx_u8__39_comb;
  wire [7:0] p1_idx_u8__41_comb;
  wire [7:0] p1_idx_u8__43_comb;
  wire [7:0] p1_idx_u8__45_comb;
  wire [7:0] p1_idx_u8__47_comb;
  wire [7:0] p1_idx_u8__49_comb;
  wire [7:0] p1_idx_u8__51_comb;
  wire [7:0] p1_idx_u8__53_comb;
  wire [7:0] p1_idx_u8__55_comb;
  wire [7:0] p1_idx_u8__57_comb;
  wire [7:0] p1_idx_u8__59_comb;
  wire [7:0] p1_idx_u8__61_comb;
  wire [9:0] p1_array_concat_8163_comb[0:55];
  wire [9:0] p1_row7_comb[0:7];
  wire [5:0] p1_add_8168_comb;
  wire [4:0] p1_add_8211_comb;
  wire [7:0] p1_actual_index__15_comb;
  wire [3:0] p1_add_8377_comb;
  wire [7:0] p1_actual_index__17_comb;
  wire [6:0] p1_add_8379_comb;
  wire [7:0] p1_actual_index__19_comb;
  wire [5:0] p1_add_8381_comb;
  wire [7:0] p1_actual_index__21_comb;
  wire [6:0] p1_add_8383_comb;
  wire [7:0] p1_actual_index__23_comb;
  wire [4:0] p1_add_8385_comb;
  wire [7:0] p1_actual_index__25_comb;
  wire [6:0] p1_add_8387_comb;
  wire [7:0] p1_actual_index__27_comb;
  wire [5:0] p1_add_8389_comb;
  wire [7:0] p1_actual_index__29_comb;
  wire [6:0] p1_add_8391_comb;
  wire [7:0] p1_actual_index__31_comb;
  wire [2:0] p1_add_8393_comb;
  wire [7:0] p1_actual_index__33_comb;
  wire [6:0] p1_add_8395_comb;
  wire [7:0] p1_actual_index__35_comb;
  wire [5:0] p1_add_8397_comb;
  wire [7:0] p1_actual_index__37_comb;
  wire [6:0] p1_add_8399_comb;
  wire [7:0] p1_actual_index__39_comb;
  wire [4:0] p1_add_8401_comb;
  wire [7:0] p1_actual_index__41_comb;
  wire [6:0] p1_add_8403_comb;
  wire [7:0] p1_actual_index__43_comb;
  wire [5:0] p1_add_8405_comb;
  wire [7:0] p1_actual_index__45_comb;
  wire [6:0] p1_add_8407_comb;
  wire [7:0] p1_actual_index__47_comb;
  wire [3:0] p1_add_8409_comb;
  wire [7:0] p1_actual_index__49_comb;
  wire [6:0] p1_add_8411_comb;
  wire [7:0] p1_actual_index__51_comb;
  wire [5:0] p1_add_8413_comb;
  wire [7:0] p1_actual_index__53_comb;
  wire [6:0] p1_add_8415_comb;
  wire [7:0] p1_actual_index__55_comb;
  wire [4:0] p1_add_8417_comb;
  wire [7:0] p1_actual_index__57_comb;
  wire [6:0] p1_add_8419_comb;
  wire [7:0] p1_actual_index__59_comb;
  wire [5:0] p1_add_8421_comb;
  wire [7:0] p1_actual_index__61_comb;
  wire [6:0] p1_add_8423_comb;
  wire [9:0] p1_flat_comb[0:63];
  wire [7:0] p1_actual_index__14_comb;
  wire [7:0] p1_actual_index__2_comb;
  wire [7:0] p1_actual_index__4_comb;
  wire [7:0] p1_actual_index__6_comb;
  wire [7:0] p1_actual_index__10_comb;
  wire [7:0] p1_actual_index__12_comb;
  wire [7:0] p1_actual_index__8_comb;
  wire [7:0] p1_actual_index__16_comb;
  wire [7:0] p1_actual_index__18_comb;
  wire [7:0] p1_actual_index__20_comb;
  wire [7:0] p1_actual_index__22_comb;
  wire [7:0] p1_actual_index__24_comb;
  wire [7:0] p1_actual_index__26_comb;
  wire [7:0] p1_actual_index__28_comb;
  wire [7:0] p1_actual_index__30_comb;
  wire [7:0] p1_actual_index__32_comb;
  wire [7:0] p1_actual_index__34_comb;
  wire [7:0] p1_actual_index__36_comb;
  wire [7:0] p1_actual_index__38_comb;
  wire [7:0] p1_actual_index__40_comb;
  wire [7:0] p1_actual_index__42_comb;
  wire [7:0] p1_actual_index__44_comb;
  wire [7:0] p1_actual_index__46_comb;
  wire [7:0] p1_actual_index__48_comb;
  wire [7:0] p1_actual_index__50_comb;
  wire [7:0] p1_actual_index__52_comb;
  wire [7:0] p1_actual_index__54_comb;
  wire [7:0] p1_actual_index__56_comb;
  wire [7:0] p1_actual_index__58_comb;
  wire [7:0] p1_actual_index__60_comb;
  wire [7:0] p1_actual_index__62_comb;
  wire [9:0] p1_value_comb;
  wire [9:0] p1_and_8187_comb;
  wire [9:0] p1_and_8318_comb;
  wire [9:0] p1_and_8320_comb;
  wire [9:0] p1_and_8315_comb;
  wire [9:0] p1_and_8308_comb;
  wire [9:0] p1_and_8301_comb;
  wire [9:0] p1_and_8290_comb;
  wire [9:0] p1_and_8281_comb;
  wire [9:0] p1_and_8271_comb;
  wire [9:0] p1_and_8244_comb;
  wire [9:0] p1_and_8235_comb;
  wire [9:0] p1_and_8227_comb;
  wire [9:0] p1_and_8195_comb;
  wire [7:0] p1_bin_value_comb;
  wire p1_eq_8198_comb;
  wire [9:0] p1_and_8199_comb;
  wire p1_ne_8323_comb;
  wire p1_ne_8324_comb;
  wire p1_ne_8322_comb;
  wire p1_ne_8317_comb;
  wire p1_ne_8310_comb;
  wire p1_ne_8303_comb;
  wire p1_ne_8292_comb;
  wire p1_ne_8283_comb;
  wire [9:0] p1_and_8247_comb;
  wire p1_ne_8254_comb;
  wire p1_ne_8246_comb;
  wire p1_ne_8237_comb;
  wire p1_ne_8207_comb;
  wire [7:0] p1_flipped_comb;
  wire [1:0] p1_idx_u8__1_squeezed_comb;
  wire p1_eq_8210_comb;
  wire p1_not_8325_comb;
  wire p1_eq_8255_comb;
  wire [1:0] p1_sel_8218_comb;
  wire [1:0] p1_sign_ext_8219_comb;
  wire p1_and_8848_comb;
  wire [7:0] p1_code_list_comb;
  assign p1_row0_comb[0] = p0_matrix[3'h0][0];
  assign p1_row0_comb[1] = p0_matrix[3'h0][1];
  assign p1_row0_comb[2] = p0_matrix[3'h0][2];
  assign p1_row0_comb[3] = p0_matrix[3'h0][3];
  assign p1_row0_comb[4] = p0_matrix[3'h0][4];
  assign p1_row0_comb[5] = p0_matrix[3'h0][5];
  assign p1_row0_comb[6] = p0_matrix[3'h0][6];
  assign p1_row0_comb[7] = p0_matrix[3'h0][7];
  assign p1_row1_comb[0] = p0_matrix[3'h1][0];
  assign p1_row1_comb[1] = p0_matrix[3'h1][1];
  assign p1_row1_comb[2] = p0_matrix[3'h1][2];
  assign p1_row1_comb[3] = p0_matrix[3'h1][3];
  assign p1_row1_comb[4] = p0_matrix[3'h1][4];
  assign p1_row1_comb[5] = p0_matrix[3'h1][5];
  assign p1_row1_comb[6] = p0_matrix[3'h1][6];
  assign p1_row1_comb[7] = p0_matrix[3'h1][7];
  assign p1_array_concat_8141_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_8141_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_8141_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_8141_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_8141_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_8141_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_8141_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_8141_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_8141_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_8141_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_8141_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_8141_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_8141_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_8141_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_8141_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_8141_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_8144_comb[0] = p1_array_concat_8141_comb[0];
  assign p1_array_concat_8144_comb[1] = p1_array_concat_8141_comb[1];
  assign p1_array_concat_8144_comb[2] = p1_array_concat_8141_comb[2];
  assign p1_array_concat_8144_comb[3] = p1_array_concat_8141_comb[3];
  assign p1_array_concat_8144_comb[4] = p1_array_concat_8141_comb[4];
  assign p1_array_concat_8144_comb[5] = p1_array_concat_8141_comb[5];
  assign p1_array_concat_8144_comb[6] = p1_array_concat_8141_comb[6];
  assign p1_array_concat_8144_comb[7] = p1_array_concat_8141_comb[7];
  assign p1_array_concat_8144_comb[8] = p1_array_concat_8141_comb[8];
  assign p1_array_concat_8144_comb[9] = p1_array_concat_8141_comb[9];
  assign p1_array_concat_8144_comb[10] = p1_array_concat_8141_comb[10];
  assign p1_array_concat_8144_comb[11] = p1_array_concat_8141_comb[11];
  assign p1_array_concat_8144_comb[12] = p1_array_concat_8141_comb[12];
  assign p1_array_concat_8144_comb[13] = p1_array_concat_8141_comb[13];
  assign p1_array_concat_8144_comb[14] = p1_array_concat_8141_comb[14];
  assign p1_array_concat_8144_comb[15] = p1_array_concat_8141_comb[15];
  assign p1_array_concat_8144_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_8144_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_8144_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_8144_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_8144_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_8144_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_8144_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_8144_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_idx_u8__4_squeezed_comb = 3'h4;
  assign p1_array_concat_8147_comb[0] = p1_array_concat_8144_comb[0];
  assign p1_array_concat_8147_comb[1] = p1_array_concat_8144_comb[1];
  assign p1_array_concat_8147_comb[2] = p1_array_concat_8144_comb[2];
  assign p1_array_concat_8147_comb[3] = p1_array_concat_8144_comb[3];
  assign p1_array_concat_8147_comb[4] = p1_array_concat_8144_comb[4];
  assign p1_array_concat_8147_comb[5] = p1_array_concat_8144_comb[5];
  assign p1_array_concat_8147_comb[6] = p1_array_concat_8144_comb[6];
  assign p1_array_concat_8147_comb[7] = p1_array_concat_8144_comb[7];
  assign p1_array_concat_8147_comb[8] = p1_array_concat_8144_comb[8];
  assign p1_array_concat_8147_comb[9] = p1_array_concat_8144_comb[9];
  assign p1_array_concat_8147_comb[10] = p1_array_concat_8144_comb[10];
  assign p1_array_concat_8147_comb[11] = p1_array_concat_8144_comb[11];
  assign p1_array_concat_8147_comb[12] = p1_array_concat_8144_comb[12];
  assign p1_array_concat_8147_comb[13] = p1_array_concat_8144_comb[13];
  assign p1_array_concat_8147_comb[14] = p1_array_concat_8144_comb[14];
  assign p1_array_concat_8147_comb[15] = p1_array_concat_8144_comb[15];
  assign p1_array_concat_8147_comb[16] = p1_array_concat_8144_comb[16];
  assign p1_array_concat_8147_comb[17] = p1_array_concat_8144_comb[17];
  assign p1_array_concat_8147_comb[18] = p1_array_concat_8144_comb[18];
  assign p1_array_concat_8147_comb[19] = p1_array_concat_8144_comb[19];
  assign p1_array_concat_8147_comb[20] = p1_array_concat_8144_comb[20];
  assign p1_array_concat_8147_comb[21] = p1_array_concat_8144_comb[21];
  assign p1_array_concat_8147_comb[22] = p1_array_concat_8144_comb[22];
  assign p1_array_concat_8147_comb[23] = p1_array_concat_8144_comb[23];
  assign p1_array_concat_8147_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_8147_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_8147_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_8147_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_8147_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_8147_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_8147_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_8147_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[p1_idx_u8__4_squeezed_comb][0];
  assign p1_row4_comb[1] = p0_matrix[p1_idx_u8__4_squeezed_comb][1];
  assign p1_row4_comb[2] = p0_matrix[p1_idx_u8__4_squeezed_comb][2];
  assign p1_row4_comb[3] = p0_matrix[p1_idx_u8__4_squeezed_comb][3];
  assign p1_row4_comb[4] = p0_matrix[p1_idx_u8__4_squeezed_comb][4];
  assign p1_row4_comb[5] = p0_matrix[p1_idx_u8__4_squeezed_comb][5];
  assign p1_row4_comb[6] = p0_matrix[p1_idx_u8__4_squeezed_comb][6];
  assign p1_row4_comb[7] = p0_matrix[p1_idx_u8__4_squeezed_comb][7];
  assign p1_idx_u8__5_squeezed_comb = 3'h5;
  assign p1_array_concat_8150_comb[0] = p1_array_concat_8147_comb[0];
  assign p1_array_concat_8150_comb[1] = p1_array_concat_8147_comb[1];
  assign p1_array_concat_8150_comb[2] = p1_array_concat_8147_comb[2];
  assign p1_array_concat_8150_comb[3] = p1_array_concat_8147_comb[3];
  assign p1_array_concat_8150_comb[4] = p1_array_concat_8147_comb[4];
  assign p1_array_concat_8150_comb[5] = p1_array_concat_8147_comb[5];
  assign p1_array_concat_8150_comb[6] = p1_array_concat_8147_comb[6];
  assign p1_array_concat_8150_comb[7] = p1_array_concat_8147_comb[7];
  assign p1_array_concat_8150_comb[8] = p1_array_concat_8147_comb[8];
  assign p1_array_concat_8150_comb[9] = p1_array_concat_8147_comb[9];
  assign p1_array_concat_8150_comb[10] = p1_array_concat_8147_comb[10];
  assign p1_array_concat_8150_comb[11] = p1_array_concat_8147_comb[11];
  assign p1_array_concat_8150_comb[12] = p1_array_concat_8147_comb[12];
  assign p1_array_concat_8150_comb[13] = p1_array_concat_8147_comb[13];
  assign p1_array_concat_8150_comb[14] = p1_array_concat_8147_comb[14];
  assign p1_array_concat_8150_comb[15] = p1_array_concat_8147_comb[15];
  assign p1_array_concat_8150_comb[16] = p1_array_concat_8147_comb[16];
  assign p1_array_concat_8150_comb[17] = p1_array_concat_8147_comb[17];
  assign p1_array_concat_8150_comb[18] = p1_array_concat_8147_comb[18];
  assign p1_array_concat_8150_comb[19] = p1_array_concat_8147_comb[19];
  assign p1_array_concat_8150_comb[20] = p1_array_concat_8147_comb[20];
  assign p1_array_concat_8150_comb[21] = p1_array_concat_8147_comb[21];
  assign p1_array_concat_8150_comb[22] = p1_array_concat_8147_comb[22];
  assign p1_array_concat_8150_comb[23] = p1_array_concat_8147_comb[23];
  assign p1_array_concat_8150_comb[24] = p1_array_concat_8147_comb[24];
  assign p1_array_concat_8150_comb[25] = p1_array_concat_8147_comb[25];
  assign p1_array_concat_8150_comb[26] = p1_array_concat_8147_comb[26];
  assign p1_array_concat_8150_comb[27] = p1_array_concat_8147_comb[27];
  assign p1_array_concat_8150_comb[28] = p1_array_concat_8147_comb[28];
  assign p1_array_concat_8150_comb[29] = p1_array_concat_8147_comb[29];
  assign p1_array_concat_8150_comb[30] = p1_array_concat_8147_comb[30];
  assign p1_array_concat_8150_comb[31] = p1_array_concat_8147_comb[31];
  assign p1_array_concat_8150_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_8150_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_8150_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_8150_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_8150_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_8150_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_8150_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_8150_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[p1_idx_u8__5_squeezed_comb][0];
  assign p1_row5_comb[1] = p0_matrix[p1_idx_u8__5_squeezed_comb][1];
  assign p1_row5_comb[2] = p0_matrix[p1_idx_u8__5_squeezed_comb][2];
  assign p1_row5_comb[3] = p0_matrix[p1_idx_u8__5_squeezed_comb][3];
  assign p1_row5_comb[4] = p0_matrix[p1_idx_u8__5_squeezed_comb][4];
  assign p1_row5_comb[5] = p0_matrix[p1_idx_u8__5_squeezed_comb][5];
  assign p1_row5_comb[6] = p0_matrix[p1_idx_u8__5_squeezed_comb][6];
  assign p1_row5_comb[7] = p0_matrix[p1_idx_u8__5_squeezed_comb][7];
  assign p1_idx_u8__6_squeezed_comb = 3'h6;
  assign p1_idx_u8__1_comb = 8'h01;
  assign p1_idx_u8__3_comb = 8'h03;
  assign p1_idx_u8__5_comb = 8'h05;
  assign p1_idx_u8__7_comb = 8'h07;
  assign p1_idx_u8__9_comb = 8'h09;
  assign p1_idx_u8__11_comb = 8'h0b;
  assign p1_idx_u8__13_comb = 8'h0d;
  assign p1_array_concat_8156_comb[0] = p1_array_concat_8150_comb[0];
  assign p1_array_concat_8156_comb[1] = p1_array_concat_8150_comb[1];
  assign p1_array_concat_8156_comb[2] = p1_array_concat_8150_comb[2];
  assign p1_array_concat_8156_comb[3] = p1_array_concat_8150_comb[3];
  assign p1_array_concat_8156_comb[4] = p1_array_concat_8150_comb[4];
  assign p1_array_concat_8156_comb[5] = p1_array_concat_8150_comb[5];
  assign p1_array_concat_8156_comb[6] = p1_array_concat_8150_comb[6];
  assign p1_array_concat_8156_comb[7] = p1_array_concat_8150_comb[7];
  assign p1_array_concat_8156_comb[8] = p1_array_concat_8150_comb[8];
  assign p1_array_concat_8156_comb[9] = p1_array_concat_8150_comb[9];
  assign p1_array_concat_8156_comb[10] = p1_array_concat_8150_comb[10];
  assign p1_array_concat_8156_comb[11] = p1_array_concat_8150_comb[11];
  assign p1_array_concat_8156_comb[12] = p1_array_concat_8150_comb[12];
  assign p1_array_concat_8156_comb[13] = p1_array_concat_8150_comb[13];
  assign p1_array_concat_8156_comb[14] = p1_array_concat_8150_comb[14];
  assign p1_array_concat_8156_comb[15] = p1_array_concat_8150_comb[15];
  assign p1_array_concat_8156_comb[16] = p1_array_concat_8150_comb[16];
  assign p1_array_concat_8156_comb[17] = p1_array_concat_8150_comb[17];
  assign p1_array_concat_8156_comb[18] = p1_array_concat_8150_comb[18];
  assign p1_array_concat_8156_comb[19] = p1_array_concat_8150_comb[19];
  assign p1_array_concat_8156_comb[20] = p1_array_concat_8150_comb[20];
  assign p1_array_concat_8156_comb[21] = p1_array_concat_8150_comb[21];
  assign p1_array_concat_8156_comb[22] = p1_array_concat_8150_comb[22];
  assign p1_array_concat_8156_comb[23] = p1_array_concat_8150_comb[23];
  assign p1_array_concat_8156_comb[24] = p1_array_concat_8150_comb[24];
  assign p1_array_concat_8156_comb[25] = p1_array_concat_8150_comb[25];
  assign p1_array_concat_8156_comb[26] = p1_array_concat_8150_comb[26];
  assign p1_array_concat_8156_comb[27] = p1_array_concat_8150_comb[27];
  assign p1_array_concat_8156_comb[28] = p1_array_concat_8150_comb[28];
  assign p1_array_concat_8156_comb[29] = p1_array_concat_8150_comb[29];
  assign p1_array_concat_8156_comb[30] = p1_array_concat_8150_comb[30];
  assign p1_array_concat_8156_comb[31] = p1_array_concat_8150_comb[31];
  assign p1_array_concat_8156_comb[32] = p1_array_concat_8150_comb[32];
  assign p1_array_concat_8156_comb[33] = p1_array_concat_8150_comb[33];
  assign p1_array_concat_8156_comb[34] = p1_array_concat_8150_comb[34];
  assign p1_array_concat_8156_comb[35] = p1_array_concat_8150_comb[35];
  assign p1_array_concat_8156_comb[36] = p1_array_concat_8150_comb[36];
  assign p1_array_concat_8156_comb[37] = p1_array_concat_8150_comb[37];
  assign p1_array_concat_8156_comb[38] = p1_array_concat_8150_comb[38];
  assign p1_array_concat_8156_comb[39] = p1_array_concat_8150_comb[39];
  assign p1_array_concat_8156_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_8156_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_8156_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_8156_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_8156_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_8156_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_8156_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_8156_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[p1_idx_u8__6_squeezed_comb][0];
  assign p1_row6_comb[1] = p0_matrix[p1_idx_u8__6_squeezed_comb][1];
  assign p1_row6_comb[2] = p0_matrix[p1_idx_u8__6_squeezed_comb][2];
  assign p1_row6_comb[3] = p0_matrix[p1_idx_u8__6_squeezed_comb][3];
  assign p1_row6_comb[4] = p0_matrix[p1_idx_u8__6_squeezed_comb][4];
  assign p1_row6_comb[5] = p0_matrix[p1_idx_u8__6_squeezed_comb][5];
  assign p1_row6_comb[6] = p0_matrix[p1_idx_u8__6_squeezed_comb][6];
  assign p1_row6_comb[7] = p0_matrix[p1_idx_u8__6_squeezed_comb][7];
  assign p1_idx_u8__7_squeezed_comb = 3'h7;
  assign p1_add_8159_comb = p0_start_pix[7:1] + 7'h07;
  assign p1_actual_index__1_comb = p0_start_pix + p1_idx_u8__1_comb;
  assign p1_add_8274_comb = p0_start_pix[7:1] + 7'h01;
  assign p1_actual_index__3_comb = p0_start_pix + p1_idx_u8__3_comb;
  assign p1_add_8257_comb = p0_start_pix[7:2] + 6'h01;
  assign p1_actual_index__5_comb = p0_start_pix + p1_idx_u8__5_comb;
  assign p1_add_8241_comb = p0_start_pix[7:1] + 7'h03;
  assign p1_actual_index__7_comb = p0_start_pix + p1_idx_u8__7_comb;
  assign p1_actual_index__9_comb = p0_start_pix + p1_idx_u8__9_comb;
  assign p1_add_8192_comb = p0_start_pix[7:1] + 7'h05;
  assign p1_actual_index__11_comb = p0_start_pix + p1_idx_u8__11_comb;
  assign p1_actual_index__13_comb = p0_start_pix + p1_idx_u8__13_comb;
  assign p1_idx_u8__15_comb = 8'h0f;
  assign p1_idx_u8__17_comb = 8'h11;
  assign p1_idx_u8__19_comb = 8'h13;
  assign p1_idx_u8__21_comb = 8'h15;
  assign p1_idx_u8__23_comb = 8'h17;
  assign p1_idx_u8__25_comb = 8'h19;
  assign p1_idx_u8__27_comb = 8'h1b;
  assign p1_idx_u8__29_comb = 8'h1d;
  assign p1_idx_u8__31_comb = 8'h1f;
  assign p1_idx_u8__33_comb = 8'h21;
  assign p1_idx_u8__35_comb = 8'h23;
  assign p1_idx_u8__37_comb = 8'h25;
  assign p1_idx_u8__39_comb = 8'h27;
  assign p1_idx_u8__41_comb = 8'h29;
  assign p1_idx_u8__43_comb = 8'h2b;
  assign p1_idx_u8__45_comb = 8'h2d;
  assign p1_idx_u8__47_comb = 8'h2f;
  assign p1_idx_u8__49_comb = 8'h31;
  assign p1_idx_u8__51_comb = 8'h33;
  assign p1_idx_u8__53_comb = 8'h35;
  assign p1_idx_u8__55_comb = 8'h37;
  assign p1_idx_u8__57_comb = 8'h39;
  assign p1_idx_u8__59_comb = 8'h3b;
  assign p1_idx_u8__61_comb = 8'h3d;
  assign p1_array_concat_8163_comb[0] = p1_array_concat_8156_comb[0];
  assign p1_array_concat_8163_comb[1] = p1_array_concat_8156_comb[1];
  assign p1_array_concat_8163_comb[2] = p1_array_concat_8156_comb[2];
  assign p1_array_concat_8163_comb[3] = p1_array_concat_8156_comb[3];
  assign p1_array_concat_8163_comb[4] = p1_array_concat_8156_comb[4];
  assign p1_array_concat_8163_comb[5] = p1_array_concat_8156_comb[5];
  assign p1_array_concat_8163_comb[6] = p1_array_concat_8156_comb[6];
  assign p1_array_concat_8163_comb[7] = p1_array_concat_8156_comb[7];
  assign p1_array_concat_8163_comb[8] = p1_array_concat_8156_comb[8];
  assign p1_array_concat_8163_comb[9] = p1_array_concat_8156_comb[9];
  assign p1_array_concat_8163_comb[10] = p1_array_concat_8156_comb[10];
  assign p1_array_concat_8163_comb[11] = p1_array_concat_8156_comb[11];
  assign p1_array_concat_8163_comb[12] = p1_array_concat_8156_comb[12];
  assign p1_array_concat_8163_comb[13] = p1_array_concat_8156_comb[13];
  assign p1_array_concat_8163_comb[14] = p1_array_concat_8156_comb[14];
  assign p1_array_concat_8163_comb[15] = p1_array_concat_8156_comb[15];
  assign p1_array_concat_8163_comb[16] = p1_array_concat_8156_comb[16];
  assign p1_array_concat_8163_comb[17] = p1_array_concat_8156_comb[17];
  assign p1_array_concat_8163_comb[18] = p1_array_concat_8156_comb[18];
  assign p1_array_concat_8163_comb[19] = p1_array_concat_8156_comb[19];
  assign p1_array_concat_8163_comb[20] = p1_array_concat_8156_comb[20];
  assign p1_array_concat_8163_comb[21] = p1_array_concat_8156_comb[21];
  assign p1_array_concat_8163_comb[22] = p1_array_concat_8156_comb[22];
  assign p1_array_concat_8163_comb[23] = p1_array_concat_8156_comb[23];
  assign p1_array_concat_8163_comb[24] = p1_array_concat_8156_comb[24];
  assign p1_array_concat_8163_comb[25] = p1_array_concat_8156_comb[25];
  assign p1_array_concat_8163_comb[26] = p1_array_concat_8156_comb[26];
  assign p1_array_concat_8163_comb[27] = p1_array_concat_8156_comb[27];
  assign p1_array_concat_8163_comb[28] = p1_array_concat_8156_comb[28];
  assign p1_array_concat_8163_comb[29] = p1_array_concat_8156_comb[29];
  assign p1_array_concat_8163_comb[30] = p1_array_concat_8156_comb[30];
  assign p1_array_concat_8163_comb[31] = p1_array_concat_8156_comb[31];
  assign p1_array_concat_8163_comb[32] = p1_array_concat_8156_comb[32];
  assign p1_array_concat_8163_comb[33] = p1_array_concat_8156_comb[33];
  assign p1_array_concat_8163_comb[34] = p1_array_concat_8156_comb[34];
  assign p1_array_concat_8163_comb[35] = p1_array_concat_8156_comb[35];
  assign p1_array_concat_8163_comb[36] = p1_array_concat_8156_comb[36];
  assign p1_array_concat_8163_comb[37] = p1_array_concat_8156_comb[37];
  assign p1_array_concat_8163_comb[38] = p1_array_concat_8156_comb[38];
  assign p1_array_concat_8163_comb[39] = p1_array_concat_8156_comb[39];
  assign p1_array_concat_8163_comb[40] = p1_array_concat_8156_comb[40];
  assign p1_array_concat_8163_comb[41] = p1_array_concat_8156_comb[41];
  assign p1_array_concat_8163_comb[42] = p1_array_concat_8156_comb[42];
  assign p1_array_concat_8163_comb[43] = p1_array_concat_8156_comb[43];
  assign p1_array_concat_8163_comb[44] = p1_array_concat_8156_comb[44];
  assign p1_array_concat_8163_comb[45] = p1_array_concat_8156_comb[45];
  assign p1_array_concat_8163_comb[46] = p1_array_concat_8156_comb[46];
  assign p1_array_concat_8163_comb[47] = p1_array_concat_8156_comb[47];
  assign p1_array_concat_8163_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_8163_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_8163_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_8163_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_8163_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_8163_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_8163_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_8163_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[p1_idx_u8__7_squeezed_comb][0];
  assign p1_row7_comb[1] = p0_matrix[p1_idx_u8__7_squeezed_comb][1];
  assign p1_row7_comb[2] = p0_matrix[p1_idx_u8__7_squeezed_comb][2];
  assign p1_row7_comb[3] = p0_matrix[p1_idx_u8__7_squeezed_comb][3];
  assign p1_row7_comb[4] = p0_matrix[p1_idx_u8__7_squeezed_comb][4];
  assign p1_row7_comb[5] = p0_matrix[p1_idx_u8__7_squeezed_comb][5];
  assign p1_row7_comb[6] = p0_matrix[p1_idx_u8__7_squeezed_comb][6];
  assign p1_row7_comb[7] = p0_matrix[p1_idx_u8__7_squeezed_comb][7];
  assign p1_add_8168_comb = p0_start_pix[7:2] + 6'h03;
  assign p1_add_8211_comb = p0_start_pix[7:3] + 5'h01;
  assign p1_actual_index__15_comb = p0_start_pix + p1_idx_u8__15_comb;
  assign p1_add_8377_comb = p0_start_pix[7:4] + 4'h1;
  assign p1_actual_index__17_comb = p0_start_pix + p1_idx_u8__17_comb;
  assign p1_add_8379_comb = p0_start_pix[7:1] + 7'h09;
  assign p1_actual_index__19_comb = p0_start_pix + p1_idx_u8__19_comb;
  assign p1_add_8381_comb = p0_start_pix[7:2] + 6'h05;
  assign p1_actual_index__21_comb = p0_start_pix + p1_idx_u8__21_comb;
  assign p1_add_8383_comb = p0_start_pix[7:1] + 7'h0b;
  assign p1_actual_index__23_comb = p0_start_pix + p1_idx_u8__23_comb;
  assign p1_add_8385_comb = p0_start_pix[7:3] + 5'h03;
  assign p1_actual_index__25_comb = p0_start_pix + p1_idx_u8__25_comb;
  assign p1_add_8387_comb = p0_start_pix[7:1] + 7'h0d;
  assign p1_actual_index__27_comb = p0_start_pix + p1_idx_u8__27_comb;
  assign p1_add_8389_comb = p0_start_pix[7:2] + 6'h07;
  assign p1_actual_index__29_comb = p0_start_pix + p1_idx_u8__29_comb;
  assign p1_add_8391_comb = p0_start_pix[7:1] + 7'h0f;
  assign p1_actual_index__31_comb = p0_start_pix + p1_idx_u8__31_comb;
  assign p1_add_8393_comb = p0_start_pix[7:5] + 3'h1;
  assign p1_actual_index__33_comb = p0_start_pix + p1_idx_u8__33_comb;
  assign p1_add_8395_comb = p0_start_pix[7:1] + 7'h11;
  assign p1_actual_index__35_comb = p0_start_pix + p1_idx_u8__35_comb;
  assign p1_add_8397_comb = p0_start_pix[7:2] + 6'h09;
  assign p1_actual_index__37_comb = p0_start_pix + p1_idx_u8__37_comb;
  assign p1_add_8399_comb = p0_start_pix[7:1] + 7'h13;
  assign p1_actual_index__39_comb = p0_start_pix + p1_idx_u8__39_comb;
  assign p1_add_8401_comb = p0_start_pix[7:3] + 5'h05;
  assign p1_actual_index__41_comb = p0_start_pix + p1_idx_u8__41_comb;
  assign p1_add_8403_comb = p0_start_pix[7:1] + 7'h15;
  assign p1_actual_index__43_comb = p0_start_pix + p1_idx_u8__43_comb;
  assign p1_add_8405_comb = p0_start_pix[7:2] + 6'h0b;
  assign p1_actual_index__45_comb = p0_start_pix + p1_idx_u8__45_comb;
  assign p1_add_8407_comb = p0_start_pix[7:1] + 7'h17;
  assign p1_actual_index__47_comb = p0_start_pix + p1_idx_u8__47_comb;
  assign p1_add_8409_comb = p0_start_pix[7:4] + 4'h3;
  assign p1_actual_index__49_comb = p0_start_pix + p1_idx_u8__49_comb;
  assign p1_add_8411_comb = p0_start_pix[7:1] + 7'h19;
  assign p1_actual_index__51_comb = p0_start_pix + p1_idx_u8__51_comb;
  assign p1_add_8413_comb = p0_start_pix[7:2] + 6'h0d;
  assign p1_actual_index__53_comb = p0_start_pix + p1_idx_u8__53_comb;
  assign p1_add_8415_comb = p0_start_pix[7:1] + 7'h1b;
  assign p1_actual_index__55_comb = p0_start_pix + p1_idx_u8__55_comb;
  assign p1_add_8417_comb = p0_start_pix[7:3] + 5'h07;
  assign p1_actual_index__57_comb = p0_start_pix + p1_idx_u8__57_comb;
  assign p1_add_8419_comb = p0_start_pix[7:1] + 7'h1d;
  assign p1_actual_index__59_comb = p0_start_pix + p1_idx_u8__59_comb;
  assign p1_add_8421_comb = p0_start_pix[7:2] + 6'h0f;
  assign p1_actual_index__61_comb = p0_start_pix + p1_idx_u8__61_comb;
  assign p1_add_8423_comb = p0_start_pix[7:1] + 7'h1f;
  assign p1_flat_comb[0] = p1_array_concat_8163_comb[0];
  assign p1_flat_comb[1] = p1_array_concat_8163_comb[1];
  assign p1_flat_comb[2] = p1_array_concat_8163_comb[2];
  assign p1_flat_comb[3] = p1_array_concat_8163_comb[3];
  assign p1_flat_comb[4] = p1_array_concat_8163_comb[4];
  assign p1_flat_comb[5] = p1_array_concat_8163_comb[5];
  assign p1_flat_comb[6] = p1_array_concat_8163_comb[6];
  assign p1_flat_comb[7] = p1_array_concat_8163_comb[7];
  assign p1_flat_comb[8] = p1_array_concat_8163_comb[8];
  assign p1_flat_comb[9] = p1_array_concat_8163_comb[9];
  assign p1_flat_comb[10] = p1_array_concat_8163_comb[10];
  assign p1_flat_comb[11] = p1_array_concat_8163_comb[11];
  assign p1_flat_comb[12] = p1_array_concat_8163_comb[12];
  assign p1_flat_comb[13] = p1_array_concat_8163_comb[13];
  assign p1_flat_comb[14] = p1_array_concat_8163_comb[14];
  assign p1_flat_comb[15] = p1_array_concat_8163_comb[15];
  assign p1_flat_comb[16] = p1_array_concat_8163_comb[16];
  assign p1_flat_comb[17] = p1_array_concat_8163_comb[17];
  assign p1_flat_comb[18] = p1_array_concat_8163_comb[18];
  assign p1_flat_comb[19] = p1_array_concat_8163_comb[19];
  assign p1_flat_comb[20] = p1_array_concat_8163_comb[20];
  assign p1_flat_comb[21] = p1_array_concat_8163_comb[21];
  assign p1_flat_comb[22] = p1_array_concat_8163_comb[22];
  assign p1_flat_comb[23] = p1_array_concat_8163_comb[23];
  assign p1_flat_comb[24] = p1_array_concat_8163_comb[24];
  assign p1_flat_comb[25] = p1_array_concat_8163_comb[25];
  assign p1_flat_comb[26] = p1_array_concat_8163_comb[26];
  assign p1_flat_comb[27] = p1_array_concat_8163_comb[27];
  assign p1_flat_comb[28] = p1_array_concat_8163_comb[28];
  assign p1_flat_comb[29] = p1_array_concat_8163_comb[29];
  assign p1_flat_comb[30] = p1_array_concat_8163_comb[30];
  assign p1_flat_comb[31] = p1_array_concat_8163_comb[31];
  assign p1_flat_comb[32] = p1_array_concat_8163_comb[32];
  assign p1_flat_comb[33] = p1_array_concat_8163_comb[33];
  assign p1_flat_comb[34] = p1_array_concat_8163_comb[34];
  assign p1_flat_comb[35] = p1_array_concat_8163_comb[35];
  assign p1_flat_comb[36] = p1_array_concat_8163_comb[36];
  assign p1_flat_comb[37] = p1_array_concat_8163_comb[37];
  assign p1_flat_comb[38] = p1_array_concat_8163_comb[38];
  assign p1_flat_comb[39] = p1_array_concat_8163_comb[39];
  assign p1_flat_comb[40] = p1_array_concat_8163_comb[40];
  assign p1_flat_comb[41] = p1_array_concat_8163_comb[41];
  assign p1_flat_comb[42] = p1_array_concat_8163_comb[42];
  assign p1_flat_comb[43] = p1_array_concat_8163_comb[43];
  assign p1_flat_comb[44] = p1_array_concat_8163_comb[44];
  assign p1_flat_comb[45] = p1_array_concat_8163_comb[45];
  assign p1_flat_comb[46] = p1_array_concat_8163_comb[46];
  assign p1_flat_comb[47] = p1_array_concat_8163_comb[47];
  assign p1_flat_comb[48] = p1_array_concat_8163_comb[48];
  assign p1_flat_comb[49] = p1_array_concat_8163_comb[49];
  assign p1_flat_comb[50] = p1_array_concat_8163_comb[50];
  assign p1_flat_comb[51] = p1_array_concat_8163_comb[51];
  assign p1_flat_comb[52] = p1_array_concat_8163_comb[52];
  assign p1_flat_comb[53] = p1_array_concat_8163_comb[53];
  assign p1_flat_comb[54] = p1_array_concat_8163_comb[54];
  assign p1_flat_comb[55] = p1_array_concat_8163_comb[55];
  assign p1_flat_comb[56] = p1_row7_comb[0];
  assign p1_flat_comb[57] = p1_row7_comb[1];
  assign p1_flat_comb[58] = p1_row7_comb[2];
  assign p1_flat_comb[59] = p1_row7_comb[3];
  assign p1_flat_comb[60] = p1_row7_comb[4];
  assign p1_flat_comb[61] = p1_row7_comb[5];
  assign p1_flat_comb[62] = p1_row7_comb[6];
  assign p1_flat_comb[63] = p1_row7_comb[7];
  assign p1_actual_index__14_comb = {p1_add_8159_comb, p0_start_pix[0]};
  assign p1_actual_index__2_comb = {p1_add_8274_comb, p0_start_pix[0]};
  assign p1_actual_index__4_comb = {p1_add_8257_comb, p0_start_pix[1:0]};
  assign p1_actual_index__6_comb = {p1_add_8241_comb, p0_start_pix[0]};
  assign p1_actual_index__10_comb = {p1_add_8192_comb, p0_start_pix[0]};
  assign p1_actual_index__12_comb = {p1_add_8168_comb, p0_start_pix[1:0]};
  assign p1_actual_index__8_comb = {p1_add_8211_comb, p0_start_pix[2:0]};
  assign p1_actual_index__16_comb = {p1_add_8377_comb, p0_start_pix[3:0]};
  assign p1_actual_index__18_comb = {p1_add_8379_comb, p0_start_pix[0]};
  assign p1_actual_index__20_comb = {p1_add_8381_comb, p0_start_pix[1:0]};
  assign p1_actual_index__22_comb = {p1_add_8383_comb, p0_start_pix[0]};
  assign p1_actual_index__24_comb = {p1_add_8385_comb, p0_start_pix[2:0]};
  assign p1_actual_index__26_comb = {p1_add_8387_comb, p0_start_pix[0]};
  assign p1_actual_index__28_comb = {p1_add_8389_comb, p0_start_pix[1:0]};
  assign p1_actual_index__30_comb = {p1_add_8391_comb, p0_start_pix[0]};
  assign p1_actual_index__32_comb = {p1_add_8393_comb, p0_start_pix[4:0]};
  assign p1_actual_index__34_comb = {p1_add_8395_comb, p0_start_pix[0]};
  assign p1_actual_index__36_comb = {p1_add_8397_comb, p0_start_pix[1:0]};
  assign p1_actual_index__38_comb = {p1_add_8399_comb, p0_start_pix[0]};
  assign p1_actual_index__40_comb = {p1_add_8401_comb, p0_start_pix[2:0]};
  assign p1_actual_index__42_comb = {p1_add_8403_comb, p0_start_pix[0]};
  assign p1_actual_index__44_comb = {p1_add_8405_comb, p0_start_pix[1:0]};
  assign p1_actual_index__46_comb = {p1_add_8407_comb, p0_start_pix[0]};
  assign p1_actual_index__48_comb = {p1_add_8409_comb, p0_start_pix[3:0]};
  assign p1_actual_index__50_comb = {p1_add_8411_comb, p0_start_pix[0]};
  assign p1_actual_index__52_comb = {p1_add_8413_comb, p0_start_pix[1:0]};
  assign p1_actual_index__54_comb = {p1_add_8415_comb, p0_start_pix[0]};
  assign p1_actual_index__56_comb = {p1_add_8417_comb, p0_start_pix[2:0]};
  assign p1_actual_index__58_comb = {p1_add_8419_comb, p0_start_pix[0]};
  assign p1_actual_index__60_comb = {p1_add_8421_comb, p0_start_pix[1:0]};
  assign p1_actual_index__62_comb = {p1_add_8423_comb, p0_start_pix[0]};
  assign p1_value_comb = p0_matrix[3'h0][3'h0];
  assign p1_and_8187_comb = p1_flat_comb[p1_actual_index__14_comb > 8'h3f ? 6'h3f : p1_actual_index__14_comb[5:0]] & {10{~(p1_add_8159_comb[5] | p1_add_8159_comb[6])}};
  assign p1_and_8318_comb = p1_flat_comb[p0_start_pix > 8'h3f ? 6'h3f : p0_start_pix[5:0]] & {10{~(p0_start_pix[6] | p0_start_pix[7])}};
  assign p1_and_8320_comb = p1_flat_comb[p1_actual_index__1_comb > 8'h3f ? 6'h3f : p1_actual_index__1_comb[5:0]] & {10{~(p1_actual_index__1_comb[6] | p1_actual_index__1_comb[7])}};
  assign p1_and_8315_comb = p1_flat_comb[p1_actual_index__2_comb > 8'h3f ? 6'h3f : p1_actual_index__2_comb[5:0]] & {10{~(p1_add_8274_comb[5] | p1_add_8274_comb[6])}};
  assign p1_and_8308_comb = p1_flat_comb[p1_actual_index__3_comb > 8'h3f ? 6'h3f : p1_actual_index__3_comb[5:0]] & {10{~(p1_actual_index__3_comb[6] | p1_actual_index__3_comb[7])}};
  assign p1_and_8301_comb = p1_flat_comb[p1_actual_index__4_comb > 8'h3f ? 6'h3f : p1_actual_index__4_comb[5:0]] & {10{~(p1_add_8257_comb[4] | p1_add_8257_comb[5])}};
  assign p1_and_8290_comb = p1_flat_comb[p1_actual_index__5_comb > 8'h3f ? 6'h3f : p1_actual_index__5_comb[5:0]] & {10{~(p1_actual_index__5_comb[6] | p1_actual_index__5_comb[7])}};
  assign p1_and_8281_comb = p1_flat_comb[p1_actual_index__6_comb > 8'h3f ? 6'h3f : p1_actual_index__6_comb[5:0]] & {10{~(p1_add_8241_comb[5] | p1_add_8241_comb[6])}};
  assign p1_and_8271_comb = p1_flat_comb[p1_actual_index__7_comb > 8'h3f ? 6'h3f : p1_actual_index__7_comb[5:0]] & {10{~(p1_actual_index__7_comb[6] | p1_actual_index__7_comb[7])}};
  assign p1_and_8244_comb = p1_flat_comb[p1_actual_index__9_comb > 8'h3f ? 6'h3f : p1_actual_index__9_comb[5:0]] & {10{~(p1_actual_index__9_comb[6] | p1_actual_index__9_comb[7])}};
  assign p1_and_8235_comb = p1_flat_comb[p1_actual_index__10_comb > 8'h3f ? 6'h3f : p1_actual_index__10_comb[5:0]] & {10{~(p1_add_8192_comb[5] | p1_add_8192_comb[6])}};
  assign p1_and_8227_comb = p1_flat_comb[p1_actual_index__11_comb > 8'h3f ? 6'h3f : p1_actual_index__11_comb[5:0]] & {10{~(p1_actual_index__11_comb[6] | p1_actual_index__11_comb[7])}};
  assign p1_and_8195_comb = p1_flat_comb[p1_actual_index__13_comb > 8'h3f ? 6'h3f : p1_actual_index__13_comb[5:0]] & {10{~(p1_actual_index__13_comb[6] | p1_actual_index__13_comb[7])}};
  assign p1_bin_value_comb = p1_value_comb[7:0];
  assign p1_eq_8198_comb = p1_and_8187_comb == 10'h000;
  assign p1_and_8199_comb = p1_flat_comb[p1_actual_index__12_comb > 8'h3f ? 6'h3f : p1_actual_index__12_comb[5:0]] & {10{~(p1_add_8168_comb[4] | p1_add_8168_comb[5])}};
  assign p1_ne_8323_comb = p1_and_8318_comb != 10'h000;
  assign p1_ne_8324_comb = p1_and_8320_comb != 10'h000;
  assign p1_ne_8322_comb = p1_and_8315_comb != 10'h000;
  assign p1_ne_8317_comb = p1_and_8308_comb != 10'h000;
  assign p1_ne_8310_comb = p1_and_8301_comb != 10'h000;
  assign p1_ne_8303_comb = p1_and_8290_comb != 10'h000;
  assign p1_ne_8292_comb = p1_and_8281_comb != 10'h000;
  assign p1_ne_8283_comb = p1_and_8271_comb != 10'h000;
  assign p1_and_8247_comb = p1_flat_comb[p1_actual_index__8_comb > 8'h3f ? 6'h3f : p1_actual_index__8_comb[5:0]] & {10{~(p1_add_8211_comb[3] | p1_add_8211_comb[4])}};
  assign p1_ne_8254_comb = p1_and_8244_comb != 10'h000;
  assign p1_ne_8246_comb = p1_and_8235_comb != 10'h000;
  assign p1_ne_8237_comb = p1_and_8227_comb != 10'h000;
  assign p1_ne_8207_comb = p1_and_8195_comb != 10'h000;
  assign p1_flipped_comb = ~p1_bin_value_comb;
  assign p1_idx_u8__1_squeezed_comb = 2'h1;
  assign p1_eq_8210_comb = p1_and_8199_comb == 10'h000;
  assign p1_not_8325_comb = ~p1_ne_8323_comb;
  assign p1_eq_8255_comb = p1_and_8247_comb == 10'h000;
  assign p1_sel_8218_comb = p1_ne_8207_comb ? p1_idx_u8__1_squeezed_comb : {1'h1, p1_eq_8198_comb};
  assign p1_sign_ext_8219_comb = {2{p1_eq_8210_comb}};
  assign p1_and_8848_comb = p1_not_8325_comb & ~p1_ne_8324_comb & ~p1_ne_8322_comb & ~p1_ne_8317_comb & ~p1_ne_8310_comb & ~p1_ne_8303_comb & ~p1_ne_8292_comb & ~p1_ne_8283_comb & p1_eq_8255_comb & ~p1_ne_8254_comb & ~p1_ne_8246_comb & ~p1_ne_8237_comb & p1_eq_8210_comb & ~p1_ne_8207_comb & p1_eq_8198_comb & (p1_flat_comb[p1_actual_index__15_comb > 8'h3f ? 6'h3f : p1_actual_index__15_comb[5:0]] & {10{~(p1_actual_index__15_comb[6] | p1_actual_index__15_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__16_comb > 8'h3f ? 6'h3f : p1_actual_index__16_comb[5:0]] & {10{~(p1_add_8377_comb[2] | p1_add_8377_comb[3])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__17_comb > 8'h3f ? 6'h3f : p1_actual_index__17_comb[5:0]] & {10{~(p1_actual_index__17_comb[6] | p1_actual_index__17_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__18_comb > 8'h3f ? 6'h3f : p1_actual_index__18_comb[5:0]] & {10{~(p1_add_8379_comb[5] | p1_add_8379_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__19_comb > 8'h3f ? 6'h3f : p1_actual_index__19_comb[5:0]] & {10{~(p1_actual_index__19_comb[6] | p1_actual_index__19_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__20_comb > 8'h3f ? 6'h3f : p1_actual_index__20_comb[5:0]] & {10{~(p1_add_8381_comb[4] | p1_add_8381_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__21_comb > 8'h3f ? 6'h3f : p1_actual_index__21_comb[5:0]] & {10{~(p1_actual_index__21_comb[6] | p1_actual_index__21_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__22_comb > 8'h3f ? 6'h3f : p1_actual_index__22_comb[5:0]] & {10{~(p1_add_8383_comb[5] | p1_add_8383_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__23_comb > 8'h3f ? 6'h3f : p1_actual_index__23_comb[5:0]] & {10{~(p1_actual_index__23_comb[6] | p1_actual_index__23_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__24_comb > 8'h3f ? 6'h3f : p1_actual_index__24_comb[5:0]] & {10{~(p1_add_8385_comb[3] | p1_add_8385_comb[4])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__25_comb > 8'h3f ? 6'h3f : p1_actual_index__25_comb[5:0]] & {10{~(p1_actual_index__25_comb[6] | p1_actual_index__25_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__26_comb > 8'h3f ? 6'h3f : p1_actual_index__26_comb[5:0]] & {10{~(p1_add_8387_comb[5] | p1_add_8387_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__27_comb > 8'h3f ? 6'h3f : p1_actual_index__27_comb[5:0]] & {10{~(p1_actual_index__27_comb[6] | p1_actual_index__27_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__28_comb > 8'h3f ? 6'h3f : p1_actual_index__28_comb[5:0]] & {10{~(p1_add_8389_comb[4] | p1_add_8389_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__29_comb > 8'h3f ? 6'h3f : p1_actual_index__29_comb[5:0]] & {10{~(p1_actual_index__29_comb[6] | p1_actual_index__29_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__30_comb > 8'h3f ? 6'h3f : p1_actual_index__30_comb[5:0]] & {10{~(p1_add_8391_comb[5] | p1_add_8391_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__31_comb > 8'h3f ? 6'h3f : p1_actual_index__31_comb[5:0]] & {10{~(p1_actual_index__31_comb[6] | p1_actual_index__31_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__32_comb > 8'h3f ? 6'h3f : p1_actual_index__32_comb[5:0]] & {10{~(p1_add_8393_comb[1] | p1_add_8393_comb[2])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__33_comb > 8'h3f ? 6'h3f : p1_actual_index__33_comb[5:0]] & {10{~(p1_actual_index__33_comb[6] | p1_actual_index__33_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__34_comb > 8'h3f ? 6'h3f : p1_actual_index__34_comb[5:0]] & {10{~(p1_add_8395_comb[5] | p1_add_8395_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__35_comb > 8'h3f ? 6'h3f : p1_actual_index__35_comb[5:0]] & {10{~(p1_actual_index__35_comb[6] | p1_actual_index__35_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__36_comb > 8'h3f ? 6'h3f : p1_actual_index__36_comb[5:0]] & {10{~(p1_add_8397_comb[4] | p1_add_8397_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__37_comb > 8'h3f ? 6'h3f : p1_actual_index__37_comb[5:0]] & {10{~(p1_actual_index__37_comb[6] | p1_actual_index__37_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__38_comb > 8'h3f ? 6'h3f : p1_actual_index__38_comb[5:0]] & {10{~(p1_add_8399_comb[5] | p1_add_8399_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__39_comb > 8'h3f ? 6'h3f : p1_actual_index__39_comb[5:0]] & {10{~(p1_actual_index__39_comb[6] | p1_actual_index__39_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__40_comb > 8'h3f ? 6'h3f : p1_actual_index__40_comb[5:0]] & {10{~(p1_add_8401_comb[3] | p1_add_8401_comb[4])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__41_comb > 8'h3f ? 6'h3f : p1_actual_index__41_comb[5:0]] & {10{~(p1_actual_index__41_comb[6] | p1_actual_index__41_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__42_comb > 8'h3f ? 6'h3f : p1_actual_index__42_comb[5:0]] & {10{~(p1_add_8403_comb[5] | p1_add_8403_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__43_comb > 8'h3f ? 6'h3f : p1_actual_index__43_comb[5:0]] & {10{~(p1_actual_index__43_comb[6] | p1_actual_index__43_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__44_comb > 8'h3f ? 6'h3f : p1_actual_index__44_comb[5:0]] & {10{~(p1_add_8405_comb[4] | p1_add_8405_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__45_comb > 8'h3f ? 6'h3f : p1_actual_index__45_comb[5:0]] & {10{~(p1_actual_index__45_comb[6] | p1_actual_index__45_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__46_comb > 8'h3f ? 6'h3f : p1_actual_index__46_comb[5:0]] & {10{~(p1_add_8407_comb[5] | p1_add_8407_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__47_comb > 8'h3f ? 6'h3f : p1_actual_index__47_comb[5:0]] & {10{~(p1_actual_index__47_comb[6] | p1_actual_index__47_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__48_comb > 8'h3f ? 6'h3f : p1_actual_index__48_comb[5:0]] & {10{~(p1_add_8409_comb[2] | p1_add_8409_comb[3])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__49_comb > 8'h3f ? 6'h3f : p1_actual_index__49_comb[5:0]] & {10{~(p1_actual_index__49_comb[6] | p1_actual_index__49_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__50_comb > 8'h3f ? 6'h3f : p1_actual_index__50_comb[5:0]] & {10{~(p1_add_8411_comb[5] | p1_add_8411_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__51_comb > 8'h3f ? 6'h3f : p1_actual_index__51_comb[5:0]] & {10{~(p1_actual_index__51_comb[6] | p1_actual_index__51_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__52_comb > 8'h3f ? 6'h3f : p1_actual_index__52_comb[5:0]] & {10{~(p1_add_8413_comb[4] | p1_add_8413_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__53_comb > 8'h3f ? 6'h3f : p1_actual_index__53_comb[5:0]] & {10{~(p1_actual_index__53_comb[6] | p1_actual_index__53_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__54_comb > 8'h3f ? 6'h3f : p1_actual_index__54_comb[5:0]] & {10{~(p1_add_8415_comb[5] | p1_add_8415_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__55_comb > 8'h3f ? 6'h3f : p1_actual_index__55_comb[5:0]] & {10{~(p1_actual_index__55_comb[6] | p1_actual_index__55_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__56_comb > 8'h3f ? 6'h3f : p1_actual_index__56_comb[5:0]] & {10{~(p1_add_8417_comb[3] | p1_add_8417_comb[4])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__57_comb > 8'h3f ? 6'h3f : p1_actual_index__57_comb[5:0]] & {10{~(p1_actual_index__57_comb[6] | p1_actual_index__57_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__58_comb > 8'h3f ? 6'h3f : p1_actual_index__58_comb[5:0]] & {10{~(p1_add_8419_comb[5] | p1_add_8419_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__59_comb > 8'h3f ? 6'h3f : p1_actual_index__59_comb[5:0]] & {10{~(p1_actual_index__59_comb[6] | p1_actual_index__59_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__60_comb > 8'h3f ? 6'h3f : p1_actual_index__60_comb[5:0]] & {10{~(p1_add_8421_comb[4] | p1_add_8421_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__61_comb > 8'h3f ? 6'h3f : p1_actual_index__61_comb[5:0]] & {10{~(p1_actual_index__61_comb[6] | p1_actual_index__61_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__62_comb > 8'h3f ? 6'h3f : p1_actual_index__62_comb[5:0]] & {10{~(p1_add_8423_comb[5] | p1_add_8423_comb[6])}}) == 10'h000;
  assign p1_code_list_comb = ($signed(p1_value_comb) <= $signed(10'h000) ? p1_flipped_comb : p1_bin_value_comb) & {8{p1_value_comb != 10'h000}};

  // Registers for pipe stage 1:
  reg p1_is_luminance;
  reg [9:0] p1_and_8187;
  reg [9:0] p1_and_8195;
  reg [9:0] p1_and_8199;
  reg [1:0] p1_sel_8218;
  reg [1:0] p1_sign_ext_8219;
  reg [9:0] p1_and_8227;
  reg [9:0] p1_and_8235;
  reg p1_ne_8237;
  reg [9:0] p1_and_8244;
  reg p1_ne_8246;
  reg [9:0] p1_and_8247;
  reg p1_ne_8254;
  reg p1_eq_8255;
  reg [9:0] p1_and_8271;
  reg [9:0] p1_and_8281;
  reg p1_ne_8283;
  reg [9:0] p1_and_8290;
  reg p1_ne_8292;
  reg [9:0] p1_and_8301;
  reg p1_ne_8303;
  reg [9:0] p1_and_8308;
  reg p1_ne_8310;
  reg [9:0] p1_and_8315;
  reg p1_ne_8317;
  reg [9:0] p1_and_8318;
  reg [9:0] p1_and_8320;
  reg p1_ne_8322;
  reg p1_ne_8323;
  reg p1_ne_8324;
  reg p1_not_8325;
  reg p1_and_8848;
  reg [7:0] p1_code_list;
  always @ (posedge clk) begin
    p1_is_luminance <= p0_is_luminance;
    p1_and_8187 <= p1_and_8187_comb;
    p1_and_8195 <= p1_and_8195_comb;
    p1_and_8199 <= p1_and_8199_comb;
    p1_sel_8218 <= p1_sel_8218_comb;
    p1_sign_ext_8219 <= p1_sign_ext_8219_comb;
    p1_and_8227 <= p1_and_8227_comb;
    p1_and_8235 <= p1_and_8235_comb;
    p1_ne_8237 <= p1_ne_8237_comb;
    p1_and_8244 <= p1_and_8244_comb;
    p1_ne_8246 <= p1_ne_8246_comb;
    p1_and_8247 <= p1_and_8247_comb;
    p1_ne_8254 <= p1_ne_8254_comb;
    p1_eq_8255 <= p1_eq_8255_comb;
    p1_and_8271 <= p1_and_8271_comb;
    p1_and_8281 <= p1_and_8281_comb;
    p1_ne_8283 <= p1_ne_8283_comb;
    p1_and_8290 <= p1_and_8290_comb;
    p1_ne_8292 <= p1_ne_8292_comb;
    p1_and_8301 <= p1_and_8301_comb;
    p1_ne_8303 <= p1_ne_8303_comb;
    p1_and_8308 <= p1_and_8308_comb;
    p1_ne_8310 <= p1_ne_8310_comb;
    p1_and_8315 <= p1_and_8315_comb;
    p1_ne_8317 <= p1_ne_8317_comb;
    p1_and_8318 <= p1_and_8318_comb;
    p1_and_8320 <= p1_and_8320_comb;
    p1_ne_8322 <= p1_ne_8322_comb;
    p1_ne_8323 <= p1_ne_8323_comb;
    p1_ne_8324 <= p1_ne_8324_comb;
    p1_not_8325 <= p1_not_8325_comb;
    p1_and_8848 <= p1_and_8848_comb;
    p1_code_list <= p1_code_list_comb;
  end

  // ===== Pipe stage 2:
  wire [2:0] p2_and_8935_comb;
  wire [3:0] p2_sel_8944_comb;
  wire [3:0] p2_sel_8948_comb;
  assign p2_and_8935_comb = (p1_ne_8254 ? 3'h1 : (p1_ne_8246 ? 3'h2 : (p1_ne_8237 ? 3'h3 : {1'h1, p1_sel_8218 & p1_sign_ext_8219}))) & {3{p1_eq_8255}};
  assign p2_sel_8944_comb = p1_ne_8310 ? 4'h4 : (p1_ne_8303 ? 4'h5 : (p1_ne_8292 ? 4'h6 : (p1_ne_8283 ? 4'h7 : {1'h1, p2_and_8935_comb})));
  assign p2_sel_8948_comb = p1_ne_8322 ? 4'h2 : (p1_ne_8317 ? 4'h3 : p2_sel_8944_comb);

  // Registers for pipe stage 2:
  reg p2_is_luminance;
  reg [9:0] p2_and_8187;
  reg [9:0] p2_and_8195;
  reg [9:0] p2_and_8199;
  reg [9:0] p2_and_8227;
  reg [9:0] p2_and_8235;
  reg [9:0] p2_and_8244;
  reg [9:0] p2_and_8247;
  reg [9:0] p2_and_8271;
  reg [9:0] p2_and_8281;
  reg [9:0] p2_and_8290;
  reg [9:0] p2_and_8301;
  reg [9:0] p2_and_8308;
  reg [9:0] p2_and_8315;
  reg [9:0] p2_and_8318;
  reg [9:0] p2_and_8320;
  reg p2_ne_8323;
  reg p2_ne_8324;
  reg [3:0] p2_sel_8948;
  reg p2_not_8325;
  reg p2_and_8848;
  reg [7:0] p2_code_list;
  always @ (posedge clk) begin
    p2_is_luminance <= p1_is_luminance;
    p2_and_8187 <= p1_and_8187;
    p2_and_8195 <= p1_and_8195;
    p2_and_8199 <= p1_and_8199;
    p2_and_8227 <= p1_and_8227;
    p2_and_8235 <= p1_and_8235;
    p2_and_8244 <= p1_and_8244;
    p2_and_8247 <= p1_and_8247;
    p2_and_8271 <= p1_and_8271;
    p2_and_8281 <= p1_and_8281;
    p2_and_8290 <= p1_and_8290;
    p2_and_8301 <= p1_and_8301;
    p2_and_8308 <= p1_and_8308;
    p2_and_8315 <= p1_and_8315;
    p2_and_8318 <= p1_and_8318;
    p2_and_8320 <= p1_and_8320;
    p2_ne_8323 <= p1_ne_8323;
    p2_ne_8324 <= p1_ne_8324;
    p2_sel_8948 <= p2_sel_8948_comb;
    p2_not_8325 <= p1_not_8325;
    p2_and_8848 <= p1_and_8848;
    p2_code_list <= p1_code_list;
  end

  // ===== Pipe stage 3:
  wire [3:0] p3_sel_8994_comb;
  wire [3:0] p3_run_comb;
  wire [9:0] p3_value__1_comb;
  wire [7:0] p3_bin_value__2_comb;
  wire [7:0] p3_value_abs_comb;
  wire [1:0] p3_idx_u8__1_squeezed__1_comb;
  wire [1:0] p3_idx_u8__2_squeezed_comb;
  wire [1:0] p3_idx_u8__3_squeezed_comb;
  wire p3_eq_9030_comb;
  wire [7:0] p3_flipped__1_comb;
  wire [2:0] p3_idx_u8__4_squeezed__1_comb;
  wire [7:0] p3_code_list__1_comb;
  wire [2:0] p3_sel_9020_comb;
  wire [2:0] p3_idx_u8__5_squeezed__1_comb;
  wire p3_or_reduce_9023_comb;
  wire [2:0] p3_sel_9024_comb;
  wire p3_or_reduce_9025_comb;
  wire p3_bit_slice_9026_comb;
  wire p3_ne_9028_comb;
  wire p3_or_9032_comb;
  wire [7:0] p3_sel_9043_comb;
  wire [3:0] p3_sel_9044_comb;
  assign p3_sel_8994_comb = p2_ne_8324 ? 4'h1 : p2_sel_8948;
  assign p3_run_comb = p3_sel_8994_comb & {4{p2_not_8325}};
  assign p3_value__1_comb = p3_run_comb == 4'h0 ? p2_and_8318 : (p3_run_comb == 4'h1 ? p2_and_8320 : (p3_run_comb == 4'h2 ? p2_and_8315 : (p3_run_comb == 4'h3 ? p2_and_8308 : (p3_run_comb == 4'h4 ? p2_and_8301 : (p3_run_comb == 4'h5 ? p2_and_8290 : (p3_run_comb == 4'h6 ? p2_and_8281 : (p3_run_comb == 4'h7 ? p2_and_8271 : (p3_run_comb == 4'h8 ? p2_and_8247 : (p3_run_comb == 4'h9 ? p2_and_8244 : (p3_run_comb == 4'ha ? p2_and_8235 : (p3_run_comb == 4'hb ? p2_and_8227 : (p3_run_comb == 4'hc ? p2_and_8199 : (p3_run_comb == 4'hd ? p2_and_8195 : (p3_run_comb == 4'he ? p2_and_8187 : 10'h000))))))))))))));
  assign p3_bin_value__2_comb = p3_value__1_comb[7:0];
  assign p3_value_abs_comb = p3_value__1_comb[9] ? -p3_bin_value__2_comb : p3_bin_value__2_comb;
  assign p3_idx_u8__1_squeezed__1_comb = 2'h1;
  assign p3_idx_u8__2_squeezed_comb = 2'h2;
  assign p3_idx_u8__3_squeezed_comb = 2'h3;
  assign p3_eq_9030_comb = p3_run_comb == 4'hf;
  assign p3_flipped__1_comb = ~p3_bin_value__2_comb;
  assign p3_idx_u8__4_squeezed__1_comb = 3'h4;
  assign p3_code_list__1_comb = $signed(p3_value__1_comb) <= $signed(10'h000) ? p3_flipped__1_comb : p3_bin_value__2_comb;
  assign p3_sel_9020_comb = |p3_value_abs_comb[7:3] ? p3_idx_u8__4_squeezed__1_comb : {1'h0, |p3_value_abs_comb[7:2] ? p3_idx_u8__3_squeezed_comb : (|p3_value_abs_comb[7:1] ? p3_idx_u8__2_squeezed_comb : p3_idx_u8__1_squeezed__1_comb)};
  assign p3_idx_u8__5_squeezed__1_comb = 3'h5;
  assign p3_or_reduce_9023_comb = |p3_value_abs_comb[7:5];
  assign p3_sel_9024_comb = |p3_value_abs_comb[7:4] ? p3_idx_u8__5_squeezed__1_comb : p3_sel_9020_comb;
  assign p3_or_reduce_9025_comb = |p3_value_abs_comb[7:6];
  assign p3_bit_slice_9026_comb = p3_value_abs_comb[7];
  assign p3_ne_9028_comb = p3_value_abs_comb != 8'h00;
  assign p3_or_9032_comb = p2_and_8848 | p3_eq_9030_comb;
  assign p3_sel_9043_comb = p2_and_8848 ? p2_code_list : p3_code_list__1_comb & {8{~p3_eq_9030_comb}};
  assign p3_sel_9044_comb = p2_and_8848 ? 4'hf : p3_sel_8994_comb & {4{~(p3_eq_9030_comb | p2_ne_8323)}};

  // Registers for pipe stage 3:
  reg p3_is_luminance;
  reg [3:0] p3_run;
  reg p3_or_reduce_9023;
  reg [2:0] p3_sel_9024;
  reg p3_or_reduce_9025;
  reg p3_bit_slice_9026;
  reg p3_ne_9028;
  reg p3_or_9032;
  reg [7:0] p3_sel_9043;
  reg [3:0] p3_sel_9044;
  always @ (posedge clk) begin
    p3_is_luminance <= p2_is_luminance;
    p3_run <= p3_run_comb;
    p3_or_reduce_9023 <= p3_or_reduce_9023_comb;
    p3_sel_9024 <= p3_sel_9024_comb;
    p3_or_reduce_9025 <= p3_or_reduce_9025_comb;
    p3_bit_slice_9026 <= p3_bit_slice_9026_comb;
    p3_ne_9028 <= p3_ne_9028_comb;
    p3_or_9032 <= p3_or_9032_comb;
    p3_sel_9043 <= p3_sel_9043_comb;
    p3_sel_9044 <= p3_sel_9044_comb;
  end

  // ===== Pipe stage 4:
  wire [2:0] p4_idx_u8__6_squeezed__1_comb;
  wire [2:0] p4_idx_u8__7_squeezed__1_comb;
  wire [3:0] p4_idx_u8__8_squeezed_comb;
  wire [7:0] p4_size_comb;
  wire [7:0] p4_run_size_str_u8_comb;
  wire [4:0] p4_huffman_length_squeezed_comb;
  wire [4:0] p4_idx_u8__2_squeezed__1_comb;
  wire [15:0] p4_huffman_code_full_comb;
  wire [35:0] p4_tuple_9097_comb;
  assign p4_idx_u8__6_squeezed__1_comb = 3'h6;
  assign p4_idx_u8__7_squeezed__1_comb = 3'h7;
  assign p4_idx_u8__8_squeezed_comb = 4'h8;
  assign p4_size_comb = {4'h0, p3_bit_slice_9026 ? p4_idx_u8__8_squeezed_comb : {1'h0, p3_or_reduce_9025 ? p4_idx_u8__7_squeezed__1_comb : (p3_or_reduce_9023 ? p4_idx_u8__6_squeezed__1_comb : p3_sel_9024)}} & {8{p3_ne_9028}};
  assign p4_run_size_str_u8_comb = {p3_run, 4'h0} | p4_size_comb;
  assign p4_huffman_length_squeezed_comb = p3_is_luminance ? literal_9081[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_9079[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_idx_u8__2_squeezed__1_comb = 5'h02;
  assign p4_huffman_code_full_comb = p3_is_luminance ? literal_9083[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_9082[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_tuple_9097_comb = {p4_huffman_code_full_comb & {16{~p3_or_9032}}, {3'h0, p3_or_9032 ? p4_idx_u8__2_squeezed__1_comb : p4_huffman_length_squeezed_comb}, p3_sel_9043, p3_sel_9044};

  // Registers for pipe stage 4:
  reg [35:0] p4_tuple_9097;
  always @ (posedge clk) begin
    p4_tuple_9097 <= p4_tuple_9097_comb;
  end
  assign out = p4_tuple_9097;
endmodule
