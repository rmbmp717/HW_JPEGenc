module Huffman_ACenc(
  input wire clk,
  input wire [511:0] matrix,
  input wire is_luminance,
  output wire [31:0] out
);
  wire [7:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[7:0];
  assign matrix_unflattened[0][1] = matrix[15:8];
  assign matrix_unflattened[0][2] = matrix[23:16];
  assign matrix_unflattened[0][3] = matrix[31:24];
  assign matrix_unflattened[0][4] = matrix[39:32];
  assign matrix_unflattened[0][5] = matrix[47:40];
  assign matrix_unflattened[0][6] = matrix[55:48];
  assign matrix_unflattened[0][7] = matrix[63:56];
  assign matrix_unflattened[1][0] = matrix[71:64];
  assign matrix_unflattened[1][1] = matrix[79:72];
  assign matrix_unflattened[1][2] = matrix[87:80];
  assign matrix_unflattened[1][3] = matrix[95:88];
  assign matrix_unflattened[1][4] = matrix[103:96];
  assign matrix_unflattened[1][5] = matrix[111:104];
  assign matrix_unflattened[1][6] = matrix[119:112];
  assign matrix_unflattened[1][7] = matrix[127:120];
  assign matrix_unflattened[2][0] = matrix[135:128];
  assign matrix_unflattened[2][1] = matrix[143:136];
  assign matrix_unflattened[2][2] = matrix[151:144];
  assign matrix_unflattened[2][3] = matrix[159:152];
  assign matrix_unflattened[2][4] = matrix[167:160];
  assign matrix_unflattened[2][5] = matrix[175:168];
  assign matrix_unflattened[2][6] = matrix[183:176];
  assign matrix_unflattened[2][7] = matrix[191:184];
  assign matrix_unflattened[3][0] = matrix[199:192];
  assign matrix_unflattened[3][1] = matrix[207:200];
  assign matrix_unflattened[3][2] = matrix[215:208];
  assign matrix_unflattened[3][3] = matrix[223:216];
  assign matrix_unflattened[3][4] = matrix[231:224];
  assign matrix_unflattened[3][5] = matrix[239:232];
  assign matrix_unflattened[3][6] = matrix[247:240];
  assign matrix_unflattened[3][7] = matrix[255:248];
  assign matrix_unflattened[4][0] = matrix[263:256];
  assign matrix_unflattened[4][1] = matrix[271:264];
  assign matrix_unflattened[4][2] = matrix[279:272];
  assign matrix_unflattened[4][3] = matrix[287:280];
  assign matrix_unflattened[4][4] = matrix[295:288];
  assign matrix_unflattened[4][5] = matrix[303:296];
  assign matrix_unflattened[4][6] = matrix[311:304];
  assign matrix_unflattened[4][7] = matrix[319:312];
  assign matrix_unflattened[5][0] = matrix[327:320];
  assign matrix_unflattened[5][1] = matrix[335:328];
  assign matrix_unflattened[5][2] = matrix[343:336];
  assign matrix_unflattened[5][3] = matrix[351:344];
  assign matrix_unflattened[5][4] = matrix[359:352];
  assign matrix_unflattened[5][5] = matrix[367:360];
  assign matrix_unflattened[5][6] = matrix[375:368];
  assign matrix_unflattened[5][7] = matrix[383:376];
  assign matrix_unflattened[6][0] = matrix[391:384];
  assign matrix_unflattened[6][1] = matrix[399:392];
  assign matrix_unflattened[6][2] = matrix[407:400];
  assign matrix_unflattened[6][3] = matrix[415:408];
  assign matrix_unflattened[6][4] = matrix[423:416];
  assign matrix_unflattened[6][5] = matrix[431:424];
  assign matrix_unflattened[6][6] = matrix[439:432];
  assign matrix_unflattened[6][7] = matrix[447:440];
  assign matrix_unflattened[7][0] = matrix[455:448];
  assign matrix_unflattened[7][1] = matrix[463:456];
  assign matrix_unflattened[7][2] = matrix[471:464];
  assign matrix_unflattened[7][3] = matrix[479:472];
  assign matrix_unflattened[7][4] = matrix[487:480];
  assign matrix_unflattened[7][5] = matrix[495:488];
  assign matrix_unflattened[7][6] = matrix[503:496];
  assign matrix_unflattened[7][7] = matrix[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_matrix[0:7][0:7];
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_array_index_4701_comb;
  wire [7:0] p1_array_index_4705_comb;
  wire p1_eq_4708_comb;
  wire [7:0] p1_array_index_4709_comb;
  wire p1_ne_4711_comb;
  wire p1_eq_4714_comb;
  wire [7:0] p1_array_index_4721_comb;
  wire [7:0] p1_array_index_4727_comb;
  wire p1_ne_4729_comb;
  wire [7:0] p1_array_index_4734_comb;
  wire p1_ne_4736_comb;
  wire [2:0] p1_sel_4737_comb;
  wire [7:0] p1_array_index_4739_comb;
  wire p1_ne_4741_comb;
  wire p1_eq_4744_comb;
  wire [7:0] p1_array_index_4751_comb;
  wire [7:0] p1_array_index_4757_comb;
  wire p1_ne_4759_comb;
  wire [7:0] p1_array_index_4764_comb;
  wire p1_ne_4766_comb;
  wire [3:0] p1_sel_4767_comb;
  wire [7:0] p1_array_index_4771_comb;
  wire p1_ne_4773_comb;
  wire [7:0] p1_array_index_4778_comb;
  wire p1_ne_4780_comb;
  wire [7:0] p1_array_index_4785_comb;
  wire p1_ne_4787_comb;
  wire [7:0] p1_array_index_4790_comb;
  wire p1_ne_4792_comb;
  wire p1_ne_4797_comb;
  wire [3:0] p1_sel_4798_comb;
  wire [7:0] p1_array_index_4800_comb;
  wire p1_ne_4803_comb;
  wire [7:0] p1_array_index_4807_comb;
  wire [7:0] p1_value_comb;
  wire [7:0] p1_flipped_comb;
  wire [7:0] p1_code_list_comb;
  wire [7:0] p1_sign_ext_5067_comb;
  wire [15:0] p1_concat_5068_comb;
  wire [31:0] p1_tuple_5071_comb;
  assign p1_array_index_4701_comb = p0_matrix[3'h1][3'h7];
  assign p1_array_index_4705_comb = p0_matrix[3'h1][3'h6];
  assign p1_eq_4708_comb = p1_array_index_4701_comb == 8'h00;
  assign p1_array_index_4709_comb = p0_matrix[3'h1][3'h5];
  assign p1_ne_4711_comb = p1_array_index_4705_comb != 8'h00;
  assign p1_eq_4714_comb = p1_array_index_4709_comb == 8'h00;
  assign p1_array_index_4721_comb = p0_matrix[3'h1][3'h4];
  assign p1_array_index_4727_comb = p0_matrix[3'h1][3'h3];
  assign p1_ne_4729_comb = p1_array_index_4721_comb != 8'h00;
  assign p1_array_index_4734_comb = p0_matrix[3'h1][3'h2];
  assign p1_ne_4736_comb = p1_array_index_4727_comb != 8'h00;
  assign p1_sel_4737_comb = p1_ne_4729_comb ? 3'h3 : {1'h1, (p1_ne_4711_comb ? 2'h1 : {1'h1, p1_eq_4708_comb}) & {2{p1_eq_4714_comb}}};
  assign p1_array_index_4739_comb = p0_matrix[3'h1][3'h1];
  assign p1_ne_4741_comb = p1_array_index_4734_comb != 8'h00;
  assign p1_eq_4744_comb = p1_array_index_4739_comb == 8'h00;
  assign p1_array_index_4751_comb = p0_matrix[3'h1][3'h0];
  assign p1_array_index_4757_comb = p0_matrix[3'h0][3'h7];
  assign p1_ne_4759_comb = p1_array_index_4751_comb != 8'h00;
  assign p1_array_index_4764_comb = p0_matrix[3'h0][3'h6];
  assign p1_ne_4766_comb = p1_array_index_4757_comb != 8'h00;
  assign p1_sel_4767_comb = p1_ne_4759_comb ? 4'h7 : {1'h1, (p1_ne_4741_comb ? 3'h1 : (p1_ne_4736_comb ? 3'h2 : p1_sel_4737_comb)) & {3{p1_eq_4744_comb}}};
  assign p1_array_index_4771_comb = p0_matrix[3'h0][3'h5];
  assign p1_ne_4773_comb = p1_array_index_4764_comb != 8'h00;
  assign p1_array_index_4778_comb = p0_matrix[3'h0][3'h4];
  assign p1_ne_4780_comb = p1_array_index_4771_comb != 8'h00;
  assign p1_array_index_4785_comb = p0_matrix[3'h0][3'h3];
  assign p1_ne_4787_comb = p1_array_index_4778_comb != 8'h00;
  assign p1_array_index_4790_comb = p0_matrix[3'h0][3'h2];
  assign p1_ne_4792_comb = p1_array_index_4785_comb != 8'h00;
  assign p1_ne_4797_comb = p1_array_index_4790_comb != 8'h00;
  assign p1_sel_4798_comb = p1_ne_4792_comb ? 4'h2 : (p1_ne_4787_comb ? 4'h3 : (p1_ne_4780_comb ? 4'h4 : (p1_ne_4773_comb ? 4'h5 : (p1_ne_4766_comb ? 4'h6 : p1_sel_4767_comb))));
  assign p1_array_index_4800_comb = p0_matrix[3'h0][3'h1];
  assign p1_ne_4803_comb = p1_array_index_4800_comb != 8'h00;
  assign p1_array_index_4807_comb = p0_matrix[3'h2][3'h0];
  assign p1_value_comb = {p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h00 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h01 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h02 ? p1_array_index_4790_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h03 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h04 ? p1_array_index_4785_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h05 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h06 ? p1_array_index_4778_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h07 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h08 ? p1_array_index_4771_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h09 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h0a ? p1_array_index_4764_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h0b ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h0c ? p1_array_index_4757_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h0d ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h0e ? p1_array_index_4751_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h0f ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h10 ? p1_array_index_4739_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h11 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h12 ? p1_array_index_4734_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h13 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h14 ? p1_array_index_4727_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h15 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h16 ? p1_array_index_4721_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h17 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h18 ? p1_array_index_4709_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h19 ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h1a ? p1_array_index_4705_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h1b ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h1c ? p1_array_index_4701_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h1d ? p1_array_index_4800_comb : ({p1_ne_4797_comb ? 4'h1 : p1_sel_4798_comb, p1_ne_4803_comb} == 5'h1e ? p1_array_index_4807_comb : p1_array_index_4800_comb))))))))))))))))))))))))))))));
  assign p1_flipped_comb = ~p1_value_comb;
  assign p1_code_list_comb = ~((|p1_value_comb[7:1]) | p1_value_comb[0]) ? p1_flipped_comb : p1_value_comb;
  assign p1_sign_ext_5067_comb = {8{~(~p1_ne_4803_comb & ~p1_ne_4797_comb & ~p1_ne_4792_comb & ~p1_ne_4787_comb & ~p1_ne_4780_comb & ~p1_ne_4773_comb & ~p1_ne_4766_comb & ~p1_ne_4759_comb & p1_eq_4744_comb & ~p1_ne_4741_comb & ~p1_ne_4736_comb & ~p1_ne_4729_comb & p1_eq_4714_comb & ~p1_ne_4711_comb & p1_eq_4708_comb & p1_array_index_4807_comb == 8'h00 & p0_matrix[3'h2][3'h1] == 8'h00 & p0_matrix[3'h2][3'h2] == 8'h00 & p0_matrix[3'h2][3'h3] == 8'h00 & p0_matrix[3'h2][3'h4] == 8'h00 & p0_matrix[3'h2][3'h5] == 8'h00 & p0_matrix[3'h2][3'h6] == 8'h00 & p0_matrix[3'h2][3'h7] == 8'h00 & p0_matrix[3'h3][3'h0] == 8'h00 & p0_matrix[3'h3][3'h1] == 8'h00 & p0_matrix[3'h3][3'h2] == 8'h00 & p0_matrix[3'h3][3'h3] == 8'h00 & p0_matrix[3'h3][3'h4] == 8'h00 & p0_matrix[3'h3][3'h5] == 8'h00 & p0_matrix[3'h3][3'h6] == 8'h00 & p0_matrix[3'h3][3'h7] == 8'h00 & p0_matrix[3'h4][3'h0] == 8'h00 & p0_matrix[3'h4][3'h1] == 8'h00 & p0_matrix[3'h4][3'h2] == 8'h00 & p0_matrix[3'h4][3'h3] == 8'h00 & p0_matrix[3'h4][3'h4] == 8'h00 & p0_matrix[3'h4][3'h5] == 8'h00 & p0_matrix[3'h4][3'h6] == 8'h00 & p0_matrix[3'h4][3'h7] == 8'h00 & p0_matrix[3'h5][3'h0] == 8'h00 & p0_matrix[3'h5][3'h1] == 8'h00 & p0_matrix[3'h5][3'h2] == 8'h00 & p0_matrix[3'h5][3'h3] == 8'h00 & p0_matrix[3'h5][3'h4] == 8'h00 & p0_matrix[3'h5][3'h5] == 8'h00 & p0_matrix[3'h5][3'h6] == 8'h00 & p0_matrix[3'h5][3'h7] == 8'h00 & p0_matrix[3'h6][3'h0] == 8'h00 & p0_matrix[3'h6][3'h1] == 8'h00 & p0_matrix[3'h6][3'h2] == 8'h00 & p0_matrix[3'h6][3'h3] == 8'h00 & p0_matrix[3'h6][3'h4] == 8'h00 & p0_matrix[3'h6][3'h5] == 8'h00 & p0_matrix[3'h6][3'h6] == 8'h00 & p0_matrix[3'h6][3'h7] == 8'h00 & p0_matrix[3'h7][3'h0] == 8'h00 & p0_matrix[3'h7][3'h1] == 8'h00 & p0_matrix[3'h7][3'h2] == 8'h00 & p0_matrix[3'h7][3'h3] == 8'h00 & p0_matrix[3'h7][3'h4] == 8'h00 & p0_matrix[3'h7][3'h5] == 8'h00 & p0_matrix[3'h7][3'h6] == 8'h00 & p0_matrix[3'h7][3'h7] == 8'h00)}};
  assign p1_concat_5068_comb = {15'h0000, ~(~p1_ne_4803_comb & ~p1_ne_4797_comb & ~p1_ne_4792_comb & ~p1_ne_4787_comb & ~p1_ne_4780_comb & ~p1_ne_4773_comb & ~p1_ne_4766_comb & ~p1_ne_4759_comb & p1_eq_4744_comb & ~p1_ne_4741_comb & ~p1_ne_4736_comb & ~p1_ne_4729_comb & p1_eq_4714_comb & ~p1_ne_4711_comb & p1_eq_4708_comb & p1_array_index_4807_comb == 8'h00 & p0_matrix[3'h2][3'h1] == 8'h00 & p0_matrix[3'h2][3'h2] == 8'h00 & p0_matrix[3'h2][3'h3] == 8'h00 & p0_matrix[3'h2][3'h4] == 8'h00 & p0_matrix[3'h2][3'h5] == 8'h00 & p0_matrix[3'h2][3'h6] == 8'h00 & p0_matrix[3'h2][3'h7] == 8'h00 & p0_matrix[3'h3][3'h0] == 8'h00 & p0_matrix[3'h3][3'h1] == 8'h00 & p0_matrix[3'h3][3'h2] == 8'h00 & p0_matrix[3'h3][3'h3] == 8'h00 & p0_matrix[3'h3][3'h4] == 8'h00 & p0_matrix[3'h3][3'h5] == 8'h00 & p0_matrix[3'h3][3'h6] == 8'h00 & p0_matrix[3'h3][3'h7] == 8'h00 & p0_matrix[3'h4][3'h0] == 8'h00 & p0_matrix[3'h4][3'h1] == 8'h00 & p0_matrix[3'h4][3'h2] == 8'h00 & p0_matrix[3'h4][3'h3] == 8'h00 & p0_matrix[3'h4][3'h4] == 8'h00 & p0_matrix[3'h4][3'h5] == 8'h00 & p0_matrix[3'h4][3'h6] == 8'h00 & p0_matrix[3'h4][3'h7] == 8'h00 & p0_matrix[3'h5][3'h0] == 8'h00 & p0_matrix[3'h5][3'h1] == 8'h00 & p0_matrix[3'h5][3'h2] == 8'h00 & p0_matrix[3'h5][3'h3] == 8'h00 & p0_matrix[3'h5][3'h4] == 8'h00 & p0_matrix[3'h5][3'h5] == 8'h00 & p0_matrix[3'h5][3'h6] == 8'h00 & p0_matrix[3'h5][3'h7] == 8'h00 & p0_matrix[3'h6][3'h0] == 8'h00 & p0_matrix[3'h6][3'h1] == 8'h00 & p0_matrix[3'h6][3'h2] == 8'h00 & p0_matrix[3'h6][3'h3] == 8'h00 & p0_matrix[3'h6][3'h4] == 8'h00 & p0_matrix[3'h6][3'h5] == 8'h00 & p0_matrix[3'h6][3'h6] == 8'h00 & p0_matrix[3'h6][3'h7] == 8'h00 & p0_matrix[3'h7][3'h0] == 8'h00 & p0_matrix[3'h7][3'h1] == 8'h00 & p0_matrix[3'h7][3'h2] == 8'h00 & p0_matrix[3'h7][3'h3] == 8'h00 & p0_matrix[3'h7][3'h4] == 8'h00 & p0_matrix[3'h7][3'h5] == 8'h00 & p0_matrix[3'h7][3'h6] == 8'h00 & p0_matrix[3'h7][3'h7] == 8'h00)};
  assign p1_tuple_5071_comb = {p1_concat_5068_comb, 8'h02, p1_code_list_comb & p1_sign_ext_5067_comb};

  // Registers for pipe stage 1:
  reg [31:0] p1_tuple_5071;
  always @ (posedge clk) begin
    p1_tuple_5071 <= p1_tuple_5071_comb;
  end
  assign out = p1_tuple_5071;
endmodule
