module Huffman_ACenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire [7:0] start_pix,
  input wire [7:0] pre_start_pix,
  input wire is_luminance,
  output wire [65:0] out
);
  wire [4:0] literal_12664[0:251];
  assign literal_12664[0] = 5'h02;
  assign literal_12664[1] = 5'h02;
  assign literal_12664[2] = 5'h03;
  assign literal_12664[3] = 5'h04;
  assign literal_12664[4] = 5'h05;
  assign literal_12664[5] = 5'h07;
  assign literal_12664[6] = 5'h08;
  assign literal_12664[7] = 5'h0e;
  assign literal_12664[8] = 5'h10;
  assign literal_12664[9] = 5'h10;
  assign literal_12664[10] = 5'h10;
  assign literal_12664[11] = 5'h00;
  assign literal_12664[12] = 5'h00;
  assign literal_12664[13] = 5'h00;
  assign literal_12664[14] = 5'h00;
  assign literal_12664[15] = 5'h00;
  assign literal_12664[16] = 5'h00;
  assign literal_12664[17] = 5'h03;
  assign literal_12664[18] = 5'h06;
  assign literal_12664[19] = 5'h07;
  assign literal_12664[20] = 5'h09;
  assign literal_12664[21] = 5'h0b;
  assign literal_12664[22] = 5'h0d;
  assign literal_12664[23] = 5'h10;
  assign literal_12664[24] = 5'h10;
  assign literal_12664[25] = 5'h10;
  assign literal_12664[26] = 5'h10;
  assign literal_12664[27] = 5'h00;
  assign literal_12664[28] = 5'h00;
  assign literal_12664[29] = 5'h00;
  assign literal_12664[30] = 5'h00;
  assign literal_12664[31] = 5'h00;
  assign literal_12664[32] = 5'h00;
  assign literal_12664[33] = 5'h05;
  assign literal_12664[34] = 5'h07;
  assign literal_12664[35] = 5'h0a;
  assign literal_12664[36] = 5'h0c;
  assign literal_12664[37] = 5'h0d;
  assign literal_12664[38] = 5'h10;
  assign literal_12664[39] = 5'h10;
  assign literal_12664[40] = 5'h10;
  assign literal_12664[41] = 5'h10;
  assign literal_12664[42] = 5'h10;
  assign literal_12664[43] = 5'h00;
  assign literal_12664[44] = 5'h00;
  assign literal_12664[45] = 5'h00;
  assign literal_12664[46] = 5'h00;
  assign literal_12664[47] = 5'h00;
  assign literal_12664[48] = 5'h00;
  assign literal_12664[49] = 5'h06;
  assign literal_12664[50] = 5'h08;
  assign literal_12664[51] = 5'h0b;
  assign literal_12664[52] = 5'h0c;
  assign literal_12664[53] = 5'h0f;
  assign literal_12664[54] = 5'h10;
  assign literal_12664[55] = 5'h10;
  assign literal_12664[56] = 5'h10;
  assign literal_12664[57] = 5'h10;
  assign literal_12664[58] = 5'h10;
  assign literal_12664[59] = 5'h00;
  assign literal_12664[60] = 5'h00;
  assign literal_12664[61] = 5'h00;
  assign literal_12664[62] = 5'h00;
  assign literal_12664[63] = 5'h00;
  assign literal_12664[64] = 5'h00;
  assign literal_12664[65] = 5'h06;
  assign literal_12664[66] = 5'h0a;
  assign literal_12664[67] = 5'h0c;
  assign literal_12664[68] = 5'h0f;
  assign literal_12664[69] = 5'h10;
  assign literal_12664[70] = 5'h10;
  assign literal_12664[71] = 5'h10;
  assign literal_12664[72] = 5'h10;
  assign literal_12664[73] = 5'h10;
  assign literal_12664[74] = 5'h10;
  assign literal_12664[75] = 5'h00;
  assign literal_12664[76] = 5'h00;
  assign literal_12664[77] = 5'h00;
  assign literal_12664[78] = 5'h00;
  assign literal_12664[79] = 5'h00;
  assign literal_12664[80] = 5'h00;
  assign literal_12664[81] = 5'h07;
  assign literal_12664[82] = 5'h0b;
  assign literal_12664[83] = 5'h0d;
  assign literal_12664[84] = 5'h10;
  assign literal_12664[85] = 5'h10;
  assign literal_12664[86] = 5'h10;
  assign literal_12664[87] = 5'h10;
  assign literal_12664[88] = 5'h10;
  assign literal_12664[89] = 5'h10;
  assign literal_12664[90] = 5'h10;
  assign literal_12664[91] = 5'h00;
  assign literal_12664[92] = 5'h00;
  assign literal_12664[93] = 5'h00;
  assign literal_12664[94] = 5'h00;
  assign literal_12664[95] = 5'h00;
  assign literal_12664[96] = 5'h00;
  assign literal_12664[97] = 5'h07;
  assign literal_12664[98] = 5'h0b;
  assign literal_12664[99] = 5'h0d;
  assign literal_12664[100] = 5'h10;
  assign literal_12664[101] = 5'h10;
  assign literal_12664[102] = 5'h10;
  assign literal_12664[103] = 5'h10;
  assign literal_12664[104] = 5'h10;
  assign literal_12664[105] = 5'h10;
  assign literal_12664[106] = 5'h10;
  assign literal_12664[107] = 5'h00;
  assign literal_12664[108] = 5'h00;
  assign literal_12664[109] = 5'h00;
  assign literal_12664[110] = 5'h00;
  assign literal_12664[111] = 5'h00;
  assign literal_12664[112] = 5'h00;
  assign literal_12664[113] = 5'h08;
  assign literal_12664[114] = 5'h0b;
  assign literal_12664[115] = 5'h0e;
  assign literal_12664[116] = 5'h10;
  assign literal_12664[117] = 5'h10;
  assign literal_12664[118] = 5'h10;
  assign literal_12664[119] = 5'h10;
  assign literal_12664[120] = 5'h10;
  assign literal_12664[121] = 5'h10;
  assign literal_12664[122] = 5'h10;
  assign literal_12664[123] = 5'h00;
  assign literal_12664[124] = 5'h00;
  assign literal_12664[125] = 5'h00;
  assign literal_12664[126] = 5'h00;
  assign literal_12664[127] = 5'h00;
  assign literal_12664[128] = 5'h00;
  assign literal_12664[129] = 5'h08;
  assign literal_12664[130] = 5'h0c;
  assign literal_12664[131] = 5'h10;
  assign literal_12664[132] = 5'h10;
  assign literal_12664[133] = 5'h10;
  assign literal_12664[134] = 5'h10;
  assign literal_12664[135] = 5'h10;
  assign literal_12664[136] = 5'h10;
  assign literal_12664[137] = 5'h10;
  assign literal_12664[138] = 5'h10;
  assign literal_12664[139] = 5'h00;
  assign literal_12664[140] = 5'h00;
  assign literal_12664[141] = 5'h00;
  assign literal_12664[142] = 5'h00;
  assign literal_12664[143] = 5'h00;
  assign literal_12664[144] = 5'h00;
  assign literal_12664[145] = 5'h08;
  assign literal_12664[146] = 5'h0d;
  assign literal_12664[147] = 5'h10;
  assign literal_12664[148] = 5'h10;
  assign literal_12664[149] = 5'h10;
  assign literal_12664[150] = 5'h10;
  assign literal_12664[151] = 5'h10;
  assign literal_12664[152] = 5'h10;
  assign literal_12664[153] = 5'h10;
  assign literal_12664[154] = 5'h10;
  assign literal_12664[155] = 5'h00;
  assign literal_12664[156] = 5'h00;
  assign literal_12664[157] = 5'h00;
  assign literal_12664[158] = 5'h00;
  assign literal_12664[159] = 5'h00;
  assign literal_12664[160] = 5'h00;
  assign literal_12664[161] = 5'h09;
  assign literal_12664[162] = 5'h0d;
  assign literal_12664[163] = 5'h10;
  assign literal_12664[164] = 5'h10;
  assign literal_12664[165] = 5'h10;
  assign literal_12664[166] = 5'h10;
  assign literal_12664[167] = 5'h10;
  assign literal_12664[168] = 5'h10;
  assign literal_12664[169] = 5'h10;
  assign literal_12664[170] = 5'h10;
  assign literal_12664[171] = 5'h00;
  assign literal_12664[172] = 5'h00;
  assign literal_12664[173] = 5'h00;
  assign literal_12664[174] = 5'h00;
  assign literal_12664[175] = 5'h00;
  assign literal_12664[176] = 5'h00;
  assign literal_12664[177] = 5'h09;
  assign literal_12664[178] = 5'h0d;
  assign literal_12664[179] = 5'h10;
  assign literal_12664[180] = 5'h10;
  assign literal_12664[181] = 5'h10;
  assign literal_12664[182] = 5'h10;
  assign literal_12664[183] = 5'h10;
  assign literal_12664[184] = 5'h10;
  assign literal_12664[185] = 5'h10;
  assign literal_12664[186] = 5'h10;
  assign literal_12664[187] = 5'h00;
  assign literal_12664[188] = 5'h00;
  assign literal_12664[189] = 5'h00;
  assign literal_12664[190] = 5'h00;
  assign literal_12664[191] = 5'h00;
  assign literal_12664[192] = 5'h00;
  assign literal_12664[193] = 5'h0a;
  assign literal_12664[194] = 5'h0d;
  assign literal_12664[195] = 5'h10;
  assign literal_12664[196] = 5'h10;
  assign literal_12664[197] = 5'h10;
  assign literal_12664[198] = 5'h10;
  assign literal_12664[199] = 5'h10;
  assign literal_12664[200] = 5'h10;
  assign literal_12664[201] = 5'h10;
  assign literal_12664[202] = 5'h10;
  assign literal_12664[203] = 5'h00;
  assign literal_12664[204] = 5'h00;
  assign literal_12664[205] = 5'h00;
  assign literal_12664[206] = 5'h00;
  assign literal_12664[207] = 5'h00;
  assign literal_12664[208] = 5'h00;
  assign literal_12664[209] = 5'h0a;
  assign literal_12664[210] = 5'h0e;
  assign literal_12664[211] = 5'h10;
  assign literal_12664[212] = 5'h10;
  assign literal_12664[213] = 5'h10;
  assign literal_12664[214] = 5'h10;
  assign literal_12664[215] = 5'h10;
  assign literal_12664[216] = 5'h10;
  assign literal_12664[217] = 5'h10;
  assign literal_12664[218] = 5'h10;
  assign literal_12664[219] = 5'h00;
  assign literal_12664[220] = 5'h00;
  assign literal_12664[221] = 5'h00;
  assign literal_12664[222] = 5'h00;
  assign literal_12664[223] = 5'h00;
  assign literal_12664[224] = 5'h00;
  assign literal_12664[225] = 5'h0a;
  assign literal_12664[226] = 5'h0f;
  assign literal_12664[227] = 5'h10;
  assign literal_12664[228] = 5'h10;
  assign literal_12664[229] = 5'h10;
  assign literal_12664[230] = 5'h10;
  assign literal_12664[231] = 5'h10;
  assign literal_12664[232] = 5'h10;
  assign literal_12664[233] = 5'h10;
  assign literal_12664[234] = 5'h10;
  assign literal_12664[235] = 5'h00;
  assign literal_12664[236] = 5'h00;
  assign literal_12664[237] = 5'h00;
  assign literal_12664[238] = 5'h00;
  assign literal_12664[239] = 5'h00;
  assign literal_12664[240] = 5'h09;
  assign literal_12664[241] = 5'h0b;
  assign literal_12664[242] = 5'h10;
  assign literal_12664[243] = 5'h10;
  assign literal_12664[244] = 5'h10;
  assign literal_12664[245] = 5'h10;
  assign literal_12664[246] = 5'h10;
  assign literal_12664[247] = 5'h10;
  assign literal_12664[248] = 5'h10;
  assign literal_12664[249] = 5'h10;
  assign literal_12664[250] = 5'h10;
  assign literal_12664[251] = 5'h00;
  wire [4:0] literal_12666[0:251];
  assign literal_12666[0] = 5'h04;
  assign literal_12666[1] = 5'h02;
  assign literal_12666[2] = 5'h02;
  assign literal_12666[3] = 5'h03;
  assign literal_12666[4] = 5'h04;
  assign literal_12666[5] = 5'h05;
  assign literal_12666[6] = 5'h07;
  assign literal_12666[7] = 5'h09;
  assign literal_12666[8] = 5'h10;
  assign literal_12666[9] = 5'h10;
  assign literal_12666[10] = 5'h10;
  assign literal_12666[11] = 5'h00;
  assign literal_12666[12] = 5'h00;
  assign literal_12666[13] = 5'h00;
  assign literal_12666[14] = 5'h00;
  assign literal_12666[15] = 5'h00;
  assign literal_12666[16] = 5'h00;
  assign literal_12666[17] = 5'h04;
  assign literal_12666[18] = 5'h05;
  assign literal_12666[19] = 5'h07;
  assign literal_12666[20] = 5'h09;
  assign literal_12666[21] = 5'h0a;
  assign literal_12666[22] = 5'h0b;
  assign literal_12666[23] = 5'h10;
  assign literal_12666[24] = 5'h10;
  assign literal_12666[25] = 5'h10;
  assign literal_12666[26] = 5'h10;
  assign literal_12666[27] = 5'h00;
  assign literal_12666[28] = 5'h00;
  assign literal_12666[29] = 5'h00;
  assign literal_12666[30] = 5'h00;
  assign literal_12666[31] = 5'h00;
  assign literal_12666[32] = 5'h00;
  assign literal_12666[33] = 5'h05;
  assign literal_12666[34] = 5'h08;
  assign literal_12666[35] = 5'h0a;
  assign literal_12666[36] = 5'h0c;
  assign literal_12666[37] = 5'h0e;
  assign literal_12666[38] = 5'h10;
  assign literal_12666[39] = 5'h10;
  assign literal_12666[40] = 5'h10;
  assign literal_12666[41] = 5'h10;
  assign literal_12666[42] = 5'h10;
  assign literal_12666[43] = 5'h00;
  assign literal_12666[44] = 5'h00;
  assign literal_12666[45] = 5'h00;
  assign literal_12666[46] = 5'h00;
  assign literal_12666[47] = 5'h00;
  assign literal_12666[48] = 5'h00;
  assign literal_12666[49] = 5'h06;
  assign literal_12666[50] = 5'h09;
  assign literal_12666[51] = 5'h0b;
  assign literal_12666[52] = 5'h0e;
  assign literal_12666[53] = 5'h10;
  assign literal_12666[54] = 5'h10;
  assign literal_12666[55] = 5'h10;
  assign literal_12666[56] = 5'h10;
  assign literal_12666[57] = 5'h10;
  assign literal_12666[58] = 5'h10;
  assign literal_12666[59] = 5'h00;
  assign literal_12666[60] = 5'h00;
  assign literal_12666[61] = 5'h00;
  assign literal_12666[62] = 5'h00;
  assign literal_12666[63] = 5'h00;
  assign literal_12666[64] = 5'h00;
  assign literal_12666[65] = 5'h06;
  assign literal_12666[66] = 5'h0a;
  assign literal_12666[67] = 5'h0e;
  assign literal_12666[68] = 5'h10;
  assign literal_12666[69] = 5'h10;
  assign literal_12666[70] = 5'h10;
  assign literal_12666[71] = 5'h10;
  assign literal_12666[72] = 5'h10;
  assign literal_12666[73] = 5'h10;
  assign literal_12666[74] = 5'h10;
  assign literal_12666[75] = 5'h00;
  assign literal_12666[76] = 5'h00;
  assign literal_12666[77] = 5'h00;
  assign literal_12666[78] = 5'h00;
  assign literal_12666[79] = 5'h00;
  assign literal_12666[80] = 5'h00;
  assign literal_12666[81] = 5'h07;
  assign literal_12666[82] = 5'h0a;
  assign literal_12666[83] = 5'h0e;
  assign literal_12666[84] = 5'h10;
  assign literal_12666[85] = 5'h10;
  assign literal_12666[86] = 5'h10;
  assign literal_12666[87] = 5'h10;
  assign literal_12666[88] = 5'h10;
  assign literal_12666[89] = 5'h10;
  assign literal_12666[90] = 5'h10;
  assign literal_12666[91] = 5'h00;
  assign literal_12666[92] = 5'h00;
  assign literal_12666[93] = 5'h00;
  assign literal_12666[94] = 5'h00;
  assign literal_12666[95] = 5'h00;
  assign literal_12666[96] = 5'h00;
  assign literal_12666[97] = 5'h07;
  assign literal_12666[98] = 5'h0c;
  assign literal_12666[99] = 5'h0f;
  assign literal_12666[100] = 5'h10;
  assign literal_12666[101] = 5'h10;
  assign literal_12666[102] = 5'h10;
  assign literal_12666[103] = 5'h10;
  assign literal_12666[104] = 5'h10;
  assign literal_12666[105] = 5'h10;
  assign literal_12666[106] = 5'h10;
  assign literal_12666[107] = 5'h00;
  assign literal_12666[108] = 5'h00;
  assign literal_12666[109] = 5'h00;
  assign literal_12666[110] = 5'h00;
  assign literal_12666[111] = 5'h00;
  assign literal_12666[112] = 5'h00;
  assign literal_12666[113] = 5'h08;
  assign literal_12666[114] = 5'h0c;
  assign literal_12666[115] = 5'h10;
  assign literal_12666[116] = 5'h10;
  assign literal_12666[117] = 5'h10;
  assign literal_12666[118] = 5'h10;
  assign literal_12666[119] = 5'h10;
  assign literal_12666[120] = 5'h10;
  assign literal_12666[121] = 5'h10;
  assign literal_12666[122] = 5'h10;
  assign literal_12666[123] = 5'h00;
  assign literal_12666[124] = 5'h00;
  assign literal_12666[125] = 5'h00;
  assign literal_12666[126] = 5'h00;
  assign literal_12666[127] = 5'h00;
  assign literal_12666[128] = 5'h00;
  assign literal_12666[129] = 5'h09;
  assign literal_12666[130] = 5'h0d;
  assign literal_12666[131] = 5'h10;
  assign literal_12666[132] = 5'h10;
  assign literal_12666[133] = 5'h10;
  assign literal_12666[134] = 5'h10;
  assign literal_12666[135] = 5'h10;
  assign literal_12666[136] = 5'h10;
  assign literal_12666[137] = 5'h10;
  assign literal_12666[138] = 5'h10;
  assign literal_12666[139] = 5'h00;
  assign literal_12666[140] = 5'h00;
  assign literal_12666[141] = 5'h00;
  assign literal_12666[142] = 5'h00;
  assign literal_12666[143] = 5'h00;
  assign literal_12666[144] = 5'h00;
  assign literal_12666[145] = 5'h09;
  assign literal_12666[146] = 5'h0e;
  assign literal_12666[147] = 5'h10;
  assign literal_12666[148] = 5'h10;
  assign literal_12666[149] = 5'h10;
  assign literal_12666[150] = 5'h10;
  assign literal_12666[151] = 5'h10;
  assign literal_12666[152] = 5'h10;
  assign literal_12666[153] = 5'h10;
  assign literal_12666[154] = 5'h10;
  assign literal_12666[155] = 5'h00;
  assign literal_12666[156] = 5'h00;
  assign literal_12666[157] = 5'h00;
  assign literal_12666[158] = 5'h00;
  assign literal_12666[159] = 5'h00;
  assign literal_12666[160] = 5'h00;
  assign literal_12666[161] = 5'h09;
  assign literal_12666[162] = 5'h0e;
  assign literal_12666[163] = 5'h10;
  assign literal_12666[164] = 5'h10;
  assign literal_12666[165] = 5'h10;
  assign literal_12666[166] = 5'h10;
  assign literal_12666[167] = 5'h10;
  assign literal_12666[168] = 5'h10;
  assign literal_12666[169] = 5'h10;
  assign literal_12666[170] = 5'h10;
  assign literal_12666[171] = 5'h00;
  assign literal_12666[172] = 5'h00;
  assign literal_12666[173] = 5'h00;
  assign literal_12666[174] = 5'h00;
  assign literal_12666[175] = 5'h00;
  assign literal_12666[176] = 5'h00;
  assign literal_12666[177] = 5'h0a;
  assign literal_12666[178] = 5'h0f;
  assign literal_12666[179] = 5'h10;
  assign literal_12666[180] = 5'h10;
  assign literal_12666[181] = 5'h10;
  assign literal_12666[182] = 5'h10;
  assign literal_12666[183] = 5'h10;
  assign literal_12666[184] = 5'h10;
  assign literal_12666[185] = 5'h10;
  assign literal_12666[186] = 5'h10;
  assign literal_12666[187] = 5'h00;
  assign literal_12666[188] = 5'h00;
  assign literal_12666[189] = 5'h00;
  assign literal_12666[190] = 5'h00;
  assign literal_12666[191] = 5'h00;
  assign literal_12666[192] = 5'h00;
  assign literal_12666[193] = 5'h0a;
  assign literal_12666[194] = 5'h10;
  assign literal_12666[195] = 5'h10;
  assign literal_12666[196] = 5'h10;
  assign literal_12666[197] = 5'h10;
  assign literal_12666[198] = 5'h10;
  assign literal_12666[199] = 5'h10;
  assign literal_12666[200] = 5'h10;
  assign literal_12666[201] = 5'h10;
  assign literal_12666[202] = 5'h10;
  assign literal_12666[203] = 5'h00;
  assign literal_12666[204] = 5'h00;
  assign literal_12666[205] = 5'h00;
  assign literal_12666[206] = 5'h00;
  assign literal_12666[207] = 5'h00;
  assign literal_12666[208] = 5'h00;
  assign literal_12666[209] = 5'h0a;
  assign literal_12666[210] = 5'h10;
  assign literal_12666[211] = 5'h10;
  assign literal_12666[212] = 5'h10;
  assign literal_12666[213] = 5'h10;
  assign literal_12666[214] = 5'h10;
  assign literal_12666[215] = 5'h10;
  assign literal_12666[216] = 5'h10;
  assign literal_12666[217] = 5'h10;
  assign literal_12666[218] = 5'h10;
  assign literal_12666[219] = 5'h00;
  assign literal_12666[220] = 5'h00;
  assign literal_12666[221] = 5'h00;
  assign literal_12666[222] = 5'h00;
  assign literal_12666[223] = 5'h00;
  assign literal_12666[224] = 5'h00;
  assign literal_12666[225] = 5'h0b;
  assign literal_12666[226] = 5'h10;
  assign literal_12666[227] = 5'h10;
  assign literal_12666[228] = 5'h10;
  assign literal_12666[229] = 5'h10;
  assign literal_12666[230] = 5'h10;
  assign literal_12666[231] = 5'h10;
  assign literal_12666[232] = 5'h10;
  assign literal_12666[233] = 5'h10;
  assign literal_12666[234] = 5'h10;
  assign literal_12666[235] = 5'h00;
  assign literal_12666[236] = 5'h00;
  assign literal_12666[237] = 5'h00;
  assign literal_12666[238] = 5'h00;
  assign literal_12666[239] = 5'h00;
  assign literal_12666[240] = 5'h0c;
  assign literal_12666[241] = 5'h0d;
  assign literal_12666[242] = 5'h10;
  assign literal_12666[243] = 5'h10;
  assign literal_12666[244] = 5'h10;
  assign literal_12666[245] = 5'h10;
  assign literal_12666[246] = 5'h10;
  assign literal_12666[247] = 5'h10;
  assign literal_12666[248] = 5'h10;
  assign literal_12666[249] = 5'h10;
  assign literal_12666[250] = 5'h10;
  assign literal_12666[251] = 5'h00;
  wire [15:0] literal_12671[0:251];
  assign literal_12671[0] = 16'h0001;
  assign literal_12671[1] = 16'h0000;
  assign literal_12671[2] = 16'h0004;
  assign literal_12671[3] = 16'h000c;
  assign literal_12671[4] = 16'h001a;
  assign literal_12671[5] = 16'h0076;
  assign literal_12671[6] = 16'h00f6;
  assign literal_12671[7] = 16'h3fe0;
  assign literal_12671[8] = 16'hff96;
  assign literal_12671[9] = 16'hff97;
  assign literal_12671[10] = 16'hff98;
  assign literal_12671[11] = 16'h0000;
  assign literal_12671[12] = 16'h0000;
  assign literal_12671[13] = 16'h0000;
  assign literal_12671[14] = 16'h0000;
  assign literal_12671[15] = 16'h0000;
  assign literal_12671[16] = 16'h0000;
  assign literal_12671[17] = 16'h0005;
  assign literal_12671[18] = 16'h0038;
  assign literal_12671[19] = 16'h0078;
  assign literal_12671[20] = 16'h01f9;
  assign literal_12671[21] = 16'h07f2;
  assign literal_12671[22] = 16'h1fe8;
  assign literal_12671[23] = 16'hff93;
  assign literal_12671[24] = 16'hff99;
  assign literal_12671[25] = 16'hff9a;
  assign literal_12671[26] = 16'hff9e;
  assign literal_12671[27] = 16'h0000;
  assign literal_12671[28] = 16'h0000;
  assign literal_12671[29] = 16'h0000;
  assign literal_12671[30] = 16'h0000;
  assign literal_12671[31] = 16'h0000;
  assign literal_12671[32] = 16'h0000;
  assign literal_12671[33] = 16'h001b;
  assign literal_12671[34] = 16'h007a;
  assign literal_12671[35] = 16'h03f7;
  assign literal_12671[36] = 16'h0ff0;
  assign literal_12671[37] = 16'h1feb;
  assign literal_12671[38] = 16'hff9b;
  assign literal_12671[39] = 16'hff9f;
  assign literal_12671[40] = 16'hffa8;
  assign literal_12671[41] = 16'hffa9;
  assign literal_12671[42] = 16'hfff1;
  assign literal_12671[43] = 16'h0000;
  assign literal_12671[44] = 16'h0000;
  assign literal_12671[45] = 16'h0000;
  assign literal_12671[46] = 16'h0000;
  assign literal_12671[47] = 16'h0000;
  assign literal_12671[48] = 16'h0000;
  assign literal_12671[49] = 16'h0039;
  assign literal_12671[50] = 16'h00fa;
  assign literal_12671[51] = 16'h07f7;
  assign literal_12671[52] = 16'h0ff1;
  assign literal_12671[53] = 16'h7fc6;
  assign literal_12671[54] = 16'hff9c;
  assign literal_12671[55] = 16'hffa3;
  assign literal_12671[56] = 16'hffd7;
  assign literal_12671[57] = 16'hffe4;
  assign literal_12671[58] = 16'hfff2;
  assign literal_12671[59] = 16'h0000;
  assign literal_12671[60] = 16'h0000;
  assign literal_12671[61] = 16'h0000;
  assign literal_12671[62] = 16'h0000;
  assign literal_12671[63] = 16'h0000;
  assign literal_12671[64] = 16'h0000;
  assign literal_12671[65] = 16'h003a;
  assign literal_12671[66] = 16'h03f8;
  assign literal_12671[67] = 16'h0ff2;
  assign literal_12671[68] = 16'h7fc8;
  assign literal_12671[69] = 16'hff9d;
  assign literal_12671[70] = 16'hffbf;
  assign literal_12671[71] = 16'hffcb;
  assign literal_12671[72] = 16'hffd8;
  assign literal_12671[73] = 16'hffe5;
  assign literal_12671[74] = 16'hfff3;
  assign literal_12671[75] = 16'h0000;
  assign literal_12671[76] = 16'h0000;
  assign literal_12671[77] = 16'h0000;
  assign literal_12671[78] = 16'h0000;
  assign literal_12671[79] = 16'h0000;
  assign literal_12671[80] = 16'h0000;
  assign literal_12671[81] = 16'h0077;
  assign literal_12671[82] = 16'h07f3;
  assign literal_12671[83] = 16'h1fea;
  assign literal_12671[84] = 16'hff94;
  assign literal_12671[85] = 16'hffa2;
  assign literal_12671[86] = 16'hffc0;
  assign literal_12671[87] = 16'hffcc;
  assign literal_12671[88] = 16'hffd9;
  assign literal_12671[89] = 16'hffe6;
  assign literal_12671[90] = 16'hfff4;
  assign literal_12671[91] = 16'h0000;
  assign literal_12671[92] = 16'h0000;
  assign literal_12671[93] = 16'h0000;
  assign literal_12671[94] = 16'h0000;
  assign literal_12671[95] = 16'h0000;
  assign literal_12671[96] = 16'h0000;
  assign literal_12671[97] = 16'h0079;
  assign literal_12671[98] = 16'h07f4;
  assign literal_12671[99] = 16'h1fed;
  assign literal_12671[100] = 16'hffa0;
  assign literal_12671[101] = 16'hffb5;
  assign literal_12671[102] = 16'hffc1;
  assign literal_12671[103] = 16'hffcd;
  assign literal_12671[104] = 16'hffda;
  assign literal_12671[105] = 16'hffe7;
  assign literal_12671[106] = 16'hfff5;
  assign literal_12671[107] = 16'h0000;
  assign literal_12671[108] = 16'h0000;
  assign literal_12671[109] = 16'h0000;
  assign literal_12671[110] = 16'h0000;
  assign literal_12671[111] = 16'h0000;
  assign literal_12671[112] = 16'h0000;
  assign literal_12671[113] = 16'h00f7;
  assign literal_12671[114] = 16'h07f5;
  assign literal_12671[115] = 16'h3fe1;
  assign literal_12671[116] = 16'hffa1;
  assign literal_12671[117] = 16'hffb6;
  assign literal_12671[118] = 16'hffc2;
  assign literal_12671[119] = 16'hffce;
  assign literal_12671[120] = 16'hffdb;
  assign literal_12671[121] = 16'hffe8;
  assign literal_12671[122] = 16'hfff6;
  assign literal_12671[123] = 16'h0000;
  assign literal_12671[124] = 16'h0000;
  assign literal_12671[125] = 16'h0000;
  assign literal_12671[126] = 16'h0000;
  assign literal_12671[127] = 16'h0000;
  assign literal_12671[128] = 16'h0000;
  assign literal_12671[129] = 16'h00f8;
  assign literal_12671[130] = 16'h0ff3;
  assign literal_12671[131] = 16'hff92;
  assign literal_12671[132] = 16'hffad;
  assign literal_12671[133] = 16'hffb7;
  assign literal_12671[134] = 16'hffc3;
  assign literal_12671[135] = 16'hffcf;
  assign literal_12671[136] = 16'hffdc;
  assign literal_12671[137] = 16'hffe9;
  assign literal_12671[138] = 16'hfff7;
  assign literal_12671[139] = 16'h0000;
  assign literal_12671[140] = 16'h0000;
  assign literal_12671[141] = 16'h0000;
  assign literal_12671[142] = 16'h0000;
  assign literal_12671[143] = 16'h0000;
  assign literal_12671[144] = 16'h0000;
  assign literal_12671[145] = 16'h00f9;
  assign literal_12671[146] = 16'h1fe9;
  assign literal_12671[147] = 16'hff95;
  assign literal_12671[148] = 16'hffae;
  assign literal_12671[149] = 16'hffb8;
  assign literal_12671[150] = 16'hffc4;
  assign literal_12671[151] = 16'hffd0;
  assign literal_12671[152] = 16'hffdd;
  assign literal_12671[153] = 16'hffea;
  assign literal_12671[154] = 16'hfff8;
  assign literal_12671[155] = 16'h0000;
  assign literal_12671[156] = 16'h0000;
  assign literal_12671[157] = 16'h0000;
  assign literal_12671[158] = 16'h0000;
  assign literal_12671[159] = 16'h0000;
  assign literal_12671[160] = 16'h0000;
  assign literal_12671[161] = 16'h01f6;
  assign literal_12671[162] = 16'h1fec;
  assign literal_12671[163] = 16'hffa5;
  assign literal_12671[164] = 16'hffaf;
  assign literal_12671[165] = 16'hffb9;
  assign literal_12671[166] = 16'hffc5;
  assign literal_12671[167] = 16'hffd1;
  assign literal_12671[168] = 16'hffde;
  assign literal_12671[169] = 16'hffeb;
  assign literal_12671[170] = 16'hfff9;
  assign literal_12671[171] = 16'h0000;
  assign literal_12671[172] = 16'h0000;
  assign literal_12671[173] = 16'h0000;
  assign literal_12671[174] = 16'h0000;
  assign literal_12671[175] = 16'h0000;
  assign literal_12671[176] = 16'h0000;
  assign literal_12671[177] = 16'h01f7;
  assign literal_12671[178] = 16'h1fee;
  assign literal_12671[179] = 16'hffa6;
  assign literal_12671[180] = 16'hffb0;
  assign literal_12671[181] = 16'hffba;
  assign literal_12671[182] = 16'hffc6;
  assign literal_12671[183] = 16'hffd2;
  assign literal_12671[184] = 16'hffdf;
  assign literal_12671[185] = 16'hffec;
  assign literal_12671[186] = 16'hfffa;
  assign literal_12671[187] = 16'h0000;
  assign literal_12671[188] = 16'h0000;
  assign literal_12671[189] = 16'h0000;
  assign literal_12671[190] = 16'h0000;
  assign literal_12671[191] = 16'h0000;
  assign literal_12671[192] = 16'h0000;
  assign literal_12671[193] = 16'h03f4;
  assign literal_12671[194] = 16'h1fef;
  assign literal_12671[195] = 16'hffa7;
  assign literal_12671[196] = 16'hffb1;
  assign literal_12671[197] = 16'hffbb;
  assign literal_12671[198] = 16'hffc7;
  assign literal_12671[199] = 16'hffd3;
  assign literal_12671[200] = 16'hffe0;
  assign literal_12671[201] = 16'hffed;
  assign literal_12671[202] = 16'hfffb;
  assign literal_12671[203] = 16'h0000;
  assign literal_12671[204] = 16'h0000;
  assign literal_12671[205] = 16'h0000;
  assign literal_12671[206] = 16'h0000;
  assign literal_12671[207] = 16'h0000;
  assign literal_12671[208] = 16'h0000;
  assign literal_12671[209] = 16'h03f5;
  assign literal_12671[210] = 16'h3fe2;
  assign literal_12671[211] = 16'hffaa;
  assign literal_12671[212] = 16'hffb2;
  assign literal_12671[213] = 16'hffbc;
  assign literal_12671[214] = 16'hffc8;
  assign literal_12671[215] = 16'hffd4;
  assign literal_12671[216] = 16'hffe1;
  assign literal_12671[217] = 16'hffee;
  assign literal_12671[218] = 16'hfffc;
  assign literal_12671[219] = 16'h0000;
  assign literal_12671[220] = 16'h0000;
  assign literal_12671[221] = 16'h0000;
  assign literal_12671[222] = 16'h0000;
  assign literal_12671[223] = 16'h0000;
  assign literal_12671[224] = 16'h0000;
  assign literal_12671[225] = 16'h03f6;
  assign literal_12671[226] = 16'h7fc7;
  assign literal_12671[227] = 16'hffab;
  assign literal_12671[228] = 16'hffb3;
  assign literal_12671[229] = 16'hffbd;
  assign literal_12671[230] = 16'hffc9;
  assign literal_12671[231] = 16'hffd5;
  assign literal_12671[232] = 16'hffe2;
  assign literal_12671[233] = 16'hffef;
  assign literal_12671[234] = 16'hfffd;
  assign literal_12671[235] = 16'h0000;
  assign literal_12671[236] = 16'h0000;
  assign literal_12671[237] = 16'h0000;
  assign literal_12671[238] = 16'h0000;
  assign literal_12671[239] = 16'h0000;
  assign literal_12671[240] = 16'h01f8;
  assign literal_12671[241] = 16'h07f6;
  assign literal_12671[242] = 16'hffa4;
  assign literal_12671[243] = 16'hffac;
  assign literal_12671[244] = 16'hffb4;
  assign literal_12671[245] = 16'hffbe;
  assign literal_12671[246] = 16'hffca;
  assign literal_12671[247] = 16'hffd6;
  assign literal_12671[248] = 16'hffe3;
  assign literal_12671[249] = 16'hfff0;
  assign literal_12671[250] = 16'hfffe;
  assign literal_12671[251] = 16'h0000;
  wire [15:0] literal_12672[0:251];
  assign literal_12672[0] = 16'h000c;
  assign literal_12672[1] = 16'h0000;
  assign literal_12672[2] = 16'h0001;
  assign literal_12672[3] = 16'h0004;
  assign literal_12672[4] = 16'h000b;
  assign literal_12672[5] = 16'h001a;
  assign literal_12672[6] = 16'h0079;
  assign literal_12672[7] = 16'h01f9;
  assign literal_12672[8] = 16'hff9c;
  assign literal_12672[9] = 16'hff9f;
  assign literal_12672[10] = 16'hffa0;
  assign literal_12672[11] = 16'h0000;
  assign literal_12672[12] = 16'h0000;
  assign literal_12672[13] = 16'h0000;
  assign literal_12672[14] = 16'h0000;
  assign literal_12672[15] = 16'h0000;
  assign literal_12672[16] = 16'h0000;
  assign literal_12672[17] = 16'h000a;
  assign literal_12672[18] = 16'h001c;
  assign literal_12672[19] = 16'h007a;
  assign literal_12672[20] = 16'h01f5;
  assign literal_12672[21] = 16'h03f4;
  assign literal_12672[22] = 16'h07f8;
  assign literal_12672[23] = 16'hff95;
  assign literal_12672[24] = 16'hffa1;
  assign literal_12672[25] = 16'hffa2;
  assign literal_12672[26] = 16'hffad;
  assign literal_12672[27] = 16'h0000;
  assign literal_12672[28] = 16'h0000;
  assign literal_12672[29] = 16'h0000;
  assign literal_12672[30] = 16'h0000;
  assign literal_12672[31] = 16'h0000;
  assign literal_12672[32] = 16'h0000;
  assign literal_12672[33] = 16'h001b;
  assign literal_12672[34] = 16'h00f8;
  assign literal_12672[35] = 16'h03f7;
  assign literal_12672[36] = 16'h0ff4;
  assign literal_12672[37] = 16'h3fdc;
  assign literal_12672[38] = 16'hff9d;
  assign literal_12672[39] = 16'hff90;
  assign literal_12672[40] = 16'hffac;
  assign literal_12672[41] = 16'hffe3;
  assign literal_12672[42] = 16'hfff1;
  assign literal_12672[43] = 16'h0000;
  assign literal_12672[44] = 16'h0000;
  assign literal_12672[45] = 16'h0000;
  assign literal_12672[46] = 16'h0000;
  assign literal_12672[47] = 16'h0000;
  assign literal_12672[48] = 16'h0000;
  assign literal_12672[49] = 16'h003a;
  assign literal_12672[50] = 16'h01f6;
  assign literal_12672[51] = 16'h07f7;
  assign literal_12672[52] = 16'h3fde;
  assign literal_12672[53] = 16'hff8e;
  assign literal_12672[54] = 16'hff94;
  assign literal_12672[55] = 16'hffc9;
  assign literal_12672[56] = 16'hffd6;
  assign literal_12672[57] = 16'hffe4;
  assign literal_12672[58] = 16'hfff2;
  assign literal_12672[59] = 16'h0000;
  assign literal_12672[60] = 16'h0000;
  assign literal_12672[61] = 16'h0000;
  assign literal_12672[62] = 16'h0000;
  assign literal_12672[63] = 16'h0000;
  assign literal_12672[64] = 16'h0000;
  assign literal_12672[65] = 16'h003b;
  assign literal_12672[66] = 16'h03f6;
  assign literal_12672[67] = 16'h3fdd;
  assign literal_12672[68] = 16'hff8f;
  assign literal_12672[69] = 16'hffa5;
  assign literal_12672[70] = 16'hffa6;
  assign literal_12672[71] = 16'hffca;
  assign literal_12672[72] = 16'hffd7;
  assign literal_12672[73] = 16'hffe5;
  assign literal_12672[74] = 16'hfff3;
  assign literal_12672[75] = 16'h0000;
  assign literal_12672[76] = 16'h0000;
  assign literal_12672[77] = 16'h0000;
  assign literal_12672[78] = 16'h0000;
  assign literal_12672[79] = 16'h0000;
  assign literal_12672[80] = 16'h0000;
  assign literal_12672[81] = 16'h0078;
  assign literal_12672[82] = 16'h03f9;
  assign literal_12672[83] = 16'h3fdf;
  assign literal_12672[84] = 16'hff96;
  assign literal_12672[85] = 16'hffab;
  assign literal_12672[86] = 16'hffa9;
  assign literal_12672[87] = 16'hffcb;
  assign literal_12672[88] = 16'hffd8;
  assign literal_12672[89] = 16'hffe6;
  assign literal_12672[90] = 16'hfff4;
  assign literal_12672[91] = 16'h0000;
  assign literal_12672[92] = 16'h0000;
  assign literal_12672[93] = 16'h0000;
  assign literal_12672[94] = 16'h0000;
  assign literal_12672[95] = 16'h0000;
  assign literal_12672[96] = 16'h0000;
  assign literal_12672[97] = 16'h007b;
  assign literal_12672[98] = 16'h0ff2;
  assign literal_12672[99] = 16'h7fc5;
  assign literal_12672[100] = 16'hff97;
  assign literal_12672[101] = 16'hffb5;
  assign literal_12672[102] = 16'hffbf;
  assign literal_12672[103] = 16'hffcc;
  assign literal_12672[104] = 16'hffd9;
  assign literal_12672[105] = 16'hffe7;
  assign literal_12672[106] = 16'hfff5;
  assign literal_12672[107] = 16'h0000;
  assign literal_12672[108] = 16'h0000;
  assign literal_12672[109] = 16'h0000;
  assign literal_12672[110] = 16'h0000;
  assign literal_12672[111] = 16'h0000;
  assign literal_12672[112] = 16'h0000;
  assign literal_12672[113] = 16'h00f9;
  assign literal_12672[114] = 16'h0ff5;
  assign literal_12672[115] = 16'hff8c;
  assign literal_12672[116] = 16'hff98;
  assign literal_12672[117] = 16'hffb6;
  assign literal_12672[118] = 16'hffc0;
  assign literal_12672[119] = 16'hffcd;
  assign literal_12672[120] = 16'hffda;
  assign literal_12672[121] = 16'hffe8;
  assign literal_12672[122] = 16'hfff6;
  assign literal_12672[123] = 16'h0000;
  assign literal_12672[124] = 16'h0000;
  assign literal_12672[125] = 16'h0000;
  assign literal_12672[126] = 16'h0000;
  assign literal_12672[127] = 16'h0000;
  assign literal_12672[128] = 16'h0000;
  assign literal_12672[129] = 16'h01f4;
  assign literal_12672[130] = 16'h1fec;
  assign literal_12672[131] = 16'hff9e;
  assign literal_12672[132] = 16'hffa3;
  assign literal_12672[133] = 16'hffb7;
  assign literal_12672[134] = 16'hffc1;
  assign literal_12672[135] = 16'hffce;
  assign literal_12672[136] = 16'hffdb;
  assign literal_12672[137] = 16'hffe9;
  assign literal_12672[138] = 16'hfff7;
  assign literal_12672[139] = 16'h0000;
  assign literal_12672[140] = 16'h0000;
  assign literal_12672[141] = 16'h0000;
  assign literal_12672[142] = 16'h0000;
  assign literal_12672[143] = 16'h0000;
  assign literal_12672[144] = 16'h0000;
  assign literal_12672[145] = 16'h01f7;
  assign literal_12672[146] = 16'h3fe0;
  assign literal_12672[147] = 16'hff91;
  assign literal_12672[148] = 16'hffa4;
  assign literal_12672[149] = 16'hffb8;
  assign literal_12672[150] = 16'hffc2;
  assign literal_12672[151] = 16'hffcf;
  assign literal_12672[152] = 16'hffdc;
  assign literal_12672[153] = 16'hffea;
  assign literal_12672[154] = 16'hfff8;
  assign literal_12672[155] = 16'h0000;
  assign literal_12672[156] = 16'h0000;
  assign literal_12672[157] = 16'h0000;
  assign literal_12672[158] = 16'h0000;
  assign literal_12672[159] = 16'h0000;
  assign literal_12672[160] = 16'h0000;
  assign literal_12672[161] = 16'h01f8;
  assign literal_12672[162] = 16'h3fe1;
  assign literal_12672[163] = 16'hff92;
  assign literal_12672[164] = 16'hffa7;
  assign literal_12672[165] = 16'hffb9;
  assign literal_12672[166] = 16'hffc3;
  assign literal_12672[167] = 16'hffd0;
  assign literal_12672[168] = 16'hffdd;
  assign literal_12672[169] = 16'hffeb;
  assign literal_12672[170] = 16'hfff9;
  assign literal_12672[171] = 16'h0000;
  assign literal_12672[172] = 16'h0000;
  assign literal_12672[173] = 16'h0000;
  assign literal_12672[174] = 16'h0000;
  assign literal_12672[175] = 16'h0000;
  assign literal_12672[176] = 16'h0000;
  assign literal_12672[177] = 16'h03f5;
  assign literal_12672[178] = 16'h7fc4;
  assign literal_12672[179] = 16'hff93;
  assign literal_12672[180] = 16'hffa8;
  assign literal_12672[181] = 16'hffba;
  assign literal_12672[182] = 16'hffc4;
  assign literal_12672[183] = 16'hffd1;
  assign literal_12672[184] = 16'hffde;
  assign literal_12672[185] = 16'hffec;
  assign literal_12672[186] = 16'hfffa;
  assign literal_12672[187] = 16'h0000;
  assign literal_12672[188] = 16'h0000;
  assign literal_12672[189] = 16'h0000;
  assign literal_12672[190] = 16'h0000;
  assign literal_12672[191] = 16'h0000;
  assign literal_12672[192] = 16'h0000;
  assign literal_12672[193] = 16'h03f8;
  assign literal_12672[194] = 16'hff8d;
  assign literal_12672[195] = 16'hff99;
  assign literal_12672[196] = 16'hffb1;
  assign literal_12672[197] = 16'hffbb;
  assign literal_12672[198] = 16'hffc5;
  assign literal_12672[199] = 16'hffd2;
  assign literal_12672[200] = 16'hffdf;
  assign literal_12672[201] = 16'hffed;
  assign literal_12672[202] = 16'hfffb;
  assign literal_12672[203] = 16'h0000;
  assign literal_12672[204] = 16'h0000;
  assign literal_12672[205] = 16'h0000;
  assign literal_12672[206] = 16'h0000;
  assign literal_12672[207] = 16'h0000;
  assign literal_12672[208] = 16'h0000;
  assign literal_12672[209] = 16'h03fa;
  assign literal_12672[210] = 16'hff9a;
  assign literal_12672[211] = 16'hffaa;
  assign literal_12672[212] = 16'hffb2;
  assign literal_12672[213] = 16'hffbc;
  assign literal_12672[214] = 16'hffc6;
  assign literal_12672[215] = 16'hffd3;
  assign literal_12672[216] = 16'hffe0;
  assign literal_12672[217] = 16'hffee;
  assign literal_12672[218] = 16'hfffc;
  assign literal_12672[219] = 16'h0000;
  assign literal_12672[220] = 16'h0000;
  assign literal_12672[221] = 16'h0000;
  assign literal_12672[222] = 16'h0000;
  assign literal_12672[223] = 16'h0000;
  assign literal_12672[224] = 16'h0000;
  assign literal_12672[225] = 16'h07f6;
  assign literal_12672[226] = 16'hff9b;
  assign literal_12672[227] = 16'hffaf;
  assign literal_12672[228] = 16'hffb3;
  assign literal_12672[229] = 16'hffbd;
  assign literal_12672[230] = 16'hffc7;
  assign literal_12672[231] = 16'hffd4;
  assign literal_12672[232] = 16'hffe1;
  assign literal_12672[233] = 16'hffef;
  assign literal_12672[234] = 16'hfffd;
  assign literal_12672[235] = 16'h0000;
  assign literal_12672[236] = 16'h0000;
  assign literal_12672[237] = 16'h0000;
  assign literal_12672[238] = 16'h0000;
  assign literal_12672[239] = 16'h0000;
  assign literal_12672[240] = 16'h0ff3;
  assign literal_12672[241] = 16'h1fed;
  assign literal_12672[242] = 16'hffae;
  assign literal_12672[243] = 16'hffb0;
  assign literal_12672[244] = 16'hffb4;
  assign literal_12672[245] = 16'hffbe;
  assign literal_12672[246] = 16'hffc8;
  assign literal_12672[247] = 16'hffd5;
  assign literal_12672[248] = 16'hffe2;
  assign literal_12672[249] = 16'hfff0;
  assign literal_12672[250] = 16'hfffe;
  assign literal_12672[251] = 16'h0000;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire p1_next_pix__1_squeezed_squeezed_const_msb_bits_comb;
  wire p1_next_pix__1_squeezed_squeezed_const_msb_bits__5_comb;
  wire [8:0] p1_concat_11197_comb;
  wire [7:0] p1_concat_11199_comb;
  wire [8:0] p1_add_11202_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__16_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__15_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__14_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__13_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__12_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__11_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__10_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__9_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__8_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__7_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__6_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__5_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__4_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__3_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__1_comb;
  wire [2:0] p1_run_0_squeezed_const_msb_bits__2_comb;
  wire [7:0] p1_add_11333_comb;
  wire [9:0] p1_array_index_11336_comb;
  wire [9:0] p1_array_index_11337_comb;
  wire [9:0] p1_array_index_11338_comb;
  wire [9:0] p1_array_index_11339_comb;
  wire [9:0] p1_array_index_11340_comb;
  wire [9:0] p1_array_index_11341_comb;
  wire [9:0] p1_array_index_11342_comb;
  wire [9:0] p1_array_index_11343_comb;
  wire [9:0] p1_array_index_11344_comb;
  wire [9:0] p1_array_index_11345_comb;
  wire [9:0] p1_array_index_11346_comb;
  wire [9:0] p1_array_index_11347_comb;
  wire [9:0] p1_array_index_11348_comb;
  wire [9:0] p1_array_index_11349_comb;
  wire [9:0] p1_array_index_11350_comb;
  wire [9:0] p1_array_index_11351_comb;
  wire [9:0] p1_array_index_11352_comb;
  wire [9:0] p1_array_index_11353_comb;
  wire [9:0] p1_array_index_11354_comb;
  wire [9:0] p1_array_index_11355_comb;
  wire [9:0] p1_array_index_11356_comb;
  wire [9:0] p1_array_index_11357_comb;
  wire [9:0] p1_array_index_11358_comb;
  wire [9:0] p1_array_index_11359_comb;
  wire [9:0] p1_array_index_11360_comb;
  wire [9:0] p1_array_index_11361_comb;
  wire [9:0] p1_array_index_11362_comb;
  wire [9:0] p1_array_index_11363_comb;
  wire [9:0] p1_array_index_11364_comb;
  wire [9:0] p1_array_index_11365_comb;
  wire [9:0] p1_array_index_11366_comb;
  wire [9:0] p1_array_index_11367_comb;
  wire [9:0] p1_array_index_11368_comb;
  wire [9:0] p1_array_index_11369_comb;
  wire [9:0] p1_array_index_11370_comb;
  wire [9:0] p1_array_index_11371_comb;
  wire [9:0] p1_array_index_11372_comb;
  wire [9:0] p1_array_index_11373_comb;
  wire [9:0] p1_array_index_11374_comb;
  wire [9:0] p1_array_index_11375_comb;
  wire [9:0] p1_array_index_11376_comb;
  wire [9:0] p1_array_index_11377_comb;
  wire [9:0] p1_array_index_11378_comb;
  wire [9:0] p1_array_index_11379_comb;
  wire [9:0] p1_array_index_11380_comb;
  wire [9:0] p1_array_index_11381_comb;
  wire [9:0] p1_array_index_11382_comb;
  wire [9:0] p1_array_index_11383_comb;
  wire [9:0] p1_array_index_11384_comb;
  wire [9:0] p1_array_index_11385_comb;
  wire [9:0] p1_array_index_11386_comb;
  wire [9:0] p1_array_index_11387_comb;
  wire [9:0] p1_array_index_11388_comb;
  wire [9:0] p1_array_index_11389_comb;
  wire [9:0] p1_array_index_11390_comb;
  wire [9:0] p1_array_index_11391_comb;
  wire [9:0] p1_array_index_11392_comb;
  wire [9:0] p1_array_index_11393_comb;
  wire [9:0] p1_array_index_11394_comb;
  wire [9:0] p1_array_index_11395_comb;
  wire [9:0] p1_array_index_11396_comb;
  wire [9:0] p1_array_index_11397_comb;
  wire [9:0] p1_array_index_11398_comb;
  wire [9:0] p1_array_index_11399_comb;
  wire [8:0] p1_add_11401_comb;
  wire p1_next_pix__1_squeezed_squeezed_const_msb_bits__6_comb;
  wire [6:0] p1_concat_11409_comb;
  wire [6:0] p1_add_11421_comb;
  wire [8:0] p1_add_11431_comb;
  wire [1:0] p1_concat_11434_comb;
  wire p1_next_pix__1_squeezed_squeezed_const_msb_bits__7_comb;
  wire [7:0] p1_add_11439_comb;
  wire [1:0] p1_sel_11444_comb;
  wire [1:0] p1_sign_ext_11445_comb;
  wire [8:0] p1_add_11447_comb;
  wire [5:0] p1_add_11474_comb;
  wire [8:0] p1_add_11485_comb;
  wire [7:0] p1_add_11493_comb;
  wire [8:0] p1_add_11501_comb;
  wire [6:0] p1_add_11510_comb;
  wire [8:0] p1_add_11520_comb;
  wire [7:0] p1_add_11529_comb;
  wire [8:0] p1_add_11546_comb;
  wire [2:0] p1_sel_11479_comb;
  wire [2:0] p1_sel_11488_comb;
  wire p1_nor_11490_comb;
  wire [2:0] p1_sel_11498_comb;
  wire p1_or_11517_comb;
  wire p1_or_11527_comb;
  wire p1_or_11536_comb;
  wire p1_or_11544_comb;
  wire p1_or_11552_comb;
  wire p1_or_11556_comb;
  wire p1_or_11560_comb;
  wire p1_nor_11563_comb;
  assign p1_next_pix__1_squeezed_squeezed_const_msb_bits_comb = 1'h0;
  assign p1_next_pix__1_squeezed_squeezed_const_msb_bits__5_comb = 1'h0;
  assign p1_concat_11197_comb = {p1_next_pix__1_squeezed_squeezed_const_msb_bits_comb, p0_start_pix};
  assign p1_concat_11199_comb = {p1_next_pix__1_squeezed_squeezed_const_msb_bits__5_comb, p0_start_pix[7:1]};
  assign p1_add_11202_comb = p1_concat_11197_comb + 9'h00f;
  assign p1_run_0_squeezed_const_msb_bits__16_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__15_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__14_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__13_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__12_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__11_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__10_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__9_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__8_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__7_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__6_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__5_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__4_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__3_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__1_comb = 3'h0;
  assign p1_run_0_squeezed_const_msb_bits__2_comb = 3'h0;
  assign p1_add_11333_comb = p1_concat_11199_comb + 8'h07;
  assign p1_array_index_11336_comb = p0_matrix[3'h7][3'h7];
  assign p1_array_index_11337_comb = p0_matrix[3'h7][3'h6];
  assign p1_array_index_11338_comb = p0_matrix[3'h7][3'h5];
  assign p1_array_index_11339_comb = p0_matrix[3'h7][3'h4];
  assign p1_array_index_11340_comb = p0_matrix[3'h7][3'h3];
  assign p1_array_index_11341_comb = p0_matrix[3'h7][3'h2];
  assign p1_array_index_11342_comb = p0_matrix[3'h7][3'h1];
  assign p1_array_index_11343_comb = p0_matrix[3'h7][p1_run_0_squeezed_const_msb_bits__16_comb];
  assign p1_array_index_11344_comb = p0_matrix[3'h6][3'h7];
  assign p1_array_index_11345_comb = p0_matrix[3'h6][3'h6];
  assign p1_array_index_11346_comb = p0_matrix[3'h6][3'h5];
  assign p1_array_index_11347_comb = p0_matrix[3'h6][3'h4];
  assign p1_array_index_11348_comb = p0_matrix[3'h6][3'h3];
  assign p1_array_index_11349_comb = p0_matrix[3'h6][3'h2];
  assign p1_array_index_11350_comb = p0_matrix[3'h6][3'h1];
  assign p1_array_index_11351_comb = p0_matrix[3'h6][p1_run_0_squeezed_const_msb_bits__15_comb];
  assign p1_array_index_11352_comb = p0_matrix[3'h5][3'h7];
  assign p1_array_index_11353_comb = p0_matrix[3'h5][3'h6];
  assign p1_array_index_11354_comb = p0_matrix[3'h5][3'h5];
  assign p1_array_index_11355_comb = p0_matrix[3'h5][3'h4];
  assign p1_array_index_11356_comb = p0_matrix[3'h5][3'h3];
  assign p1_array_index_11357_comb = p0_matrix[3'h5][3'h2];
  assign p1_array_index_11358_comb = p0_matrix[3'h5][3'h1];
  assign p1_array_index_11359_comb = p0_matrix[3'h5][p1_run_0_squeezed_const_msb_bits__14_comb];
  assign p1_array_index_11360_comb = p0_matrix[3'h4][3'h7];
  assign p1_array_index_11361_comb = p0_matrix[3'h4][3'h6];
  assign p1_array_index_11362_comb = p0_matrix[3'h4][3'h5];
  assign p1_array_index_11363_comb = p0_matrix[3'h4][3'h4];
  assign p1_array_index_11364_comb = p0_matrix[3'h4][3'h3];
  assign p1_array_index_11365_comb = p0_matrix[3'h4][3'h2];
  assign p1_array_index_11366_comb = p0_matrix[3'h4][3'h1];
  assign p1_array_index_11367_comb = p0_matrix[3'h4][p1_run_0_squeezed_const_msb_bits__13_comb];
  assign p1_array_index_11368_comb = p0_matrix[3'h3][3'h7];
  assign p1_array_index_11369_comb = p0_matrix[3'h3][3'h6];
  assign p1_array_index_11370_comb = p0_matrix[3'h3][3'h5];
  assign p1_array_index_11371_comb = p0_matrix[3'h3][3'h4];
  assign p1_array_index_11372_comb = p0_matrix[3'h3][3'h3];
  assign p1_array_index_11373_comb = p0_matrix[3'h3][3'h2];
  assign p1_array_index_11374_comb = p0_matrix[3'h3][3'h1];
  assign p1_array_index_11375_comb = p0_matrix[3'h3][p1_run_0_squeezed_const_msb_bits__12_comb];
  assign p1_array_index_11376_comb = p0_matrix[3'h2][3'h7];
  assign p1_array_index_11377_comb = p0_matrix[3'h2][3'h6];
  assign p1_array_index_11378_comb = p0_matrix[3'h2][3'h5];
  assign p1_array_index_11379_comb = p0_matrix[3'h2][3'h4];
  assign p1_array_index_11380_comb = p0_matrix[3'h2][3'h3];
  assign p1_array_index_11381_comb = p0_matrix[3'h2][3'h2];
  assign p1_array_index_11382_comb = p0_matrix[3'h2][3'h1];
  assign p1_array_index_11383_comb = p0_matrix[3'h2][p1_run_0_squeezed_const_msb_bits__11_comb];
  assign p1_array_index_11384_comb = p0_matrix[3'h1][3'h7];
  assign p1_array_index_11385_comb = p0_matrix[3'h1][3'h6];
  assign p1_array_index_11386_comb = p0_matrix[3'h1][3'h5];
  assign p1_array_index_11387_comb = p0_matrix[3'h1][3'h4];
  assign p1_array_index_11388_comb = p0_matrix[3'h1][3'h3];
  assign p1_array_index_11389_comb = p0_matrix[3'h1][3'h2];
  assign p1_array_index_11390_comb = p0_matrix[3'h1][3'h1];
  assign p1_array_index_11391_comb = p0_matrix[3'h1][p1_run_0_squeezed_const_msb_bits__10_comb];
  assign p1_array_index_11392_comb = p0_matrix[p1_run_0_squeezed_const_msb_bits__9_comb][3'h7];
  assign p1_array_index_11393_comb = p0_matrix[p1_run_0_squeezed_const_msb_bits__8_comb][3'h6];
  assign p1_array_index_11394_comb = p0_matrix[p1_run_0_squeezed_const_msb_bits__7_comb][3'h5];
  assign p1_array_index_11395_comb = p0_matrix[p1_run_0_squeezed_const_msb_bits__6_comb][3'h4];
  assign p1_array_index_11396_comb = p0_matrix[p1_run_0_squeezed_const_msb_bits__5_comb][3'h3];
  assign p1_array_index_11397_comb = p0_matrix[p1_run_0_squeezed_const_msb_bits__4_comb][3'h2];
  assign p1_array_index_11398_comb = p0_matrix[p1_run_0_squeezed_const_msb_bits__3_comb][3'h1];
  assign p1_array_index_11399_comb = p0_matrix[p1_run_0_squeezed_const_msb_bits__1_comb][p1_run_0_squeezed_const_msb_bits__2_comb];
  assign p1_add_11401_comb = p1_concat_11197_comb + 9'h00d;
  assign p1_next_pix__1_squeezed_squeezed_const_msb_bits__6_comb = 1'h0;
  assign p1_concat_11409_comb = {p1_next_pix__1_squeezed_squeezed_const_msb_bits__6_comb, p0_start_pix[7:2]};
  assign p1_add_11421_comb = p1_concat_11409_comb + 7'h03;
  assign p1_add_11431_comb = p1_concat_11197_comb + 9'h00b;
  assign p1_concat_11434_comb = {1'h1, ~((|p1_add_11202_comb[8:6]) | ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11202_comb} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000)};
  assign p1_next_pix__1_squeezed_squeezed_const_msb_bits__7_comb = 1'h0;
  assign p1_add_11439_comb = p1_concat_11199_comb + 8'h05;
  assign p1_sel_11444_comb = (|p1_add_11333_comb[7:5]) | ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11333_comb, p0_start_pix[0]} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000 ? 2'h1 : p1_concat_11434_comb;
  assign p1_sign_ext_11445_comb = {2{~((|p1_add_11401_comb[8:6]) | ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11401_comb} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000)}};
  assign p1_add_11447_comb = p1_concat_11197_comb + 9'h009;
  assign p1_add_11474_comb = {p1_next_pix__1_squeezed_squeezed_const_msb_bits__7_comb, p0_start_pix[7:3]} + 6'h01;
  assign p1_add_11485_comb = p1_concat_11197_comb + 9'h007;
  assign p1_add_11493_comb = p1_concat_11199_comb + 8'h03;
  assign p1_add_11501_comb = p1_concat_11197_comb + 9'h005;
  assign p1_add_11510_comb = p1_concat_11409_comb + 7'h01;
  assign p1_add_11520_comb = p1_concat_11197_comb + 9'h003;
  assign p1_add_11529_comb = p1_concat_11199_comb + 8'h01;
  assign p1_add_11546_comb = p1_concat_11197_comb + 9'h001;
  assign p1_sel_11479_comb = (|p1_add_11421_comb[6:4]) | ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11421_comb, p0_start_pix[1:0]} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000 ? 3'h3 : {1'h1, p1_sel_11444_comb & p1_sign_ext_11445_comb};
  assign p1_sel_11488_comb = (|p1_add_11431_comb[8:6]) | ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11431_comb} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000 ? 3'h2 : p1_sel_11479_comb;
  assign p1_nor_11490_comb = ~((|p1_add_11447_comb[8:6]) | ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11447_comb} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000);
  assign p1_sel_11498_comb = (|p1_add_11439_comb[7:5]) | ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11439_comb, p0_start_pix[0]} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000 ? 3'h1 : p1_sel_11488_comb;
  assign p1_or_11517_comb = (|p1_add_11474_comb[5:3]) | ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11474_comb, p0_start_pix[2:0]} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_11527_comb = (|p1_add_11485_comb[8:6]) | ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11485_comb} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_11536_comb = (|p1_add_11493_comb[7:5]) | ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11493_comb, p0_start_pix[0]} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_11544_comb = (|p1_add_11501_comb[8:6]) | ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11501_comb} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_11552_comb = (|p1_add_11510_comb[6:4]) | ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11510_comb, p0_start_pix[1:0]} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_11556_comb = (|p1_add_11520_comb[8:6]) | ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11520_comb} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_11560_comb = (|p1_add_11529_comb[7:5]) | ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11529_comb, p0_start_pix[0]} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_nor_11563_comb = ~(p1_add_11546_comb > 9'h03e | ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0000 ? p1_array_index_11336_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0001 ? p1_array_index_11337_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0002 ? p1_array_index_11338_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0003 ? p1_array_index_11339_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0004 ? p1_array_index_11340_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0005 ? p1_array_index_11341_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0006 ? p1_array_index_11342_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0007 ? p1_array_index_11343_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0008 ? p1_array_index_11344_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0009 ? p1_array_index_11345_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_000a ? p1_array_index_11346_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_000b ? p1_array_index_11347_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_000c ? p1_array_index_11348_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_000d ? p1_array_index_11349_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_000e ? p1_array_index_11350_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_000f ? p1_array_index_11351_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0010 ? p1_array_index_11352_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0011 ? p1_array_index_11353_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0012 ? p1_array_index_11354_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0013 ? p1_array_index_11355_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0014 ? p1_array_index_11356_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0015 ? p1_array_index_11357_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0016 ? p1_array_index_11358_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0017 ? p1_array_index_11359_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0018 ? p1_array_index_11360_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0019 ? p1_array_index_11361_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_001a ? p1_array_index_11362_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_001b ? p1_array_index_11363_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_001c ? p1_array_index_11364_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_001d ? p1_array_index_11365_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_001e ? p1_array_index_11366_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_001f ? p1_array_index_11367_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0020 ? p1_array_index_11368_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0021 ? p1_array_index_11369_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0022 ? p1_array_index_11370_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0023 ? p1_array_index_11371_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0024 ? p1_array_index_11372_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0025 ? p1_array_index_11373_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0026 ? p1_array_index_11374_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0027 ? p1_array_index_11375_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0028 ? p1_array_index_11376_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0029 ? p1_array_index_11377_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_002a ? p1_array_index_11378_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_002b ? p1_array_index_11379_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_002c ? p1_array_index_11380_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_002d ? p1_array_index_11381_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_002e ? p1_array_index_11382_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_002f ? p1_array_index_11383_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0030 ? p1_array_index_11384_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0031 ? p1_array_index_11385_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0032 ? p1_array_index_11386_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0033 ? p1_array_index_11387_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0034 ? p1_array_index_11388_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0035 ? p1_array_index_11389_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0036 ? p1_array_index_11390_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0037 ? p1_array_index_11391_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0038 ? p1_array_index_11392_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_0039 ? p1_array_index_11393_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_003a ? p1_array_index_11394_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_003b ? p1_array_index_11395_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_003c ? p1_array_index_11396_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_003d ? p1_array_index_11397_comb : ({23'h00_0000, p1_add_11546_comb} == 32'h0000_003e ? p1_array_index_11398_comb : p1_array_index_11399_comb))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000);

  // Registers for pipe stage 1:
  reg [7:0] p1_start_pix;
  reg p1_is_luminance;
  reg [9:0] p1_array_index_11336;
  reg [9:0] p1_array_index_11337;
  reg [9:0] p1_array_index_11338;
  reg [9:0] p1_array_index_11339;
  reg [9:0] p1_array_index_11340;
  reg [9:0] p1_array_index_11341;
  reg [9:0] p1_array_index_11342;
  reg [9:0] p1_array_index_11343;
  reg [9:0] p1_array_index_11344;
  reg [9:0] p1_array_index_11345;
  reg [9:0] p1_array_index_11346;
  reg [9:0] p1_array_index_11347;
  reg [9:0] p1_array_index_11348;
  reg [9:0] p1_array_index_11349;
  reg [9:0] p1_array_index_11350;
  reg [9:0] p1_array_index_11351;
  reg [9:0] p1_array_index_11352;
  reg [9:0] p1_array_index_11353;
  reg [9:0] p1_array_index_11354;
  reg [9:0] p1_array_index_11355;
  reg [9:0] p1_array_index_11356;
  reg [9:0] p1_array_index_11357;
  reg [9:0] p1_array_index_11358;
  reg [9:0] p1_array_index_11359;
  reg [9:0] p1_array_index_11360;
  reg [9:0] p1_array_index_11361;
  reg [9:0] p1_array_index_11362;
  reg [9:0] p1_array_index_11363;
  reg [9:0] p1_array_index_11364;
  reg [9:0] p1_array_index_11365;
  reg [9:0] p1_array_index_11366;
  reg [9:0] p1_array_index_11367;
  reg [9:0] p1_array_index_11368;
  reg [9:0] p1_array_index_11369;
  reg [9:0] p1_array_index_11370;
  reg [9:0] p1_array_index_11371;
  reg [9:0] p1_array_index_11372;
  reg [9:0] p1_array_index_11373;
  reg [9:0] p1_array_index_11374;
  reg [9:0] p1_array_index_11375;
  reg [9:0] p1_array_index_11376;
  reg [9:0] p1_array_index_11377;
  reg [9:0] p1_array_index_11378;
  reg [9:0] p1_array_index_11379;
  reg [9:0] p1_array_index_11380;
  reg [9:0] p1_array_index_11381;
  reg [9:0] p1_array_index_11382;
  reg [9:0] p1_array_index_11383;
  reg [9:0] p1_array_index_11384;
  reg [9:0] p1_array_index_11385;
  reg [9:0] p1_array_index_11386;
  reg [9:0] p1_array_index_11387;
  reg [9:0] p1_array_index_11388;
  reg [9:0] p1_array_index_11389;
  reg [9:0] p1_array_index_11390;
  reg [9:0] p1_array_index_11391;
  reg [9:0] p1_array_index_11392;
  reg [9:0] p1_array_index_11393;
  reg [9:0] p1_array_index_11394;
  reg [9:0] p1_array_index_11395;
  reg [9:0] p1_array_index_11396;
  reg [9:0] p1_array_index_11397;
  reg [9:0] p1_array_index_11398;
  reg [9:0] p1_array_index_11399;
  reg p1_nor_11490;
  reg [2:0] p1_sel_11498;
  reg p1_or_11517;
  reg p1_or_11527;
  reg p1_or_11536;
  reg p1_or_11544;
  reg p1_or_11552;
  reg p1_or_11556;
  reg p1_or_11560;
  reg p1_nor_11563;
  always @ (posedge clk) begin
    p1_start_pix <= p0_start_pix;
    p1_is_luminance <= p0_is_luminance;
    p1_array_index_11336 <= p1_array_index_11336_comb;
    p1_array_index_11337 <= p1_array_index_11337_comb;
    p1_array_index_11338 <= p1_array_index_11338_comb;
    p1_array_index_11339 <= p1_array_index_11339_comb;
    p1_array_index_11340 <= p1_array_index_11340_comb;
    p1_array_index_11341 <= p1_array_index_11341_comb;
    p1_array_index_11342 <= p1_array_index_11342_comb;
    p1_array_index_11343 <= p1_array_index_11343_comb;
    p1_array_index_11344 <= p1_array_index_11344_comb;
    p1_array_index_11345 <= p1_array_index_11345_comb;
    p1_array_index_11346 <= p1_array_index_11346_comb;
    p1_array_index_11347 <= p1_array_index_11347_comb;
    p1_array_index_11348 <= p1_array_index_11348_comb;
    p1_array_index_11349 <= p1_array_index_11349_comb;
    p1_array_index_11350 <= p1_array_index_11350_comb;
    p1_array_index_11351 <= p1_array_index_11351_comb;
    p1_array_index_11352 <= p1_array_index_11352_comb;
    p1_array_index_11353 <= p1_array_index_11353_comb;
    p1_array_index_11354 <= p1_array_index_11354_comb;
    p1_array_index_11355 <= p1_array_index_11355_comb;
    p1_array_index_11356 <= p1_array_index_11356_comb;
    p1_array_index_11357 <= p1_array_index_11357_comb;
    p1_array_index_11358 <= p1_array_index_11358_comb;
    p1_array_index_11359 <= p1_array_index_11359_comb;
    p1_array_index_11360 <= p1_array_index_11360_comb;
    p1_array_index_11361 <= p1_array_index_11361_comb;
    p1_array_index_11362 <= p1_array_index_11362_comb;
    p1_array_index_11363 <= p1_array_index_11363_comb;
    p1_array_index_11364 <= p1_array_index_11364_comb;
    p1_array_index_11365 <= p1_array_index_11365_comb;
    p1_array_index_11366 <= p1_array_index_11366_comb;
    p1_array_index_11367 <= p1_array_index_11367_comb;
    p1_array_index_11368 <= p1_array_index_11368_comb;
    p1_array_index_11369 <= p1_array_index_11369_comb;
    p1_array_index_11370 <= p1_array_index_11370_comb;
    p1_array_index_11371 <= p1_array_index_11371_comb;
    p1_array_index_11372 <= p1_array_index_11372_comb;
    p1_array_index_11373 <= p1_array_index_11373_comb;
    p1_array_index_11374 <= p1_array_index_11374_comb;
    p1_array_index_11375 <= p1_array_index_11375_comb;
    p1_array_index_11376 <= p1_array_index_11376_comb;
    p1_array_index_11377 <= p1_array_index_11377_comb;
    p1_array_index_11378 <= p1_array_index_11378_comb;
    p1_array_index_11379 <= p1_array_index_11379_comb;
    p1_array_index_11380 <= p1_array_index_11380_comb;
    p1_array_index_11381 <= p1_array_index_11381_comb;
    p1_array_index_11382 <= p1_array_index_11382_comb;
    p1_array_index_11383 <= p1_array_index_11383_comb;
    p1_array_index_11384 <= p1_array_index_11384_comb;
    p1_array_index_11385 <= p1_array_index_11385_comb;
    p1_array_index_11386 <= p1_array_index_11386_comb;
    p1_array_index_11387 <= p1_array_index_11387_comb;
    p1_array_index_11388 <= p1_array_index_11388_comb;
    p1_array_index_11389 <= p1_array_index_11389_comb;
    p1_array_index_11390 <= p1_array_index_11390_comb;
    p1_array_index_11391 <= p1_array_index_11391_comb;
    p1_array_index_11392 <= p1_array_index_11392_comb;
    p1_array_index_11393 <= p1_array_index_11393_comb;
    p1_array_index_11394 <= p1_array_index_11394_comb;
    p1_array_index_11395 <= p1_array_index_11395_comb;
    p1_array_index_11396 <= p1_array_index_11396_comb;
    p1_array_index_11397 <= p1_array_index_11397_comb;
    p1_array_index_11398 <= p1_array_index_11398_comb;
    p1_array_index_11399 <= p1_array_index_11399_comb;
    p1_nor_11490 <= p1_nor_11490_comb;
    p1_sel_11498 <= p1_sel_11498_comb;
    p1_or_11517 <= p1_or_11517_comb;
    p1_or_11527 <= p1_or_11527_comb;
    p1_or_11536 <= p1_or_11536_comb;
    p1_or_11544 <= p1_or_11544_comb;
    p1_or_11552 <= p1_or_11552_comb;
    p1_or_11556 <= p1_or_11556_comb;
    p1_or_11560 <= p1_or_11560_comb;
    p1_nor_11563 <= p1_nor_11563_comb;
  end

  // ===== Pipe stage 2:
  wire [3:0] p2_sel_11725_comb;
  wire p2_next_pix__1_squeezed_squeezed_const_msb_bits__4_comb;
  wire [4:0] p2_concat_11736_comb;
  wire [4:0] p2_zero_num__1_comb;
  wire [4:0] p2_add_11743_comb;
  wire p2_eq_11744_comb;
  assign p2_sel_11725_comb = p1_or_11536 ? 4'h5 : (p1_or_11527 ? 4'h6 : (p1_or_11517 ? 4'h7 : {1'h1, p1_sel_11498 & {3{p1_nor_11490}}}));
  assign p2_next_pix__1_squeezed_squeezed_const_msb_bits__4_comb = 1'h0;
  assign p2_concat_11736_comb = {p2_next_pix__1_squeezed_squeezed_const_msb_bits__4_comb, p1_or_11560 ? 4'h1 : (p1_or_11556 ? 4'h2 : (p1_or_11552 ? 4'h3 : (p1_or_11544 ? 4'h4 : p2_sel_11725_comb)))};
  assign p2_zero_num__1_comb = p2_concat_11736_comb & {5{p1_nor_11563}};
  assign p2_add_11743_comb = p2_zero_num__1_comb + 5'h01;
  assign p2_eq_11744_comb = ({24'h00_0000, p1_start_pix} == 32'h0000_0000 ? p1_array_index_11336 : ({24'h00_0000, p1_start_pix} == 32'h0000_0001 ? p1_array_index_11337 : ({24'h00_0000, p1_start_pix} == 32'h0000_0002 ? p1_array_index_11338 : ({24'h00_0000, p1_start_pix} == 32'h0000_0003 ? p1_array_index_11339 : ({24'h00_0000, p1_start_pix} == 32'h0000_0004 ? p1_array_index_11340 : ({24'h00_0000, p1_start_pix} == 32'h0000_0005 ? p1_array_index_11341 : ({24'h00_0000, p1_start_pix} == 32'h0000_0006 ? p1_array_index_11342 : ({24'h00_0000, p1_start_pix} == 32'h0000_0007 ? p1_array_index_11343 : ({24'h00_0000, p1_start_pix} == 32'h0000_0008 ? p1_array_index_11344 : ({24'h00_0000, p1_start_pix} == 32'h0000_0009 ? p1_array_index_11345 : ({24'h00_0000, p1_start_pix} == 32'h0000_000a ? p1_array_index_11346 : ({24'h00_0000, p1_start_pix} == 32'h0000_000b ? p1_array_index_11347 : ({24'h00_0000, p1_start_pix} == 32'h0000_000c ? p1_array_index_11348 : ({24'h00_0000, p1_start_pix} == 32'h0000_000d ? p1_array_index_11349 : ({24'h00_0000, p1_start_pix} == 32'h0000_000e ? p1_array_index_11350 : ({24'h00_0000, p1_start_pix} == 32'h0000_000f ? p1_array_index_11351 : ({24'h00_0000, p1_start_pix} == 32'h0000_0010 ? p1_array_index_11352 : ({24'h00_0000, p1_start_pix} == 32'h0000_0011 ? p1_array_index_11353 : ({24'h00_0000, p1_start_pix} == 32'h0000_0012 ? p1_array_index_11354 : ({24'h00_0000, p1_start_pix} == 32'h0000_0013 ? p1_array_index_11355 : ({24'h00_0000, p1_start_pix} == 32'h0000_0014 ? p1_array_index_11356 : ({24'h00_0000, p1_start_pix} == 32'h0000_0015 ? p1_array_index_11357 : ({24'h00_0000, p1_start_pix} == 32'h0000_0016 ? p1_array_index_11358 : ({24'h00_0000, p1_start_pix} == 32'h0000_0017 ? p1_array_index_11359 : ({24'h00_0000, p1_start_pix} == 32'h0000_0018 ? p1_array_index_11360 : ({24'h00_0000, p1_start_pix} == 32'h0000_0019 ? p1_array_index_11361 : ({24'h00_0000, p1_start_pix} == 32'h0000_001a ? p1_array_index_11362 : ({24'h00_0000, p1_start_pix} == 32'h0000_001b ? p1_array_index_11363 : ({24'h00_0000, p1_start_pix} == 32'h0000_001c ? p1_array_index_11364 : ({24'h00_0000, p1_start_pix} == 32'h0000_001d ? p1_array_index_11365 : ({24'h00_0000, p1_start_pix} == 32'h0000_001e ? p1_array_index_11366 : ({24'h00_0000, p1_start_pix} == 32'h0000_001f ? p1_array_index_11367 : ({24'h00_0000, p1_start_pix} == 32'h0000_0020 ? p1_array_index_11368 : ({24'h00_0000, p1_start_pix} == 32'h0000_0021 ? p1_array_index_11369 : ({24'h00_0000, p1_start_pix} == 32'h0000_0022 ? p1_array_index_11370 : ({24'h00_0000, p1_start_pix} == 32'h0000_0023 ? p1_array_index_11371 : ({24'h00_0000, p1_start_pix} == 32'h0000_0024 ? p1_array_index_11372 : ({24'h00_0000, p1_start_pix} == 32'h0000_0025 ? p1_array_index_11373 : ({24'h00_0000, p1_start_pix} == 32'h0000_0026 ? p1_array_index_11374 : ({24'h00_0000, p1_start_pix} == 32'h0000_0027 ? p1_array_index_11375 : ({24'h00_0000, p1_start_pix} == 32'h0000_0028 ? p1_array_index_11376 : ({24'h00_0000, p1_start_pix} == 32'h0000_0029 ? p1_array_index_11377 : ({24'h00_0000, p1_start_pix} == 32'h0000_002a ? p1_array_index_11378 : ({24'h00_0000, p1_start_pix} == 32'h0000_002b ? p1_array_index_11379 : ({24'h00_0000, p1_start_pix} == 32'h0000_002c ? p1_array_index_11380 : ({24'h00_0000, p1_start_pix} == 32'h0000_002d ? p1_array_index_11381 : ({24'h00_0000, p1_start_pix} == 32'h0000_002e ? p1_array_index_11382 : ({24'h00_0000, p1_start_pix} == 32'h0000_002f ? p1_array_index_11383 : ({24'h00_0000, p1_start_pix} == 32'h0000_0030 ? p1_array_index_11384 : ({24'h00_0000, p1_start_pix} == 32'h0000_0031 ? p1_array_index_11385 : ({24'h00_0000, p1_start_pix} == 32'h0000_0032 ? p1_array_index_11386 : ({24'h00_0000, p1_start_pix} == 32'h0000_0033 ? p1_array_index_11387 : ({24'h00_0000, p1_start_pix} == 32'h0000_0034 ? p1_array_index_11388 : ({24'h00_0000, p1_start_pix} == 32'h0000_0035 ? p1_array_index_11389 : ({24'h00_0000, p1_start_pix} == 32'h0000_0036 ? p1_array_index_11390 : ({24'h00_0000, p1_start_pix} == 32'h0000_0037 ? p1_array_index_11391 : ({24'h00_0000, p1_start_pix} == 32'h0000_0038 ? p1_array_index_11392 : ({24'h00_0000, p1_start_pix} == 32'h0000_0039 ? p1_array_index_11393 : ({24'h00_0000, p1_start_pix} == 32'h0000_003a ? p1_array_index_11394 : ({24'h00_0000, p1_start_pix} == 32'h0000_003b ? p1_array_index_11395 : ({24'h00_0000, p1_start_pix} == 32'h0000_003c ? p1_array_index_11396 : ({24'h00_0000, p1_start_pix} == 32'h0000_003d ? p1_array_index_11397 : ({24'h00_0000, p1_start_pix} == 32'h0000_003e ? p1_array_index_11398 : p1_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) == 10'h000;

  // Registers for pipe stage 2:
  reg [7:0] p2_start_pix;
  reg p2_is_luminance;
  reg [9:0] p2_array_index_11336;
  reg [9:0] p2_array_index_11337;
  reg [9:0] p2_array_index_11338;
  reg [9:0] p2_array_index_11339;
  reg [9:0] p2_array_index_11340;
  reg [9:0] p2_array_index_11341;
  reg [9:0] p2_array_index_11342;
  reg [9:0] p2_array_index_11343;
  reg [9:0] p2_array_index_11344;
  reg [9:0] p2_array_index_11345;
  reg [9:0] p2_array_index_11346;
  reg [9:0] p2_array_index_11347;
  reg [9:0] p2_array_index_11348;
  reg [9:0] p2_array_index_11349;
  reg [9:0] p2_array_index_11350;
  reg [9:0] p2_array_index_11351;
  reg [9:0] p2_array_index_11352;
  reg [9:0] p2_array_index_11353;
  reg [9:0] p2_array_index_11354;
  reg [9:0] p2_array_index_11355;
  reg [9:0] p2_array_index_11356;
  reg [9:0] p2_array_index_11357;
  reg [9:0] p2_array_index_11358;
  reg [9:0] p2_array_index_11359;
  reg [9:0] p2_array_index_11360;
  reg [9:0] p2_array_index_11361;
  reg [9:0] p2_array_index_11362;
  reg [9:0] p2_array_index_11363;
  reg [9:0] p2_array_index_11364;
  reg [9:0] p2_array_index_11365;
  reg [9:0] p2_array_index_11366;
  reg [9:0] p2_array_index_11367;
  reg [9:0] p2_array_index_11368;
  reg [9:0] p2_array_index_11369;
  reg [9:0] p2_array_index_11370;
  reg [9:0] p2_array_index_11371;
  reg [9:0] p2_array_index_11372;
  reg [9:0] p2_array_index_11373;
  reg [9:0] p2_array_index_11374;
  reg [9:0] p2_array_index_11375;
  reg [9:0] p2_array_index_11376;
  reg [9:0] p2_array_index_11377;
  reg [9:0] p2_array_index_11378;
  reg [9:0] p2_array_index_11379;
  reg [9:0] p2_array_index_11380;
  reg [9:0] p2_array_index_11381;
  reg [9:0] p2_array_index_11382;
  reg [9:0] p2_array_index_11383;
  reg [9:0] p2_array_index_11384;
  reg [9:0] p2_array_index_11385;
  reg [9:0] p2_array_index_11386;
  reg [9:0] p2_array_index_11387;
  reg [9:0] p2_array_index_11388;
  reg [9:0] p2_array_index_11389;
  reg [9:0] p2_array_index_11390;
  reg [9:0] p2_array_index_11391;
  reg [9:0] p2_array_index_11392;
  reg [9:0] p2_array_index_11393;
  reg [9:0] p2_array_index_11394;
  reg [9:0] p2_array_index_11395;
  reg [9:0] p2_array_index_11396;
  reg [9:0] p2_array_index_11397;
  reg [9:0] p2_array_index_11398;
  reg [9:0] p2_array_index_11399;
  reg [4:0] p2_add_11743;
  reg p2_eq_11744;
  always @ (posedge clk) begin
    p2_start_pix <= p1_start_pix;
    p2_is_luminance <= p1_is_luminance;
    p2_array_index_11336 <= p1_array_index_11336;
    p2_array_index_11337 <= p1_array_index_11337;
    p2_array_index_11338 <= p1_array_index_11338;
    p2_array_index_11339 <= p1_array_index_11339;
    p2_array_index_11340 <= p1_array_index_11340;
    p2_array_index_11341 <= p1_array_index_11341;
    p2_array_index_11342 <= p1_array_index_11342;
    p2_array_index_11343 <= p1_array_index_11343;
    p2_array_index_11344 <= p1_array_index_11344;
    p2_array_index_11345 <= p1_array_index_11345;
    p2_array_index_11346 <= p1_array_index_11346;
    p2_array_index_11347 <= p1_array_index_11347;
    p2_array_index_11348 <= p1_array_index_11348;
    p2_array_index_11349 <= p1_array_index_11349;
    p2_array_index_11350 <= p1_array_index_11350;
    p2_array_index_11351 <= p1_array_index_11351;
    p2_array_index_11352 <= p1_array_index_11352;
    p2_array_index_11353 <= p1_array_index_11353;
    p2_array_index_11354 <= p1_array_index_11354;
    p2_array_index_11355 <= p1_array_index_11355;
    p2_array_index_11356 <= p1_array_index_11356;
    p2_array_index_11357 <= p1_array_index_11357;
    p2_array_index_11358 <= p1_array_index_11358;
    p2_array_index_11359 <= p1_array_index_11359;
    p2_array_index_11360 <= p1_array_index_11360;
    p2_array_index_11361 <= p1_array_index_11361;
    p2_array_index_11362 <= p1_array_index_11362;
    p2_array_index_11363 <= p1_array_index_11363;
    p2_array_index_11364 <= p1_array_index_11364;
    p2_array_index_11365 <= p1_array_index_11365;
    p2_array_index_11366 <= p1_array_index_11366;
    p2_array_index_11367 <= p1_array_index_11367;
    p2_array_index_11368 <= p1_array_index_11368;
    p2_array_index_11369 <= p1_array_index_11369;
    p2_array_index_11370 <= p1_array_index_11370;
    p2_array_index_11371 <= p1_array_index_11371;
    p2_array_index_11372 <= p1_array_index_11372;
    p2_array_index_11373 <= p1_array_index_11373;
    p2_array_index_11374 <= p1_array_index_11374;
    p2_array_index_11375 <= p1_array_index_11375;
    p2_array_index_11376 <= p1_array_index_11376;
    p2_array_index_11377 <= p1_array_index_11377;
    p2_array_index_11378 <= p1_array_index_11378;
    p2_array_index_11379 <= p1_array_index_11379;
    p2_array_index_11380 <= p1_array_index_11380;
    p2_array_index_11381 <= p1_array_index_11381;
    p2_array_index_11382 <= p1_array_index_11382;
    p2_array_index_11383 <= p1_array_index_11383;
    p2_array_index_11384 <= p1_array_index_11384;
    p2_array_index_11385 <= p1_array_index_11385;
    p2_array_index_11386 <= p1_array_index_11386;
    p2_array_index_11387 <= p1_array_index_11387;
    p2_array_index_11388 <= p1_array_index_11388;
    p2_array_index_11389 <= p1_array_index_11389;
    p2_array_index_11390 <= p1_array_index_11390;
    p2_array_index_11391 <= p1_array_index_11391;
    p2_array_index_11392 <= p1_array_index_11392;
    p2_array_index_11393 <= p1_array_index_11393;
    p2_array_index_11394 <= p1_array_index_11394;
    p2_array_index_11395 <= p1_array_index_11395;
    p2_array_index_11396 <= p1_array_index_11396;
    p2_array_index_11397 <= p1_array_index_11397;
    p2_array_index_11398 <= p1_array_index_11398;
    p2_array_index_11399 <= p1_array_index_11399;
    p2_add_11743 <= p2_add_11743_comb;
    p2_eq_11744 <= p2_eq_11744_comb;
  end

  // ===== Pipe stage 3:
  wire [2:0] p3_run_0_squeezed_const_msb_bits_comb;
  wire [7:0] p3_value_pix_num_comb;
  wire [7:0] p3_start_pix_1__1_comb;
  wire [7:0] p3_add_11885_comb;
  wire [9:0] p3_value__1_comb;
  wire [7:0] p3_actual_index__65_comb;
  wire [6:0] p3_add_11988_comb;
  wire [7:0] p3_actual_index__67_comb;
  wire [5:0] p3_add_11990_comb;
  wire [7:0] p3_actual_index__69_comb;
  wire [6:0] p3_add_11992_comb;
  wire [7:0] p3_actual_index__71_comb;
  wire [4:0] p3_add_11994_comb;
  wire [7:0] p3_actual_index__73_comb;
  wire [6:0] p3_add_11996_comb;
  wire [7:0] p3_actual_index__75_comb;
  wire [5:0] p3_add_11998_comb;
  wire [7:0] p3_actual_index__77_comb;
  wire [6:0] p3_add_12000_comb;
  wire [7:0] p3_actual_index__79_comb;
  wire [3:0] p3_add_12002_comb;
  wire [7:0] p3_actual_index__81_comb;
  wire [6:0] p3_add_12004_comb;
  wire [7:0] p3_actual_index__83_comb;
  wire [5:0] p3_add_12006_comb;
  wire [7:0] p3_actual_index__85_comb;
  wire [6:0] p3_add_12008_comb;
  wire [7:0] p3_actual_index__87_comb;
  wire [4:0] p3_add_12010_comb;
  wire [7:0] p3_actual_index__89_comb;
  wire [6:0] p3_add_12012_comb;
  wire [7:0] p3_actual_index__91_comb;
  wire [5:0] p3_add_12014_comb;
  wire [7:0] p3_actual_index__93_comb;
  wire [6:0] p3_add_12016_comb;
  wire [7:0] p3_actual_index__95_comb;
  wire [2:0] p3_add_12018_comb;
  wire [7:0] p3_actual_index__97_comb;
  wire [6:0] p3_add_12020_comb;
  wire [7:0] p3_actual_index__99_comb;
  wire [5:0] p3_add_12022_comb;
  wire [7:0] p3_actual_index__101_comb;
  wire [6:0] p3_add_12024_comb;
  wire [7:0] p3_actual_index__103_comb;
  wire [4:0] p3_add_12026_comb;
  wire [7:0] p3_actual_index__105_comb;
  wire [6:0] p3_add_12028_comb;
  wire [7:0] p3_actual_index__107_comb;
  wire [5:0] p3_add_12030_comb;
  wire [7:0] p3_actual_index__109_comb;
  wire [6:0] p3_add_12032_comb;
  wire [7:0] p3_actual_index__111_comb;
  wire [3:0] p3_add_12034_comb;
  wire [7:0] p3_actual_index__113_comb;
  wire [6:0] p3_add_12036_comb;
  wire [7:0] p3_actual_index__115_comb;
  wire [5:0] p3_add_12038_comb;
  wire [7:0] p3_actual_index__117_comb;
  wire [6:0] p3_add_12040_comb;
  wire [7:0] p3_actual_index__119_comb;
  wire [4:0] p3_add_12042_comb;
  wire [7:0] p3_actual_index__121_comb;
  wire [6:0] p3_add_12044_comb;
  wire [7:0] p3_actual_index__123_comb;
  wire [5:0] p3_add_12046_comb;
  wire [7:0] p3_actual_index__125_comb;
  wire [6:0] p3_add_12048_comb;
  wire [7:0] p3_actual_index__127_comb;
  wire [7:0] p3_bin_value__1_comb;
  wire [7:0] p3_bin_value_comb;
  wire [7:0] p3_actual_index__66_comb;
  wire [7:0] p3_actual_index__68_comb;
  wire [7:0] p3_actual_index__70_comb;
  wire [7:0] p3_actual_index__72_comb;
  wire [7:0] p3_actual_index__74_comb;
  wire [7:0] p3_actual_index__76_comb;
  wire [7:0] p3_actual_index__78_comb;
  wire [7:0] p3_actual_index__80_comb;
  wire [7:0] p3_actual_index__82_comb;
  wire [7:0] p3_actual_index__84_comb;
  wire [7:0] p3_actual_index__86_comb;
  wire [7:0] p3_actual_index__88_comb;
  wire [7:0] p3_actual_index__90_comb;
  wire [7:0] p3_actual_index__92_comb;
  wire [7:0] p3_actual_index__94_comb;
  wire [7:0] p3_actual_index__96_comb;
  wire [7:0] p3_actual_index__98_comb;
  wire [7:0] p3_actual_index__100_comb;
  wire [7:0] p3_actual_index__102_comb;
  wire [7:0] p3_actual_index__104_comb;
  wire [7:0] p3_actual_index__106_comb;
  wire [7:0] p3_actual_index__108_comb;
  wire [7:0] p3_actual_index__110_comb;
  wire [7:0] p3_actual_index__112_comb;
  wire [7:0] p3_actual_index__114_comb;
  wire [7:0] p3_actual_index__116_comb;
  wire [7:0] p3_actual_index__118_comb;
  wire [7:0] p3_actual_index__120_comb;
  wire [7:0] p3_actual_index__122_comb;
  wire [7:0] p3_actual_index__124_comb;
  wire [7:0] p3_actual_index__126_comb;
  wire [7:0] p3_value_abs_comb;
  wire [9:0] p3_value_comb;
  wire p3_and_12599_comb;
  wire p3_next_pix__1_squeezed_squeezed_const_msb_bits__1_comb;
  wire [7:0] p3_flipped_comb;
  wire [7:0] p3_Code_list_comb;
  wire p3_or_reduce_11910_comb;
  wire [2:0] p3_sel_11911_comb;
  wire p3_or_reduce_11914_comb;
  wire p3_bit_slice_11983_comb;
  wire [4:0] p3_value_pix_num_squeezed_comb;
  wire p3_or_reduce_11986_comb;
  wire p3_bit_slice_12183_comb;
  wire p3_eq_12184_comb;
  wire [7:0] p3_code_list_comb;
  assign p3_run_0_squeezed_const_msb_bits_comb = 3'h0;
  assign p3_value_pix_num_comb = {p3_run_0_squeezed_const_msb_bits_comb, p2_add_11743} & {8{p2_eq_11744}};
  assign p3_start_pix_1__1_comb = p2_start_pix > 8'h40 ? 8'h40 : p2_start_pix;
  assign p3_add_11885_comb = p2_start_pix + p3_value_pix_num_comb;
  assign p3_value__1_comb = p3_add_11885_comb == 8'h00 ? p2_array_index_11336 : (p3_add_11885_comb == 8'h01 ? p2_array_index_11337 : (p3_add_11885_comb == 8'h02 ? p2_array_index_11338 : (p3_add_11885_comb == 8'h03 ? p2_array_index_11339 : (p3_add_11885_comb == 8'h04 ? p2_array_index_11340 : (p3_add_11885_comb == 8'h05 ? p2_array_index_11341 : (p3_add_11885_comb == 8'h06 ? p2_array_index_11342 : (p3_add_11885_comb == 8'h07 ? p2_array_index_11343 : (p3_add_11885_comb == 8'h08 ? p2_array_index_11344 : (p3_add_11885_comb == 8'h09 ? p2_array_index_11345 : (p3_add_11885_comb == 8'h0a ? p2_array_index_11346 : (p3_add_11885_comb == 8'h0b ? p2_array_index_11347 : (p3_add_11885_comb == 8'h0c ? p2_array_index_11348 : (p3_add_11885_comb == 8'h0d ? p2_array_index_11349 : (p3_add_11885_comb == 8'h0e ? p2_array_index_11350 : (p3_add_11885_comb == 8'h0f ? p2_array_index_11351 : (p3_add_11885_comb == 8'h10 ? p2_array_index_11352 : (p3_add_11885_comb == 8'h11 ? p2_array_index_11353 : (p3_add_11885_comb == 8'h12 ? p2_array_index_11354 : (p3_add_11885_comb == 8'h13 ? p2_array_index_11355 : (p3_add_11885_comb == 8'h14 ? p2_array_index_11356 : (p3_add_11885_comb == 8'h15 ? p2_array_index_11357 : (p3_add_11885_comb == 8'h16 ? p2_array_index_11358 : (p3_add_11885_comb == 8'h17 ? p2_array_index_11359 : (p3_add_11885_comb == 8'h18 ? p2_array_index_11360 : (p3_add_11885_comb == 8'h19 ? p2_array_index_11361 : (p3_add_11885_comb == 8'h1a ? p2_array_index_11362 : (p3_add_11885_comb == 8'h1b ? p2_array_index_11363 : (p3_add_11885_comb == 8'h1c ? p2_array_index_11364 : (p3_add_11885_comb == 8'h1d ? p2_array_index_11365 : (p3_add_11885_comb == 8'h1e ? p2_array_index_11366 : (p3_add_11885_comb == 8'h1f ? p2_array_index_11367 : (p3_add_11885_comb == 8'h20 ? p2_array_index_11368 : (p3_add_11885_comb == 8'h21 ? p2_array_index_11369 : (p3_add_11885_comb == 8'h22 ? p2_array_index_11370 : (p3_add_11885_comb == 8'h23 ? p2_array_index_11371 : (p3_add_11885_comb == 8'h24 ? p2_array_index_11372 : (p3_add_11885_comb == 8'h25 ? p2_array_index_11373 : (p3_add_11885_comb == 8'h26 ? p2_array_index_11374 : (p3_add_11885_comb == 8'h27 ? p2_array_index_11375 : (p3_add_11885_comb == 8'h28 ? p2_array_index_11376 : (p3_add_11885_comb == 8'h29 ? p2_array_index_11377 : (p3_add_11885_comb == 8'h2a ? p2_array_index_11378 : (p3_add_11885_comb == 8'h2b ? p2_array_index_11379 : (p3_add_11885_comb == 8'h2c ? p2_array_index_11380 : (p3_add_11885_comb == 8'h2d ? p2_array_index_11381 : (p3_add_11885_comb == 8'h2e ? p2_array_index_11382 : (p3_add_11885_comb == 8'h2f ? p2_array_index_11383 : (p3_add_11885_comb == 8'h30 ? p2_array_index_11384 : (p3_add_11885_comb == 8'h31 ? p2_array_index_11385 : (p3_add_11885_comb == 8'h32 ? p2_array_index_11386 : (p3_add_11885_comb == 8'h33 ? p2_array_index_11387 : (p3_add_11885_comb == 8'h34 ? p2_array_index_11388 : (p3_add_11885_comb == 8'h35 ? p2_array_index_11389 : (p3_add_11885_comb == 8'h36 ? p2_array_index_11390 : (p3_add_11885_comb == 8'h37 ? p2_array_index_11391 : (p3_add_11885_comb == 8'h38 ? p2_array_index_11392 : (p3_add_11885_comb == 8'h39 ? p2_array_index_11393 : (p3_add_11885_comb == 8'h3a ? p2_array_index_11394 : (p3_add_11885_comb == 8'h3b ? p2_array_index_11395 : (p3_add_11885_comb == 8'h3c ? p2_array_index_11396 : (p3_add_11885_comb == 8'h3d ? p2_array_index_11397 : (p3_add_11885_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign p3_actual_index__65_comb = p3_start_pix_1__1_comb + 8'h01;
  assign p3_add_11988_comb = p3_start_pix_1__1_comb[7:1] + 7'h01;
  assign p3_actual_index__67_comb = p3_start_pix_1__1_comb + 8'h03;
  assign p3_add_11990_comb = p3_start_pix_1__1_comb[7:2] + 6'h01;
  assign p3_actual_index__69_comb = p3_start_pix_1__1_comb + 8'h05;
  assign p3_add_11992_comb = p3_start_pix_1__1_comb[7:1] + 7'h03;
  assign p3_actual_index__71_comb = p3_start_pix_1__1_comb + 8'h07;
  assign p3_add_11994_comb = p3_start_pix_1__1_comb[7:3] + 5'h01;
  assign p3_actual_index__73_comb = p3_start_pix_1__1_comb + 8'h09;
  assign p3_add_11996_comb = p3_start_pix_1__1_comb[7:1] + 7'h05;
  assign p3_actual_index__75_comb = p3_start_pix_1__1_comb + 8'h0b;
  assign p3_add_11998_comb = p3_start_pix_1__1_comb[7:2] + 6'h03;
  assign p3_actual_index__77_comb = p3_start_pix_1__1_comb + 8'h0d;
  assign p3_add_12000_comb = p3_start_pix_1__1_comb[7:1] + 7'h07;
  assign p3_actual_index__79_comb = p3_start_pix_1__1_comb + 8'h0f;
  assign p3_add_12002_comb = p3_start_pix_1__1_comb[7:4] + 4'h1;
  assign p3_actual_index__81_comb = p3_start_pix_1__1_comb + 8'h11;
  assign p3_add_12004_comb = p3_start_pix_1__1_comb[7:1] + 7'h09;
  assign p3_actual_index__83_comb = p3_start_pix_1__1_comb + 8'h13;
  assign p3_add_12006_comb = p3_start_pix_1__1_comb[7:2] + 6'h05;
  assign p3_actual_index__85_comb = p3_start_pix_1__1_comb + 8'h15;
  assign p3_add_12008_comb = p3_start_pix_1__1_comb[7:1] + 7'h0b;
  assign p3_actual_index__87_comb = p3_start_pix_1__1_comb + 8'h17;
  assign p3_add_12010_comb = p3_start_pix_1__1_comb[7:3] + 5'h03;
  assign p3_actual_index__89_comb = p3_start_pix_1__1_comb + 8'h19;
  assign p3_add_12012_comb = p3_start_pix_1__1_comb[7:1] + 7'h0d;
  assign p3_actual_index__91_comb = p3_start_pix_1__1_comb + 8'h1b;
  assign p3_add_12014_comb = p3_start_pix_1__1_comb[7:2] + 6'h07;
  assign p3_actual_index__93_comb = p3_start_pix_1__1_comb + 8'h1d;
  assign p3_add_12016_comb = p3_start_pix_1__1_comb[7:1] + 7'h0f;
  assign p3_actual_index__95_comb = p3_start_pix_1__1_comb + 8'h1f;
  assign p3_add_12018_comb = p3_start_pix_1__1_comb[7:5] + 3'h1;
  assign p3_actual_index__97_comb = p3_start_pix_1__1_comb + 8'h21;
  assign p3_add_12020_comb = p3_start_pix_1__1_comb[7:1] + 7'h11;
  assign p3_actual_index__99_comb = p3_start_pix_1__1_comb + 8'h23;
  assign p3_add_12022_comb = p3_start_pix_1__1_comb[7:2] + 6'h09;
  assign p3_actual_index__101_comb = p3_start_pix_1__1_comb + 8'h25;
  assign p3_add_12024_comb = p3_start_pix_1__1_comb[7:1] + 7'h13;
  assign p3_actual_index__103_comb = p3_start_pix_1__1_comb + 8'h27;
  assign p3_add_12026_comb = p3_start_pix_1__1_comb[7:3] + 5'h05;
  assign p3_actual_index__105_comb = p3_start_pix_1__1_comb + 8'h29;
  assign p3_add_12028_comb = p3_start_pix_1__1_comb[7:1] + 7'h15;
  assign p3_actual_index__107_comb = p3_start_pix_1__1_comb + 8'h2b;
  assign p3_add_12030_comb = p3_start_pix_1__1_comb[7:2] + 6'h0b;
  assign p3_actual_index__109_comb = p3_start_pix_1__1_comb + 8'h2d;
  assign p3_add_12032_comb = p3_start_pix_1__1_comb[7:1] + 7'h17;
  assign p3_actual_index__111_comb = p3_start_pix_1__1_comb + 8'h2f;
  assign p3_add_12034_comb = p3_start_pix_1__1_comb[7:4] + 4'h3;
  assign p3_actual_index__113_comb = p3_start_pix_1__1_comb + 8'h31;
  assign p3_add_12036_comb = p3_start_pix_1__1_comb[7:1] + 7'h19;
  assign p3_actual_index__115_comb = p3_start_pix_1__1_comb + 8'h33;
  assign p3_add_12038_comb = p3_start_pix_1__1_comb[7:2] + 6'h0d;
  assign p3_actual_index__117_comb = p3_start_pix_1__1_comb + 8'h35;
  assign p3_add_12040_comb = p3_start_pix_1__1_comb[7:1] + 7'h1b;
  assign p3_actual_index__119_comb = p3_start_pix_1__1_comb + 8'h37;
  assign p3_add_12042_comb = p3_start_pix_1__1_comb[7:3] + 5'h07;
  assign p3_actual_index__121_comb = p3_start_pix_1__1_comb + 8'h39;
  assign p3_add_12044_comb = p3_start_pix_1__1_comb[7:1] + 7'h1d;
  assign p3_actual_index__123_comb = p3_start_pix_1__1_comb + 8'h3b;
  assign p3_add_12046_comb = p3_start_pix_1__1_comb[7:2] + 6'h0f;
  assign p3_actual_index__125_comb = p3_start_pix_1__1_comb + 8'h3d;
  assign p3_add_12048_comb = p3_start_pix_1__1_comb[7:1] + 7'h1f;
  assign p3_actual_index__127_comb = p3_start_pix_1__1_comb + 8'h3f;
  assign p3_bin_value__1_comb = p3_value__1_comb[7:0];
  assign p3_bin_value_comb = -p3_bin_value__1_comb;
  assign p3_actual_index__66_comb = {p3_add_11988_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__68_comb = {p3_add_11990_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__70_comb = {p3_add_11992_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__72_comb = {p3_add_11994_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__74_comb = {p3_add_11996_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__76_comb = {p3_add_11998_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__78_comb = {p3_add_12000_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__80_comb = {p3_add_12002_comb, p3_start_pix_1__1_comb[3:0]};
  assign p3_actual_index__82_comb = {p3_add_12004_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__84_comb = {p3_add_12006_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__86_comb = {p3_add_12008_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__88_comb = {p3_add_12010_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__90_comb = {p3_add_12012_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__92_comb = {p3_add_12014_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__94_comb = {p3_add_12016_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__96_comb = {p3_add_12018_comb, p3_start_pix_1__1_comb[4:0]};
  assign p3_actual_index__98_comb = {p3_add_12020_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__100_comb = {p3_add_12022_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__102_comb = {p3_add_12024_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__104_comb = {p3_add_12026_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__106_comb = {p3_add_12028_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__108_comb = {p3_add_12030_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__110_comb = {p3_add_12032_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__112_comb = {p3_add_12034_comb, p3_start_pix_1__1_comb[3:0]};
  assign p3_actual_index__114_comb = {p3_add_12036_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__116_comb = {p3_add_12038_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__118_comb = {p3_add_12040_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__120_comb = {p3_add_12042_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__122_comb = {p3_add_12044_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__124_comb = {p3_add_12046_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__126_comb = {p3_add_12048_comb, p3_start_pix_1__1_comb[0]};
  assign p3_value_abs_comb = p3_value__1_comb[9] ? p3_bin_value_comb : p3_bin_value__1_comb;
  assign p3_value_comb = p2_start_pix == 8'h00 ? p2_array_index_11336 : (p2_start_pix == 8'h01 ? p2_array_index_11337 : (p2_start_pix == 8'h02 ? p2_array_index_11338 : (p2_start_pix == 8'h03 ? p2_array_index_11339 : (p2_start_pix == 8'h04 ? p2_array_index_11340 : (p2_start_pix == 8'h05 ? p2_array_index_11341 : (p2_start_pix == 8'h06 ? p2_array_index_11342 : (p2_start_pix == 8'h07 ? p2_array_index_11343 : (p2_start_pix == 8'h08 ? p2_array_index_11344 : (p2_start_pix == 8'h09 ? p2_array_index_11345 : (p2_start_pix == 8'h0a ? p2_array_index_11346 : (p2_start_pix == 8'h0b ? p2_array_index_11347 : (p2_start_pix == 8'h0c ? p2_array_index_11348 : (p2_start_pix == 8'h0d ? p2_array_index_11349 : (p2_start_pix == 8'h0e ? p2_array_index_11350 : (p2_start_pix == 8'h0f ? p2_array_index_11351 : (p2_start_pix == 8'h10 ? p2_array_index_11352 : (p2_start_pix == 8'h11 ? p2_array_index_11353 : (p2_start_pix == 8'h12 ? p2_array_index_11354 : (p2_start_pix == 8'h13 ? p2_array_index_11355 : (p2_start_pix == 8'h14 ? p2_array_index_11356 : (p2_start_pix == 8'h15 ? p2_array_index_11357 : (p2_start_pix == 8'h16 ? p2_array_index_11358 : (p2_start_pix == 8'h17 ? p2_array_index_11359 : (p2_start_pix == 8'h18 ? p2_array_index_11360 : (p2_start_pix == 8'h19 ? p2_array_index_11361 : (p2_start_pix == 8'h1a ? p2_array_index_11362 : (p2_start_pix == 8'h1b ? p2_array_index_11363 : (p2_start_pix == 8'h1c ? p2_array_index_11364 : (p2_start_pix == 8'h1d ? p2_array_index_11365 : (p2_start_pix == 8'h1e ? p2_array_index_11366 : (p2_start_pix == 8'h1f ? p2_array_index_11367 : (p2_start_pix == 8'h20 ? p2_array_index_11368 : (p2_start_pix == 8'h21 ? p2_array_index_11369 : (p2_start_pix == 8'h22 ? p2_array_index_11370 : (p2_start_pix == 8'h23 ? p2_array_index_11371 : (p2_start_pix == 8'h24 ? p2_array_index_11372 : (p2_start_pix == 8'h25 ? p2_array_index_11373 : (p2_start_pix == 8'h26 ? p2_array_index_11374 : (p2_start_pix == 8'h27 ? p2_array_index_11375 : (p2_start_pix == 8'h28 ? p2_array_index_11376 : (p2_start_pix == 8'h29 ? p2_array_index_11377 : (p2_start_pix == 8'h2a ? p2_array_index_11378 : (p2_start_pix == 8'h2b ? p2_array_index_11379 : (p2_start_pix == 8'h2c ? p2_array_index_11380 : (p2_start_pix == 8'h2d ? p2_array_index_11381 : (p2_start_pix == 8'h2e ? p2_array_index_11382 : (p2_start_pix == 8'h2f ? p2_array_index_11383 : (p2_start_pix == 8'h30 ? p2_array_index_11384 : (p2_start_pix == 8'h31 ? p2_array_index_11385 : (p2_start_pix == 8'h32 ? p2_array_index_11386 : (p2_start_pix == 8'h33 ? p2_array_index_11387 : (p2_start_pix == 8'h34 ? p2_array_index_11388 : (p2_start_pix == 8'h35 ? p2_array_index_11389 : (p2_start_pix == 8'h36 ? p2_array_index_11390 : (p2_start_pix == 8'h37 ? p2_array_index_11391 : (p2_start_pix == 8'h38 ? p2_array_index_11392 : (p2_start_pix == 8'h39 ? p2_array_index_11393 : (p2_start_pix == 8'h3a ? p2_array_index_11394 : (p2_start_pix == 8'h3b ? p2_array_index_11395 : (p2_start_pix == 8'h3c ? p2_array_index_11396 : (p2_start_pix == 8'h3d ? p2_array_index_11397 : (p2_start_pix == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign p3_and_12599_comb = (p3_value_comb & {10{~p3_start_pix_1__1_comb[6]}}) == 10'h000 & ((p3_actual_index__65_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__65_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__65_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__65_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__65_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__65_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__65_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__65_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__65_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__65_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__65_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__65_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__65_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__65_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__65_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__65_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__65_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__65_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__65_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__65_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__65_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__65_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__65_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__65_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__65_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__65_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__65_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__65_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__65_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__65_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__65_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__65_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__65_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__65_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__65_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__65_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__65_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__65_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__65_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__65_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__65_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__65_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__65_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__65_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__65_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__65_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__65_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__65_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__65_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__65_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__65_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__65_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__65_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__65_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__65_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__65_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__65_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__65_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__65_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__65_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__65_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__65_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__65_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__65_comb[6] | p3_actual_index__65_comb[7])}}) == 10'h000 & ((p3_actual_index__66_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__66_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__66_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__66_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__66_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__66_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__66_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__66_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__66_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__66_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__66_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__66_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__66_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__66_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__66_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__66_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__66_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__66_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__66_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__66_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__66_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__66_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__66_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__66_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__66_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__66_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__66_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__66_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__66_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__66_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__66_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__66_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__66_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__66_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__66_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__66_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__66_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__66_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__66_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__66_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__66_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__66_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__66_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__66_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__66_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__66_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__66_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__66_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__66_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__66_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__66_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__66_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__66_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__66_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__66_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__66_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__66_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__66_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__66_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__66_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__66_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__66_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__66_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_11988_comb[5] | p3_add_11988_comb[6])}}) == 10'h000 & ((p3_actual_index__67_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__67_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__67_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__67_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__67_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__67_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__67_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__67_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__67_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__67_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__67_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__67_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__67_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__67_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__67_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__67_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__67_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__67_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__67_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__67_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__67_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__67_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__67_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__67_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__67_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__67_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__67_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__67_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__67_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__67_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__67_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__67_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__67_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__67_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__67_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__67_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__67_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__67_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__67_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__67_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__67_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__67_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__67_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__67_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__67_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__67_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__67_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__67_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__67_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__67_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__67_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__67_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__67_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__67_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__67_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__67_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__67_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__67_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__67_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__67_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__67_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__67_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__67_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__67_comb[6] | p3_actual_index__67_comb[7])}}) == 10'h000 & ((p3_actual_index__68_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__68_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__68_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__68_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__68_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__68_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__68_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__68_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__68_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__68_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__68_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__68_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__68_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__68_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__68_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__68_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__68_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__68_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__68_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__68_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__68_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__68_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__68_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__68_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__68_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__68_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__68_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__68_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__68_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__68_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__68_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__68_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__68_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__68_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__68_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__68_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__68_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__68_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__68_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__68_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__68_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__68_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__68_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__68_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__68_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__68_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__68_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__68_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__68_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__68_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__68_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__68_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__68_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__68_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__68_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__68_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__68_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__68_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__68_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__68_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__68_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__68_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__68_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_11990_comb[4] | p3_add_11990_comb[5])}}) == 10'h000 & ((p3_actual_index__69_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__69_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__69_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__69_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__69_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__69_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__69_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__69_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__69_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__69_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__69_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__69_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__69_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__69_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__69_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__69_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__69_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__69_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__69_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__69_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__69_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__69_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__69_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__69_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__69_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__69_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__69_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__69_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__69_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__69_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__69_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__69_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__69_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__69_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__69_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__69_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__69_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__69_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__69_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__69_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__69_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__69_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__69_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__69_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__69_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__69_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__69_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__69_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__69_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__69_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__69_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__69_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__69_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__69_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__69_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__69_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__69_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__69_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__69_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__69_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__69_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__69_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__69_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__69_comb[6] | p3_actual_index__69_comb[7])}}) == 10'h000 & ((p3_actual_index__70_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__70_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__70_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__70_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__70_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__70_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__70_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__70_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__70_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__70_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__70_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__70_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__70_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__70_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__70_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__70_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__70_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__70_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__70_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__70_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__70_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__70_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__70_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__70_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__70_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__70_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__70_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__70_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__70_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__70_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__70_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__70_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__70_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__70_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__70_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__70_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__70_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__70_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__70_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__70_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__70_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__70_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__70_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__70_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__70_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__70_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__70_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__70_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__70_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__70_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__70_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__70_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__70_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__70_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__70_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__70_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__70_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__70_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__70_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__70_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__70_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__70_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__70_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_11992_comb[5] | p3_add_11992_comb[6])}}) == 10'h000 & ((p3_actual_index__71_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__71_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__71_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__71_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__71_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__71_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__71_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__71_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__71_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__71_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__71_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__71_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__71_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__71_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__71_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__71_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__71_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__71_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__71_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__71_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__71_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__71_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__71_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__71_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__71_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__71_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__71_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__71_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__71_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__71_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__71_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__71_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__71_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__71_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__71_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__71_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__71_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__71_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__71_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__71_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__71_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__71_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__71_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__71_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__71_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__71_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__71_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__71_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__71_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__71_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__71_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__71_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__71_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__71_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__71_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__71_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__71_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__71_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__71_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__71_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__71_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__71_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__71_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__71_comb[6] | p3_actual_index__71_comb[7])}}) == 10'h000 & ((p3_actual_index__72_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__72_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__72_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__72_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__72_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__72_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__72_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__72_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__72_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__72_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__72_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__72_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__72_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__72_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__72_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__72_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__72_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__72_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__72_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__72_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__72_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__72_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__72_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__72_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__72_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__72_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__72_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__72_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__72_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__72_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__72_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__72_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__72_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__72_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__72_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__72_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__72_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__72_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__72_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__72_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__72_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__72_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__72_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__72_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__72_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__72_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__72_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__72_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__72_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__72_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__72_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__72_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__72_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__72_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__72_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__72_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__72_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__72_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__72_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__72_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__72_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__72_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__72_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_11994_comb[3] | p3_add_11994_comb[4])}}) == 10'h000 & ((p3_actual_index__73_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__73_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__73_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__73_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__73_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__73_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__73_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__73_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__73_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__73_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__73_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__73_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__73_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__73_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__73_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__73_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__73_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__73_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__73_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__73_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__73_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__73_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__73_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__73_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__73_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__73_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__73_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__73_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__73_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__73_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__73_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__73_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__73_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__73_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__73_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__73_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__73_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__73_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__73_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__73_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__73_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__73_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__73_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__73_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__73_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__73_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__73_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__73_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__73_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__73_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__73_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__73_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__73_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__73_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__73_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__73_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__73_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__73_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__73_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__73_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__73_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__73_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__73_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__73_comb[6] | p3_actual_index__73_comb[7])}}) == 10'h000 & ((p3_actual_index__74_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__74_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__74_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__74_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__74_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__74_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__74_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__74_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__74_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__74_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__74_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__74_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__74_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__74_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__74_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__74_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__74_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__74_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__74_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__74_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__74_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__74_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__74_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__74_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__74_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__74_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__74_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__74_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__74_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__74_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__74_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__74_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__74_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__74_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__74_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__74_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__74_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__74_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__74_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__74_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__74_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__74_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__74_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__74_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__74_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__74_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__74_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__74_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__74_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__74_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__74_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__74_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__74_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__74_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__74_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__74_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__74_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__74_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__74_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__74_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__74_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__74_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__74_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_11996_comb[5] | p3_add_11996_comb[6])}}) == 10'h000 & ((p3_actual_index__75_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__75_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__75_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__75_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__75_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__75_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__75_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__75_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__75_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__75_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__75_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__75_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__75_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__75_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__75_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__75_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__75_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__75_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__75_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__75_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__75_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__75_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__75_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__75_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__75_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__75_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__75_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__75_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__75_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__75_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__75_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__75_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__75_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__75_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__75_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__75_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__75_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__75_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__75_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__75_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__75_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__75_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__75_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__75_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__75_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__75_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__75_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__75_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__75_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__75_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__75_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__75_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__75_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__75_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__75_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__75_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__75_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__75_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__75_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__75_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__75_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__75_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__75_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__75_comb[6] | p3_actual_index__75_comb[7])}}) == 10'h000 & ((p3_actual_index__76_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__76_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__76_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__76_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__76_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__76_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__76_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__76_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__76_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__76_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__76_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__76_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__76_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__76_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__76_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__76_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__76_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__76_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__76_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__76_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__76_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__76_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__76_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__76_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__76_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__76_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__76_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__76_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__76_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__76_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__76_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__76_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__76_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__76_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__76_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__76_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__76_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__76_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__76_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__76_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__76_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__76_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__76_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__76_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__76_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__76_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__76_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__76_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__76_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__76_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__76_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__76_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__76_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__76_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__76_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__76_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__76_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__76_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__76_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__76_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__76_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__76_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__76_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_11998_comb[4] | p3_add_11998_comb[5])}}) == 10'h000 & ((p3_actual_index__77_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__77_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__77_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__77_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__77_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__77_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__77_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__77_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__77_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__77_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__77_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__77_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__77_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__77_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__77_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__77_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__77_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__77_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__77_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__77_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__77_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__77_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__77_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__77_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__77_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__77_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__77_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__77_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__77_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__77_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__77_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__77_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__77_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__77_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__77_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__77_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__77_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__77_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__77_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__77_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__77_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__77_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__77_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__77_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__77_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__77_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__77_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__77_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__77_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__77_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__77_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__77_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__77_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__77_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__77_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__77_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__77_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__77_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__77_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__77_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__77_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__77_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__77_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__77_comb[6] | p3_actual_index__77_comb[7])}}) == 10'h000 & ((p3_actual_index__78_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__78_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__78_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__78_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__78_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__78_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__78_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__78_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__78_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__78_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__78_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__78_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__78_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__78_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__78_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__78_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__78_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__78_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__78_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__78_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__78_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__78_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__78_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__78_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__78_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__78_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__78_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__78_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__78_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__78_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__78_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__78_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__78_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__78_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__78_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__78_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__78_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__78_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__78_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__78_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__78_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__78_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__78_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__78_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__78_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__78_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__78_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__78_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__78_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__78_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__78_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__78_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__78_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__78_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__78_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__78_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__78_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__78_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__78_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__78_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__78_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__78_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__78_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12000_comb[5] | p3_add_12000_comb[6])}}) == 10'h000 & ((p3_actual_index__79_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__79_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__79_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__79_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__79_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__79_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__79_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__79_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__79_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__79_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__79_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__79_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__79_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__79_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__79_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__79_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__79_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__79_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__79_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__79_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__79_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__79_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__79_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__79_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__79_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__79_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__79_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__79_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__79_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__79_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__79_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__79_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__79_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__79_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__79_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__79_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__79_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__79_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__79_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__79_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__79_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__79_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__79_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__79_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__79_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__79_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__79_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__79_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__79_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__79_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__79_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__79_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__79_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__79_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__79_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__79_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__79_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__79_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__79_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__79_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__79_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__79_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__79_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__79_comb[6] | p3_actual_index__79_comb[7])}}) == 10'h000 & ((p3_actual_index__80_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__80_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__80_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__80_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__80_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__80_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__80_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__80_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__80_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__80_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__80_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__80_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__80_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__80_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__80_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__80_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__80_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__80_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__80_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__80_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__80_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__80_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__80_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__80_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__80_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__80_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__80_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__80_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__80_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__80_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__80_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__80_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__80_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__80_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__80_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__80_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__80_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__80_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__80_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__80_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__80_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__80_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__80_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__80_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__80_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__80_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__80_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__80_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__80_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__80_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__80_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__80_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__80_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__80_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__80_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__80_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__80_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__80_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__80_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__80_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__80_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__80_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__80_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12002_comb[2] | p3_add_12002_comb[3])}}) == 10'h000 & ((p3_actual_index__81_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__81_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__81_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__81_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__81_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__81_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__81_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__81_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__81_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__81_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__81_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__81_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__81_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__81_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__81_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__81_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__81_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__81_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__81_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__81_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__81_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__81_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__81_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__81_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__81_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__81_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__81_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__81_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__81_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__81_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__81_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__81_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__81_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__81_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__81_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__81_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__81_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__81_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__81_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__81_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__81_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__81_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__81_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__81_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__81_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__81_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__81_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__81_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__81_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__81_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__81_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__81_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__81_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__81_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__81_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__81_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__81_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__81_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__81_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__81_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__81_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__81_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__81_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__81_comb[6] | p3_actual_index__81_comb[7])}}) == 10'h000 & ((p3_actual_index__82_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__82_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__82_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__82_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__82_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__82_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__82_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__82_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__82_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__82_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__82_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__82_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__82_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__82_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__82_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__82_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__82_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__82_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__82_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__82_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__82_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__82_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__82_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__82_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__82_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__82_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__82_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__82_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__82_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__82_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__82_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__82_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__82_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__82_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__82_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__82_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__82_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__82_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__82_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__82_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__82_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__82_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__82_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__82_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__82_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__82_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__82_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__82_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__82_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__82_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__82_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__82_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__82_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__82_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__82_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__82_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__82_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__82_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__82_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__82_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__82_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__82_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__82_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12004_comb[5] | p3_add_12004_comb[6])}}) == 10'h000 & ((p3_actual_index__83_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__83_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__83_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__83_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__83_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__83_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__83_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__83_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__83_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__83_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__83_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__83_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__83_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__83_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__83_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__83_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__83_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__83_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__83_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__83_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__83_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__83_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__83_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__83_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__83_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__83_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__83_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__83_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__83_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__83_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__83_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__83_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__83_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__83_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__83_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__83_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__83_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__83_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__83_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__83_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__83_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__83_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__83_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__83_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__83_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__83_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__83_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__83_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__83_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__83_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__83_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__83_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__83_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__83_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__83_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__83_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__83_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__83_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__83_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__83_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__83_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__83_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__83_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__83_comb[6] | p3_actual_index__83_comb[7])}}) == 10'h000 & ((p3_actual_index__84_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__84_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__84_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__84_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__84_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__84_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__84_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__84_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__84_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__84_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__84_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__84_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__84_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__84_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__84_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__84_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__84_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__84_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__84_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__84_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__84_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__84_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__84_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__84_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__84_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__84_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__84_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__84_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__84_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__84_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__84_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__84_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__84_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__84_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__84_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__84_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__84_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__84_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__84_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__84_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__84_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__84_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__84_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__84_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__84_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__84_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__84_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__84_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__84_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__84_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__84_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__84_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__84_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__84_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__84_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__84_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__84_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__84_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__84_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__84_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__84_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__84_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__84_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12006_comb[4] | p3_add_12006_comb[5])}}) == 10'h000 & ((p3_actual_index__85_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__85_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__85_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__85_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__85_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__85_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__85_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__85_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__85_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__85_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__85_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__85_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__85_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__85_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__85_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__85_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__85_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__85_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__85_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__85_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__85_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__85_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__85_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__85_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__85_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__85_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__85_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__85_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__85_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__85_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__85_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__85_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__85_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__85_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__85_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__85_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__85_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__85_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__85_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__85_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__85_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__85_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__85_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__85_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__85_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__85_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__85_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__85_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__85_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__85_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__85_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__85_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__85_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__85_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__85_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__85_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__85_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__85_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__85_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__85_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__85_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__85_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__85_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__85_comb[6] | p3_actual_index__85_comb[7])}}) == 10'h000 & ((p3_actual_index__86_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__86_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__86_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__86_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__86_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__86_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__86_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__86_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__86_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__86_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__86_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__86_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__86_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__86_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__86_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__86_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__86_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__86_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__86_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__86_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__86_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__86_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__86_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__86_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__86_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__86_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__86_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__86_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__86_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__86_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__86_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__86_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__86_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__86_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__86_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__86_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__86_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__86_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__86_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__86_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__86_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__86_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__86_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__86_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__86_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__86_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__86_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__86_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__86_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__86_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__86_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__86_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__86_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__86_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__86_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__86_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__86_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__86_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__86_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__86_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__86_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__86_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__86_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12008_comb[5] | p3_add_12008_comb[6])}}) == 10'h000 & ((p3_actual_index__87_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__87_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__87_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__87_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__87_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__87_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__87_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__87_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__87_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__87_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__87_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__87_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__87_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__87_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__87_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__87_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__87_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__87_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__87_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__87_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__87_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__87_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__87_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__87_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__87_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__87_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__87_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__87_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__87_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__87_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__87_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__87_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__87_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__87_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__87_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__87_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__87_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__87_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__87_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__87_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__87_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__87_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__87_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__87_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__87_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__87_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__87_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__87_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__87_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__87_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__87_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__87_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__87_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__87_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__87_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__87_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__87_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__87_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__87_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__87_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__87_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__87_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__87_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__87_comb[6] | p3_actual_index__87_comb[7])}}) == 10'h000 & ((p3_actual_index__88_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__88_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__88_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__88_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__88_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__88_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__88_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__88_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__88_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__88_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__88_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__88_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__88_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__88_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__88_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__88_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__88_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__88_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__88_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__88_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__88_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__88_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__88_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__88_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__88_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__88_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__88_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__88_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__88_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__88_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__88_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__88_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__88_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__88_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__88_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__88_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__88_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__88_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__88_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__88_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__88_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__88_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__88_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__88_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__88_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__88_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__88_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__88_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__88_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__88_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__88_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__88_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__88_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__88_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__88_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__88_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__88_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__88_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__88_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__88_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__88_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__88_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__88_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12010_comb[3] | p3_add_12010_comb[4])}}) == 10'h000 & ((p3_actual_index__89_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__89_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__89_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__89_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__89_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__89_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__89_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__89_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__89_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__89_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__89_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__89_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__89_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__89_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__89_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__89_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__89_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__89_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__89_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__89_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__89_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__89_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__89_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__89_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__89_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__89_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__89_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__89_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__89_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__89_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__89_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__89_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__89_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__89_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__89_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__89_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__89_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__89_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__89_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__89_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__89_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__89_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__89_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__89_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__89_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__89_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__89_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__89_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__89_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__89_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__89_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__89_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__89_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__89_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__89_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__89_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__89_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__89_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__89_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__89_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__89_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__89_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__89_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__89_comb[6] | p3_actual_index__89_comb[7])}}) == 10'h000 & ((p3_actual_index__90_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__90_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__90_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__90_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__90_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__90_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__90_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__90_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__90_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__90_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__90_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__90_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__90_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__90_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__90_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__90_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__90_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__90_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__90_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__90_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__90_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__90_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__90_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__90_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__90_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__90_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__90_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__90_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__90_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__90_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__90_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__90_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__90_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__90_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__90_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__90_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__90_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__90_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__90_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__90_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__90_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__90_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__90_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__90_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__90_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__90_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__90_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__90_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__90_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__90_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__90_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__90_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__90_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__90_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__90_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__90_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__90_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__90_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__90_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__90_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__90_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__90_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__90_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12012_comb[5] | p3_add_12012_comb[6])}}) == 10'h000 & ((p3_actual_index__91_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__91_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__91_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__91_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__91_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__91_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__91_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__91_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__91_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__91_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__91_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__91_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__91_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__91_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__91_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__91_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__91_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__91_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__91_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__91_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__91_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__91_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__91_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__91_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__91_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__91_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__91_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__91_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__91_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__91_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__91_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__91_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__91_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__91_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__91_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__91_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__91_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__91_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__91_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__91_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__91_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__91_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__91_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__91_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__91_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__91_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__91_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__91_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__91_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__91_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__91_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__91_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__91_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__91_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__91_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__91_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__91_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__91_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__91_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__91_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__91_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__91_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__91_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__91_comb[6] | p3_actual_index__91_comb[7])}}) == 10'h000 & ((p3_actual_index__92_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__92_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__92_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__92_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__92_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__92_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__92_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__92_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__92_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__92_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__92_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__92_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__92_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__92_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__92_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__92_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__92_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__92_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__92_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__92_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__92_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__92_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__92_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__92_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__92_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__92_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__92_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__92_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__92_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__92_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__92_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__92_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__92_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__92_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__92_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__92_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__92_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__92_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__92_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__92_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__92_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__92_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__92_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__92_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__92_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__92_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__92_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__92_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__92_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__92_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__92_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__92_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__92_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__92_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__92_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__92_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__92_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__92_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__92_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__92_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__92_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__92_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__92_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12014_comb[4] | p3_add_12014_comb[5])}}) == 10'h000 & ((p3_actual_index__93_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__93_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__93_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__93_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__93_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__93_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__93_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__93_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__93_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__93_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__93_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__93_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__93_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__93_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__93_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__93_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__93_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__93_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__93_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__93_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__93_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__93_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__93_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__93_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__93_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__93_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__93_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__93_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__93_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__93_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__93_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__93_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__93_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__93_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__93_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__93_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__93_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__93_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__93_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__93_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__93_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__93_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__93_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__93_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__93_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__93_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__93_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__93_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__93_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__93_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__93_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__93_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__93_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__93_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__93_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__93_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__93_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__93_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__93_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__93_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__93_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__93_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__93_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__93_comb[6] | p3_actual_index__93_comb[7])}}) == 10'h000 & ((p3_actual_index__94_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__94_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__94_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__94_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__94_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__94_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__94_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__94_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__94_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__94_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__94_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__94_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__94_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__94_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__94_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__94_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__94_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__94_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__94_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__94_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__94_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__94_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__94_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__94_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__94_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__94_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__94_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__94_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__94_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__94_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__94_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__94_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__94_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__94_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__94_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__94_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__94_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__94_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__94_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__94_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__94_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__94_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__94_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__94_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__94_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__94_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__94_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__94_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__94_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__94_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__94_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__94_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__94_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__94_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__94_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__94_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__94_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__94_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__94_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__94_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__94_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__94_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__94_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12016_comb[5] | p3_add_12016_comb[6])}}) == 10'h000 & ((p3_actual_index__95_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__95_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__95_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__95_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__95_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__95_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__95_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__95_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__95_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__95_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__95_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__95_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__95_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__95_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__95_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__95_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__95_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__95_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__95_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__95_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__95_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__95_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__95_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__95_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__95_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__95_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__95_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__95_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__95_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__95_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__95_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__95_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__95_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__95_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__95_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__95_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__95_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__95_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__95_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__95_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__95_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__95_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__95_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__95_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__95_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__95_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__95_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__95_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__95_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__95_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__95_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__95_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__95_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__95_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__95_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__95_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__95_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__95_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__95_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__95_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__95_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__95_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__95_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__95_comb[6] | p3_actual_index__95_comb[7])}}) == 10'h000 & ((p3_actual_index__96_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__96_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__96_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__96_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__96_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__96_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__96_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__96_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__96_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__96_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__96_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__96_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__96_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__96_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__96_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__96_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__96_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__96_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__96_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__96_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__96_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__96_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__96_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__96_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__96_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__96_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__96_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__96_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__96_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__96_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__96_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__96_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__96_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__96_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__96_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__96_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__96_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__96_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__96_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__96_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__96_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__96_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__96_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__96_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__96_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__96_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__96_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__96_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__96_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__96_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__96_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__96_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__96_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__96_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__96_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__96_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__96_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__96_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__96_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__96_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__96_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__96_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__96_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12018_comb[1] | p3_add_12018_comb[2])}}) == 10'h000 & ((p3_actual_index__97_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__97_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__97_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__97_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__97_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__97_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__97_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__97_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__97_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__97_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__97_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__97_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__97_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__97_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__97_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__97_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__97_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__97_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__97_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__97_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__97_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__97_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__97_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__97_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__97_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__97_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__97_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__97_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__97_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__97_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__97_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__97_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__97_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__97_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__97_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__97_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__97_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__97_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__97_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__97_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__97_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__97_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__97_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__97_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__97_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__97_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__97_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__97_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__97_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__97_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__97_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__97_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__97_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__97_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__97_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__97_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__97_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__97_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__97_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__97_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__97_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__97_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__97_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__97_comb[6] | p3_actual_index__97_comb[7])}}) == 10'h000 & ((p3_actual_index__98_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__98_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__98_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__98_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__98_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__98_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__98_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__98_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__98_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__98_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__98_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__98_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__98_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__98_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__98_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__98_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__98_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__98_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__98_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__98_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__98_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__98_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__98_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__98_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__98_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__98_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__98_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__98_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__98_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__98_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__98_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__98_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__98_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__98_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__98_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__98_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__98_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__98_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__98_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__98_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__98_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__98_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__98_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__98_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__98_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__98_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__98_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__98_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__98_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__98_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__98_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__98_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__98_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__98_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__98_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__98_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__98_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__98_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__98_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__98_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__98_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__98_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__98_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12020_comb[5] | p3_add_12020_comb[6])}}) == 10'h000 & ((p3_actual_index__99_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__99_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__99_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__99_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__99_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__99_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__99_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__99_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__99_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__99_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__99_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__99_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__99_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__99_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__99_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__99_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__99_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__99_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__99_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__99_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__99_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__99_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__99_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__99_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__99_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__99_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__99_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__99_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__99_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__99_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__99_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__99_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__99_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__99_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__99_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__99_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__99_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__99_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__99_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__99_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__99_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__99_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__99_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__99_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__99_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__99_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__99_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__99_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__99_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__99_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__99_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__99_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__99_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__99_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__99_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__99_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__99_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__99_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__99_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__99_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__99_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__99_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__99_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__99_comb[6] | p3_actual_index__99_comb[7])}}) == 10'h000 & ((p3_actual_index__100_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__100_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__100_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__100_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__100_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__100_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__100_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__100_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__100_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__100_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__100_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__100_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__100_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__100_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__100_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__100_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__100_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__100_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__100_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__100_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__100_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__100_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__100_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__100_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__100_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__100_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__100_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__100_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__100_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__100_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__100_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__100_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__100_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__100_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__100_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__100_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__100_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__100_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__100_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__100_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__100_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__100_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__100_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__100_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__100_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__100_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__100_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__100_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__100_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__100_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__100_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__100_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__100_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__100_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__100_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__100_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__100_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__100_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__100_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__100_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__100_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__100_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__100_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12022_comb[4] | p3_add_12022_comb[5])}}) == 10'h000 & ((p3_actual_index__101_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__101_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__101_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__101_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__101_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__101_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__101_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__101_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__101_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__101_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__101_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__101_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__101_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__101_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__101_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__101_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__101_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__101_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__101_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__101_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__101_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__101_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__101_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__101_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__101_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__101_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__101_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__101_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__101_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__101_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__101_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__101_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__101_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__101_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__101_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__101_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__101_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__101_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__101_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__101_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__101_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__101_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__101_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__101_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__101_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__101_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__101_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__101_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__101_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__101_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__101_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__101_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__101_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__101_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__101_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__101_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__101_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__101_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__101_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__101_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__101_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__101_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__101_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__101_comb[6] | p3_actual_index__101_comb[7])}}) == 10'h000 & ((p3_actual_index__102_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__102_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__102_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__102_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__102_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__102_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__102_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__102_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__102_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__102_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__102_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__102_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__102_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__102_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__102_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__102_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__102_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__102_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__102_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__102_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__102_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__102_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__102_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__102_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__102_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__102_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__102_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__102_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__102_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__102_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__102_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__102_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__102_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__102_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__102_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__102_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__102_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__102_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__102_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__102_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__102_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__102_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__102_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__102_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__102_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__102_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__102_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__102_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__102_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__102_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__102_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__102_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__102_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__102_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__102_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__102_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__102_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__102_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__102_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__102_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__102_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__102_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__102_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12024_comb[5] | p3_add_12024_comb[6])}}) == 10'h000 & ((p3_actual_index__103_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__103_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__103_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__103_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__103_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__103_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__103_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__103_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__103_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__103_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__103_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__103_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__103_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__103_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__103_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__103_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__103_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__103_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__103_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__103_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__103_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__103_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__103_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__103_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__103_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__103_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__103_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__103_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__103_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__103_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__103_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__103_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__103_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__103_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__103_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__103_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__103_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__103_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__103_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__103_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__103_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__103_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__103_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__103_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__103_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__103_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__103_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__103_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__103_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__103_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__103_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__103_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__103_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__103_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__103_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__103_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__103_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__103_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__103_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__103_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__103_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__103_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__103_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__103_comb[6] | p3_actual_index__103_comb[7])}}) == 10'h000 & ((p3_actual_index__104_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__104_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__104_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__104_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__104_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__104_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__104_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__104_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__104_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__104_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__104_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__104_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__104_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__104_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__104_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__104_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__104_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__104_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__104_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__104_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__104_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__104_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__104_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__104_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__104_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__104_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__104_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__104_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__104_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__104_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__104_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__104_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__104_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__104_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__104_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__104_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__104_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__104_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__104_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__104_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__104_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__104_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__104_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__104_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__104_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__104_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__104_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__104_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__104_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__104_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__104_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__104_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__104_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__104_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__104_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__104_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__104_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__104_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__104_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__104_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__104_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__104_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__104_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12026_comb[3] | p3_add_12026_comb[4])}}) == 10'h000 & ((p3_actual_index__105_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__105_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__105_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__105_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__105_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__105_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__105_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__105_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__105_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__105_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__105_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__105_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__105_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__105_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__105_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__105_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__105_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__105_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__105_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__105_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__105_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__105_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__105_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__105_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__105_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__105_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__105_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__105_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__105_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__105_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__105_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__105_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__105_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__105_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__105_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__105_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__105_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__105_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__105_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__105_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__105_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__105_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__105_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__105_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__105_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__105_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__105_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__105_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__105_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__105_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__105_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__105_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__105_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__105_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__105_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__105_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__105_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__105_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__105_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__105_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__105_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__105_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__105_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__105_comb[6] | p3_actual_index__105_comb[7])}}) == 10'h000 & ((p3_actual_index__106_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__106_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__106_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__106_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__106_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__106_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__106_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__106_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__106_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__106_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__106_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__106_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__106_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__106_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__106_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__106_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__106_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__106_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__106_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__106_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__106_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__106_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__106_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__106_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__106_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__106_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__106_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__106_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__106_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__106_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__106_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__106_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__106_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__106_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__106_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__106_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__106_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__106_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__106_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__106_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__106_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__106_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__106_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__106_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__106_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__106_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__106_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__106_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__106_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__106_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__106_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__106_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__106_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__106_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__106_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__106_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__106_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__106_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__106_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__106_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__106_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__106_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__106_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12028_comb[5] | p3_add_12028_comb[6])}}) == 10'h000 & ((p3_actual_index__107_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__107_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__107_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__107_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__107_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__107_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__107_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__107_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__107_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__107_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__107_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__107_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__107_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__107_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__107_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__107_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__107_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__107_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__107_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__107_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__107_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__107_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__107_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__107_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__107_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__107_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__107_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__107_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__107_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__107_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__107_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__107_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__107_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__107_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__107_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__107_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__107_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__107_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__107_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__107_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__107_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__107_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__107_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__107_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__107_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__107_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__107_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__107_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__107_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__107_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__107_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__107_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__107_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__107_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__107_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__107_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__107_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__107_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__107_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__107_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__107_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__107_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__107_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__107_comb[6] | p3_actual_index__107_comb[7])}}) == 10'h000 & ((p3_actual_index__108_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__108_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__108_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__108_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__108_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__108_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__108_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__108_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__108_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__108_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__108_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__108_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__108_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__108_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__108_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__108_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__108_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__108_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__108_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__108_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__108_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__108_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__108_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__108_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__108_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__108_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__108_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__108_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__108_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__108_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__108_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__108_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__108_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__108_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__108_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__108_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__108_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__108_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__108_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__108_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__108_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__108_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__108_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__108_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__108_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__108_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__108_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__108_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__108_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__108_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__108_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__108_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__108_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__108_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__108_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__108_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__108_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__108_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__108_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__108_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__108_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__108_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__108_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12030_comb[4] | p3_add_12030_comb[5])}}) == 10'h000 & ((p3_actual_index__109_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__109_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__109_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__109_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__109_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__109_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__109_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__109_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__109_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__109_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__109_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__109_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__109_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__109_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__109_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__109_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__109_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__109_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__109_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__109_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__109_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__109_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__109_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__109_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__109_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__109_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__109_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__109_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__109_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__109_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__109_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__109_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__109_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__109_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__109_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__109_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__109_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__109_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__109_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__109_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__109_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__109_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__109_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__109_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__109_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__109_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__109_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__109_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__109_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__109_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__109_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__109_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__109_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__109_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__109_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__109_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__109_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__109_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__109_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__109_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__109_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__109_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__109_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__109_comb[6] | p3_actual_index__109_comb[7])}}) == 10'h000 & ((p3_actual_index__110_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__110_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__110_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__110_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__110_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__110_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__110_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__110_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__110_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__110_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__110_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__110_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__110_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__110_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__110_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__110_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__110_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__110_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__110_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__110_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__110_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__110_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__110_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__110_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__110_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__110_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__110_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__110_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__110_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__110_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__110_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__110_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__110_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__110_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__110_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__110_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__110_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__110_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__110_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__110_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__110_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__110_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__110_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__110_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__110_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__110_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__110_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__110_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__110_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__110_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__110_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__110_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__110_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__110_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__110_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__110_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__110_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__110_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__110_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__110_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__110_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__110_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__110_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12032_comb[5] | p3_add_12032_comb[6])}}) == 10'h000 & ((p3_actual_index__111_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__111_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__111_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__111_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__111_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__111_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__111_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__111_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__111_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__111_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__111_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__111_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__111_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__111_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__111_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__111_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__111_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__111_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__111_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__111_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__111_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__111_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__111_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__111_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__111_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__111_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__111_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__111_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__111_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__111_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__111_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__111_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__111_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__111_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__111_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__111_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__111_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__111_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__111_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__111_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__111_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__111_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__111_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__111_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__111_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__111_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__111_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__111_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__111_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__111_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__111_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__111_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__111_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__111_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__111_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__111_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__111_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__111_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__111_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__111_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__111_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__111_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__111_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__111_comb[6] | p3_actual_index__111_comb[7])}}) == 10'h000 & ((p3_actual_index__112_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__112_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__112_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__112_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__112_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__112_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__112_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__112_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__112_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__112_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__112_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__112_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__112_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__112_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__112_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__112_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__112_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__112_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__112_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__112_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__112_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__112_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__112_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__112_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__112_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__112_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__112_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__112_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__112_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__112_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__112_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__112_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__112_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__112_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__112_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__112_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__112_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__112_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__112_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__112_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__112_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__112_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__112_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__112_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__112_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__112_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__112_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__112_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__112_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__112_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__112_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__112_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__112_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__112_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__112_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__112_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__112_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__112_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__112_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__112_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__112_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__112_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__112_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12034_comb[2] | p3_add_12034_comb[3])}}) == 10'h000 & ((p3_actual_index__113_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__113_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__113_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__113_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__113_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__113_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__113_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__113_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__113_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__113_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__113_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__113_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__113_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__113_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__113_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__113_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__113_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__113_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__113_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__113_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__113_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__113_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__113_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__113_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__113_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__113_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__113_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__113_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__113_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__113_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__113_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__113_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__113_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__113_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__113_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__113_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__113_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__113_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__113_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__113_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__113_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__113_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__113_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__113_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__113_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__113_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__113_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__113_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__113_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__113_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__113_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__113_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__113_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__113_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__113_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__113_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__113_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__113_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__113_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__113_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__113_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__113_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__113_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__113_comb[6] | p3_actual_index__113_comb[7])}}) == 10'h000 & ((p3_actual_index__114_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__114_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__114_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__114_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__114_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__114_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__114_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__114_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__114_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__114_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__114_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__114_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__114_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__114_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__114_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__114_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__114_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__114_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__114_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__114_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__114_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__114_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__114_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__114_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__114_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__114_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__114_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__114_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__114_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__114_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__114_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__114_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__114_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__114_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__114_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__114_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__114_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__114_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__114_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__114_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__114_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__114_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__114_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__114_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__114_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__114_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__114_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__114_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__114_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__114_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__114_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__114_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__114_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__114_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__114_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__114_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__114_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__114_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__114_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__114_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__114_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__114_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__114_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12036_comb[5] | p3_add_12036_comb[6])}}) == 10'h000 & ((p3_actual_index__115_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__115_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__115_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__115_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__115_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__115_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__115_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__115_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__115_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__115_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__115_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__115_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__115_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__115_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__115_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__115_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__115_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__115_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__115_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__115_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__115_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__115_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__115_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__115_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__115_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__115_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__115_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__115_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__115_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__115_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__115_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__115_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__115_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__115_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__115_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__115_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__115_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__115_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__115_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__115_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__115_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__115_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__115_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__115_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__115_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__115_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__115_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__115_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__115_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__115_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__115_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__115_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__115_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__115_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__115_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__115_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__115_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__115_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__115_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__115_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__115_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__115_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__115_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__115_comb[6] | p3_actual_index__115_comb[7])}}) == 10'h000 & ((p3_actual_index__116_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__116_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__116_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__116_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__116_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__116_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__116_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__116_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__116_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__116_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__116_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__116_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__116_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__116_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__116_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__116_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__116_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__116_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__116_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__116_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__116_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__116_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__116_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__116_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__116_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__116_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__116_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__116_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__116_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__116_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__116_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__116_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__116_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__116_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__116_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__116_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__116_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__116_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__116_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__116_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__116_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__116_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__116_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__116_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__116_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__116_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__116_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__116_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__116_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__116_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__116_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__116_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__116_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__116_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__116_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__116_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__116_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__116_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__116_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__116_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__116_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__116_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__116_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12038_comb[4] | p3_add_12038_comb[5])}}) == 10'h000 & ((p3_actual_index__117_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__117_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__117_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__117_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__117_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__117_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__117_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__117_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__117_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__117_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__117_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__117_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__117_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__117_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__117_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__117_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__117_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__117_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__117_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__117_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__117_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__117_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__117_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__117_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__117_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__117_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__117_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__117_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__117_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__117_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__117_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__117_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__117_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__117_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__117_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__117_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__117_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__117_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__117_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__117_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__117_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__117_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__117_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__117_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__117_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__117_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__117_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__117_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__117_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__117_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__117_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__117_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__117_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__117_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__117_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__117_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__117_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__117_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__117_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__117_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__117_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__117_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__117_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__117_comb[6] | p3_actual_index__117_comb[7])}}) == 10'h000 & ((p3_actual_index__118_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__118_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__118_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__118_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__118_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__118_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__118_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__118_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__118_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__118_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__118_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__118_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__118_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__118_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__118_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__118_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__118_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__118_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__118_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__118_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__118_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__118_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__118_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__118_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__118_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__118_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__118_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__118_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__118_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__118_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__118_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__118_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__118_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__118_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__118_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__118_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__118_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__118_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__118_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__118_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__118_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__118_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__118_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__118_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__118_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__118_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__118_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__118_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__118_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__118_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__118_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__118_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__118_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__118_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__118_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__118_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__118_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__118_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__118_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__118_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__118_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__118_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__118_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12040_comb[5] | p3_add_12040_comb[6])}}) == 10'h000 & ((p3_actual_index__119_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__119_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__119_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__119_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__119_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__119_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__119_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__119_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__119_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__119_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__119_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__119_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__119_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__119_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__119_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__119_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__119_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__119_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__119_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__119_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__119_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__119_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__119_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__119_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__119_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__119_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__119_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__119_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__119_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__119_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__119_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__119_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__119_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__119_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__119_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__119_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__119_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__119_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__119_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__119_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__119_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__119_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__119_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__119_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__119_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__119_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__119_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__119_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__119_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__119_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__119_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__119_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__119_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__119_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__119_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__119_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__119_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__119_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__119_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__119_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__119_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__119_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__119_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__119_comb[6] | p3_actual_index__119_comb[7])}}) == 10'h000 & ((p3_actual_index__120_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__120_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__120_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__120_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__120_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__120_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__120_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__120_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__120_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__120_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__120_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__120_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__120_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__120_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__120_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__120_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__120_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__120_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__120_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__120_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__120_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__120_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__120_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__120_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__120_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__120_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__120_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__120_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__120_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__120_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__120_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__120_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__120_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__120_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__120_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__120_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__120_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__120_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__120_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__120_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__120_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__120_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__120_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__120_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__120_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__120_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__120_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__120_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__120_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__120_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__120_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__120_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__120_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__120_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__120_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__120_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__120_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__120_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__120_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__120_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__120_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__120_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__120_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12042_comb[3] | p3_add_12042_comb[4])}}) == 10'h000 & ((p3_actual_index__121_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__121_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__121_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__121_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__121_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__121_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__121_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__121_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__121_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__121_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__121_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__121_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__121_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__121_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__121_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__121_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__121_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__121_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__121_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__121_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__121_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__121_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__121_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__121_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__121_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__121_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__121_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__121_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__121_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__121_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__121_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__121_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__121_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__121_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__121_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__121_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__121_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__121_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__121_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__121_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__121_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__121_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__121_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__121_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__121_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__121_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__121_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__121_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__121_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__121_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__121_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__121_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__121_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__121_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__121_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__121_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__121_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__121_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__121_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__121_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__121_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__121_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__121_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__121_comb[6] | p3_actual_index__121_comb[7])}}) == 10'h000 & ((p3_actual_index__122_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__122_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__122_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__122_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__122_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__122_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__122_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__122_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__122_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__122_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__122_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__122_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__122_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__122_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__122_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__122_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__122_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__122_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__122_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__122_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__122_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__122_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__122_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__122_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__122_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__122_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__122_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__122_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__122_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__122_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__122_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__122_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__122_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__122_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__122_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__122_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__122_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__122_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__122_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__122_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__122_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__122_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__122_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__122_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__122_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__122_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__122_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__122_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__122_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__122_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__122_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__122_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__122_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__122_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__122_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__122_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__122_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__122_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__122_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__122_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__122_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__122_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__122_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12044_comb[5] | p3_add_12044_comb[6])}}) == 10'h000 & ((p3_actual_index__123_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__123_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__123_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__123_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__123_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__123_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__123_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__123_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__123_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__123_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__123_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__123_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__123_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__123_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__123_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__123_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__123_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__123_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__123_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__123_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__123_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__123_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__123_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__123_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__123_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__123_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__123_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__123_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__123_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__123_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__123_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__123_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__123_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__123_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__123_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__123_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__123_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__123_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__123_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__123_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__123_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__123_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__123_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__123_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__123_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__123_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__123_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__123_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__123_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__123_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__123_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__123_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__123_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__123_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__123_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__123_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__123_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__123_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__123_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__123_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__123_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__123_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__123_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__123_comb[6] | p3_actual_index__123_comb[7])}}) == 10'h000 & ((p3_actual_index__124_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__124_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__124_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__124_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__124_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__124_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__124_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__124_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__124_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__124_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__124_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__124_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__124_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__124_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__124_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__124_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__124_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__124_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__124_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__124_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__124_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__124_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__124_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__124_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__124_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__124_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__124_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__124_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__124_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__124_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__124_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__124_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__124_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__124_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__124_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__124_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__124_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__124_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__124_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__124_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__124_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__124_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__124_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__124_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__124_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__124_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__124_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__124_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__124_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__124_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__124_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__124_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__124_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__124_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__124_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__124_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__124_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__124_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__124_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__124_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__124_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__124_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__124_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12046_comb[4] | p3_add_12046_comb[5])}}) == 10'h000 & ((p3_actual_index__125_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__125_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__125_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__125_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__125_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__125_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__125_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__125_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__125_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__125_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__125_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__125_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__125_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__125_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__125_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__125_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__125_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__125_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__125_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__125_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__125_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__125_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__125_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__125_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__125_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__125_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__125_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__125_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__125_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__125_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__125_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__125_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__125_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__125_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__125_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__125_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__125_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__125_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__125_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__125_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__125_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__125_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__125_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__125_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__125_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__125_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__125_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__125_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__125_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__125_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__125_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__125_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__125_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__125_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__125_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__125_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__125_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__125_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__125_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__125_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__125_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__125_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__125_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__125_comb[6] | p3_actual_index__125_comb[7])}}) == 10'h000 & ((p3_actual_index__126_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__126_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__126_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__126_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__126_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__126_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__126_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__126_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__126_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__126_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__126_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__126_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__126_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__126_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__126_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__126_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__126_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__126_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__126_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__126_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__126_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__126_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__126_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__126_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__126_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__126_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__126_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__126_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__126_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__126_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__126_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__126_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__126_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__126_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__126_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__126_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__126_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__126_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__126_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__126_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__126_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__126_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__126_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__126_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__126_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__126_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__126_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__126_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__126_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__126_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__126_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__126_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__126_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__126_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__126_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__126_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__126_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__126_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__126_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__126_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__126_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__126_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__126_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_add_12048_comb[5] | p3_add_12048_comb[6])}}) == 10'h000 & ((p3_actual_index__127_comb == 8'h00 ? p2_array_index_11336 : (p3_actual_index__127_comb == 8'h01 ? p2_array_index_11337 : (p3_actual_index__127_comb == 8'h02 ? p2_array_index_11338 : (p3_actual_index__127_comb == 8'h03 ? p2_array_index_11339 : (p3_actual_index__127_comb == 8'h04 ? p2_array_index_11340 : (p3_actual_index__127_comb == 8'h05 ? p2_array_index_11341 : (p3_actual_index__127_comb == 8'h06 ? p2_array_index_11342 : (p3_actual_index__127_comb == 8'h07 ? p2_array_index_11343 : (p3_actual_index__127_comb == 8'h08 ? p2_array_index_11344 : (p3_actual_index__127_comb == 8'h09 ? p2_array_index_11345 : (p3_actual_index__127_comb == 8'h0a ? p2_array_index_11346 : (p3_actual_index__127_comb == 8'h0b ? p2_array_index_11347 : (p3_actual_index__127_comb == 8'h0c ? p2_array_index_11348 : (p3_actual_index__127_comb == 8'h0d ? p2_array_index_11349 : (p3_actual_index__127_comb == 8'h0e ? p2_array_index_11350 : (p3_actual_index__127_comb == 8'h0f ? p2_array_index_11351 : (p3_actual_index__127_comb == 8'h10 ? p2_array_index_11352 : (p3_actual_index__127_comb == 8'h11 ? p2_array_index_11353 : (p3_actual_index__127_comb == 8'h12 ? p2_array_index_11354 : (p3_actual_index__127_comb == 8'h13 ? p2_array_index_11355 : (p3_actual_index__127_comb == 8'h14 ? p2_array_index_11356 : (p3_actual_index__127_comb == 8'h15 ? p2_array_index_11357 : (p3_actual_index__127_comb == 8'h16 ? p2_array_index_11358 : (p3_actual_index__127_comb == 8'h17 ? p2_array_index_11359 : (p3_actual_index__127_comb == 8'h18 ? p2_array_index_11360 : (p3_actual_index__127_comb == 8'h19 ? p2_array_index_11361 : (p3_actual_index__127_comb == 8'h1a ? p2_array_index_11362 : (p3_actual_index__127_comb == 8'h1b ? p2_array_index_11363 : (p3_actual_index__127_comb == 8'h1c ? p2_array_index_11364 : (p3_actual_index__127_comb == 8'h1d ? p2_array_index_11365 : (p3_actual_index__127_comb == 8'h1e ? p2_array_index_11366 : (p3_actual_index__127_comb == 8'h1f ? p2_array_index_11367 : (p3_actual_index__127_comb == 8'h20 ? p2_array_index_11368 : (p3_actual_index__127_comb == 8'h21 ? p2_array_index_11369 : (p3_actual_index__127_comb == 8'h22 ? p2_array_index_11370 : (p3_actual_index__127_comb == 8'h23 ? p2_array_index_11371 : (p3_actual_index__127_comb == 8'h24 ? p2_array_index_11372 : (p3_actual_index__127_comb == 8'h25 ? p2_array_index_11373 : (p3_actual_index__127_comb == 8'h26 ? p2_array_index_11374 : (p3_actual_index__127_comb == 8'h27 ? p2_array_index_11375 : (p3_actual_index__127_comb == 8'h28 ? p2_array_index_11376 : (p3_actual_index__127_comb == 8'h29 ? p2_array_index_11377 : (p3_actual_index__127_comb == 8'h2a ? p2_array_index_11378 : (p3_actual_index__127_comb == 8'h2b ? p2_array_index_11379 : (p3_actual_index__127_comb == 8'h2c ? p2_array_index_11380 : (p3_actual_index__127_comb == 8'h2d ? p2_array_index_11381 : (p3_actual_index__127_comb == 8'h2e ? p2_array_index_11382 : (p3_actual_index__127_comb == 8'h2f ? p2_array_index_11383 : (p3_actual_index__127_comb == 8'h30 ? p2_array_index_11384 : (p3_actual_index__127_comb == 8'h31 ? p2_array_index_11385 : (p3_actual_index__127_comb == 8'h32 ? p2_array_index_11386 : (p3_actual_index__127_comb == 8'h33 ? p2_array_index_11387 : (p3_actual_index__127_comb == 8'h34 ? p2_array_index_11388 : (p3_actual_index__127_comb == 8'h35 ? p2_array_index_11389 : (p3_actual_index__127_comb == 8'h36 ? p2_array_index_11390 : (p3_actual_index__127_comb == 8'h37 ? p2_array_index_11391 : (p3_actual_index__127_comb == 8'h38 ? p2_array_index_11392 : (p3_actual_index__127_comb == 8'h39 ? p2_array_index_11393 : (p3_actual_index__127_comb == 8'h3a ? p2_array_index_11394 : (p3_actual_index__127_comb == 8'h3b ? p2_array_index_11395 : (p3_actual_index__127_comb == 8'h3c ? p2_array_index_11396 : (p3_actual_index__127_comb == 8'h3d ? p2_array_index_11397 : (p3_actual_index__127_comb == 8'h3e ? p2_array_index_11398 : p2_array_index_11399))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) & {10{~(p3_actual_index__127_comb[6] | p3_actual_index__127_comb[7])}}) == 10'h000;
  assign p3_next_pix__1_squeezed_squeezed_const_msb_bits__1_comb = 1'h0;
  assign p3_flipped_comb = ~p3_bin_value_comb;
  assign p3_Code_list_comb = $signed(p3_value__1_comb) <= $signed(10'h000) ? p3_flipped_comb : p3_bin_value__1_comb;
  assign p3_or_reduce_11910_comb = |p3_value_abs_comb[7:4];
  assign p3_sel_11911_comb = |p3_value_abs_comb[7:3] ? 3'h4 : {p3_next_pix__1_squeezed_squeezed_const_msb_bits__1_comb, |p3_value_abs_comb[7:2] ? 2'h3 : (|p3_value_abs_comb[7:1] ? 2'h2 : 2'h1)};
  assign p3_or_reduce_11914_comb = |p3_value_abs_comb[7:5];
  assign p3_bit_slice_11983_comb = p3_value_pix_num_comb[4];
  assign p3_value_pix_num_squeezed_comb = p3_value_pix_num_comb[4:0];
  assign p3_or_reduce_11986_comb = |p3_value_abs_comb[7:6];
  assign p3_bit_slice_12183_comb = p3_value_abs_comb[7];
  assign p3_eq_12184_comb = p3_value_abs_comb == 8'h00;
  assign p3_code_list_comb = p3_Code_list_comb & {8{~p3_and_12599_comb}};

  // Registers for pipe stage 3:
  reg p3_is_luminance;
  reg p3_or_reduce_11910;
  reg [2:0] p3_sel_11911;
  reg p3_or_reduce_11914;
  reg p3_bit_slice_11983;
  reg [4:0] p3_value_pix_num_squeezed;
  reg [9:0] p3_value;
  reg p3_or_reduce_11986;
  reg p3_bit_slice_12183;
  reg p3_eq_12184;
  reg p3_and_12599;
  reg [7:0] p3_code_list;
  always @ (posedge clk) begin
    p3_is_luminance <= p2_is_luminance;
    p3_or_reduce_11910 <= p3_or_reduce_11910_comb;
    p3_sel_11911 <= p3_sel_11911_comb;
    p3_or_reduce_11914 <= p3_or_reduce_11914_comb;
    p3_bit_slice_11983 <= p3_bit_slice_11983_comb;
    p3_value_pix_num_squeezed <= p3_value_pix_num_squeezed_comb;
    p3_value <= p3_value_comb;
    p3_or_reduce_11986 <= p3_or_reduce_11986_comb;
    p3_bit_slice_12183 <= p3_bit_slice_12183_comb;
    p3_eq_12184 <= p3_eq_12184_comb;
    p3_and_12599 <= p3_and_12599_comb;
    p3_code_list <= p3_code_list_comb;
  end

  // ===== Pipe stage 4:
  wire [2:0] p4_run_0_squeezed_const_msb_bits__17_comb;
  wire [4:0] p4_run_0_squeezed_comb;
  wire p4_eq_12640_comb;
  wire p4_next_pix__1_squeezed_squeezed_const_msb_bits__2_comb;
  wire [7:0] p4_run_0_comb;
  wire [7:0] p4_run__1_comb;
  wire [3:0] p4_sel_12649_comb;
  wire [7:0] p4_concat_12654_comb;
  wire [4:0] p4_next_pix_0_squeezed__1_comb;
  wire [7:0] p4_Code_size_comb;
  wire [4:0] p4_next_pix_1_squeezed_squeezed_comb;
  wire [7:0] p4_run_size_str_u8_comb;
  wire [2:0] p4_sel_12673_comb;
  wire [1:0] p4_next_pix_squeezed_const_msb_bits_comb;
  wire p4_next_pix__1_squeezed_squeezed_const_msb_bits__3_comb;
  wire p4_next_pix__1_squeezed_squeezed_const_msb_bits__8_comb;
  wire [4:0] p4_next_pix__1_squeezed_squeezed_comb;
  wire [4:0] p4_Huffman_length_squeezed_comb;
  wire [5:0] p4_next_pix__1_squeezed_comb;
  wire [5:0] p4_run__1_squeezed_comb;
  wire [15:0] p4_Huffman_code_full_comb;
  wire [2:0] p4_run_0_squeezed_const_msb_bits__18_comb;
  wire [4:0] p4_huff_length_squeezed_comb;
  wire [1:0] p4_next_pix_squeezed_const_msb_bits__1_comb;
  wire [5:0] p4_next_pix_squeezed_comb;
  wire [1:0] p4_next_pix_squeezed_const_msb_bits__2_comb;
  wire [5:0] p4_run_squeezed_comb;
  wire [15:0] p4_huff_code_comb;
  wire [7:0] p4_huff_length_comb;
  wire [7:0] p4_code_size_comb;
  wire [7:0] p4_next_pix_comb;
  wire [7:0] p4_run_comb;
  wire [65:0] p4_tuple_12707_comb;
  assign p4_run_0_squeezed_const_msb_bits__17_comb = 3'h0;
  assign p4_run_0_squeezed_comb = p3_bit_slice_11983 ? 5'h0f : p3_value_pix_num_squeezed;
  assign p4_eq_12640_comb = p3_value == 10'h000;
  assign p4_next_pix__1_squeezed_squeezed_const_msb_bits__2_comb = 1'h0;
  assign p4_run_0_comb = {p4_run_0_squeezed_const_msb_bits__17_comb, p4_run_0_squeezed_comb};
  assign p4_run__1_comb = p4_run_0_comb & {8{p4_eq_12640_comb}};
  assign p4_sel_12649_comb = p3_bit_slice_12183 ? 4'h8 : {p4_next_pix__1_squeezed_squeezed_const_msb_bits__2_comb, p3_or_reduce_11986 ? 3'h7 : (p3_or_reduce_11914 ? 3'h6 : (p3_or_reduce_11910 ? 3'h5 : p3_sel_11911))};
  assign p4_concat_12654_comb = {4'h0, p4_sel_12649_comb};
  assign p4_next_pix_0_squeezed__1_comb = p3_value_pix_num_squeezed + 5'h01;
  assign p4_Code_size_comb = p4_concat_12654_comb & {8{~p3_eq_12184}};
  assign p4_next_pix_1_squeezed_squeezed_comb = p4_eq_12640_comb ? p4_next_pix_0_squeezed__1_comb : 5'h01;
  assign p4_run_size_str_u8_comb = {p4_run__1_comb[3:0], 4'h0} | p4_Code_size_comb;
  assign p4_sel_12673_comb = p3_is_luminance ? 3'h4 : 3'h1;
  assign p4_next_pix_squeezed_const_msb_bits_comb = 2'h0;
  assign p4_next_pix__1_squeezed_squeezed_const_msb_bits__3_comb = 1'h0;
  assign p4_next_pix__1_squeezed_squeezed_const_msb_bits__8_comb = 1'h0;
  assign p4_next_pix__1_squeezed_squeezed_comb = p4_next_pix_1_squeezed_squeezed_comb > 5'h10 ? 5'h10 : p4_next_pix_1_squeezed_squeezed_comb;
  assign p4_Huffman_length_squeezed_comb = p3_is_luminance ? literal_12666[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_12664[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_next_pix__1_squeezed_comb = {p4_next_pix__1_squeezed_squeezed_const_msb_bits__8_comb, p4_next_pix__1_squeezed_squeezed_comb};
  assign p4_run__1_squeezed_comb = p4_run__1_comb[5:0];
  assign p4_Huffman_code_full_comb = p3_is_luminance ? literal_12672[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_12671[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_run_0_squeezed_const_msb_bits__18_comb = 3'h0;
  assign p4_huff_length_squeezed_comb = p3_and_12599 ? {p4_next_pix_squeezed_const_msb_bits_comb, p3_is_luminance ? 2'h2 : 2'h1, p4_next_pix__1_squeezed_squeezed_const_msb_bits__3_comb} : p4_Huffman_length_squeezed_comb;
  assign p4_next_pix_squeezed_const_msb_bits__1_comb = 2'h0;
  assign p4_next_pix_squeezed_comb = p3_and_12599 ? 6'h3f : p4_next_pix__1_squeezed_comb;
  assign p4_next_pix_squeezed_const_msb_bits__2_comb = 2'h0;
  assign p4_run_squeezed_comb = p3_and_12599 ? 6'h3f : p4_run__1_squeezed_comb;
  assign p4_huff_code_comb = p3_and_12599 ? {12'h000, {{1{p4_sel_12673_comb[2]}}, p4_sel_12673_comb}} : p4_Huffman_code_full_comb;
  assign p4_huff_length_comb = {p4_run_0_squeezed_const_msb_bits__18_comb, p4_huff_length_squeezed_comb};
  assign p4_code_size_comb = p4_concat_12654_comb & {8{~(p3_and_12599 | p3_eq_12184)}};
  assign p4_next_pix_comb = {p4_next_pix_squeezed_const_msb_bits__1_comb, p4_next_pix_squeezed_comb};
  assign p4_run_comb = {p4_next_pix_squeezed_const_msb_bits__2_comb, p4_run_squeezed_comb};
  assign p4_tuple_12707_comb = {p4_huff_code_comb, p4_huff_length_comb, p3_code_list, p4_code_size_comb, p4_next_pix_comb, p4_run_comb, p3_value};

  // Registers for pipe stage 4:
  reg [65:0] p4_tuple_12707;
  always @ (posedge clk) begin
    p4_tuple_12707 <= p4_tuple_12707_comb;
  end
  assign out = p4_tuple_12707;
endmodule
