module Huffman_ACenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire [7:0] start_pix,
  input wire [7:0] pre_start_pix,
  input wire is_luminance,
  output wire [65:0] out
);
  wire [4:0] literal_11597[0:251];
  assign literal_11597[0] = 5'h02;
  assign literal_11597[1] = 5'h02;
  assign literal_11597[2] = 5'h03;
  assign literal_11597[3] = 5'h04;
  assign literal_11597[4] = 5'h05;
  assign literal_11597[5] = 5'h07;
  assign literal_11597[6] = 5'h08;
  assign literal_11597[7] = 5'h0e;
  assign literal_11597[8] = 5'h10;
  assign literal_11597[9] = 5'h10;
  assign literal_11597[10] = 5'h10;
  assign literal_11597[11] = 5'h00;
  assign literal_11597[12] = 5'h00;
  assign literal_11597[13] = 5'h00;
  assign literal_11597[14] = 5'h00;
  assign literal_11597[15] = 5'h00;
  assign literal_11597[16] = 5'h00;
  assign literal_11597[17] = 5'h03;
  assign literal_11597[18] = 5'h06;
  assign literal_11597[19] = 5'h07;
  assign literal_11597[20] = 5'h09;
  assign literal_11597[21] = 5'h0b;
  assign literal_11597[22] = 5'h0d;
  assign literal_11597[23] = 5'h10;
  assign literal_11597[24] = 5'h10;
  assign literal_11597[25] = 5'h10;
  assign literal_11597[26] = 5'h10;
  assign literal_11597[27] = 5'h00;
  assign literal_11597[28] = 5'h00;
  assign literal_11597[29] = 5'h00;
  assign literal_11597[30] = 5'h00;
  assign literal_11597[31] = 5'h00;
  assign literal_11597[32] = 5'h00;
  assign literal_11597[33] = 5'h05;
  assign literal_11597[34] = 5'h07;
  assign literal_11597[35] = 5'h0a;
  assign literal_11597[36] = 5'h0c;
  assign literal_11597[37] = 5'h0d;
  assign literal_11597[38] = 5'h10;
  assign literal_11597[39] = 5'h10;
  assign literal_11597[40] = 5'h10;
  assign literal_11597[41] = 5'h10;
  assign literal_11597[42] = 5'h10;
  assign literal_11597[43] = 5'h00;
  assign literal_11597[44] = 5'h00;
  assign literal_11597[45] = 5'h00;
  assign literal_11597[46] = 5'h00;
  assign literal_11597[47] = 5'h00;
  assign literal_11597[48] = 5'h00;
  assign literal_11597[49] = 5'h06;
  assign literal_11597[50] = 5'h08;
  assign literal_11597[51] = 5'h0b;
  assign literal_11597[52] = 5'h0c;
  assign literal_11597[53] = 5'h0f;
  assign literal_11597[54] = 5'h10;
  assign literal_11597[55] = 5'h10;
  assign literal_11597[56] = 5'h10;
  assign literal_11597[57] = 5'h10;
  assign literal_11597[58] = 5'h10;
  assign literal_11597[59] = 5'h00;
  assign literal_11597[60] = 5'h00;
  assign literal_11597[61] = 5'h00;
  assign literal_11597[62] = 5'h00;
  assign literal_11597[63] = 5'h00;
  assign literal_11597[64] = 5'h00;
  assign literal_11597[65] = 5'h06;
  assign literal_11597[66] = 5'h0a;
  assign literal_11597[67] = 5'h0c;
  assign literal_11597[68] = 5'h0f;
  assign literal_11597[69] = 5'h10;
  assign literal_11597[70] = 5'h10;
  assign literal_11597[71] = 5'h10;
  assign literal_11597[72] = 5'h10;
  assign literal_11597[73] = 5'h10;
  assign literal_11597[74] = 5'h10;
  assign literal_11597[75] = 5'h00;
  assign literal_11597[76] = 5'h00;
  assign literal_11597[77] = 5'h00;
  assign literal_11597[78] = 5'h00;
  assign literal_11597[79] = 5'h00;
  assign literal_11597[80] = 5'h00;
  assign literal_11597[81] = 5'h07;
  assign literal_11597[82] = 5'h0b;
  assign literal_11597[83] = 5'h0d;
  assign literal_11597[84] = 5'h10;
  assign literal_11597[85] = 5'h10;
  assign literal_11597[86] = 5'h10;
  assign literal_11597[87] = 5'h10;
  assign literal_11597[88] = 5'h10;
  assign literal_11597[89] = 5'h10;
  assign literal_11597[90] = 5'h10;
  assign literal_11597[91] = 5'h00;
  assign literal_11597[92] = 5'h00;
  assign literal_11597[93] = 5'h00;
  assign literal_11597[94] = 5'h00;
  assign literal_11597[95] = 5'h00;
  assign literal_11597[96] = 5'h00;
  assign literal_11597[97] = 5'h07;
  assign literal_11597[98] = 5'h0b;
  assign literal_11597[99] = 5'h0d;
  assign literal_11597[100] = 5'h10;
  assign literal_11597[101] = 5'h10;
  assign literal_11597[102] = 5'h10;
  assign literal_11597[103] = 5'h10;
  assign literal_11597[104] = 5'h10;
  assign literal_11597[105] = 5'h10;
  assign literal_11597[106] = 5'h10;
  assign literal_11597[107] = 5'h00;
  assign literal_11597[108] = 5'h00;
  assign literal_11597[109] = 5'h00;
  assign literal_11597[110] = 5'h00;
  assign literal_11597[111] = 5'h00;
  assign literal_11597[112] = 5'h00;
  assign literal_11597[113] = 5'h08;
  assign literal_11597[114] = 5'h0b;
  assign literal_11597[115] = 5'h0e;
  assign literal_11597[116] = 5'h10;
  assign literal_11597[117] = 5'h10;
  assign literal_11597[118] = 5'h10;
  assign literal_11597[119] = 5'h10;
  assign literal_11597[120] = 5'h10;
  assign literal_11597[121] = 5'h10;
  assign literal_11597[122] = 5'h10;
  assign literal_11597[123] = 5'h00;
  assign literal_11597[124] = 5'h00;
  assign literal_11597[125] = 5'h00;
  assign literal_11597[126] = 5'h00;
  assign literal_11597[127] = 5'h00;
  assign literal_11597[128] = 5'h00;
  assign literal_11597[129] = 5'h08;
  assign literal_11597[130] = 5'h0c;
  assign literal_11597[131] = 5'h10;
  assign literal_11597[132] = 5'h10;
  assign literal_11597[133] = 5'h10;
  assign literal_11597[134] = 5'h10;
  assign literal_11597[135] = 5'h10;
  assign literal_11597[136] = 5'h10;
  assign literal_11597[137] = 5'h10;
  assign literal_11597[138] = 5'h10;
  assign literal_11597[139] = 5'h00;
  assign literal_11597[140] = 5'h00;
  assign literal_11597[141] = 5'h00;
  assign literal_11597[142] = 5'h00;
  assign literal_11597[143] = 5'h00;
  assign literal_11597[144] = 5'h00;
  assign literal_11597[145] = 5'h08;
  assign literal_11597[146] = 5'h0d;
  assign literal_11597[147] = 5'h10;
  assign literal_11597[148] = 5'h10;
  assign literal_11597[149] = 5'h10;
  assign literal_11597[150] = 5'h10;
  assign literal_11597[151] = 5'h10;
  assign literal_11597[152] = 5'h10;
  assign literal_11597[153] = 5'h10;
  assign literal_11597[154] = 5'h10;
  assign literal_11597[155] = 5'h00;
  assign literal_11597[156] = 5'h00;
  assign literal_11597[157] = 5'h00;
  assign literal_11597[158] = 5'h00;
  assign literal_11597[159] = 5'h00;
  assign literal_11597[160] = 5'h00;
  assign literal_11597[161] = 5'h09;
  assign literal_11597[162] = 5'h0d;
  assign literal_11597[163] = 5'h10;
  assign literal_11597[164] = 5'h10;
  assign literal_11597[165] = 5'h10;
  assign literal_11597[166] = 5'h10;
  assign literal_11597[167] = 5'h10;
  assign literal_11597[168] = 5'h10;
  assign literal_11597[169] = 5'h10;
  assign literal_11597[170] = 5'h10;
  assign literal_11597[171] = 5'h00;
  assign literal_11597[172] = 5'h00;
  assign literal_11597[173] = 5'h00;
  assign literal_11597[174] = 5'h00;
  assign literal_11597[175] = 5'h00;
  assign literal_11597[176] = 5'h00;
  assign literal_11597[177] = 5'h09;
  assign literal_11597[178] = 5'h0d;
  assign literal_11597[179] = 5'h10;
  assign literal_11597[180] = 5'h10;
  assign literal_11597[181] = 5'h10;
  assign literal_11597[182] = 5'h10;
  assign literal_11597[183] = 5'h10;
  assign literal_11597[184] = 5'h10;
  assign literal_11597[185] = 5'h10;
  assign literal_11597[186] = 5'h10;
  assign literal_11597[187] = 5'h00;
  assign literal_11597[188] = 5'h00;
  assign literal_11597[189] = 5'h00;
  assign literal_11597[190] = 5'h00;
  assign literal_11597[191] = 5'h00;
  assign literal_11597[192] = 5'h00;
  assign literal_11597[193] = 5'h0a;
  assign literal_11597[194] = 5'h0d;
  assign literal_11597[195] = 5'h10;
  assign literal_11597[196] = 5'h10;
  assign literal_11597[197] = 5'h10;
  assign literal_11597[198] = 5'h10;
  assign literal_11597[199] = 5'h10;
  assign literal_11597[200] = 5'h10;
  assign literal_11597[201] = 5'h10;
  assign literal_11597[202] = 5'h10;
  assign literal_11597[203] = 5'h00;
  assign literal_11597[204] = 5'h00;
  assign literal_11597[205] = 5'h00;
  assign literal_11597[206] = 5'h00;
  assign literal_11597[207] = 5'h00;
  assign literal_11597[208] = 5'h00;
  assign literal_11597[209] = 5'h0a;
  assign literal_11597[210] = 5'h0e;
  assign literal_11597[211] = 5'h10;
  assign literal_11597[212] = 5'h10;
  assign literal_11597[213] = 5'h10;
  assign literal_11597[214] = 5'h10;
  assign literal_11597[215] = 5'h10;
  assign literal_11597[216] = 5'h10;
  assign literal_11597[217] = 5'h10;
  assign literal_11597[218] = 5'h10;
  assign literal_11597[219] = 5'h00;
  assign literal_11597[220] = 5'h00;
  assign literal_11597[221] = 5'h00;
  assign literal_11597[222] = 5'h00;
  assign literal_11597[223] = 5'h00;
  assign literal_11597[224] = 5'h00;
  assign literal_11597[225] = 5'h0a;
  assign literal_11597[226] = 5'h0f;
  assign literal_11597[227] = 5'h10;
  assign literal_11597[228] = 5'h10;
  assign literal_11597[229] = 5'h10;
  assign literal_11597[230] = 5'h10;
  assign literal_11597[231] = 5'h10;
  assign literal_11597[232] = 5'h10;
  assign literal_11597[233] = 5'h10;
  assign literal_11597[234] = 5'h10;
  assign literal_11597[235] = 5'h00;
  assign literal_11597[236] = 5'h00;
  assign literal_11597[237] = 5'h00;
  assign literal_11597[238] = 5'h00;
  assign literal_11597[239] = 5'h00;
  assign literal_11597[240] = 5'h09;
  assign literal_11597[241] = 5'h0b;
  assign literal_11597[242] = 5'h10;
  assign literal_11597[243] = 5'h10;
  assign literal_11597[244] = 5'h10;
  assign literal_11597[245] = 5'h10;
  assign literal_11597[246] = 5'h10;
  assign literal_11597[247] = 5'h10;
  assign literal_11597[248] = 5'h10;
  assign literal_11597[249] = 5'h10;
  assign literal_11597[250] = 5'h10;
  assign literal_11597[251] = 5'h00;
  wire [4:0] literal_11599[0:251];
  assign literal_11599[0] = 5'h04;
  assign literal_11599[1] = 5'h02;
  assign literal_11599[2] = 5'h02;
  assign literal_11599[3] = 5'h03;
  assign literal_11599[4] = 5'h04;
  assign literal_11599[5] = 5'h05;
  assign literal_11599[6] = 5'h07;
  assign literal_11599[7] = 5'h09;
  assign literal_11599[8] = 5'h10;
  assign literal_11599[9] = 5'h10;
  assign literal_11599[10] = 5'h10;
  assign literal_11599[11] = 5'h00;
  assign literal_11599[12] = 5'h00;
  assign literal_11599[13] = 5'h00;
  assign literal_11599[14] = 5'h00;
  assign literal_11599[15] = 5'h00;
  assign literal_11599[16] = 5'h00;
  assign literal_11599[17] = 5'h04;
  assign literal_11599[18] = 5'h05;
  assign literal_11599[19] = 5'h07;
  assign literal_11599[20] = 5'h09;
  assign literal_11599[21] = 5'h0a;
  assign literal_11599[22] = 5'h0b;
  assign literal_11599[23] = 5'h10;
  assign literal_11599[24] = 5'h10;
  assign literal_11599[25] = 5'h10;
  assign literal_11599[26] = 5'h10;
  assign literal_11599[27] = 5'h00;
  assign literal_11599[28] = 5'h00;
  assign literal_11599[29] = 5'h00;
  assign literal_11599[30] = 5'h00;
  assign literal_11599[31] = 5'h00;
  assign literal_11599[32] = 5'h00;
  assign literal_11599[33] = 5'h05;
  assign literal_11599[34] = 5'h08;
  assign literal_11599[35] = 5'h0a;
  assign literal_11599[36] = 5'h0c;
  assign literal_11599[37] = 5'h0e;
  assign literal_11599[38] = 5'h10;
  assign literal_11599[39] = 5'h10;
  assign literal_11599[40] = 5'h10;
  assign literal_11599[41] = 5'h10;
  assign literal_11599[42] = 5'h10;
  assign literal_11599[43] = 5'h00;
  assign literal_11599[44] = 5'h00;
  assign literal_11599[45] = 5'h00;
  assign literal_11599[46] = 5'h00;
  assign literal_11599[47] = 5'h00;
  assign literal_11599[48] = 5'h00;
  assign literal_11599[49] = 5'h06;
  assign literal_11599[50] = 5'h09;
  assign literal_11599[51] = 5'h0b;
  assign literal_11599[52] = 5'h0e;
  assign literal_11599[53] = 5'h10;
  assign literal_11599[54] = 5'h10;
  assign literal_11599[55] = 5'h10;
  assign literal_11599[56] = 5'h10;
  assign literal_11599[57] = 5'h10;
  assign literal_11599[58] = 5'h10;
  assign literal_11599[59] = 5'h00;
  assign literal_11599[60] = 5'h00;
  assign literal_11599[61] = 5'h00;
  assign literal_11599[62] = 5'h00;
  assign literal_11599[63] = 5'h00;
  assign literal_11599[64] = 5'h00;
  assign literal_11599[65] = 5'h06;
  assign literal_11599[66] = 5'h0a;
  assign literal_11599[67] = 5'h0e;
  assign literal_11599[68] = 5'h10;
  assign literal_11599[69] = 5'h10;
  assign literal_11599[70] = 5'h10;
  assign literal_11599[71] = 5'h10;
  assign literal_11599[72] = 5'h10;
  assign literal_11599[73] = 5'h10;
  assign literal_11599[74] = 5'h10;
  assign literal_11599[75] = 5'h00;
  assign literal_11599[76] = 5'h00;
  assign literal_11599[77] = 5'h00;
  assign literal_11599[78] = 5'h00;
  assign literal_11599[79] = 5'h00;
  assign literal_11599[80] = 5'h00;
  assign literal_11599[81] = 5'h07;
  assign literal_11599[82] = 5'h0a;
  assign literal_11599[83] = 5'h0e;
  assign literal_11599[84] = 5'h10;
  assign literal_11599[85] = 5'h10;
  assign literal_11599[86] = 5'h10;
  assign literal_11599[87] = 5'h10;
  assign literal_11599[88] = 5'h10;
  assign literal_11599[89] = 5'h10;
  assign literal_11599[90] = 5'h10;
  assign literal_11599[91] = 5'h00;
  assign literal_11599[92] = 5'h00;
  assign literal_11599[93] = 5'h00;
  assign literal_11599[94] = 5'h00;
  assign literal_11599[95] = 5'h00;
  assign literal_11599[96] = 5'h00;
  assign literal_11599[97] = 5'h07;
  assign literal_11599[98] = 5'h0c;
  assign literal_11599[99] = 5'h0f;
  assign literal_11599[100] = 5'h10;
  assign literal_11599[101] = 5'h10;
  assign literal_11599[102] = 5'h10;
  assign literal_11599[103] = 5'h10;
  assign literal_11599[104] = 5'h10;
  assign literal_11599[105] = 5'h10;
  assign literal_11599[106] = 5'h10;
  assign literal_11599[107] = 5'h00;
  assign literal_11599[108] = 5'h00;
  assign literal_11599[109] = 5'h00;
  assign literal_11599[110] = 5'h00;
  assign literal_11599[111] = 5'h00;
  assign literal_11599[112] = 5'h00;
  assign literal_11599[113] = 5'h08;
  assign literal_11599[114] = 5'h0c;
  assign literal_11599[115] = 5'h10;
  assign literal_11599[116] = 5'h10;
  assign literal_11599[117] = 5'h10;
  assign literal_11599[118] = 5'h10;
  assign literal_11599[119] = 5'h10;
  assign literal_11599[120] = 5'h10;
  assign literal_11599[121] = 5'h10;
  assign literal_11599[122] = 5'h10;
  assign literal_11599[123] = 5'h00;
  assign literal_11599[124] = 5'h00;
  assign literal_11599[125] = 5'h00;
  assign literal_11599[126] = 5'h00;
  assign literal_11599[127] = 5'h00;
  assign literal_11599[128] = 5'h00;
  assign literal_11599[129] = 5'h09;
  assign literal_11599[130] = 5'h0d;
  assign literal_11599[131] = 5'h10;
  assign literal_11599[132] = 5'h10;
  assign literal_11599[133] = 5'h10;
  assign literal_11599[134] = 5'h10;
  assign literal_11599[135] = 5'h10;
  assign literal_11599[136] = 5'h10;
  assign literal_11599[137] = 5'h10;
  assign literal_11599[138] = 5'h10;
  assign literal_11599[139] = 5'h00;
  assign literal_11599[140] = 5'h00;
  assign literal_11599[141] = 5'h00;
  assign literal_11599[142] = 5'h00;
  assign literal_11599[143] = 5'h00;
  assign literal_11599[144] = 5'h00;
  assign literal_11599[145] = 5'h09;
  assign literal_11599[146] = 5'h0e;
  assign literal_11599[147] = 5'h10;
  assign literal_11599[148] = 5'h10;
  assign literal_11599[149] = 5'h10;
  assign literal_11599[150] = 5'h10;
  assign literal_11599[151] = 5'h10;
  assign literal_11599[152] = 5'h10;
  assign literal_11599[153] = 5'h10;
  assign literal_11599[154] = 5'h10;
  assign literal_11599[155] = 5'h00;
  assign literal_11599[156] = 5'h00;
  assign literal_11599[157] = 5'h00;
  assign literal_11599[158] = 5'h00;
  assign literal_11599[159] = 5'h00;
  assign literal_11599[160] = 5'h00;
  assign literal_11599[161] = 5'h09;
  assign literal_11599[162] = 5'h0e;
  assign literal_11599[163] = 5'h10;
  assign literal_11599[164] = 5'h10;
  assign literal_11599[165] = 5'h10;
  assign literal_11599[166] = 5'h10;
  assign literal_11599[167] = 5'h10;
  assign literal_11599[168] = 5'h10;
  assign literal_11599[169] = 5'h10;
  assign literal_11599[170] = 5'h10;
  assign literal_11599[171] = 5'h00;
  assign literal_11599[172] = 5'h00;
  assign literal_11599[173] = 5'h00;
  assign literal_11599[174] = 5'h00;
  assign literal_11599[175] = 5'h00;
  assign literal_11599[176] = 5'h00;
  assign literal_11599[177] = 5'h0a;
  assign literal_11599[178] = 5'h0f;
  assign literal_11599[179] = 5'h10;
  assign literal_11599[180] = 5'h10;
  assign literal_11599[181] = 5'h10;
  assign literal_11599[182] = 5'h10;
  assign literal_11599[183] = 5'h10;
  assign literal_11599[184] = 5'h10;
  assign literal_11599[185] = 5'h10;
  assign literal_11599[186] = 5'h10;
  assign literal_11599[187] = 5'h00;
  assign literal_11599[188] = 5'h00;
  assign literal_11599[189] = 5'h00;
  assign literal_11599[190] = 5'h00;
  assign literal_11599[191] = 5'h00;
  assign literal_11599[192] = 5'h00;
  assign literal_11599[193] = 5'h0a;
  assign literal_11599[194] = 5'h10;
  assign literal_11599[195] = 5'h10;
  assign literal_11599[196] = 5'h10;
  assign literal_11599[197] = 5'h10;
  assign literal_11599[198] = 5'h10;
  assign literal_11599[199] = 5'h10;
  assign literal_11599[200] = 5'h10;
  assign literal_11599[201] = 5'h10;
  assign literal_11599[202] = 5'h10;
  assign literal_11599[203] = 5'h00;
  assign literal_11599[204] = 5'h00;
  assign literal_11599[205] = 5'h00;
  assign literal_11599[206] = 5'h00;
  assign literal_11599[207] = 5'h00;
  assign literal_11599[208] = 5'h00;
  assign literal_11599[209] = 5'h0a;
  assign literal_11599[210] = 5'h10;
  assign literal_11599[211] = 5'h10;
  assign literal_11599[212] = 5'h10;
  assign literal_11599[213] = 5'h10;
  assign literal_11599[214] = 5'h10;
  assign literal_11599[215] = 5'h10;
  assign literal_11599[216] = 5'h10;
  assign literal_11599[217] = 5'h10;
  assign literal_11599[218] = 5'h10;
  assign literal_11599[219] = 5'h00;
  assign literal_11599[220] = 5'h00;
  assign literal_11599[221] = 5'h00;
  assign literal_11599[222] = 5'h00;
  assign literal_11599[223] = 5'h00;
  assign literal_11599[224] = 5'h00;
  assign literal_11599[225] = 5'h0b;
  assign literal_11599[226] = 5'h10;
  assign literal_11599[227] = 5'h10;
  assign literal_11599[228] = 5'h10;
  assign literal_11599[229] = 5'h10;
  assign literal_11599[230] = 5'h10;
  assign literal_11599[231] = 5'h10;
  assign literal_11599[232] = 5'h10;
  assign literal_11599[233] = 5'h10;
  assign literal_11599[234] = 5'h10;
  assign literal_11599[235] = 5'h00;
  assign literal_11599[236] = 5'h00;
  assign literal_11599[237] = 5'h00;
  assign literal_11599[238] = 5'h00;
  assign literal_11599[239] = 5'h00;
  assign literal_11599[240] = 5'h0c;
  assign literal_11599[241] = 5'h0d;
  assign literal_11599[242] = 5'h10;
  assign literal_11599[243] = 5'h10;
  assign literal_11599[244] = 5'h10;
  assign literal_11599[245] = 5'h10;
  assign literal_11599[246] = 5'h10;
  assign literal_11599[247] = 5'h10;
  assign literal_11599[248] = 5'h10;
  assign literal_11599[249] = 5'h10;
  assign literal_11599[250] = 5'h10;
  assign literal_11599[251] = 5'h00;
  wire [15:0] literal_11602[0:251];
  assign literal_11602[0] = 16'h0001;
  assign literal_11602[1] = 16'h0000;
  assign literal_11602[2] = 16'h0004;
  assign literal_11602[3] = 16'h000c;
  assign literal_11602[4] = 16'h001a;
  assign literal_11602[5] = 16'h0076;
  assign literal_11602[6] = 16'h00f6;
  assign literal_11602[7] = 16'h3fe0;
  assign literal_11602[8] = 16'hff96;
  assign literal_11602[9] = 16'hff97;
  assign literal_11602[10] = 16'hff98;
  assign literal_11602[11] = 16'h0000;
  assign literal_11602[12] = 16'h0000;
  assign literal_11602[13] = 16'h0000;
  assign literal_11602[14] = 16'h0000;
  assign literal_11602[15] = 16'h0000;
  assign literal_11602[16] = 16'h0000;
  assign literal_11602[17] = 16'h0005;
  assign literal_11602[18] = 16'h0038;
  assign literal_11602[19] = 16'h0078;
  assign literal_11602[20] = 16'h01f9;
  assign literal_11602[21] = 16'h07f2;
  assign literal_11602[22] = 16'h1fe8;
  assign literal_11602[23] = 16'hff93;
  assign literal_11602[24] = 16'hff99;
  assign literal_11602[25] = 16'hff9a;
  assign literal_11602[26] = 16'hff9e;
  assign literal_11602[27] = 16'h0000;
  assign literal_11602[28] = 16'h0000;
  assign literal_11602[29] = 16'h0000;
  assign literal_11602[30] = 16'h0000;
  assign literal_11602[31] = 16'h0000;
  assign literal_11602[32] = 16'h0000;
  assign literal_11602[33] = 16'h001b;
  assign literal_11602[34] = 16'h007a;
  assign literal_11602[35] = 16'h03f7;
  assign literal_11602[36] = 16'h0ff0;
  assign literal_11602[37] = 16'h1feb;
  assign literal_11602[38] = 16'hff9b;
  assign literal_11602[39] = 16'hff9f;
  assign literal_11602[40] = 16'hffa8;
  assign literal_11602[41] = 16'hffa9;
  assign literal_11602[42] = 16'hfff1;
  assign literal_11602[43] = 16'h0000;
  assign literal_11602[44] = 16'h0000;
  assign literal_11602[45] = 16'h0000;
  assign literal_11602[46] = 16'h0000;
  assign literal_11602[47] = 16'h0000;
  assign literal_11602[48] = 16'h0000;
  assign literal_11602[49] = 16'h0039;
  assign literal_11602[50] = 16'h00fa;
  assign literal_11602[51] = 16'h07f7;
  assign literal_11602[52] = 16'h0ff1;
  assign literal_11602[53] = 16'h7fc6;
  assign literal_11602[54] = 16'hff9c;
  assign literal_11602[55] = 16'hffa3;
  assign literal_11602[56] = 16'hffd7;
  assign literal_11602[57] = 16'hffe4;
  assign literal_11602[58] = 16'hfff2;
  assign literal_11602[59] = 16'h0000;
  assign literal_11602[60] = 16'h0000;
  assign literal_11602[61] = 16'h0000;
  assign literal_11602[62] = 16'h0000;
  assign literal_11602[63] = 16'h0000;
  assign literal_11602[64] = 16'h0000;
  assign literal_11602[65] = 16'h003a;
  assign literal_11602[66] = 16'h03f8;
  assign literal_11602[67] = 16'h0ff2;
  assign literal_11602[68] = 16'h7fc8;
  assign literal_11602[69] = 16'hff9d;
  assign literal_11602[70] = 16'hffbf;
  assign literal_11602[71] = 16'hffcb;
  assign literal_11602[72] = 16'hffd8;
  assign literal_11602[73] = 16'hffe5;
  assign literal_11602[74] = 16'hfff3;
  assign literal_11602[75] = 16'h0000;
  assign literal_11602[76] = 16'h0000;
  assign literal_11602[77] = 16'h0000;
  assign literal_11602[78] = 16'h0000;
  assign literal_11602[79] = 16'h0000;
  assign literal_11602[80] = 16'h0000;
  assign literal_11602[81] = 16'h0077;
  assign literal_11602[82] = 16'h07f3;
  assign literal_11602[83] = 16'h1fea;
  assign literal_11602[84] = 16'hff94;
  assign literal_11602[85] = 16'hffa2;
  assign literal_11602[86] = 16'hffc0;
  assign literal_11602[87] = 16'hffcc;
  assign literal_11602[88] = 16'hffd9;
  assign literal_11602[89] = 16'hffe6;
  assign literal_11602[90] = 16'hfff4;
  assign literal_11602[91] = 16'h0000;
  assign literal_11602[92] = 16'h0000;
  assign literal_11602[93] = 16'h0000;
  assign literal_11602[94] = 16'h0000;
  assign literal_11602[95] = 16'h0000;
  assign literal_11602[96] = 16'h0000;
  assign literal_11602[97] = 16'h0079;
  assign literal_11602[98] = 16'h07f4;
  assign literal_11602[99] = 16'h1fed;
  assign literal_11602[100] = 16'hffa0;
  assign literal_11602[101] = 16'hffb5;
  assign literal_11602[102] = 16'hffc1;
  assign literal_11602[103] = 16'hffcd;
  assign literal_11602[104] = 16'hffda;
  assign literal_11602[105] = 16'hffe7;
  assign literal_11602[106] = 16'hfff5;
  assign literal_11602[107] = 16'h0000;
  assign literal_11602[108] = 16'h0000;
  assign literal_11602[109] = 16'h0000;
  assign literal_11602[110] = 16'h0000;
  assign literal_11602[111] = 16'h0000;
  assign literal_11602[112] = 16'h0000;
  assign literal_11602[113] = 16'h00f7;
  assign literal_11602[114] = 16'h07f5;
  assign literal_11602[115] = 16'h3fe1;
  assign literal_11602[116] = 16'hffa1;
  assign literal_11602[117] = 16'hffb6;
  assign literal_11602[118] = 16'hffc2;
  assign literal_11602[119] = 16'hffce;
  assign literal_11602[120] = 16'hffdb;
  assign literal_11602[121] = 16'hffe8;
  assign literal_11602[122] = 16'hfff6;
  assign literal_11602[123] = 16'h0000;
  assign literal_11602[124] = 16'h0000;
  assign literal_11602[125] = 16'h0000;
  assign literal_11602[126] = 16'h0000;
  assign literal_11602[127] = 16'h0000;
  assign literal_11602[128] = 16'h0000;
  assign literal_11602[129] = 16'h00f8;
  assign literal_11602[130] = 16'h0ff3;
  assign literal_11602[131] = 16'hff92;
  assign literal_11602[132] = 16'hffad;
  assign literal_11602[133] = 16'hffb7;
  assign literal_11602[134] = 16'hffc3;
  assign literal_11602[135] = 16'hffcf;
  assign literal_11602[136] = 16'hffdc;
  assign literal_11602[137] = 16'hffe9;
  assign literal_11602[138] = 16'hfff7;
  assign literal_11602[139] = 16'h0000;
  assign literal_11602[140] = 16'h0000;
  assign literal_11602[141] = 16'h0000;
  assign literal_11602[142] = 16'h0000;
  assign literal_11602[143] = 16'h0000;
  assign literal_11602[144] = 16'h0000;
  assign literal_11602[145] = 16'h00f9;
  assign literal_11602[146] = 16'h1fe9;
  assign literal_11602[147] = 16'hff95;
  assign literal_11602[148] = 16'hffae;
  assign literal_11602[149] = 16'hffb8;
  assign literal_11602[150] = 16'hffc4;
  assign literal_11602[151] = 16'hffd0;
  assign literal_11602[152] = 16'hffdd;
  assign literal_11602[153] = 16'hffea;
  assign literal_11602[154] = 16'hfff8;
  assign literal_11602[155] = 16'h0000;
  assign literal_11602[156] = 16'h0000;
  assign literal_11602[157] = 16'h0000;
  assign literal_11602[158] = 16'h0000;
  assign literal_11602[159] = 16'h0000;
  assign literal_11602[160] = 16'h0000;
  assign literal_11602[161] = 16'h01f6;
  assign literal_11602[162] = 16'h1fec;
  assign literal_11602[163] = 16'hffa5;
  assign literal_11602[164] = 16'hffaf;
  assign literal_11602[165] = 16'hffb9;
  assign literal_11602[166] = 16'hffc5;
  assign literal_11602[167] = 16'hffd1;
  assign literal_11602[168] = 16'hffde;
  assign literal_11602[169] = 16'hffeb;
  assign literal_11602[170] = 16'hfff9;
  assign literal_11602[171] = 16'h0000;
  assign literal_11602[172] = 16'h0000;
  assign literal_11602[173] = 16'h0000;
  assign literal_11602[174] = 16'h0000;
  assign literal_11602[175] = 16'h0000;
  assign literal_11602[176] = 16'h0000;
  assign literal_11602[177] = 16'h01f7;
  assign literal_11602[178] = 16'h1fee;
  assign literal_11602[179] = 16'hffa6;
  assign literal_11602[180] = 16'hffb0;
  assign literal_11602[181] = 16'hffba;
  assign literal_11602[182] = 16'hffc6;
  assign literal_11602[183] = 16'hffd2;
  assign literal_11602[184] = 16'hffdf;
  assign literal_11602[185] = 16'hffec;
  assign literal_11602[186] = 16'hfffa;
  assign literal_11602[187] = 16'h0000;
  assign literal_11602[188] = 16'h0000;
  assign literal_11602[189] = 16'h0000;
  assign literal_11602[190] = 16'h0000;
  assign literal_11602[191] = 16'h0000;
  assign literal_11602[192] = 16'h0000;
  assign literal_11602[193] = 16'h03f4;
  assign literal_11602[194] = 16'h1fef;
  assign literal_11602[195] = 16'hffa7;
  assign literal_11602[196] = 16'hffb1;
  assign literal_11602[197] = 16'hffbb;
  assign literal_11602[198] = 16'hffc7;
  assign literal_11602[199] = 16'hffd3;
  assign literal_11602[200] = 16'hffe0;
  assign literal_11602[201] = 16'hffed;
  assign literal_11602[202] = 16'hfffb;
  assign literal_11602[203] = 16'h0000;
  assign literal_11602[204] = 16'h0000;
  assign literal_11602[205] = 16'h0000;
  assign literal_11602[206] = 16'h0000;
  assign literal_11602[207] = 16'h0000;
  assign literal_11602[208] = 16'h0000;
  assign literal_11602[209] = 16'h03f5;
  assign literal_11602[210] = 16'h3fe2;
  assign literal_11602[211] = 16'hffaa;
  assign literal_11602[212] = 16'hffb2;
  assign literal_11602[213] = 16'hffbc;
  assign literal_11602[214] = 16'hffc8;
  assign literal_11602[215] = 16'hffd4;
  assign literal_11602[216] = 16'hffe1;
  assign literal_11602[217] = 16'hffee;
  assign literal_11602[218] = 16'hfffc;
  assign literal_11602[219] = 16'h0000;
  assign literal_11602[220] = 16'h0000;
  assign literal_11602[221] = 16'h0000;
  assign literal_11602[222] = 16'h0000;
  assign literal_11602[223] = 16'h0000;
  assign literal_11602[224] = 16'h0000;
  assign literal_11602[225] = 16'h03f6;
  assign literal_11602[226] = 16'h7fc7;
  assign literal_11602[227] = 16'hffab;
  assign literal_11602[228] = 16'hffb3;
  assign literal_11602[229] = 16'hffbd;
  assign literal_11602[230] = 16'hffc9;
  assign literal_11602[231] = 16'hffd5;
  assign literal_11602[232] = 16'hffe2;
  assign literal_11602[233] = 16'hffef;
  assign literal_11602[234] = 16'hfffd;
  assign literal_11602[235] = 16'h0000;
  assign literal_11602[236] = 16'h0000;
  assign literal_11602[237] = 16'h0000;
  assign literal_11602[238] = 16'h0000;
  assign literal_11602[239] = 16'h0000;
  assign literal_11602[240] = 16'h01f8;
  assign literal_11602[241] = 16'h07f6;
  assign literal_11602[242] = 16'hffa4;
  assign literal_11602[243] = 16'hffac;
  assign literal_11602[244] = 16'hffb4;
  assign literal_11602[245] = 16'hffbe;
  assign literal_11602[246] = 16'hffca;
  assign literal_11602[247] = 16'hffd6;
  assign literal_11602[248] = 16'hffe3;
  assign literal_11602[249] = 16'hfff0;
  assign literal_11602[250] = 16'hfffe;
  assign literal_11602[251] = 16'h0000;
  wire [15:0] literal_11603[0:251];
  assign literal_11603[0] = 16'h000c;
  assign literal_11603[1] = 16'h0000;
  assign literal_11603[2] = 16'h0001;
  assign literal_11603[3] = 16'h0004;
  assign literal_11603[4] = 16'h000b;
  assign literal_11603[5] = 16'h001a;
  assign literal_11603[6] = 16'h0079;
  assign literal_11603[7] = 16'h01f9;
  assign literal_11603[8] = 16'hff9c;
  assign literal_11603[9] = 16'hff9f;
  assign literal_11603[10] = 16'hffa0;
  assign literal_11603[11] = 16'h0000;
  assign literal_11603[12] = 16'h0000;
  assign literal_11603[13] = 16'h0000;
  assign literal_11603[14] = 16'h0000;
  assign literal_11603[15] = 16'h0000;
  assign literal_11603[16] = 16'h0000;
  assign literal_11603[17] = 16'h000a;
  assign literal_11603[18] = 16'h001c;
  assign literal_11603[19] = 16'h007a;
  assign literal_11603[20] = 16'h01f5;
  assign literal_11603[21] = 16'h03f4;
  assign literal_11603[22] = 16'h07f8;
  assign literal_11603[23] = 16'hff95;
  assign literal_11603[24] = 16'hffa1;
  assign literal_11603[25] = 16'hffa2;
  assign literal_11603[26] = 16'hffad;
  assign literal_11603[27] = 16'h0000;
  assign literal_11603[28] = 16'h0000;
  assign literal_11603[29] = 16'h0000;
  assign literal_11603[30] = 16'h0000;
  assign literal_11603[31] = 16'h0000;
  assign literal_11603[32] = 16'h0000;
  assign literal_11603[33] = 16'h001b;
  assign literal_11603[34] = 16'h00f8;
  assign literal_11603[35] = 16'h03f7;
  assign literal_11603[36] = 16'h0ff4;
  assign literal_11603[37] = 16'h3fdc;
  assign literal_11603[38] = 16'hff9d;
  assign literal_11603[39] = 16'hff90;
  assign literal_11603[40] = 16'hffac;
  assign literal_11603[41] = 16'hffe3;
  assign literal_11603[42] = 16'hfff1;
  assign literal_11603[43] = 16'h0000;
  assign literal_11603[44] = 16'h0000;
  assign literal_11603[45] = 16'h0000;
  assign literal_11603[46] = 16'h0000;
  assign literal_11603[47] = 16'h0000;
  assign literal_11603[48] = 16'h0000;
  assign literal_11603[49] = 16'h003a;
  assign literal_11603[50] = 16'h01f6;
  assign literal_11603[51] = 16'h07f7;
  assign literal_11603[52] = 16'h3fde;
  assign literal_11603[53] = 16'hff8e;
  assign literal_11603[54] = 16'hff94;
  assign literal_11603[55] = 16'hffc9;
  assign literal_11603[56] = 16'hffd6;
  assign literal_11603[57] = 16'hffe4;
  assign literal_11603[58] = 16'hfff2;
  assign literal_11603[59] = 16'h0000;
  assign literal_11603[60] = 16'h0000;
  assign literal_11603[61] = 16'h0000;
  assign literal_11603[62] = 16'h0000;
  assign literal_11603[63] = 16'h0000;
  assign literal_11603[64] = 16'h0000;
  assign literal_11603[65] = 16'h003b;
  assign literal_11603[66] = 16'h03f6;
  assign literal_11603[67] = 16'h3fdd;
  assign literal_11603[68] = 16'hff8f;
  assign literal_11603[69] = 16'hffa5;
  assign literal_11603[70] = 16'hffa6;
  assign literal_11603[71] = 16'hffca;
  assign literal_11603[72] = 16'hffd7;
  assign literal_11603[73] = 16'hffe5;
  assign literal_11603[74] = 16'hfff3;
  assign literal_11603[75] = 16'h0000;
  assign literal_11603[76] = 16'h0000;
  assign literal_11603[77] = 16'h0000;
  assign literal_11603[78] = 16'h0000;
  assign literal_11603[79] = 16'h0000;
  assign literal_11603[80] = 16'h0000;
  assign literal_11603[81] = 16'h0078;
  assign literal_11603[82] = 16'h03f9;
  assign literal_11603[83] = 16'h3fdf;
  assign literal_11603[84] = 16'hff96;
  assign literal_11603[85] = 16'hffab;
  assign literal_11603[86] = 16'hffa9;
  assign literal_11603[87] = 16'hffcb;
  assign literal_11603[88] = 16'hffd8;
  assign literal_11603[89] = 16'hffe6;
  assign literal_11603[90] = 16'hfff4;
  assign literal_11603[91] = 16'h0000;
  assign literal_11603[92] = 16'h0000;
  assign literal_11603[93] = 16'h0000;
  assign literal_11603[94] = 16'h0000;
  assign literal_11603[95] = 16'h0000;
  assign literal_11603[96] = 16'h0000;
  assign literal_11603[97] = 16'h007b;
  assign literal_11603[98] = 16'h0ff2;
  assign literal_11603[99] = 16'h7fc5;
  assign literal_11603[100] = 16'hff97;
  assign literal_11603[101] = 16'hffb5;
  assign literal_11603[102] = 16'hffbf;
  assign literal_11603[103] = 16'hffcc;
  assign literal_11603[104] = 16'hffd9;
  assign literal_11603[105] = 16'hffe7;
  assign literal_11603[106] = 16'hfff5;
  assign literal_11603[107] = 16'h0000;
  assign literal_11603[108] = 16'h0000;
  assign literal_11603[109] = 16'h0000;
  assign literal_11603[110] = 16'h0000;
  assign literal_11603[111] = 16'h0000;
  assign literal_11603[112] = 16'h0000;
  assign literal_11603[113] = 16'h00f9;
  assign literal_11603[114] = 16'h0ff5;
  assign literal_11603[115] = 16'hff8c;
  assign literal_11603[116] = 16'hff98;
  assign literal_11603[117] = 16'hffb6;
  assign literal_11603[118] = 16'hffc0;
  assign literal_11603[119] = 16'hffcd;
  assign literal_11603[120] = 16'hffda;
  assign literal_11603[121] = 16'hffe8;
  assign literal_11603[122] = 16'hfff6;
  assign literal_11603[123] = 16'h0000;
  assign literal_11603[124] = 16'h0000;
  assign literal_11603[125] = 16'h0000;
  assign literal_11603[126] = 16'h0000;
  assign literal_11603[127] = 16'h0000;
  assign literal_11603[128] = 16'h0000;
  assign literal_11603[129] = 16'h01f4;
  assign literal_11603[130] = 16'h1fec;
  assign literal_11603[131] = 16'hff9e;
  assign literal_11603[132] = 16'hffa3;
  assign literal_11603[133] = 16'hffb7;
  assign literal_11603[134] = 16'hffc1;
  assign literal_11603[135] = 16'hffce;
  assign literal_11603[136] = 16'hffdb;
  assign literal_11603[137] = 16'hffe9;
  assign literal_11603[138] = 16'hfff7;
  assign literal_11603[139] = 16'h0000;
  assign literal_11603[140] = 16'h0000;
  assign literal_11603[141] = 16'h0000;
  assign literal_11603[142] = 16'h0000;
  assign literal_11603[143] = 16'h0000;
  assign literal_11603[144] = 16'h0000;
  assign literal_11603[145] = 16'h01f7;
  assign literal_11603[146] = 16'h3fe0;
  assign literal_11603[147] = 16'hff91;
  assign literal_11603[148] = 16'hffa4;
  assign literal_11603[149] = 16'hffb8;
  assign literal_11603[150] = 16'hffc2;
  assign literal_11603[151] = 16'hffcf;
  assign literal_11603[152] = 16'hffdc;
  assign literal_11603[153] = 16'hffea;
  assign literal_11603[154] = 16'hfff8;
  assign literal_11603[155] = 16'h0000;
  assign literal_11603[156] = 16'h0000;
  assign literal_11603[157] = 16'h0000;
  assign literal_11603[158] = 16'h0000;
  assign literal_11603[159] = 16'h0000;
  assign literal_11603[160] = 16'h0000;
  assign literal_11603[161] = 16'h01f8;
  assign literal_11603[162] = 16'h3fe1;
  assign literal_11603[163] = 16'hff92;
  assign literal_11603[164] = 16'hffa7;
  assign literal_11603[165] = 16'hffb9;
  assign literal_11603[166] = 16'hffc3;
  assign literal_11603[167] = 16'hffd0;
  assign literal_11603[168] = 16'hffdd;
  assign literal_11603[169] = 16'hffeb;
  assign literal_11603[170] = 16'hfff9;
  assign literal_11603[171] = 16'h0000;
  assign literal_11603[172] = 16'h0000;
  assign literal_11603[173] = 16'h0000;
  assign literal_11603[174] = 16'h0000;
  assign literal_11603[175] = 16'h0000;
  assign literal_11603[176] = 16'h0000;
  assign literal_11603[177] = 16'h03f5;
  assign literal_11603[178] = 16'h7fc4;
  assign literal_11603[179] = 16'hff93;
  assign literal_11603[180] = 16'hffa8;
  assign literal_11603[181] = 16'hffba;
  assign literal_11603[182] = 16'hffc4;
  assign literal_11603[183] = 16'hffd1;
  assign literal_11603[184] = 16'hffde;
  assign literal_11603[185] = 16'hffec;
  assign literal_11603[186] = 16'hfffa;
  assign literal_11603[187] = 16'h0000;
  assign literal_11603[188] = 16'h0000;
  assign literal_11603[189] = 16'h0000;
  assign literal_11603[190] = 16'h0000;
  assign literal_11603[191] = 16'h0000;
  assign literal_11603[192] = 16'h0000;
  assign literal_11603[193] = 16'h03f8;
  assign literal_11603[194] = 16'hff8d;
  assign literal_11603[195] = 16'hff99;
  assign literal_11603[196] = 16'hffb1;
  assign literal_11603[197] = 16'hffbb;
  assign literal_11603[198] = 16'hffc5;
  assign literal_11603[199] = 16'hffd2;
  assign literal_11603[200] = 16'hffdf;
  assign literal_11603[201] = 16'hffed;
  assign literal_11603[202] = 16'hfffb;
  assign literal_11603[203] = 16'h0000;
  assign literal_11603[204] = 16'h0000;
  assign literal_11603[205] = 16'h0000;
  assign literal_11603[206] = 16'h0000;
  assign literal_11603[207] = 16'h0000;
  assign literal_11603[208] = 16'h0000;
  assign literal_11603[209] = 16'h03fa;
  assign literal_11603[210] = 16'hff9a;
  assign literal_11603[211] = 16'hffaa;
  assign literal_11603[212] = 16'hffb2;
  assign literal_11603[213] = 16'hffbc;
  assign literal_11603[214] = 16'hffc6;
  assign literal_11603[215] = 16'hffd3;
  assign literal_11603[216] = 16'hffe0;
  assign literal_11603[217] = 16'hffee;
  assign literal_11603[218] = 16'hfffc;
  assign literal_11603[219] = 16'h0000;
  assign literal_11603[220] = 16'h0000;
  assign literal_11603[221] = 16'h0000;
  assign literal_11603[222] = 16'h0000;
  assign literal_11603[223] = 16'h0000;
  assign literal_11603[224] = 16'h0000;
  assign literal_11603[225] = 16'h07f6;
  assign literal_11603[226] = 16'hff9b;
  assign literal_11603[227] = 16'hffaf;
  assign literal_11603[228] = 16'hffb3;
  assign literal_11603[229] = 16'hffbd;
  assign literal_11603[230] = 16'hffc7;
  assign literal_11603[231] = 16'hffd4;
  assign literal_11603[232] = 16'hffe1;
  assign literal_11603[233] = 16'hffef;
  assign literal_11603[234] = 16'hfffd;
  assign literal_11603[235] = 16'h0000;
  assign literal_11603[236] = 16'h0000;
  assign literal_11603[237] = 16'h0000;
  assign literal_11603[238] = 16'h0000;
  assign literal_11603[239] = 16'h0000;
  assign literal_11603[240] = 16'h0ff3;
  assign literal_11603[241] = 16'h1fed;
  assign literal_11603[242] = 16'hffae;
  assign literal_11603[243] = 16'hffb0;
  assign literal_11603[244] = 16'hffb4;
  assign literal_11603[245] = 16'hffbe;
  assign literal_11603[246] = 16'hffc8;
  assign literal_11603[247] = 16'hffd5;
  assign literal_11603[248] = 16'hffe2;
  assign literal_11603[249] = 16'hfff0;
  assign literal_11603[250] = 16'hfffe;
  assign literal_11603[251] = 16'h0000;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [2:0] p1_run_0_squeezed_const_msb_bits_comb;
  wire [9:0] p1_row0_comb[0:7];
  wire [9:0] p1_row1_comb[0:7];
  wire [9:0] p1_array_concat_10569_comb[0:15];
  wire [9:0] p1_row2_comb[0:7];
  wire [9:0] p1_array_concat_10572_comb[0:23];
  wire [9:0] p1_row3_comb[0:7];
  wire [9:0] p1_array_concat_10575_comb[0:31];
  wire [9:0] p1_row4_comb[0:7];
  wire [9:0] p1_array_concat_10578_comb[0:39];
  wire [9:0] p1_row5_comb[0:7];
  wire p1_next_pix__1_squeezed_squeezed_const_msb_bits__5_comb;
  wire p1_next_pix__1_squeezed_squeezed_const_msb_bits_comb;
  wire [9:0] p1_array_concat_10584_comb[0:47];
  wire [9:0] p1_row6_comb[0:7];
  wire [7:0] p1_concat_10587_comb;
  wire [8:0] p1_concat_10589_comb;
  wire [9:0] p1_array_concat_10591_comb[0:55];
  wire [9:0] p1_row7_comb[0:7];
  wire [7:0] p1_add_10593_comb;
  wire [8:0] p1_add_10595_comb;
  wire [9:0] p1_flat_ac_comb[0:63];
  wire p1_next_pix__1_squeezed_squeezed_const_msb_bits__6_comb;
  wire p1_next_pix__1_squeezed_squeezed_const_msb_bits__7_comb;
  wire [8:0] p1_concat_10600_comb;
  wire [8:0] p1_add_10604_comb;
  wire [6:0] p1_concat_10605_comb;
  wire [6:0] p1_add_10615_comb;
  wire [7:0] p1_add_10630_comb;
  wire [5:0] p1_add_10659_comb;
  wire [7:0] p1_add_10671_comb;
  wire [6:0] p1_add_10684_comb;
  wire [7:0] p1_add_10701_comb;
  wire [8:0] p1_concat_10625_comb;
  wire [8:0] p1_add_10631_comb;
  wire [8:0] p1_concat_10640_comb;
  wire [8:0] p1_add_10647_comb;
  wire [8:0] p1_concat_10668_comb;
  wire [8:0] p1_add_10672_comb;
  wire [8:0] p1_concat_10678_comb;
  wire [8:0] p1_add_10685_comb;
  wire [8:0] p1_concat_10694_comb;
  wire [8:0] p1_add_10702_comb;
  wire [8:0] p1_concat_10709_comb;
  wire [8:0] p1_add_10723_comb;
  wire [1:0] p1_and_10646_comb;
  wire p1_or_10655_comb;
  wire p1_or_10663_comb;
  wire p1_or_10669_comb;
  wire p1_nor_10670_comb;
  wire p1_or_10691_comb;
  wire p1_or_10700_comb;
  wire p1_or_10708_comb;
  wire p1_or_10715_comb;
  wire p1_or_10722_comb;
  wire p1_or_10726_comb;
  wire p1_or_10730_comb;
  wire p1_nor_10733_comb;
  assign p1_run_0_squeezed_const_msb_bits_comb = 3'h0;
  assign p1_row0_comb[0] = p0_matrix[p1_run_0_squeezed_const_msb_bits_comb][0];
  assign p1_row0_comb[1] = p0_matrix[p1_run_0_squeezed_const_msb_bits_comb][1];
  assign p1_row0_comb[2] = p0_matrix[p1_run_0_squeezed_const_msb_bits_comb][2];
  assign p1_row0_comb[3] = p0_matrix[p1_run_0_squeezed_const_msb_bits_comb][3];
  assign p1_row0_comb[4] = p0_matrix[p1_run_0_squeezed_const_msb_bits_comb][4];
  assign p1_row0_comb[5] = p0_matrix[p1_run_0_squeezed_const_msb_bits_comb][5];
  assign p1_row0_comb[6] = p0_matrix[p1_run_0_squeezed_const_msb_bits_comb][6];
  assign p1_row0_comb[7] = p0_matrix[p1_run_0_squeezed_const_msb_bits_comb][7];
  assign p1_row1_comb[0] = p0_matrix[3'h1][0];
  assign p1_row1_comb[1] = p0_matrix[3'h1][1];
  assign p1_row1_comb[2] = p0_matrix[3'h1][2];
  assign p1_row1_comb[3] = p0_matrix[3'h1][3];
  assign p1_row1_comb[4] = p0_matrix[3'h1][4];
  assign p1_row1_comb[5] = p0_matrix[3'h1][5];
  assign p1_row1_comb[6] = p0_matrix[3'h1][6];
  assign p1_row1_comb[7] = p0_matrix[3'h1][7];
  assign p1_array_concat_10569_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_10569_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_10569_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_10569_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_10569_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_10569_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_10569_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_10569_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_10569_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_10569_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_10569_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_10569_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_10569_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_10569_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_10569_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_10569_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_10572_comb[0] = p1_array_concat_10569_comb[0];
  assign p1_array_concat_10572_comb[1] = p1_array_concat_10569_comb[1];
  assign p1_array_concat_10572_comb[2] = p1_array_concat_10569_comb[2];
  assign p1_array_concat_10572_comb[3] = p1_array_concat_10569_comb[3];
  assign p1_array_concat_10572_comb[4] = p1_array_concat_10569_comb[4];
  assign p1_array_concat_10572_comb[5] = p1_array_concat_10569_comb[5];
  assign p1_array_concat_10572_comb[6] = p1_array_concat_10569_comb[6];
  assign p1_array_concat_10572_comb[7] = p1_array_concat_10569_comb[7];
  assign p1_array_concat_10572_comb[8] = p1_array_concat_10569_comb[8];
  assign p1_array_concat_10572_comb[9] = p1_array_concat_10569_comb[9];
  assign p1_array_concat_10572_comb[10] = p1_array_concat_10569_comb[10];
  assign p1_array_concat_10572_comb[11] = p1_array_concat_10569_comb[11];
  assign p1_array_concat_10572_comb[12] = p1_array_concat_10569_comb[12];
  assign p1_array_concat_10572_comb[13] = p1_array_concat_10569_comb[13];
  assign p1_array_concat_10572_comb[14] = p1_array_concat_10569_comb[14];
  assign p1_array_concat_10572_comb[15] = p1_array_concat_10569_comb[15];
  assign p1_array_concat_10572_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_10572_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_10572_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_10572_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_10572_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_10572_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_10572_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_10572_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_array_concat_10575_comb[0] = p1_array_concat_10572_comb[0];
  assign p1_array_concat_10575_comb[1] = p1_array_concat_10572_comb[1];
  assign p1_array_concat_10575_comb[2] = p1_array_concat_10572_comb[2];
  assign p1_array_concat_10575_comb[3] = p1_array_concat_10572_comb[3];
  assign p1_array_concat_10575_comb[4] = p1_array_concat_10572_comb[4];
  assign p1_array_concat_10575_comb[5] = p1_array_concat_10572_comb[5];
  assign p1_array_concat_10575_comb[6] = p1_array_concat_10572_comb[6];
  assign p1_array_concat_10575_comb[7] = p1_array_concat_10572_comb[7];
  assign p1_array_concat_10575_comb[8] = p1_array_concat_10572_comb[8];
  assign p1_array_concat_10575_comb[9] = p1_array_concat_10572_comb[9];
  assign p1_array_concat_10575_comb[10] = p1_array_concat_10572_comb[10];
  assign p1_array_concat_10575_comb[11] = p1_array_concat_10572_comb[11];
  assign p1_array_concat_10575_comb[12] = p1_array_concat_10572_comb[12];
  assign p1_array_concat_10575_comb[13] = p1_array_concat_10572_comb[13];
  assign p1_array_concat_10575_comb[14] = p1_array_concat_10572_comb[14];
  assign p1_array_concat_10575_comb[15] = p1_array_concat_10572_comb[15];
  assign p1_array_concat_10575_comb[16] = p1_array_concat_10572_comb[16];
  assign p1_array_concat_10575_comb[17] = p1_array_concat_10572_comb[17];
  assign p1_array_concat_10575_comb[18] = p1_array_concat_10572_comb[18];
  assign p1_array_concat_10575_comb[19] = p1_array_concat_10572_comb[19];
  assign p1_array_concat_10575_comb[20] = p1_array_concat_10572_comb[20];
  assign p1_array_concat_10575_comb[21] = p1_array_concat_10572_comb[21];
  assign p1_array_concat_10575_comb[22] = p1_array_concat_10572_comb[22];
  assign p1_array_concat_10575_comb[23] = p1_array_concat_10572_comb[23];
  assign p1_array_concat_10575_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_10575_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_10575_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_10575_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_10575_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_10575_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_10575_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_10575_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[3'h4][0];
  assign p1_row4_comb[1] = p0_matrix[3'h4][1];
  assign p1_row4_comb[2] = p0_matrix[3'h4][2];
  assign p1_row4_comb[3] = p0_matrix[3'h4][3];
  assign p1_row4_comb[4] = p0_matrix[3'h4][4];
  assign p1_row4_comb[5] = p0_matrix[3'h4][5];
  assign p1_row4_comb[6] = p0_matrix[3'h4][6];
  assign p1_row4_comb[7] = p0_matrix[3'h4][7];
  assign p1_array_concat_10578_comb[0] = p1_array_concat_10575_comb[0];
  assign p1_array_concat_10578_comb[1] = p1_array_concat_10575_comb[1];
  assign p1_array_concat_10578_comb[2] = p1_array_concat_10575_comb[2];
  assign p1_array_concat_10578_comb[3] = p1_array_concat_10575_comb[3];
  assign p1_array_concat_10578_comb[4] = p1_array_concat_10575_comb[4];
  assign p1_array_concat_10578_comb[5] = p1_array_concat_10575_comb[5];
  assign p1_array_concat_10578_comb[6] = p1_array_concat_10575_comb[6];
  assign p1_array_concat_10578_comb[7] = p1_array_concat_10575_comb[7];
  assign p1_array_concat_10578_comb[8] = p1_array_concat_10575_comb[8];
  assign p1_array_concat_10578_comb[9] = p1_array_concat_10575_comb[9];
  assign p1_array_concat_10578_comb[10] = p1_array_concat_10575_comb[10];
  assign p1_array_concat_10578_comb[11] = p1_array_concat_10575_comb[11];
  assign p1_array_concat_10578_comb[12] = p1_array_concat_10575_comb[12];
  assign p1_array_concat_10578_comb[13] = p1_array_concat_10575_comb[13];
  assign p1_array_concat_10578_comb[14] = p1_array_concat_10575_comb[14];
  assign p1_array_concat_10578_comb[15] = p1_array_concat_10575_comb[15];
  assign p1_array_concat_10578_comb[16] = p1_array_concat_10575_comb[16];
  assign p1_array_concat_10578_comb[17] = p1_array_concat_10575_comb[17];
  assign p1_array_concat_10578_comb[18] = p1_array_concat_10575_comb[18];
  assign p1_array_concat_10578_comb[19] = p1_array_concat_10575_comb[19];
  assign p1_array_concat_10578_comb[20] = p1_array_concat_10575_comb[20];
  assign p1_array_concat_10578_comb[21] = p1_array_concat_10575_comb[21];
  assign p1_array_concat_10578_comb[22] = p1_array_concat_10575_comb[22];
  assign p1_array_concat_10578_comb[23] = p1_array_concat_10575_comb[23];
  assign p1_array_concat_10578_comb[24] = p1_array_concat_10575_comb[24];
  assign p1_array_concat_10578_comb[25] = p1_array_concat_10575_comb[25];
  assign p1_array_concat_10578_comb[26] = p1_array_concat_10575_comb[26];
  assign p1_array_concat_10578_comb[27] = p1_array_concat_10575_comb[27];
  assign p1_array_concat_10578_comb[28] = p1_array_concat_10575_comb[28];
  assign p1_array_concat_10578_comb[29] = p1_array_concat_10575_comb[29];
  assign p1_array_concat_10578_comb[30] = p1_array_concat_10575_comb[30];
  assign p1_array_concat_10578_comb[31] = p1_array_concat_10575_comb[31];
  assign p1_array_concat_10578_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_10578_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_10578_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_10578_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_10578_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_10578_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_10578_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_10578_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[3'h5][0];
  assign p1_row5_comb[1] = p0_matrix[3'h5][1];
  assign p1_row5_comb[2] = p0_matrix[3'h5][2];
  assign p1_row5_comb[3] = p0_matrix[3'h5][3];
  assign p1_row5_comb[4] = p0_matrix[3'h5][4];
  assign p1_row5_comb[5] = p0_matrix[3'h5][5];
  assign p1_row5_comb[6] = p0_matrix[3'h5][6];
  assign p1_row5_comb[7] = p0_matrix[3'h5][7];
  assign p1_next_pix__1_squeezed_squeezed_const_msb_bits__5_comb = 1'h0;
  assign p1_next_pix__1_squeezed_squeezed_const_msb_bits_comb = 1'h0;
  assign p1_array_concat_10584_comb[0] = p1_array_concat_10578_comb[0];
  assign p1_array_concat_10584_comb[1] = p1_array_concat_10578_comb[1];
  assign p1_array_concat_10584_comb[2] = p1_array_concat_10578_comb[2];
  assign p1_array_concat_10584_comb[3] = p1_array_concat_10578_comb[3];
  assign p1_array_concat_10584_comb[4] = p1_array_concat_10578_comb[4];
  assign p1_array_concat_10584_comb[5] = p1_array_concat_10578_comb[5];
  assign p1_array_concat_10584_comb[6] = p1_array_concat_10578_comb[6];
  assign p1_array_concat_10584_comb[7] = p1_array_concat_10578_comb[7];
  assign p1_array_concat_10584_comb[8] = p1_array_concat_10578_comb[8];
  assign p1_array_concat_10584_comb[9] = p1_array_concat_10578_comb[9];
  assign p1_array_concat_10584_comb[10] = p1_array_concat_10578_comb[10];
  assign p1_array_concat_10584_comb[11] = p1_array_concat_10578_comb[11];
  assign p1_array_concat_10584_comb[12] = p1_array_concat_10578_comb[12];
  assign p1_array_concat_10584_comb[13] = p1_array_concat_10578_comb[13];
  assign p1_array_concat_10584_comb[14] = p1_array_concat_10578_comb[14];
  assign p1_array_concat_10584_comb[15] = p1_array_concat_10578_comb[15];
  assign p1_array_concat_10584_comb[16] = p1_array_concat_10578_comb[16];
  assign p1_array_concat_10584_comb[17] = p1_array_concat_10578_comb[17];
  assign p1_array_concat_10584_comb[18] = p1_array_concat_10578_comb[18];
  assign p1_array_concat_10584_comb[19] = p1_array_concat_10578_comb[19];
  assign p1_array_concat_10584_comb[20] = p1_array_concat_10578_comb[20];
  assign p1_array_concat_10584_comb[21] = p1_array_concat_10578_comb[21];
  assign p1_array_concat_10584_comb[22] = p1_array_concat_10578_comb[22];
  assign p1_array_concat_10584_comb[23] = p1_array_concat_10578_comb[23];
  assign p1_array_concat_10584_comb[24] = p1_array_concat_10578_comb[24];
  assign p1_array_concat_10584_comb[25] = p1_array_concat_10578_comb[25];
  assign p1_array_concat_10584_comb[26] = p1_array_concat_10578_comb[26];
  assign p1_array_concat_10584_comb[27] = p1_array_concat_10578_comb[27];
  assign p1_array_concat_10584_comb[28] = p1_array_concat_10578_comb[28];
  assign p1_array_concat_10584_comb[29] = p1_array_concat_10578_comb[29];
  assign p1_array_concat_10584_comb[30] = p1_array_concat_10578_comb[30];
  assign p1_array_concat_10584_comb[31] = p1_array_concat_10578_comb[31];
  assign p1_array_concat_10584_comb[32] = p1_array_concat_10578_comb[32];
  assign p1_array_concat_10584_comb[33] = p1_array_concat_10578_comb[33];
  assign p1_array_concat_10584_comb[34] = p1_array_concat_10578_comb[34];
  assign p1_array_concat_10584_comb[35] = p1_array_concat_10578_comb[35];
  assign p1_array_concat_10584_comb[36] = p1_array_concat_10578_comb[36];
  assign p1_array_concat_10584_comb[37] = p1_array_concat_10578_comb[37];
  assign p1_array_concat_10584_comb[38] = p1_array_concat_10578_comb[38];
  assign p1_array_concat_10584_comb[39] = p1_array_concat_10578_comb[39];
  assign p1_array_concat_10584_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_10584_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_10584_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_10584_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_10584_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_10584_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_10584_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_10584_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[3'h6][0];
  assign p1_row6_comb[1] = p0_matrix[3'h6][1];
  assign p1_row6_comb[2] = p0_matrix[3'h6][2];
  assign p1_row6_comb[3] = p0_matrix[3'h6][3];
  assign p1_row6_comb[4] = p0_matrix[3'h6][4];
  assign p1_row6_comb[5] = p0_matrix[3'h6][5];
  assign p1_row6_comb[6] = p0_matrix[3'h6][6];
  assign p1_row6_comb[7] = p0_matrix[3'h6][7];
  assign p1_concat_10587_comb = {p1_next_pix__1_squeezed_squeezed_const_msb_bits__5_comb, p0_start_pix[7:1]};
  assign p1_concat_10589_comb = {p1_next_pix__1_squeezed_squeezed_const_msb_bits_comb, p0_start_pix};
  assign p1_array_concat_10591_comb[0] = p1_array_concat_10584_comb[0];
  assign p1_array_concat_10591_comb[1] = p1_array_concat_10584_comb[1];
  assign p1_array_concat_10591_comb[2] = p1_array_concat_10584_comb[2];
  assign p1_array_concat_10591_comb[3] = p1_array_concat_10584_comb[3];
  assign p1_array_concat_10591_comb[4] = p1_array_concat_10584_comb[4];
  assign p1_array_concat_10591_comb[5] = p1_array_concat_10584_comb[5];
  assign p1_array_concat_10591_comb[6] = p1_array_concat_10584_comb[6];
  assign p1_array_concat_10591_comb[7] = p1_array_concat_10584_comb[7];
  assign p1_array_concat_10591_comb[8] = p1_array_concat_10584_comb[8];
  assign p1_array_concat_10591_comb[9] = p1_array_concat_10584_comb[9];
  assign p1_array_concat_10591_comb[10] = p1_array_concat_10584_comb[10];
  assign p1_array_concat_10591_comb[11] = p1_array_concat_10584_comb[11];
  assign p1_array_concat_10591_comb[12] = p1_array_concat_10584_comb[12];
  assign p1_array_concat_10591_comb[13] = p1_array_concat_10584_comb[13];
  assign p1_array_concat_10591_comb[14] = p1_array_concat_10584_comb[14];
  assign p1_array_concat_10591_comb[15] = p1_array_concat_10584_comb[15];
  assign p1_array_concat_10591_comb[16] = p1_array_concat_10584_comb[16];
  assign p1_array_concat_10591_comb[17] = p1_array_concat_10584_comb[17];
  assign p1_array_concat_10591_comb[18] = p1_array_concat_10584_comb[18];
  assign p1_array_concat_10591_comb[19] = p1_array_concat_10584_comb[19];
  assign p1_array_concat_10591_comb[20] = p1_array_concat_10584_comb[20];
  assign p1_array_concat_10591_comb[21] = p1_array_concat_10584_comb[21];
  assign p1_array_concat_10591_comb[22] = p1_array_concat_10584_comb[22];
  assign p1_array_concat_10591_comb[23] = p1_array_concat_10584_comb[23];
  assign p1_array_concat_10591_comb[24] = p1_array_concat_10584_comb[24];
  assign p1_array_concat_10591_comb[25] = p1_array_concat_10584_comb[25];
  assign p1_array_concat_10591_comb[26] = p1_array_concat_10584_comb[26];
  assign p1_array_concat_10591_comb[27] = p1_array_concat_10584_comb[27];
  assign p1_array_concat_10591_comb[28] = p1_array_concat_10584_comb[28];
  assign p1_array_concat_10591_comb[29] = p1_array_concat_10584_comb[29];
  assign p1_array_concat_10591_comb[30] = p1_array_concat_10584_comb[30];
  assign p1_array_concat_10591_comb[31] = p1_array_concat_10584_comb[31];
  assign p1_array_concat_10591_comb[32] = p1_array_concat_10584_comb[32];
  assign p1_array_concat_10591_comb[33] = p1_array_concat_10584_comb[33];
  assign p1_array_concat_10591_comb[34] = p1_array_concat_10584_comb[34];
  assign p1_array_concat_10591_comb[35] = p1_array_concat_10584_comb[35];
  assign p1_array_concat_10591_comb[36] = p1_array_concat_10584_comb[36];
  assign p1_array_concat_10591_comb[37] = p1_array_concat_10584_comb[37];
  assign p1_array_concat_10591_comb[38] = p1_array_concat_10584_comb[38];
  assign p1_array_concat_10591_comb[39] = p1_array_concat_10584_comb[39];
  assign p1_array_concat_10591_comb[40] = p1_array_concat_10584_comb[40];
  assign p1_array_concat_10591_comb[41] = p1_array_concat_10584_comb[41];
  assign p1_array_concat_10591_comb[42] = p1_array_concat_10584_comb[42];
  assign p1_array_concat_10591_comb[43] = p1_array_concat_10584_comb[43];
  assign p1_array_concat_10591_comb[44] = p1_array_concat_10584_comb[44];
  assign p1_array_concat_10591_comb[45] = p1_array_concat_10584_comb[45];
  assign p1_array_concat_10591_comb[46] = p1_array_concat_10584_comb[46];
  assign p1_array_concat_10591_comb[47] = p1_array_concat_10584_comb[47];
  assign p1_array_concat_10591_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_10591_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_10591_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_10591_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_10591_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_10591_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_10591_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_10591_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[3'h7][0];
  assign p1_row7_comb[1] = p0_matrix[3'h7][1];
  assign p1_row7_comb[2] = p0_matrix[3'h7][2];
  assign p1_row7_comb[3] = p0_matrix[3'h7][3];
  assign p1_row7_comb[4] = p0_matrix[3'h7][4];
  assign p1_row7_comb[5] = p0_matrix[3'h7][5];
  assign p1_row7_comb[6] = p0_matrix[3'h7][6];
  assign p1_row7_comb[7] = p0_matrix[3'h7][7];
  assign p1_add_10593_comb = p1_concat_10587_comb + 8'h07;
  assign p1_add_10595_comb = p1_concat_10589_comb + 9'h00f;
  assign p1_flat_ac_comb[0] = p1_array_concat_10591_comb[0];
  assign p1_flat_ac_comb[1] = p1_array_concat_10591_comb[1];
  assign p1_flat_ac_comb[2] = p1_array_concat_10591_comb[2];
  assign p1_flat_ac_comb[3] = p1_array_concat_10591_comb[3];
  assign p1_flat_ac_comb[4] = p1_array_concat_10591_comb[4];
  assign p1_flat_ac_comb[5] = p1_array_concat_10591_comb[5];
  assign p1_flat_ac_comb[6] = p1_array_concat_10591_comb[6];
  assign p1_flat_ac_comb[7] = p1_array_concat_10591_comb[7];
  assign p1_flat_ac_comb[8] = p1_array_concat_10591_comb[8];
  assign p1_flat_ac_comb[9] = p1_array_concat_10591_comb[9];
  assign p1_flat_ac_comb[10] = p1_array_concat_10591_comb[10];
  assign p1_flat_ac_comb[11] = p1_array_concat_10591_comb[11];
  assign p1_flat_ac_comb[12] = p1_array_concat_10591_comb[12];
  assign p1_flat_ac_comb[13] = p1_array_concat_10591_comb[13];
  assign p1_flat_ac_comb[14] = p1_array_concat_10591_comb[14];
  assign p1_flat_ac_comb[15] = p1_array_concat_10591_comb[15];
  assign p1_flat_ac_comb[16] = p1_array_concat_10591_comb[16];
  assign p1_flat_ac_comb[17] = p1_array_concat_10591_comb[17];
  assign p1_flat_ac_comb[18] = p1_array_concat_10591_comb[18];
  assign p1_flat_ac_comb[19] = p1_array_concat_10591_comb[19];
  assign p1_flat_ac_comb[20] = p1_array_concat_10591_comb[20];
  assign p1_flat_ac_comb[21] = p1_array_concat_10591_comb[21];
  assign p1_flat_ac_comb[22] = p1_array_concat_10591_comb[22];
  assign p1_flat_ac_comb[23] = p1_array_concat_10591_comb[23];
  assign p1_flat_ac_comb[24] = p1_array_concat_10591_comb[24];
  assign p1_flat_ac_comb[25] = p1_array_concat_10591_comb[25];
  assign p1_flat_ac_comb[26] = p1_array_concat_10591_comb[26];
  assign p1_flat_ac_comb[27] = p1_array_concat_10591_comb[27];
  assign p1_flat_ac_comb[28] = p1_array_concat_10591_comb[28];
  assign p1_flat_ac_comb[29] = p1_array_concat_10591_comb[29];
  assign p1_flat_ac_comb[30] = p1_array_concat_10591_comb[30];
  assign p1_flat_ac_comb[31] = p1_array_concat_10591_comb[31];
  assign p1_flat_ac_comb[32] = p1_array_concat_10591_comb[32];
  assign p1_flat_ac_comb[33] = p1_array_concat_10591_comb[33];
  assign p1_flat_ac_comb[34] = p1_array_concat_10591_comb[34];
  assign p1_flat_ac_comb[35] = p1_array_concat_10591_comb[35];
  assign p1_flat_ac_comb[36] = p1_array_concat_10591_comb[36];
  assign p1_flat_ac_comb[37] = p1_array_concat_10591_comb[37];
  assign p1_flat_ac_comb[38] = p1_array_concat_10591_comb[38];
  assign p1_flat_ac_comb[39] = p1_array_concat_10591_comb[39];
  assign p1_flat_ac_comb[40] = p1_array_concat_10591_comb[40];
  assign p1_flat_ac_comb[41] = p1_array_concat_10591_comb[41];
  assign p1_flat_ac_comb[42] = p1_array_concat_10591_comb[42];
  assign p1_flat_ac_comb[43] = p1_array_concat_10591_comb[43];
  assign p1_flat_ac_comb[44] = p1_array_concat_10591_comb[44];
  assign p1_flat_ac_comb[45] = p1_array_concat_10591_comb[45];
  assign p1_flat_ac_comb[46] = p1_array_concat_10591_comb[46];
  assign p1_flat_ac_comb[47] = p1_array_concat_10591_comb[47];
  assign p1_flat_ac_comb[48] = p1_array_concat_10591_comb[48];
  assign p1_flat_ac_comb[49] = p1_array_concat_10591_comb[49];
  assign p1_flat_ac_comb[50] = p1_array_concat_10591_comb[50];
  assign p1_flat_ac_comb[51] = p1_array_concat_10591_comb[51];
  assign p1_flat_ac_comb[52] = p1_array_concat_10591_comb[52];
  assign p1_flat_ac_comb[53] = p1_array_concat_10591_comb[53];
  assign p1_flat_ac_comb[54] = p1_array_concat_10591_comb[54];
  assign p1_flat_ac_comb[55] = p1_array_concat_10591_comb[55];
  assign p1_flat_ac_comb[56] = p1_row7_comb[0];
  assign p1_flat_ac_comb[57] = p1_row7_comb[1];
  assign p1_flat_ac_comb[58] = p1_row7_comb[2];
  assign p1_flat_ac_comb[59] = p1_row7_comb[3];
  assign p1_flat_ac_comb[60] = p1_row7_comb[4];
  assign p1_flat_ac_comb[61] = p1_row7_comb[5];
  assign p1_flat_ac_comb[62] = p1_row7_comb[6];
  assign p1_flat_ac_comb[63] = p1_row7_comb[7];
  assign p1_next_pix__1_squeezed_squeezed_const_msb_bits__6_comb = 1'h0;
  assign p1_next_pix__1_squeezed_squeezed_const_msb_bits__7_comb = 1'h0;
  assign p1_concat_10600_comb = {p1_add_10593_comb, p0_start_pix[0]};
  assign p1_add_10604_comb = p1_concat_10589_comb + 9'h00d;
  assign p1_concat_10605_comb = {p1_next_pix__1_squeezed_squeezed_const_msb_bits__6_comb, p0_start_pix[7:2]};
  assign p1_add_10615_comb = p1_concat_10605_comb + 7'h03;
  assign p1_add_10630_comb = p1_concat_10587_comb + 8'h05;
  assign p1_add_10659_comb = {p1_next_pix__1_squeezed_squeezed_const_msb_bits__7_comb, p0_start_pix[7:3]} + 6'h01;
  assign p1_add_10671_comb = p1_concat_10587_comb + 8'h03;
  assign p1_add_10684_comb = p1_concat_10605_comb + 7'h01;
  assign p1_add_10701_comb = p1_concat_10587_comb + 8'h01;
  assign p1_concat_10625_comb = {p1_add_10615_comb, p0_start_pix[1:0]};
  assign p1_add_10631_comb = p1_concat_10589_comb + 9'h00b;
  assign p1_concat_10640_comb = {p1_add_10630_comb, p0_start_pix[0]};
  assign p1_add_10647_comb = p1_concat_10589_comb + 9'h009;
  assign p1_concat_10668_comb = {p1_add_10659_comb, p0_start_pix[2:0]};
  assign p1_add_10672_comb = p1_concat_10589_comb + 9'h007;
  assign p1_concat_10678_comb = {p1_add_10671_comb, p0_start_pix[0]};
  assign p1_add_10685_comb = p1_concat_10589_comb + 9'h005;
  assign p1_concat_10694_comb = {p1_add_10684_comb, p0_start_pix[1:0]};
  assign p1_add_10702_comb = p1_concat_10589_comb + 9'h003;
  assign p1_concat_10709_comb = {p1_add_10701_comb, p0_start_pix[0]};
  assign p1_add_10723_comb = p1_concat_10589_comb + 9'h001;
  assign p1_and_10646_comb = ((|p1_add_10593_comb[7:5]) | p1_flat_ac_comb[p1_concat_10600_comb > 9'h03f ? 6'h3f : p1_concat_10600_comb[5:0]] != 10'h000 ? 2'h1 : {1'h1, ~((|p1_add_10595_comb[8:6]) | p1_flat_ac_comb[p1_add_10595_comb > 9'h03f ? 6'h3f : p1_add_10595_comb[5:0]] != 10'h000)}) & {2{~((|p1_add_10604_comb[8:6]) | p1_flat_ac_comb[p1_add_10604_comb > 9'h03f ? 6'h3f : p1_add_10604_comb[5:0]] != 10'h000)}};
  assign p1_or_10655_comb = (|p1_add_10615_comb[6:4]) | p1_flat_ac_comb[p1_concat_10625_comb > 9'h03f ? 6'h3f : p1_concat_10625_comb[5:0]] != 10'h000;
  assign p1_or_10663_comb = (|p1_add_10631_comb[8:6]) | p1_flat_ac_comb[p1_add_10631_comb > 9'h03f ? 6'h3f : p1_add_10631_comb[5:0]] != 10'h000;
  assign p1_or_10669_comb = (|p1_add_10630_comb[7:5]) | p1_flat_ac_comb[p1_concat_10640_comb > 9'h03f ? 6'h3f : p1_concat_10640_comb[5:0]] != 10'h000;
  assign p1_nor_10670_comb = ~((|p1_add_10647_comb[8:6]) | p1_flat_ac_comb[p1_add_10647_comb > 9'h03f ? 6'h3f : p1_add_10647_comb[5:0]] != 10'h000);
  assign p1_or_10691_comb = (|p1_add_10659_comb[5:3]) | p1_flat_ac_comb[p1_concat_10668_comb > 9'h03f ? 6'h3f : p1_concat_10668_comb[5:0]] != 10'h000;
  assign p1_or_10700_comb = (|p1_add_10672_comb[8:6]) | p1_flat_ac_comb[p1_add_10672_comb > 9'h03f ? 6'h3f : p1_add_10672_comb[5:0]] != 10'h000;
  assign p1_or_10708_comb = (|p1_add_10671_comb[7:5]) | p1_flat_ac_comb[p1_concat_10678_comb > 9'h03f ? 6'h3f : p1_concat_10678_comb[5:0]] != 10'h000;
  assign p1_or_10715_comb = (|p1_add_10685_comb[8:6]) | p1_flat_ac_comb[p1_add_10685_comb > 9'h03f ? 6'h3f : p1_add_10685_comb[5:0]] != 10'h000;
  assign p1_or_10722_comb = (|p1_add_10684_comb[6:4]) | p1_flat_ac_comb[p1_concat_10694_comb > 9'h03f ? 6'h3f : p1_concat_10694_comb[5:0]] != 10'h000;
  assign p1_or_10726_comb = (|p1_add_10702_comb[8:6]) | p1_flat_ac_comb[p1_add_10702_comb > 9'h03f ? 6'h3f : p1_add_10702_comb[5:0]] != 10'h000;
  assign p1_or_10730_comb = (|p1_add_10701_comb[7:5]) | p1_flat_ac_comb[p1_concat_10709_comb > 9'h03f ? 6'h3f : p1_concat_10709_comb[5:0]] != 10'h000;
  assign p1_nor_10733_comb = ~(p1_add_10723_comb > 9'h03e | p1_flat_ac_comb[p1_add_10723_comb > 9'h03f ? 6'h3f : p1_add_10723_comb[5:0]] != 10'h000);

  // Registers for pipe stage 1:
  reg [7:0] p1_start_pix;
  reg p1_is_luminance;
  reg [9:0] p1_flat_ac[0:63];
  reg [1:0] p1_and_10646;
  reg p1_or_10655;
  reg p1_or_10663;
  reg p1_or_10669;
  reg p1_nor_10670;
  reg p1_or_10691;
  reg p1_or_10700;
  reg p1_or_10708;
  reg p1_or_10715;
  reg p1_or_10722;
  reg p1_or_10726;
  reg p1_or_10730;
  reg p1_nor_10733;
  always @ (posedge clk) begin
    p1_start_pix <= p0_start_pix;
    p1_is_luminance <= p0_is_luminance;
    p1_flat_ac[0] <= p1_flat_ac_comb[0];
    p1_flat_ac[1] <= p1_flat_ac_comb[1];
    p1_flat_ac[2] <= p1_flat_ac_comb[2];
    p1_flat_ac[3] <= p1_flat_ac_comb[3];
    p1_flat_ac[4] <= p1_flat_ac_comb[4];
    p1_flat_ac[5] <= p1_flat_ac_comb[5];
    p1_flat_ac[6] <= p1_flat_ac_comb[6];
    p1_flat_ac[7] <= p1_flat_ac_comb[7];
    p1_flat_ac[8] <= p1_flat_ac_comb[8];
    p1_flat_ac[9] <= p1_flat_ac_comb[9];
    p1_flat_ac[10] <= p1_flat_ac_comb[10];
    p1_flat_ac[11] <= p1_flat_ac_comb[11];
    p1_flat_ac[12] <= p1_flat_ac_comb[12];
    p1_flat_ac[13] <= p1_flat_ac_comb[13];
    p1_flat_ac[14] <= p1_flat_ac_comb[14];
    p1_flat_ac[15] <= p1_flat_ac_comb[15];
    p1_flat_ac[16] <= p1_flat_ac_comb[16];
    p1_flat_ac[17] <= p1_flat_ac_comb[17];
    p1_flat_ac[18] <= p1_flat_ac_comb[18];
    p1_flat_ac[19] <= p1_flat_ac_comb[19];
    p1_flat_ac[20] <= p1_flat_ac_comb[20];
    p1_flat_ac[21] <= p1_flat_ac_comb[21];
    p1_flat_ac[22] <= p1_flat_ac_comb[22];
    p1_flat_ac[23] <= p1_flat_ac_comb[23];
    p1_flat_ac[24] <= p1_flat_ac_comb[24];
    p1_flat_ac[25] <= p1_flat_ac_comb[25];
    p1_flat_ac[26] <= p1_flat_ac_comb[26];
    p1_flat_ac[27] <= p1_flat_ac_comb[27];
    p1_flat_ac[28] <= p1_flat_ac_comb[28];
    p1_flat_ac[29] <= p1_flat_ac_comb[29];
    p1_flat_ac[30] <= p1_flat_ac_comb[30];
    p1_flat_ac[31] <= p1_flat_ac_comb[31];
    p1_flat_ac[32] <= p1_flat_ac_comb[32];
    p1_flat_ac[33] <= p1_flat_ac_comb[33];
    p1_flat_ac[34] <= p1_flat_ac_comb[34];
    p1_flat_ac[35] <= p1_flat_ac_comb[35];
    p1_flat_ac[36] <= p1_flat_ac_comb[36];
    p1_flat_ac[37] <= p1_flat_ac_comb[37];
    p1_flat_ac[38] <= p1_flat_ac_comb[38];
    p1_flat_ac[39] <= p1_flat_ac_comb[39];
    p1_flat_ac[40] <= p1_flat_ac_comb[40];
    p1_flat_ac[41] <= p1_flat_ac_comb[41];
    p1_flat_ac[42] <= p1_flat_ac_comb[42];
    p1_flat_ac[43] <= p1_flat_ac_comb[43];
    p1_flat_ac[44] <= p1_flat_ac_comb[44];
    p1_flat_ac[45] <= p1_flat_ac_comb[45];
    p1_flat_ac[46] <= p1_flat_ac_comb[46];
    p1_flat_ac[47] <= p1_flat_ac_comb[47];
    p1_flat_ac[48] <= p1_flat_ac_comb[48];
    p1_flat_ac[49] <= p1_flat_ac_comb[49];
    p1_flat_ac[50] <= p1_flat_ac_comb[50];
    p1_flat_ac[51] <= p1_flat_ac_comb[51];
    p1_flat_ac[52] <= p1_flat_ac_comb[52];
    p1_flat_ac[53] <= p1_flat_ac_comb[53];
    p1_flat_ac[54] <= p1_flat_ac_comb[54];
    p1_flat_ac[55] <= p1_flat_ac_comb[55];
    p1_flat_ac[56] <= p1_flat_ac_comb[56];
    p1_flat_ac[57] <= p1_flat_ac_comb[57];
    p1_flat_ac[58] <= p1_flat_ac_comb[58];
    p1_flat_ac[59] <= p1_flat_ac_comb[59];
    p1_flat_ac[60] <= p1_flat_ac_comb[60];
    p1_flat_ac[61] <= p1_flat_ac_comb[61];
    p1_flat_ac[62] <= p1_flat_ac_comb[62];
    p1_flat_ac[63] <= p1_flat_ac_comb[63];
    p1_and_10646 <= p1_and_10646_comb;
    p1_or_10655 <= p1_or_10655_comb;
    p1_or_10663 <= p1_or_10663_comb;
    p1_or_10669 <= p1_or_10669_comb;
    p1_nor_10670 <= p1_nor_10670_comb;
    p1_or_10691 <= p1_or_10691_comb;
    p1_or_10700 <= p1_or_10700_comb;
    p1_or_10708 <= p1_or_10708_comb;
    p1_or_10715 <= p1_or_10715_comb;
    p1_or_10722 <= p1_or_10722_comb;
    p1_or_10726 <= p1_or_10726_comb;
    p1_or_10730 <= p1_or_10730_comb;
    p1_nor_10733 <= p1_nor_10733_comb;
  end

  // ===== Pipe stage 2:
  wire [2:0] p2_and_10776_comb;
  wire [3:0] p2_sel_10785_comb;
  wire p2_next_pix__1_squeezed_squeezed_const_msb_bits__4_comb;
  wire [4:0] p2_concat_10793_comb;
  wire [4:0] p2_sign_ext_10794_comb;
  wire [9:0] p2_value_comb;
  assign p2_and_10776_comb = (p1_or_10669 ? 3'h1 : (p1_or_10663 ? 3'h2 : (p1_or_10655 ? 3'h3 : {1'h1, p1_and_10646}))) & {3{p1_nor_10670}};
  assign p2_sel_10785_comb = p1_or_10715 ? 4'h4 : (p1_or_10708 ? 4'h5 : (p1_or_10700 ? 4'h6 : (p1_or_10691 ? 4'h7 : {1'h1, p2_and_10776_comb})));
  assign p2_next_pix__1_squeezed_squeezed_const_msb_bits__4_comb = 1'h0;
  assign p2_concat_10793_comb = {p2_next_pix__1_squeezed_squeezed_const_msb_bits__4_comb, p1_or_10730 ? 4'h1 : (p1_or_10726 ? 4'h2 : (p1_or_10722 ? 4'h3 : p2_sel_10785_comb))};
  assign p2_sign_ext_10794_comb = {5{p1_nor_10733}};
  assign p2_value_comb = p1_flat_ac[p1_start_pix > 8'h3f ? 6'h3f : p1_start_pix[5:0]];

  // Registers for pipe stage 2:
  reg [7:0] p2_start_pix;
  reg p2_is_luminance;
  reg [9:0] p2_flat_ac[0:63];
  reg [4:0] p2_concat_10793;
  reg [4:0] p2_sign_ext_10794;
  reg [9:0] p2_value;
  always @ (posedge clk) begin
    p2_start_pix <= p1_start_pix;
    p2_is_luminance <= p1_is_luminance;
    p2_flat_ac[0] <= p1_flat_ac[0];
    p2_flat_ac[1] <= p1_flat_ac[1];
    p2_flat_ac[2] <= p1_flat_ac[2];
    p2_flat_ac[3] <= p1_flat_ac[3];
    p2_flat_ac[4] <= p1_flat_ac[4];
    p2_flat_ac[5] <= p1_flat_ac[5];
    p2_flat_ac[6] <= p1_flat_ac[6];
    p2_flat_ac[7] <= p1_flat_ac[7];
    p2_flat_ac[8] <= p1_flat_ac[8];
    p2_flat_ac[9] <= p1_flat_ac[9];
    p2_flat_ac[10] <= p1_flat_ac[10];
    p2_flat_ac[11] <= p1_flat_ac[11];
    p2_flat_ac[12] <= p1_flat_ac[12];
    p2_flat_ac[13] <= p1_flat_ac[13];
    p2_flat_ac[14] <= p1_flat_ac[14];
    p2_flat_ac[15] <= p1_flat_ac[15];
    p2_flat_ac[16] <= p1_flat_ac[16];
    p2_flat_ac[17] <= p1_flat_ac[17];
    p2_flat_ac[18] <= p1_flat_ac[18];
    p2_flat_ac[19] <= p1_flat_ac[19];
    p2_flat_ac[20] <= p1_flat_ac[20];
    p2_flat_ac[21] <= p1_flat_ac[21];
    p2_flat_ac[22] <= p1_flat_ac[22];
    p2_flat_ac[23] <= p1_flat_ac[23];
    p2_flat_ac[24] <= p1_flat_ac[24];
    p2_flat_ac[25] <= p1_flat_ac[25];
    p2_flat_ac[26] <= p1_flat_ac[26];
    p2_flat_ac[27] <= p1_flat_ac[27];
    p2_flat_ac[28] <= p1_flat_ac[28];
    p2_flat_ac[29] <= p1_flat_ac[29];
    p2_flat_ac[30] <= p1_flat_ac[30];
    p2_flat_ac[31] <= p1_flat_ac[31];
    p2_flat_ac[32] <= p1_flat_ac[32];
    p2_flat_ac[33] <= p1_flat_ac[33];
    p2_flat_ac[34] <= p1_flat_ac[34];
    p2_flat_ac[35] <= p1_flat_ac[35];
    p2_flat_ac[36] <= p1_flat_ac[36];
    p2_flat_ac[37] <= p1_flat_ac[37];
    p2_flat_ac[38] <= p1_flat_ac[38];
    p2_flat_ac[39] <= p1_flat_ac[39];
    p2_flat_ac[40] <= p1_flat_ac[40];
    p2_flat_ac[41] <= p1_flat_ac[41];
    p2_flat_ac[42] <= p1_flat_ac[42];
    p2_flat_ac[43] <= p1_flat_ac[43];
    p2_flat_ac[44] <= p1_flat_ac[44];
    p2_flat_ac[45] <= p1_flat_ac[45];
    p2_flat_ac[46] <= p1_flat_ac[46];
    p2_flat_ac[47] <= p1_flat_ac[47];
    p2_flat_ac[48] <= p1_flat_ac[48];
    p2_flat_ac[49] <= p1_flat_ac[49];
    p2_flat_ac[50] <= p1_flat_ac[50];
    p2_flat_ac[51] <= p1_flat_ac[51];
    p2_flat_ac[52] <= p1_flat_ac[52];
    p2_flat_ac[53] <= p1_flat_ac[53];
    p2_flat_ac[54] <= p1_flat_ac[54];
    p2_flat_ac[55] <= p1_flat_ac[55];
    p2_flat_ac[56] <= p1_flat_ac[56];
    p2_flat_ac[57] <= p1_flat_ac[57];
    p2_flat_ac[58] <= p1_flat_ac[58];
    p2_flat_ac[59] <= p1_flat_ac[59];
    p2_flat_ac[60] <= p1_flat_ac[60];
    p2_flat_ac[61] <= p1_flat_ac[61];
    p2_flat_ac[62] <= p1_flat_ac[62];
    p2_flat_ac[63] <= p1_flat_ac[63];
    p2_concat_10793 <= p2_concat_10793_comb;
    p2_sign_ext_10794 <= p2_sign_ext_10794_comb;
    p2_value <= p2_value_comb;
  end

  // ===== Pipe stage 3:
  wire [4:0] p3_zero_num__1_comb;
  wire p3_ne_10811_comb;
  wire [2:0] p3_run_0_squeezed_const_msb_bits__1_comb;
  wire [4:0] p3_add_10813_comb;
  wire [7:0] p3_sign_ext_10816_comb;
  wire [7:0] p3_start_pix_1__1_comb;
  wire [7:0] p3_value_pix_num_comb;
  wire [7:0] p3_add_10818_comb;
  wire [7:0] p3_actual_index__65_comb;
  wire [6:0] p3_add_10918_comb;
  wire [7:0] p3_actual_index__67_comb;
  wire [5:0] p3_add_10920_comb;
  wire [7:0] p3_actual_index__69_comb;
  wire [6:0] p3_add_10922_comb;
  wire [7:0] p3_actual_index__71_comb;
  wire [4:0] p3_add_10924_comb;
  wire [7:0] p3_actual_index__73_comb;
  wire [6:0] p3_add_10926_comb;
  wire [7:0] p3_actual_index__75_comb;
  wire [5:0] p3_add_10928_comb;
  wire [7:0] p3_actual_index__77_comb;
  wire [6:0] p3_add_10930_comb;
  wire [7:0] p3_actual_index__79_comb;
  wire [3:0] p3_add_10932_comb;
  wire [7:0] p3_actual_index__81_comb;
  wire [6:0] p3_add_10934_comb;
  wire [7:0] p3_actual_index__83_comb;
  wire [5:0] p3_add_10936_comb;
  wire [7:0] p3_actual_index__85_comb;
  wire [6:0] p3_add_10938_comb;
  wire [7:0] p3_actual_index__87_comb;
  wire [4:0] p3_add_10940_comb;
  wire [7:0] p3_actual_index__89_comb;
  wire [6:0] p3_add_10942_comb;
  wire [7:0] p3_actual_index__91_comb;
  wire [5:0] p3_add_10944_comb;
  wire [7:0] p3_actual_index__93_comb;
  wire [6:0] p3_add_10946_comb;
  wire [7:0] p3_actual_index__95_comb;
  wire [2:0] p3_add_10948_comb;
  wire [7:0] p3_actual_index__97_comb;
  wire [6:0] p3_add_10950_comb;
  wire [7:0] p3_actual_index__99_comb;
  wire [5:0] p3_add_10952_comb;
  wire [7:0] p3_actual_index__101_comb;
  wire [6:0] p3_add_10954_comb;
  wire [7:0] p3_actual_index__103_comb;
  wire [4:0] p3_add_10956_comb;
  wire [7:0] p3_actual_index__105_comb;
  wire [6:0] p3_add_10958_comb;
  wire [7:0] p3_actual_index__107_comb;
  wire [5:0] p3_add_10960_comb;
  wire [7:0] p3_actual_index__109_comb;
  wire [6:0] p3_add_10962_comb;
  wire [7:0] p3_actual_index__111_comb;
  wire [3:0] p3_add_10964_comb;
  wire [7:0] p3_actual_index__113_comb;
  wire [6:0] p3_add_10966_comb;
  wire [7:0] p3_actual_index__115_comb;
  wire [5:0] p3_add_10968_comb;
  wire [7:0] p3_actual_index__117_comb;
  wire [6:0] p3_add_10970_comb;
  wire [7:0] p3_actual_index__119_comb;
  wire [4:0] p3_add_10972_comb;
  wire [7:0] p3_actual_index__121_comb;
  wire [6:0] p3_add_10974_comb;
  wire [7:0] p3_actual_index__123_comb;
  wire [5:0] p3_add_10976_comb;
  wire [7:0] p3_actual_index__125_comb;
  wire [6:0] p3_add_10978_comb;
  wire [7:0] p3_actual_index__127_comb;
  wire [9:0] p3_value__1_comb;
  wire [7:0] p3_bin_value__1_comb;
  wire [7:0] p3_actual_index__66_comb;
  wire [7:0] p3_actual_index__68_comb;
  wire [7:0] p3_actual_index__70_comb;
  wire [7:0] p3_actual_index__72_comb;
  wire [7:0] p3_actual_index__74_comb;
  wire [7:0] p3_actual_index__76_comb;
  wire [7:0] p3_actual_index__78_comb;
  wire [7:0] p3_actual_index__80_comb;
  wire [7:0] p3_actual_index__82_comb;
  wire [7:0] p3_actual_index__84_comb;
  wire [7:0] p3_actual_index__86_comb;
  wire [7:0] p3_actual_index__88_comb;
  wire [7:0] p3_actual_index__90_comb;
  wire [7:0] p3_actual_index__92_comb;
  wire [7:0] p3_actual_index__94_comb;
  wire [7:0] p3_actual_index__96_comb;
  wire [7:0] p3_actual_index__98_comb;
  wire [7:0] p3_actual_index__100_comb;
  wire [7:0] p3_actual_index__102_comb;
  wire [7:0] p3_actual_index__104_comb;
  wire [7:0] p3_actual_index__106_comb;
  wire [7:0] p3_actual_index__108_comb;
  wire [7:0] p3_actual_index__110_comb;
  wire [7:0] p3_actual_index__112_comb;
  wire [7:0] p3_actual_index__114_comb;
  wire [7:0] p3_actual_index__116_comb;
  wire [7:0] p3_actual_index__118_comb;
  wire [7:0] p3_actual_index__120_comb;
  wire [7:0] p3_actual_index__122_comb;
  wire [7:0] p3_actual_index__124_comb;
  wire [7:0] p3_actual_index__126_comb;
  wire [7:0] p3_bin_value_comb;
  wire [7:0] p3_value_abs_comb;
  wire [4:0] p3_next_pix_0_squeezed__1_comb;
  wire p3_and_11538_comb;
  wire [2:0] p3_run_0_squeezed_const_msb_bits__2_comb;
  wire [4:0] p3_run_0_squeezed_comb;
  wire [4:0] p3_next_pix_1_squeezed_squeezed_comb;
  wire [7:0] p3_flipped_comb;
  wire p3_next_pix__1_squeezed_squeezed_const_msb_bits__1_comb;
  wire [7:0] p3_run_0_comb;
  wire [7:0] p3_Code_list_comb;
  wire p3_or_reduce_10837_comb;
  wire [2:0] p3_concat_10838_comb;
  wire p3_or_reduce_10842_comb;
  wire p3_or_reduce_10845_comb;
  wire p3_or_reduce_10916_comb;
  wire p3_bit_slice_11116_comb;
  wire p3_eq_11117_comb;
  wire [7:0] p3_run__1_comb;
  wire [4:0] p3_next_pix__1_squeezed_squeezed_comb;
  wire [7:0] p3_code_list_comb;
  assign p3_zero_num__1_comb = p2_concat_10793 & p2_sign_ext_10794;
  assign p3_ne_10811_comb = p2_value != 10'h000;
  assign p3_run_0_squeezed_const_msb_bits__1_comb = 3'h0;
  assign p3_add_10813_comb = p3_zero_num__1_comb + 5'h01;
  assign p3_sign_ext_10816_comb = {8{~p3_ne_10811_comb}};
  assign p3_start_pix_1__1_comb = p2_start_pix > 8'h40 ? 8'h40 : p2_start_pix;
  assign p3_value_pix_num_comb = {p3_run_0_squeezed_const_msb_bits__1_comb, p3_add_10813_comb} & p3_sign_ext_10816_comb;
  assign p3_add_10818_comb = p2_start_pix + p3_value_pix_num_comb;
  assign p3_actual_index__65_comb = p3_start_pix_1__1_comb + 8'h01;
  assign p3_add_10918_comb = p3_start_pix_1__1_comb[7:1] + 7'h01;
  assign p3_actual_index__67_comb = p3_start_pix_1__1_comb + 8'h03;
  assign p3_add_10920_comb = p3_start_pix_1__1_comb[7:2] + 6'h01;
  assign p3_actual_index__69_comb = p3_start_pix_1__1_comb + 8'h05;
  assign p3_add_10922_comb = p3_start_pix_1__1_comb[7:1] + 7'h03;
  assign p3_actual_index__71_comb = p3_start_pix_1__1_comb + 8'h07;
  assign p3_add_10924_comb = p3_start_pix_1__1_comb[7:3] + 5'h01;
  assign p3_actual_index__73_comb = p3_start_pix_1__1_comb + 8'h09;
  assign p3_add_10926_comb = p3_start_pix_1__1_comb[7:1] + 7'h05;
  assign p3_actual_index__75_comb = p3_start_pix_1__1_comb + 8'h0b;
  assign p3_add_10928_comb = p3_start_pix_1__1_comb[7:2] + 6'h03;
  assign p3_actual_index__77_comb = p3_start_pix_1__1_comb + 8'h0d;
  assign p3_add_10930_comb = p3_start_pix_1__1_comb[7:1] + 7'h07;
  assign p3_actual_index__79_comb = p3_start_pix_1__1_comb + 8'h0f;
  assign p3_add_10932_comb = p3_start_pix_1__1_comb[7:4] + 4'h1;
  assign p3_actual_index__81_comb = p3_start_pix_1__1_comb + 8'h11;
  assign p3_add_10934_comb = p3_start_pix_1__1_comb[7:1] + 7'h09;
  assign p3_actual_index__83_comb = p3_start_pix_1__1_comb + 8'h13;
  assign p3_add_10936_comb = p3_start_pix_1__1_comb[7:2] + 6'h05;
  assign p3_actual_index__85_comb = p3_start_pix_1__1_comb + 8'h15;
  assign p3_add_10938_comb = p3_start_pix_1__1_comb[7:1] + 7'h0b;
  assign p3_actual_index__87_comb = p3_start_pix_1__1_comb + 8'h17;
  assign p3_add_10940_comb = p3_start_pix_1__1_comb[7:3] + 5'h03;
  assign p3_actual_index__89_comb = p3_start_pix_1__1_comb + 8'h19;
  assign p3_add_10942_comb = p3_start_pix_1__1_comb[7:1] + 7'h0d;
  assign p3_actual_index__91_comb = p3_start_pix_1__1_comb + 8'h1b;
  assign p3_add_10944_comb = p3_start_pix_1__1_comb[7:2] + 6'h07;
  assign p3_actual_index__93_comb = p3_start_pix_1__1_comb + 8'h1d;
  assign p3_add_10946_comb = p3_start_pix_1__1_comb[7:1] + 7'h0f;
  assign p3_actual_index__95_comb = p3_start_pix_1__1_comb + 8'h1f;
  assign p3_add_10948_comb = p3_start_pix_1__1_comb[7:5] + 3'h1;
  assign p3_actual_index__97_comb = p3_start_pix_1__1_comb + 8'h21;
  assign p3_add_10950_comb = p3_start_pix_1__1_comb[7:1] + 7'h11;
  assign p3_actual_index__99_comb = p3_start_pix_1__1_comb + 8'h23;
  assign p3_add_10952_comb = p3_start_pix_1__1_comb[7:2] + 6'h09;
  assign p3_actual_index__101_comb = p3_start_pix_1__1_comb + 8'h25;
  assign p3_add_10954_comb = p3_start_pix_1__1_comb[7:1] + 7'h13;
  assign p3_actual_index__103_comb = p3_start_pix_1__1_comb + 8'h27;
  assign p3_add_10956_comb = p3_start_pix_1__1_comb[7:3] + 5'h05;
  assign p3_actual_index__105_comb = p3_start_pix_1__1_comb + 8'h29;
  assign p3_add_10958_comb = p3_start_pix_1__1_comb[7:1] + 7'h15;
  assign p3_actual_index__107_comb = p3_start_pix_1__1_comb + 8'h2b;
  assign p3_add_10960_comb = p3_start_pix_1__1_comb[7:2] + 6'h0b;
  assign p3_actual_index__109_comb = p3_start_pix_1__1_comb + 8'h2d;
  assign p3_add_10962_comb = p3_start_pix_1__1_comb[7:1] + 7'h17;
  assign p3_actual_index__111_comb = p3_start_pix_1__1_comb + 8'h2f;
  assign p3_add_10964_comb = p3_start_pix_1__1_comb[7:4] + 4'h3;
  assign p3_actual_index__113_comb = p3_start_pix_1__1_comb + 8'h31;
  assign p3_add_10966_comb = p3_start_pix_1__1_comb[7:1] + 7'h19;
  assign p3_actual_index__115_comb = p3_start_pix_1__1_comb + 8'h33;
  assign p3_add_10968_comb = p3_start_pix_1__1_comb[7:2] + 6'h0d;
  assign p3_actual_index__117_comb = p3_start_pix_1__1_comb + 8'h35;
  assign p3_add_10970_comb = p3_start_pix_1__1_comb[7:1] + 7'h1b;
  assign p3_actual_index__119_comb = p3_start_pix_1__1_comb + 8'h37;
  assign p3_add_10972_comb = p3_start_pix_1__1_comb[7:3] + 5'h07;
  assign p3_actual_index__121_comb = p3_start_pix_1__1_comb + 8'h39;
  assign p3_add_10974_comb = p3_start_pix_1__1_comb[7:1] + 7'h1d;
  assign p3_actual_index__123_comb = p3_start_pix_1__1_comb + 8'h3b;
  assign p3_add_10976_comb = p3_start_pix_1__1_comb[7:2] + 6'h0f;
  assign p3_actual_index__125_comb = p3_start_pix_1__1_comb + 8'h3d;
  assign p3_add_10978_comb = p3_start_pix_1__1_comb[7:1] + 7'h1f;
  assign p3_actual_index__127_comb = p3_start_pix_1__1_comb + 8'h3f;
  assign p3_value__1_comb = p2_flat_ac[p3_add_10818_comb > 8'h3f ? 6'h3f : p3_add_10818_comb[5:0]];
  assign p3_bin_value__1_comb = p3_value__1_comb[7:0];
  assign p3_actual_index__66_comb = {p3_add_10918_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__68_comb = {p3_add_10920_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__70_comb = {p3_add_10922_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__72_comb = {p3_add_10924_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__74_comb = {p3_add_10926_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__76_comb = {p3_add_10928_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__78_comb = {p3_add_10930_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__80_comb = {p3_add_10932_comb, p3_start_pix_1__1_comb[3:0]};
  assign p3_actual_index__82_comb = {p3_add_10934_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__84_comb = {p3_add_10936_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__86_comb = {p3_add_10938_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__88_comb = {p3_add_10940_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__90_comb = {p3_add_10942_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__92_comb = {p3_add_10944_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__94_comb = {p3_add_10946_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__96_comb = {p3_add_10948_comb, p3_start_pix_1__1_comb[4:0]};
  assign p3_actual_index__98_comb = {p3_add_10950_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__100_comb = {p3_add_10952_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__102_comb = {p3_add_10954_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__104_comb = {p3_add_10956_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__106_comb = {p3_add_10958_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__108_comb = {p3_add_10960_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__110_comb = {p3_add_10962_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__112_comb = {p3_add_10964_comb, p3_start_pix_1__1_comb[3:0]};
  assign p3_actual_index__114_comb = {p3_add_10966_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__116_comb = {p3_add_10968_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__118_comb = {p3_add_10970_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__120_comb = {p3_add_10972_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__122_comb = {p3_add_10974_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__124_comb = {p3_add_10976_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__126_comb = {p3_add_10978_comb, p3_start_pix_1__1_comb[0]};
  assign p3_bin_value_comb = -p3_bin_value__1_comb;
  assign p3_value_abs_comb = p3_value__1_comb[9] ? p3_bin_value_comb : p3_bin_value__1_comb;
  assign p3_next_pix_0_squeezed__1_comb = p3_add_10813_comb + 5'h01;
  assign p3_and_11538_comb = (p2_value & {10{~p3_start_pix_1__1_comb[6]}}) == 10'h000 & (p2_flat_ac[p3_actual_index__65_comb > 8'h3f ? 6'h3f : p3_actual_index__65_comb[5:0]] & {10{~(p3_actual_index__65_comb[6] | p3_actual_index__65_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__66_comb > 8'h3f ? 6'h3f : p3_actual_index__66_comb[5:0]] & {10{~(p3_add_10918_comb[5] | p3_add_10918_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__67_comb > 8'h3f ? 6'h3f : p3_actual_index__67_comb[5:0]] & {10{~(p3_actual_index__67_comb[6] | p3_actual_index__67_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__68_comb > 8'h3f ? 6'h3f : p3_actual_index__68_comb[5:0]] & {10{~(p3_add_10920_comb[4] | p3_add_10920_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__69_comb > 8'h3f ? 6'h3f : p3_actual_index__69_comb[5:0]] & {10{~(p3_actual_index__69_comb[6] | p3_actual_index__69_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__70_comb > 8'h3f ? 6'h3f : p3_actual_index__70_comb[5:0]] & {10{~(p3_add_10922_comb[5] | p3_add_10922_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__71_comb > 8'h3f ? 6'h3f : p3_actual_index__71_comb[5:0]] & {10{~(p3_actual_index__71_comb[6] | p3_actual_index__71_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__72_comb > 8'h3f ? 6'h3f : p3_actual_index__72_comb[5:0]] & {10{~(p3_add_10924_comb[3] | p3_add_10924_comb[4])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__73_comb > 8'h3f ? 6'h3f : p3_actual_index__73_comb[5:0]] & {10{~(p3_actual_index__73_comb[6] | p3_actual_index__73_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__74_comb > 8'h3f ? 6'h3f : p3_actual_index__74_comb[5:0]] & {10{~(p3_add_10926_comb[5] | p3_add_10926_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__75_comb > 8'h3f ? 6'h3f : p3_actual_index__75_comb[5:0]] & {10{~(p3_actual_index__75_comb[6] | p3_actual_index__75_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__76_comb > 8'h3f ? 6'h3f : p3_actual_index__76_comb[5:0]] & {10{~(p3_add_10928_comb[4] | p3_add_10928_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__77_comb > 8'h3f ? 6'h3f : p3_actual_index__77_comb[5:0]] & {10{~(p3_actual_index__77_comb[6] | p3_actual_index__77_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__78_comb > 8'h3f ? 6'h3f : p3_actual_index__78_comb[5:0]] & {10{~(p3_add_10930_comb[5] | p3_add_10930_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__79_comb > 8'h3f ? 6'h3f : p3_actual_index__79_comb[5:0]] & {10{~(p3_actual_index__79_comb[6] | p3_actual_index__79_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__80_comb > 8'h3f ? 6'h3f : p3_actual_index__80_comb[5:0]] & {10{~(p3_add_10932_comb[2] | p3_add_10932_comb[3])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__81_comb > 8'h3f ? 6'h3f : p3_actual_index__81_comb[5:0]] & {10{~(p3_actual_index__81_comb[6] | p3_actual_index__81_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__82_comb > 8'h3f ? 6'h3f : p3_actual_index__82_comb[5:0]] & {10{~(p3_add_10934_comb[5] | p3_add_10934_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__83_comb > 8'h3f ? 6'h3f : p3_actual_index__83_comb[5:0]] & {10{~(p3_actual_index__83_comb[6] | p3_actual_index__83_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__84_comb > 8'h3f ? 6'h3f : p3_actual_index__84_comb[5:0]] & {10{~(p3_add_10936_comb[4] | p3_add_10936_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__85_comb > 8'h3f ? 6'h3f : p3_actual_index__85_comb[5:0]] & {10{~(p3_actual_index__85_comb[6] | p3_actual_index__85_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__86_comb > 8'h3f ? 6'h3f : p3_actual_index__86_comb[5:0]] & {10{~(p3_add_10938_comb[5] | p3_add_10938_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__87_comb > 8'h3f ? 6'h3f : p3_actual_index__87_comb[5:0]] & {10{~(p3_actual_index__87_comb[6] | p3_actual_index__87_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__88_comb > 8'h3f ? 6'h3f : p3_actual_index__88_comb[5:0]] & {10{~(p3_add_10940_comb[3] | p3_add_10940_comb[4])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__89_comb > 8'h3f ? 6'h3f : p3_actual_index__89_comb[5:0]] & {10{~(p3_actual_index__89_comb[6] | p3_actual_index__89_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__90_comb > 8'h3f ? 6'h3f : p3_actual_index__90_comb[5:0]] & {10{~(p3_add_10942_comb[5] | p3_add_10942_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__91_comb > 8'h3f ? 6'h3f : p3_actual_index__91_comb[5:0]] & {10{~(p3_actual_index__91_comb[6] | p3_actual_index__91_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__92_comb > 8'h3f ? 6'h3f : p3_actual_index__92_comb[5:0]] & {10{~(p3_add_10944_comb[4] | p3_add_10944_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__93_comb > 8'h3f ? 6'h3f : p3_actual_index__93_comb[5:0]] & {10{~(p3_actual_index__93_comb[6] | p3_actual_index__93_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__94_comb > 8'h3f ? 6'h3f : p3_actual_index__94_comb[5:0]] & {10{~(p3_add_10946_comb[5] | p3_add_10946_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__95_comb > 8'h3f ? 6'h3f : p3_actual_index__95_comb[5:0]] & {10{~(p3_actual_index__95_comb[6] | p3_actual_index__95_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__96_comb > 8'h3f ? 6'h3f : p3_actual_index__96_comb[5:0]] & {10{~(p3_add_10948_comb[1] | p3_add_10948_comb[2])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__97_comb > 8'h3f ? 6'h3f : p3_actual_index__97_comb[5:0]] & {10{~(p3_actual_index__97_comb[6] | p3_actual_index__97_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__98_comb > 8'h3f ? 6'h3f : p3_actual_index__98_comb[5:0]] & {10{~(p3_add_10950_comb[5] | p3_add_10950_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__99_comb > 8'h3f ? 6'h3f : p3_actual_index__99_comb[5:0]] & {10{~(p3_actual_index__99_comb[6] | p3_actual_index__99_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__100_comb > 8'h3f ? 6'h3f : p3_actual_index__100_comb[5:0]] & {10{~(p3_add_10952_comb[4] | p3_add_10952_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__101_comb > 8'h3f ? 6'h3f : p3_actual_index__101_comb[5:0]] & {10{~(p3_actual_index__101_comb[6] | p3_actual_index__101_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__102_comb > 8'h3f ? 6'h3f : p3_actual_index__102_comb[5:0]] & {10{~(p3_add_10954_comb[5] | p3_add_10954_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__103_comb > 8'h3f ? 6'h3f : p3_actual_index__103_comb[5:0]] & {10{~(p3_actual_index__103_comb[6] | p3_actual_index__103_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__104_comb > 8'h3f ? 6'h3f : p3_actual_index__104_comb[5:0]] & {10{~(p3_add_10956_comb[3] | p3_add_10956_comb[4])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__105_comb > 8'h3f ? 6'h3f : p3_actual_index__105_comb[5:0]] & {10{~(p3_actual_index__105_comb[6] | p3_actual_index__105_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__106_comb > 8'h3f ? 6'h3f : p3_actual_index__106_comb[5:0]] & {10{~(p3_add_10958_comb[5] | p3_add_10958_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__107_comb > 8'h3f ? 6'h3f : p3_actual_index__107_comb[5:0]] & {10{~(p3_actual_index__107_comb[6] | p3_actual_index__107_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__108_comb > 8'h3f ? 6'h3f : p3_actual_index__108_comb[5:0]] & {10{~(p3_add_10960_comb[4] | p3_add_10960_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__109_comb > 8'h3f ? 6'h3f : p3_actual_index__109_comb[5:0]] & {10{~(p3_actual_index__109_comb[6] | p3_actual_index__109_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__110_comb > 8'h3f ? 6'h3f : p3_actual_index__110_comb[5:0]] & {10{~(p3_add_10962_comb[5] | p3_add_10962_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__111_comb > 8'h3f ? 6'h3f : p3_actual_index__111_comb[5:0]] & {10{~(p3_actual_index__111_comb[6] | p3_actual_index__111_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__112_comb > 8'h3f ? 6'h3f : p3_actual_index__112_comb[5:0]] & {10{~(p3_add_10964_comb[2] | p3_add_10964_comb[3])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__113_comb > 8'h3f ? 6'h3f : p3_actual_index__113_comb[5:0]] & {10{~(p3_actual_index__113_comb[6] | p3_actual_index__113_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__114_comb > 8'h3f ? 6'h3f : p3_actual_index__114_comb[5:0]] & {10{~(p3_add_10966_comb[5] | p3_add_10966_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__115_comb > 8'h3f ? 6'h3f : p3_actual_index__115_comb[5:0]] & {10{~(p3_actual_index__115_comb[6] | p3_actual_index__115_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__116_comb > 8'h3f ? 6'h3f : p3_actual_index__116_comb[5:0]] & {10{~(p3_add_10968_comb[4] | p3_add_10968_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__117_comb > 8'h3f ? 6'h3f : p3_actual_index__117_comb[5:0]] & {10{~(p3_actual_index__117_comb[6] | p3_actual_index__117_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__118_comb > 8'h3f ? 6'h3f : p3_actual_index__118_comb[5:0]] & {10{~(p3_add_10970_comb[5] | p3_add_10970_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__119_comb > 8'h3f ? 6'h3f : p3_actual_index__119_comb[5:0]] & {10{~(p3_actual_index__119_comb[6] | p3_actual_index__119_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__120_comb > 8'h3f ? 6'h3f : p3_actual_index__120_comb[5:0]] & {10{~(p3_add_10972_comb[3] | p3_add_10972_comb[4])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__121_comb > 8'h3f ? 6'h3f : p3_actual_index__121_comb[5:0]] & {10{~(p3_actual_index__121_comb[6] | p3_actual_index__121_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__122_comb > 8'h3f ? 6'h3f : p3_actual_index__122_comb[5:0]] & {10{~(p3_add_10974_comb[5] | p3_add_10974_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__123_comb > 8'h3f ? 6'h3f : p3_actual_index__123_comb[5:0]] & {10{~(p3_actual_index__123_comb[6] | p3_actual_index__123_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__124_comb > 8'h3f ? 6'h3f : p3_actual_index__124_comb[5:0]] & {10{~(p3_add_10976_comb[4] | p3_add_10976_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__125_comb > 8'h3f ? 6'h3f : p3_actual_index__125_comb[5:0]] & {10{~(p3_actual_index__125_comb[6] | p3_actual_index__125_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__126_comb > 8'h3f ? 6'h3f : p3_actual_index__126_comb[5:0]] & {10{~(p3_add_10978_comb[5] | p3_add_10978_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__127_comb > 8'h3f ? 6'h3f : p3_actual_index__127_comb[5:0]] & {10{~(p3_actual_index__127_comb[6] | p3_actual_index__127_comb[7])}}) == 10'h000;
  assign p3_run_0_squeezed_const_msb_bits__2_comb = 3'h0;
  assign p3_run_0_squeezed_comb = p3_add_10813_comb[4] ? 5'h0f : p3_add_10813_comb;
  assign p3_next_pix_1_squeezed_squeezed_comb = p3_ne_10811_comb ? 5'h01 : p3_next_pix_0_squeezed__1_comb;
  assign p3_flipped_comb = ~p3_bin_value_comb;
  assign p3_next_pix__1_squeezed_squeezed_const_msb_bits__1_comb = 1'h0;
  assign p3_run_0_comb = {p3_run_0_squeezed_const_msb_bits__2_comb, p3_run_0_squeezed_comb};
  assign p3_Code_list_comb = $signed(p3_value__1_comb) <= $signed(10'h000) ? p3_flipped_comb : p3_bin_value__1_comb;
  assign p3_or_reduce_10837_comb = |p3_value_abs_comb[7:3];
  assign p3_concat_10838_comb = {p3_next_pix__1_squeezed_squeezed_const_msb_bits__1_comb, |p3_value_abs_comb[7:2] ? 2'h3 : (|p3_value_abs_comb[7:1] ? 2'h2 : 2'h1)};
  assign p3_or_reduce_10842_comb = |p3_value_abs_comb[7:4];
  assign p3_or_reduce_10845_comb = |p3_value_abs_comb[7:5];
  assign p3_or_reduce_10916_comb = |p3_value_abs_comb[7:6];
  assign p3_bit_slice_11116_comb = p3_value_abs_comb[7];
  assign p3_eq_11117_comb = p3_value_abs_comb == 8'h00;
  assign p3_run__1_comb = p3_run_0_comb & p3_sign_ext_10816_comb;
  assign p3_next_pix__1_squeezed_squeezed_comb = p3_next_pix_1_squeezed_squeezed_comb > 5'h10 ? 5'h10 : p3_next_pix_1_squeezed_squeezed_comb;
  assign p3_code_list_comb = p3_Code_list_comb & {8{~p3_and_11538_comb}};

  // Registers for pipe stage 3:
  reg p3_is_luminance;
  reg [9:0] p3_value;
  reg p3_or_reduce_10837;
  reg [2:0] p3_concat_10838;
  reg p3_or_reduce_10842;
  reg p3_or_reduce_10845;
  reg p3_or_reduce_10916;
  reg p3_bit_slice_11116;
  reg p3_eq_11117;
  reg [7:0] p3_run__1;
  reg p3_and_11538;
  reg [4:0] p3_next_pix__1_squeezed_squeezed;
  reg [7:0] p3_code_list;
  always @ (posedge clk) begin
    p3_is_luminance <= p2_is_luminance;
    p3_value <= p2_value;
    p3_or_reduce_10837 <= p3_or_reduce_10837_comb;
    p3_concat_10838 <= p3_concat_10838_comb;
    p3_or_reduce_10842 <= p3_or_reduce_10842_comb;
    p3_or_reduce_10845 <= p3_or_reduce_10845_comb;
    p3_or_reduce_10916 <= p3_or_reduce_10916_comb;
    p3_bit_slice_11116 <= p3_bit_slice_11116_comb;
    p3_eq_11117 <= p3_eq_11117_comb;
    p3_run__1 <= p3_run__1_comb;
    p3_and_11538 <= p3_and_11538_comb;
    p3_next_pix__1_squeezed_squeezed <= p3_next_pix__1_squeezed_squeezed_comb;
    p3_code_list <= p3_code_list_comb;
  end

  // ===== Pipe stage 4:
  wire p4_next_pix__1_squeezed_squeezed_const_msb_bits__2_comb;
  wire [3:0] p4_concat_11584_comb;
  wire [7:0] p4_concat_11591_comb;
  wire [7:0] p4_Code_size_comb;
  wire [7:0] p4_run_size_str_u8_comb;
  wire [2:0] p4_sel_11604_comb;
  wire [1:0] p4_next_pix_squeezed_const_msb_bits_comb;
  wire p4_next_pix__1_squeezed_squeezed_const_msb_bits__3_comb;
  wire p4_next_pix__1_squeezed_squeezed_const_msb_bits__8_comb;
  wire [4:0] p4_Huffman_length_squeezed_comb;
  wire [5:0] p4_next_pix__1_squeezed_comb;
  wire [5:0] p4_run__1_squeezed_comb;
  wire [15:0] p4_Huffman_code_full_comb;
  wire [2:0] p4_run_0_squeezed_const_msb_bits__3_comb;
  wire [4:0] p4_huff_length_squeezed_comb;
  wire [1:0] p4_next_pix_squeezed_const_msb_bits__1_comb;
  wire [5:0] p4_next_pix_squeezed_comb;
  wire [1:0] p4_next_pix_squeezed_const_msb_bits__2_comb;
  wire [5:0] p4_run_squeezed_comb;
  wire [15:0] p4_huff_code_comb;
  wire [7:0] p4_huff_length_comb;
  wire [7:0] p4_code_size_comb;
  wire [7:0] p4_next_pix_comb;
  wire [7:0] p4_run_comb;
  wire [65:0] p4_tuple_11637_comb;
  assign p4_next_pix__1_squeezed_squeezed_const_msb_bits__2_comb = 1'h0;
  assign p4_concat_11584_comb = {p4_next_pix__1_squeezed_squeezed_const_msb_bits__2_comb, p3_or_reduce_10916 ? 3'h7 : (p3_or_reduce_10845 ? 3'h6 : (p3_or_reduce_10842 ? 3'h5 : (p3_or_reduce_10837 ? 3'h4 : p3_concat_10838)))};
  assign p4_concat_11591_comb = {4'h0, p3_bit_slice_11116 ? 4'h8 : p4_concat_11584_comb};
  assign p4_Code_size_comb = p4_concat_11591_comb & {8{~p3_eq_11117}};
  assign p4_run_size_str_u8_comb = {p3_run__1[3:0], 4'h0} | p4_Code_size_comb;
  assign p4_sel_11604_comb = p3_is_luminance ? 3'h4 : 3'h1;
  assign p4_next_pix_squeezed_const_msb_bits_comb = 2'h0;
  assign p4_next_pix__1_squeezed_squeezed_const_msb_bits__3_comb = 1'h0;
  assign p4_next_pix__1_squeezed_squeezed_const_msb_bits__8_comb = 1'h0;
  assign p4_Huffman_length_squeezed_comb = p3_is_luminance ? literal_11599[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_11597[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_next_pix__1_squeezed_comb = {p4_next_pix__1_squeezed_squeezed_const_msb_bits__8_comb, p3_next_pix__1_squeezed_squeezed};
  assign p4_run__1_squeezed_comb = p3_run__1[5:0];
  assign p4_Huffman_code_full_comb = p3_is_luminance ? literal_11603[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_11602[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_run_0_squeezed_const_msb_bits__3_comb = 3'h0;
  assign p4_huff_length_squeezed_comb = p3_and_11538 ? {p4_next_pix_squeezed_const_msb_bits_comb, p3_is_luminance ? 2'h2 : 2'h1, p4_next_pix__1_squeezed_squeezed_const_msb_bits__3_comb} : p4_Huffman_length_squeezed_comb;
  assign p4_next_pix_squeezed_const_msb_bits__1_comb = 2'h0;
  assign p4_next_pix_squeezed_comb = p3_and_11538 ? 6'h3f : p4_next_pix__1_squeezed_comb;
  assign p4_next_pix_squeezed_const_msb_bits__2_comb = 2'h0;
  assign p4_run_squeezed_comb = p3_and_11538 ? 6'h3f : p4_run__1_squeezed_comb;
  assign p4_huff_code_comb = p3_and_11538 ? {12'h000, {{1{p4_sel_11604_comb[2]}}, p4_sel_11604_comb}} : p4_Huffman_code_full_comb;
  assign p4_huff_length_comb = {p4_run_0_squeezed_const_msb_bits__3_comb, p4_huff_length_squeezed_comb};
  assign p4_code_size_comb = p4_concat_11591_comb & {8{~(p3_and_11538 | p3_eq_11117)}};
  assign p4_next_pix_comb = {p4_next_pix_squeezed_const_msb_bits__1_comb, p4_next_pix_squeezed_comb};
  assign p4_run_comb = {p4_next_pix_squeezed_const_msb_bits__2_comb, p4_run_squeezed_comb};
  assign p4_tuple_11637_comb = {p4_huff_code_comb, p4_huff_length_comb, p3_code_list, p4_code_size_comb, p4_next_pix_comb, p4_run_comb, p3_value};

  // Registers for pipe stage 4:
  reg [65:0] p4_tuple_11637;
  always @ (posedge clk) begin
    p4_tuple_11637 <= p4_tuple_11637_comb;
  end
  assign out = p4_tuple_11637;
endmodule
