module dct_2d_s12(
  input wire clk,
  input wire [767:0] x,
  output wire [767:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [20:0] smul21b_12b_x_9b (input reg [11:0] lhs, input reg [8:0] rhs);
    reg signed [11:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [20:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul21b_12b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [19:0] smul20b_20b_x_8b (input reg [19:0] lhs, input reg [7:0] rhs);
    reg signed [19:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [19:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul20b_20b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [19:0] smul20b_20b_x_6b (input reg [19:0] lhs, input reg [5:0] rhs);
    reg signed [19:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [19:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul20b_20b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [19:0] smul20b_20b_x_7b (input reg [19:0] lhs, input reg [6:0] rhs);
    reg signed [19:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [19:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul20b_20b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [18:0] smul19b_19b_x_7b (input reg [18:0] lhs, input reg [6:0] rhs);
    reg signed [18:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [18:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul19b_19b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [23:0] umul24b_24b_x_7b (input reg [23:0] lhs, input reg [6:0] rhs);
    begin
      umul24b_24b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [11:0] x_unflattened[0:7][0:7];
  assign x_unflattened[0][0] = x[11:0];
  assign x_unflattened[0][1] = x[23:12];
  assign x_unflattened[0][2] = x[35:24];
  assign x_unflattened[0][3] = x[47:36];
  assign x_unflattened[0][4] = x[59:48];
  assign x_unflattened[0][5] = x[71:60];
  assign x_unflattened[0][6] = x[83:72];
  assign x_unflattened[0][7] = x[95:84];
  assign x_unflattened[1][0] = x[107:96];
  assign x_unflattened[1][1] = x[119:108];
  assign x_unflattened[1][2] = x[131:120];
  assign x_unflattened[1][3] = x[143:132];
  assign x_unflattened[1][4] = x[155:144];
  assign x_unflattened[1][5] = x[167:156];
  assign x_unflattened[1][6] = x[179:168];
  assign x_unflattened[1][7] = x[191:180];
  assign x_unflattened[2][0] = x[203:192];
  assign x_unflattened[2][1] = x[215:204];
  assign x_unflattened[2][2] = x[227:216];
  assign x_unflattened[2][3] = x[239:228];
  assign x_unflattened[2][4] = x[251:240];
  assign x_unflattened[2][5] = x[263:252];
  assign x_unflattened[2][6] = x[275:264];
  assign x_unflattened[2][7] = x[287:276];
  assign x_unflattened[3][0] = x[299:288];
  assign x_unflattened[3][1] = x[311:300];
  assign x_unflattened[3][2] = x[323:312];
  assign x_unflattened[3][3] = x[335:324];
  assign x_unflattened[3][4] = x[347:336];
  assign x_unflattened[3][5] = x[359:348];
  assign x_unflattened[3][6] = x[371:360];
  assign x_unflattened[3][7] = x[383:372];
  assign x_unflattened[4][0] = x[395:384];
  assign x_unflattened[4][1] = x[407:396];
  assign x_unflattened[4][2] = x[419:408];
  assign x_unflattened[4][3] = x[431:420];
  assign x_unflattened[4][4] = x[443:432];
  assign x_unflattened[4][5] = x[455:444];
  assign x_unflattened[4][6] = x[467:456];
  assign x_unflattened[4][7] = x[479:468];
  assign x_unflattened[5][0] = x[491:480];
  assign x_unflattened[5][1] = x[503:492];
  assign x_unflattened[5][2] = x[515:504];
  assign x_unflattened[5][3] = x[527:516];
  assign x_unflattened[5][4] = x[539:528];
  assign x_unflattened[5][5] = x[551:540];
  assign x_unflattened[5][6] = x[563:552];
  assign x_unflattened[5][7] = x[575:564];
  assign x_unflattened[6][0] = x[587:576];
  assign x_unflattened[6][1] = x[599:588];
  assign x_unflattened[6][2] = x[611:600];
  assign x_unflattened[6][3] = x[623:612];
  assign x_unflattened[6][4] = x[635:624];
  assign x_unflattened[6][5] = x[647:636];
  assign x_unflattened[6][6] = x[659:648];
  assign x_unflattened[6][7] = x[671:660];
  assign x_unflattened[7][0] = x[683:672];
  assign x_unflattened[7][1] = x[695:684];
  assign x_unflattened[7][2] = x[707:696];
  assign x_unflattened[7][3] = x[719:708];
  assign x_unflattened[7][4] = x[731:720];
  assign x_unflattened[7][5] = x[743:732];
  assign x_unflattened[7][6] = x[755:744];
  assign x_unflattened[7][7] = x[767:756];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [11:0] p0_x[0:7][0:7];
  always @ (posedge clk) begin
    p0_x[0][0] <= x_unflattened[0][0];
    p0_x[0][1] <= x_unflattened[0][1];
    p0_x[0][2] <= x_unflattened[0][2];
    p0_x[0][3] <= x_unflattened[0][3];
    p0_x[0][4] <= x_unflattened[0][4];
    p0_x[0][5] <= x_unflattened[0][5];
    p0_x[0][6] <= x_unflattened[0][6];
    p0_x[0][7] <= x_unflattened[0][7];
    p0_x[1][0] <= x_unflattened[1][0];
    p0_x[1][1] <= x_unflattened[1][1];
    p0_x[1][2] <= x_unflattened[1][2];
    p0_x[1][3] <= x_unflattened[1][3];
    p0_x[1][4] <= x_unflattened[1][4];
    p0_x[1][5] <= x_unflattened[1][5];
    p0_x[1][6] <= x_unflattened[1][6];
    p0_x[1][7] <= x_unflattened[1][7];
    p0_x[2][0] <= x_unflattened[2][0];
    p0_x[2][1] <= x_unflattened[2][1];
    p0_x[2][2] <= x_unflattened[2][2];
    p0_x[2][3] <= x_unflattened[2][3];
    p0_x[2][4] <= x_unflattened[2][4];
    p0_x[2][5] <= x_unflattened[2][5];
    p0_x[2][6] <= x_unflattened[2][6];
    p0_x[2][7] <= x_unflattened[2][7];
    p0_x[3][0] <= x_unflattened[3][0];
    p0_x[3][1] <= x_unflattened[3][1];
    p0_x[3][2] <= x_unflattened[3][2];
    p0_x[3][3] <= x_unflattened[3][3];
    p0_x[3][4] <= x_unflattened[3][4];
    p0_x[3][5] <= x_unflattened[3][5];
    p0_x[3][6] <= x_unflattened[3][6];
    p0_x[3][7] <= x_unflattened[3][7];
    p0_x[4][0] <= x_unflattened[4][0];
    p0_x[4][1] <= x_unflattened[4][1];
    p0_x[4][2] <= x_unflattened[4][2];
    p0_x[4][3] <= x_unflattened[4][3];
    p0_x[4][4] <= x_unflattened[4][4];
    p0_x[4][5] <= x_unflattened[4][5];
    p0_x[4][6] <= x_unflattened[4][6];
    p0_x[4][7] <= x_unflattened[4][7];
    p0_x[5][0] <= x_unflattened[5][0];
    p0_x[5][1] <= x_unflattened[5][1];
    p0_x[5][2] <= x_unflattened[5][2];
    p0_x[5][3] <= x_unflattened[5][3];
    p0_x[5][4] <= x_unflattened[5][4];
    p0_x[5][5] <= x_unflattened[5][5];
    p0_x[5][6] <= x_unflattened[5][6];
    p0_x[5][7] <= x_unflattened[5][7];
    p0_x[6][0] <= x_unflattened[6][0];
    p0_x[6][1] <= x_unflattened[6][1];
    p0_x[6][2] <= x_unflattened[6][2];
    p0_x[6][3] <= x_unflattened[6][3];
    p0_x[6][4] <= x_unflattened[6][4];
    p0_x[6][5] <= x_unflattened[6][5];
    p0_x[6][6] <= x_unflattened[6][6];
    p0_x[6][7] <= x_unflattened[6][7];
    p0_x[7][0] <= x_unflattened[7][0];
    p0_x[7][1] <= x_unflattened[7][1];
    p0_x[7][2] <= x_unflattened[7][2];
    p0_x[7][3] <= x_unflattened[7][3];
    p0_x[7][4] <= x_unflattened[7][4];
    p0_x[7][5] <= x_unflattened[7][5];
    p0_x[7][6] <= x_unflattened[7][6];
    p0_x[7][7] <= x_unflattened[7][7];
  end

  // ===== Pipe stage 1:
  wire [11:0] p1_array_index_75184_comb;
  wire [11:0] p1_array_index_75185_comb;
  wire [11:0] p1_array_index_75186_comb;
  wire [11:0] p1_array_index_75187_comb;
  wire [11:0] p1_array_index_75188_comb;
  wire [11:0] p1_array_index_75189_comb;
  wire [11:0] p1_array_index_75190_comb;
  wire [11:0] p1_array_index_75191_comb;
  wire [11:0] p1_array_index_75192_comb;
  wire [11:0] p1_array_index_75193_comb;
  wire [11:0] p1_array_index_75194_comb;
  wire [11:0] p1_array_index_75195_comb;
  wire [11:0] p1_array_index_75196_comb;
  wire [11:0] p1_array_index_75197_comb;
  wire [11:0] p1_array_index_75198_comb;
  wire [11:0] p1_array_index_75199_comb;
  wire [11:0] p1_array_index_75200_comb;
  wire [11:0] p1_array_index_75201_comb;
  wire [11:0] p1_array_index_75202_comb;
  wire [11:0] p1_array_index_75203_comb;
  wire [11:0] p1_array_index_75204_comb;
  wire [11:0] p1_array_index_75205_comb;
  wire [11:0] p1_array_index_75206_comb;
  wire [11:0] p1_array_index_75207_comb;
  wire [11:0] p1_array_index_75208_comb;
  wire [11:0] p1_array_index_75209_comb;
  wire [11:0] p1_array_index_75210_comb;
  wire [11:0] p1_array_index_75211_comb;
  wire [11:0] p1_array_index_75212_comb;
  wire [11:0] p1_array_index_75213_comb;
  wire [11:0] p1_array_index_75214_comb;
  wire [11:0] p1_array_index_75215_comb;
  wire [11:0] p1_array_index_75216_comb;
  wire [11:0] p1_array_index_75217_comb;
  wire [11:0] p1_array_index_75218_comb;
  wire [11:0] p1_array_index_75219_comb;
  wire [11:0] p1_array_index_75220_comb;
  wire [11:0] p1_array_index_75221_comb;
  wire [11:0] p1_array_index_75222_comb;
  wire [11:0] p1_array_index_75223_comb;
  wire [11:0] p1_array_index_75224_comb;
  wire [11:0] p1_array_index_75225_comb;
  wire [11:0] p1_array_index_75226_comb;
  wire [11:0] p1_array_index_75227_comb;
  wire [11:0] p1_array_index_75228_comb;
  wire [11:0] p1_array_index_75229_comb;
  wire [11:0] p1_array_index_75230_comb;
  wire [11:0] p1_array_index_75231_comb;
  wire [11:0] p1_array_index_75232_comb;
  wire [11:0] p1_array_index_75233_comb;
  wire [11:0] p1_array_index_75234_comb;
  wire [11:0] p1_array_index_75235_comb;
  wire [11:0] p1_array_index_75236_comb;
  wire [11:0] p1_array_index_75237_comb;
  wire [11:0] p1_array_index_75238_comb;
  wire [11:0] p1_array_index_75239_comb;
  wire [11:0] p1_array_index_75240_comb;
  wire [11:0] p1_array_index_75241_comb;
  wire [11:0] p1_array_index_75242_comb;
  wire [11:0] p1_array_index_75243_comb;
  wire [11:0] p1_array_index_75244_comb;
  wire [11:0] p1_array_index_75245_comb;
  wire [11:0] p1_array_index_75246_comb;
  wire [11:0] p1_array_index_75247_comb;
  wire [23:0] p1_sign_ext_75250_comb;
  wire [23:0] p1_sign_ext_75251_comb;
  wire [23:0] p1_sign_ext_75252_comb;
  wire [23:0] p1_sign_ext_75253_comb;
  wire [23:0] p1_sign_ext_75258_comb;
  wire [23:0] p1_sign_ext_75259_comb;
  wire [23:0] p1_sign_ext_75260_comb;
  wire [23:0] p1_sign_ext_75261_comb;
  wire [23:0] p1_sign_ext_75266_comb;
  wire [23:0] p1_sign_ext_75267_comb;
  wire [23:0] p1_sign_ext_75268_comb;
  wire [23:0] p1_sign_ext_75269_comb;
  wire [23:0] p1_sign_ext_75274_comb;
  wire [23:0] p1_sign_ext_75275_comb;
  wire [23:0] p1_sign_ext_75276_comb;
  wire [23:0] p1_sign_ext_75277_comb;
  wire [23:0] p1_sign_ext_75280_comb;
  wire [23:0] p1_sign_ext_75281_comb;
  wire [23:0] p1_sign_ext_75282_comb;
  wire [23:0] p1_sign_ext_75283_comb;
  wire [23:0] p1_sign_ext_75284_comb;
  wire [23:0] p1_sign_ext_75285_comb;
  wire [23:0] p1_sign_ext_75286_comb;
  wire [23:0] p1_sign_ext_75287_comb;
  wire [23:0] p1_sign_ext_75304_comb;
  wire [23:0] p1_sign_ext_75309_comb;
  wire [23:0] p1_sign_ext_75310_comb;
  wire [23:0] p1_sign_ext_75315_comb;
  wire [23:0] p1_sign_ext_75316_comb;
  wire [23:0] p1_sign_ext_75321_comb;
  wire [23:0] p1_sign_ext_75322_comb;
  wire [23:0] p1_sign_ext_75327_comb;
  wire [23:0] p1_sign_ext_75346_comb;
  wire [23:0] p1_sign_ext_75347_comb;
  wire [23:0] p1_sign_ext_75348_comb;
  wire [23:0] p1_sign_ext_75349_comb;
  wire [23:0] p1_sign_ext_75354_comb;
  wire [23:0] p1_sign_ext_75355_comb;
  wire [23:0] p1_sign_ext_75356_comb;
  wire [23:0] p1_sign_ext_75357_comb;
  wire [23:0] p1_sign_ext_75360_comb;
  wire [23:0] p1_sign_ext_75361_comb;
  wire [23:0] p1_sign_ext_75362_comb;
  wire [23:0] p1_sign_ext_75363_comb;
  wire [23:0] p1_sign_ext_75372_comb;
  wire [23:0] p1_sign_ext_75377_comb;
  wire [23:0] p1_sign_ext_75378_comb;
  wire [23:0] p1_sign_ext_75383_comb;
  wire [23:0] p1_sign_ext_75394_comb;
  wire [23:0] p1_sign_ext_75395_comb;
  wire [23:0] p1_sign_ext_75396_comb;
  wire [23:0] p1_sign_ext_75397_comb;
  wire [23:0] p1_sign_ext_75402_comb;
  wire [23:0] p1_sign_ext_75403_comb;
  wire [23:0] p1_sign_ext_75404_comb;
  wire [23:0] p1_sign_ext_75405_comb;
  wire [23:0] p1_sign_ext_75408_comb;
  wire [23:0] p1_sign_ext_75409_comb;
  wire [23:0] p1_sign_ext_75410_comb;
  wire [23:0] p1_sign_ext_75411_comb;
  wire [23:0] p1_sign_ext_75420_comb;
  wire [23:0] p1_sign_ext_75425_comb;
  wire [23:0] p1_sign_ext_75426_comb;
  wire [23:0] p1_sign_ext_75431_comb;
  wire [20:0] p1_smul_75440_comb;
  wire [20:0] p1_smul_75441_comb;
  wire [20:0] p1_smul_75450_comb;
  wire [20:0] p1_smul_75451_comb;
  wire [20:0] p1_smul_75452_comb;
  wire [20:0] p1_smul_75453_comb;
  wire [20:0] p1_smul_75462_comb;
  wire [20:0] p1_smul_75463_comb;
  wire [20:0] p1_smul_75464_comb;
  wire [20:0] p1_smul_75465_comb;
  wire [20:0] p1_smul_75474_comb;
  wire [20:0] p1_smul_75475_comb;
  wire [20:0] p1_smul_75476_comb;
  wire [20:0] p1_smul_75477_comb;
  wire [20:0] p1_smul_75486_comb;
  wire [20:0] p1_smul_75487_comb;
  wire [20:0] p1_smul_75512_comb;
  wire [20:0] p1_smul_75514_comb;
  wire [20:0] p1_smul_75517_comb;
  wire [20:0] p1_smul_75519_comb;
  wire [20:0] p1_smul_75520_comb;
  wire [20:0] p1_smul_75522_comb;
  wire [20:0] p1_smul_75525_comb;
  wire [20:0] p1_smul_75527_comb;
  wire [20:0] p1_smul_75528_comb;
  wire [20:0] p1_smul_75530_comb;
  wire [20:0] p1_smul_75533_comb;
  wire [20:0] p1_smul_75535_comb;
  wire [20:0] p1_smul_75536_comb;
  wire [20:0] p1_smul_75538_comb;
  wire [20:0] p1_smul_75541_comb;
  wire [20:0] p1_smul_75543_comb;
  wire [20:0] p1_smul_75546_comb;
  wire [20:0] p1_smul_75548_comb;
  wire [20:0] p1_smul_75549_comb;
  wire [20:0] p1_smul_75551_comb;
  wire [20:0] p1_smul_75556_comb;
  wire [20:0] p1_smul_75558_comb;
  wire [20:0] p1_smul_75559_comb;
  wire [20:0] p1_smul_75561_comb;
  wire [20:0] p1_smul_75566_comb;
  wire [20:0] p1_smul_75568_comb;
  wire [20:0] p1_smul_75569_comb;
  wire [20:0] p1_smul_75571_comb;
  wire [20:0] p1_smul_75576_comb;
  wire [20:0] p1_smul_75578_comb;
  wire [20:0] p1_smul_75579_comb;
  wire [20:0] p1_smul_75581_comb;
  wire [20:0] p1_smul_75602_comb;
  wire [20:0] p1_smul_75603_comb;
  wire [20:0] p1_smul_75604_comb;
  wire [20:0] p1_smul_75605_comb;
  wire [20:0] p1_smul_75610_comb;
  wire [20:0] p1_smul_75611_comb;
  wire [20:0] p1_smul_75612_comb;
  wire [20:0] p1_smul_75613_comb;
  wire [20:0] p1_smul_75618_comb;
  wire [20:0] p1_smul_75619_comb;
  wire [20:0] p1_smul_75620_comb;
  wire [20:0] p1_smul_75621_comb;
  wire [20:0] p1_smul_75626_comb;
  wire [20:0] p1_smul_75627_comb;
  wire [20:0] p1_smul_75628_comb;
  wire [20:0] p1_smul_75629_comb;
  wire [20:0] p1_smul_75632_comb;
  wire [20:0] p1_smul_75633_comb;
  wire [20:0] p1_smul_75642_comb;
  wire [20:0] p1_smul_75643_comb;
  wire [20:0] p1_smul_75644_comb;
  wire [20:0] p1_smul_75645_comb;
  wire [20:0] p1_smul_75654_comb;
  wire [20:0] p1_smul_75655_comb;
  wire [20:0] p1_smul_75668_comb;
  wire [20:0] p1_smul_75670_comb;
  wire [20:0] p1_smul_75673_comb;
  wire [20:0] p1_smul_75675_comb;
  wire [20:0] p1_smul_75676_comb;
  wire [20:0] p1_smul_75678_comb;
  wire [20:0] p1_smul_75681_comb;
  wire [20:0] p1_smul_75683_comb;
  wire [20:0] p1_smul_75686_comb;
  wire [20:0] p1_smul_75688_comb;
  wire [20:0] p1_smul_75689_comb;
  wire [20:0] p1_smul_75691_comb;
  wire [20:0] p1_smul_75696_comb;
  wire [20:0] p1_smul_75698_comb;
  wire [20:0] p1_smul_75699_comb;
  wire [20:0] p1_smul_75701_comb;
  wire [20:0] p1_smul_75714_comb;
  wire [20:0] p1_smul_75715_comb;
  wire [20:0] p1_smul_75716_comb;
  wire [20:0] p1_smul_75717_comb;
  wire [20:0] p1_smul_75722_comb;
  wire [20:0] p1_smul_75723_comb;
  wire [20:0] p1_smul_75724_comb;
  wire [20:0] p1_smul_75725_comb;
  wire [20:0] p1_smul_75728_comb;
  wire [20:0] p1_smul_75729_comb;
  wire [20:0] p1_smul_75738_comb;
  wire [20:0] p1_smul_75739_comb;
  wire [20:0] p1_smul_75740_comb;
  wire [20:0] p1_smul_75741_comb;
  wire [20:0] p1_smul_75750_comb;
  wire [20:0] p1_smul_75751_comb;
  wire [20:0] p1_smul_75764_comb;
  wire [20:0] p1_smul_75766_comb;
  wire [20:0] p1_smul_75769_comb;
  wire [20:0] p1_smul_75771_comb;
  wire [20:0] p1_smul_75772_comb;
  wire [20:0] p1_smul_75774_comb;
  wire [20:0] p1_smul_75777_comb;
  wire [20:0] p1_smul_75779_comb;
  wire [20:0] p1_smul_75782_comb;
  wire [20:0] p1_smul_75784_comb;
  wire [20:0] p1_smul_75785_comb;
  wire [20:0] p1_smul_75787_comb;
  wire [20:0] p1_smul_75792_comb;
  wire [20:0] p1_smul_75794_comb;
  wire [20:0] p1_smul_75795_comb;
  wire [20:0] p1_smul_75797_comb;
  wire [20:0] p1_smul_75810_comb;
  wire [20:0] p1_smul_75811_comb;
  wire [20:0] p1_smul_75812_comb;
  wire [20:0] p1_smul_75813_comb;
  wire [20:0] p1_smul_75818_comb;
  wire [20:0] p1_smul_75819_comb;
  wire [20:0] p1_smul_75820_comb;
  wire [20:0] p1_smul_75821_comb;
  wire [20:0] p1_add_75824_comb;
  wire [19:0] p1_smul_75825_comb;
  wire [19:0] p1_smul_75826_comb;
  wire [19:0] p1_smul_75827_comb;
  wire [19:0] p1_smul_75828_comb;
  wire [20:0] p1_add_75829_comb;
  wire [20:0] p1_add_75830_comb;
  wire [19:0] p1_smul_75831_comb;
  wire [19:0] p1_smul_75832_comb;
  wire [19:0] p1_smul_75833_comb;
  wire [19:0] p1_smul_75834_comb;
  wire [20:0] p1_add_75835_comb;
  wire [20:0] p1_add_75836_comb;
  wire [19:0] p1_smul_75837_comb;
  wire [19:0] p1_smul_75838_comb;
  wire [19:0] p1_smul_75839_comb;
  wire [19:0] p1_smul_75840_comb;
  wire [20:0] p1_add_75841_comb;
  wire [20:0] p1_add_75842_comb;
  wire [19:0] p1_smul_75843_comb;
  wire [19:0] p1_smul_75844_comb;
  wire [19:0] p1_smul_75845_comb;
  wire [19:0] p1_smul_75846_comb;
  wire [20:0] p1_add_75847_comb;
  wire [19:0] p1_smul_75850_comb;
  wire [19:0] p1_smul_75851_comb;
  wire [19:0] p1_smul_75856_comb;
  wire [19:0] p1_smul_75857_comb;
  wire [19:0] p1_smul_75862_comb;
  wire [19:0] p1_smul_75863_comb;
  wire [19:0] p1_smul_75868_comb;
  wire [19:0] p1_smul_75869_comb;
  wire [19:0] p1_smul_75874_comb;
  wire [19:0] p1_smul_75875_comb;
  wire [19:0] p1_smul_75880_comb;
  wire [19:0] p1_smul_75881_comb;
  wire [19:0] p1_smul_75886_comb;
  wire [19:0] p1_smul_75887_comb;
  wire [19:0] p1_smul_75892_comb;
  wire [19:0] p1_smul_75893_comb;
  wire [19:0] p1_smul_75897_comb;
  wire [19:0] p1_smul_75899_comb;
  wire [19:0] p1_smul_75900_comb;
  wire [19:0] p1_smul_75902_comb;
  wire [19:0] p1_smul_75905_comb;
  wire [19:0] p1_smul_75907_comb;
  wire [19:0] p1_smul_75908_comb;
  wire [19:0] p1_smul_75910_comb;
  wire [19:0] p1_smul_75913_comb;
  wire [19:0] p1_smul_75915_comb;
  wire [19:0] p1_smul_75916_comb;
  wire [19:0] p1_smul_75918_comb;
  wire [19:0] p1_smul_75921_comb;
  wire [19:0] p1_smul_75923_comb;
  wire [19:0] p1_smul_75924_comb;
  wire [19:0] p1_smul_75926_comb;
  wire [19:0] p1_smul_75960_comb;
  wire [19:0] p1_smul_75962_comb;
  wire [19:0] p1_smul_75965_comb;
  wire [19:0] p1_smul_75967_comb;
  wire [19:0] p1_smul_75968_comb;
  wire [19:0] p1_smul_75970_comb;
  wire [19:0] p1_smul_75973_comb;
  wire [19:0] p1_smul_75975_comb;
  wire [19:0] p1_smul_75976_comb;
  wire [19:0] p1_smul_75978_comb;
  wire [19:0] p1_smul_75981_comb;
  wire [19:0] p1_smul_75983_comb;
  wire [19:0] p1_smul_75984_comb;
  wire [19:0] p1_smul_75986_comb;
  wire [19:0] p1_smul_75989_comb;
  wire [19:0] p1_smul_75991_comb;
  wire [19:0] p1_smul_75992_comb;
  wire [19:0] p1_smul_75995_comb;
  wire [19:0] p1_smul_75998_comb;
  wire [19:0] p1_smul_76001_comb;
  wire [19:0] p1_smul_76002_comb;
  wire [19:0] p1_smul_76005_comb;
  wire [19:0] p1_smul_76008_comb;
  wire [19:0] p1_smul_76011_comb;
  wire [19:0] p1_smul_76012_comb;
  wire [19:0] p1_smul_76015_comb;
  wire [19:0] p1_smul_76018_comb;
  wire [19:0] p1_smul_76021_comb;
  wire [19:0] p1_smul_76022_comb;
  wire [19:0] p1_smul_76025_comb;
  wire [19:0] p1_smul_76028_comb;
  wire [19:0] p1_smul_76031_comb;
  wire [19:0] p1_smul_76032_comb;
  wire [19:0] p1_smul_76033_comb;
  wire [20:0] p1_add_76034_comb;
  wire [20:0] p1_add_76035_comb;
  wire [19:0] p1_smul_76036_comb;
  wire [19:0] p1_smul_76037_comb;
  wire [19:0] p1_smul_76038_comb;
  wire [19:0] p1_smul_76039_comb;
  wire [20:0] p1_add_76040_comb;
  wire [20:0] p1_add_76041_comb;
  wire [19:0] p1_smul_76042_comb;
  wire [19:0] p1_smul_76043_comb;
  wire [19:0] p1_smul_76044_comb;
  wire [19:0] p1_smul_76045_comb;
  wire [20:0] p1_add_76046_comb;
  wire [20:0] p1_add_76047_comb;
  wire [19:0] p1_smul_76048_comb;
  wire [19:0] p1_smul_76049_comb;
  wire [19:0] p1_smul_76050_comb;
  wire [19:0] p1_smul_76051_comb;
  wire [20:0] p1_add_76052_comb;
  wire [20:0] p1_add_76053_comb;
  wire [19:0] p1_smul_76054_comb;
  wire [19:0] p1_smul_76055_comb;
  wire [20:0] p1_add_76056_comb;
  wire [19:0] p1_smul_76057_comb;
  wire [19:0] p1_smul_76058_comb;
  wire [19:0] p1_smul_76059_comb;
  wire [19:0] p1_smul_76060_comb;
  wire [20:0] p1_add_76061_comb;
  wire [20:0] p1_add_76062_comb;
  wire [19:0] p1_smul_76063_comb;
  wire [19:0] p1_smul_76064_comb;
  wire [19:0] p1_smul_76065_comb;
  wire [19:0] p1_smul_76066_comb;
  wire [20:0] p1_add_76067_comb;
  wire [19:0] p1_smul_76070_comb;
  wire [19:0] p1_smul_76071_comb;
  wire [19:0] p1_smul_76076_comb;
  wire [19:0] p1_smul_76077_comb;
  wire [19:0] p1_smul_76082_comb;
  wire [19:0] p1_smul_76083_comb;
  wire [19:0] p1_smul_76088_comb;
  wire [19:0] p1_smul_76089_comb;
  wire [19:0] p1_smul_76093_comb;
  wire [19:0] p1_smul_76095_comb;
  wire [19:0] p1_smul_76096_comb;
  wire [19:0] p1_smul_76098_comb;
  wire [19:0] p1_smul_76101_comb;
  wire [19:0] p1_smul_76103_comb;
  wire [19:0] p1_smul_76104_comb;
  wire [19:0] p1_smul_76106_comb;
  wire [19:0] p1_smul_76124_comb;
  wire [19:0] p1_smul_76126_comb;
  wire [19:0] p1_smul_76129_comb;
  wire [19:0] p1_smul_76131_comb;
  wire [19:0] p1_smul_76132_comb;
  wire [19:0] p1_smul_76134_comb;
  wire [19:0] p1_smul_76137_comb;
  wire [19:0] p1_smul_76139_comb;
  wire [19:0] p1_smul_76140_comb;
  wire [19:0] p1_smul_76143_comb;
  wire [19:0] p1_smul_76146_comb;
  wire [19:0] p1_smul_76149_comb;
  wire [19:0] p1_smul_76150_comb;
  wire [19:0] p1_smul_76153_comb;
  wire [19:0] p1_smul_76156_comb;
  wire [19:0] p1_smul_76159_comb;
  wire [19:0] p1_smul_76160_comb;
  wire [19:0] p1_smul_76161_comb;
  wire [20:0] p1_add_76162_comb;
  wire [20:0] p1_add_76163_comb;
  wire [19:0] p1_smul_76164_comb;
  wire [19:0] p1_smul_76165_comb;
  wire [19:0] p1_smul_76166_comb;
  wire [19:0] p1_smul_76167_comb;
  wire [20:0] p1_add_76168_comb;
  wire [20:0] p1_add_76169_comb;
  wire [19:0] p1_smul_76170_comb;
  wire [19:0] p1_smul_76171_comb;
  wire [20:0] p1_add_76172_comb;
  wire [19:0] p1_smul_76173_comb;
  wire [19:0] p1_smul_76174_comb;
  wire [19:0] p1_smul_76175_comb;
  wire [19:0] p1_smul_76176_comb;
  wire [20:0] p1_add_76177_comb;
  wire [20:0] p1_add_76178_comb;
  wire [19:0] p1_smul_76179_comb;
  wire [19:0] p1_smul_76180_comb;
  wire [19:0] p1_smul_76181_comb;
  wire [19:0] p1_smul_76182_comb;
  wire [20:0] p1_add_76183_comb;
  wire [19:0] p1_smul_76186_comb;
  wire [19:0] p1_smul_76187_comb;
  wire [19:0] p1_smul_76192_comb;
  wire [19:0] p1_smul_76193_comb;
  wire [19:0] p1_smul_76198_comb;
  wire [19:0] p1_smul_76199_comb;
  wire [19:0] p1_smul_76204_comb;
  wire [19:0] p1_smul_76205_comb;
  wire [19:0] p1_smul_76209_comb;
  wire [19:0] p1_smul_76211_comb;
  wire [19:0] p1_smul_76212_comb;
  wire [19:0] p1_smul_76214_comb;
  wire [19:0] p1_smul_76217_comb;
  wire [19:0] p1_smul_76219_comb;
  wire [19:0] p1_smul_76220_comb;
  wire [19:0] p1_smul_76222_comb;
  wire [19:0] p1_smul_76240_comb;
  wire [19:0] p1_smul_76242_comb;
  wire [19:0] p1_smul_76245_comb;
  wire [19:0] p1_smul_76247_comb;
  wire [19:0] p1_smul_76248_comb;
  wire [19:0] p1_smul_76250_comb;
  wire [19:0] p1_smul_76253_comb;
  wire [19:0] p1_smul_76255_comb;
  wire [19:0] p1_smul_76256_comb;
  wire [19:0] p1_smul_76259_comb;
  wire [19:0] p1_smul_76262_comb;
  wire [19:0] p1_smul_76265_comb;
  wire [19:0] p1_smul_76266_comb;
  wire [19:0] p1_smul_76269_comb;
  wire [19:0] p1_smul_76272_comb;
  wire [19:0] p1_smul_76275_comb;
  wire [19:0] p1_smul_76276_comb;
  wire [19:0] p1_smul_76277_comb;
  wire [20:0] p1_add_76278_comb;
  wire [20:0] p1_add_76279_comb;
  wire [19:0] p1_smul_76280_comb;
  wire [19:0] p1_smul_76281_comb;
  wire [19:0] p1_smul_76282_comb;
  wire [19:0] p1_smul_76283_comb;
  wire [20:0] p1_add_76284_comb;
  wire [20:0] p1_add_76285_comb;
  wire [19:0] p1_smul_76286_comb;
  wire [19:0] p1_smul_76287_comb;
  wire [19:0] p1_bit_slice_76320_comb;
  wire [19:0] p1_add_76321_comb;
  wire [19:0] p1_add_76322_comb;
  wire [19:0] p1_bit_slice_76323_comb;
  wire [19:0] p1_bit_slice_76324_comb;
  wire [19:0] p1_add_76325_comb;
  wire [19:0] p1_add_76326_comb;
  wire [19:0] p1_bit_slice_76327_comb;
  wire [19:0] p1_bit_slice_76328_comb;
  wire [19:0] p1_add_76329_comb;
  wire [19:0] p1_add_76330_comb;
  wire [19:0] p1_bit_slice_76331_comb;
  wire [19:0] p1_bit_slice_76332_comb;
  wire [19:0] p1_add_76333_comb;
  wire [19:0] p1_add_76334_comb;
  wire [19:0] p1_bit_slice_76335_comb;
  wire [18:0] p1_smul_76336_comb;
  wire [18:0] p1_smul_76339_comb;
  wire [18:0] p1_smul_76340_comb;
  wire [18:0] p1_smul_76343_comb;
  wire [18:0] p1_smul_76344_comb;
  wire [18:0] p1_smul_76347_comb;
  wire [18:0] p1_smul_76348_comb;
  wire [18:0] p1_smul_76351_comb;
  wire [18:0] p1_smul_76352_comb;
  wire [18:0] p1_smul_76355_comb;
  wire [18:0] p1_smul_76356_comb;
  wire [18:0] p1_smul_76359_comb;
  wire [18:0] p1_smul_76360_comb;
  wire [18:0] p1_smul_76363_comb;
  wire [18:0] p1_smul_76364_comb;
  wire [18:0] p1_smul_76367_comb;
  wire [19:0] p1_add_76368_comb;
  wire [19:0] p1_add_76370_comb;
  wire [19:0] p1_add_76372_comb;
  wire [19:0] p1_add_76374_comb;
  wire [19:0] p1_add_76376_comb;
  wire [19:0] p1_add_76378_comb;
  wire [19:0] p1_add_76380_comb;
  wire [19:0] p1_add_76382_comb;
  wire [19:0] p1_add_76384_comb;
  wire [19:0] p1_add_76386_comb;
  wire [19:0] p1_add_76388_comb;
  wire [19:0] p1_add_76390_comb;
  wire [19:0] p1_add_76392_comb;
  wire [19:0] p1_add_76394_comb;
  wire [19:0] p1_add_76396_comb;
  wire [19:0] p1_add_76398_comb;
  wire [20:0] p1_smul_76400_comb;
  wire [20:0] p1_smul_76401_comb;
  wire [20:0] p1_smul_76402_comb;
  wire [20:0] p1_smul_76403_comb;
  wire [20:0] p1_smul_76404_comb;
  wire [20:0] p1_smul_76405_comb;
  wire [20:0] p1_smul_76406_comb;
  wire [20:0] p1_smul_76407_comb;
  wire [20:0] p1_smul_76408_comb;
  wire [20:0] p1_smul_76409_comb;
  wire [20:0] p1_smul_76410_comb;
  wire [20:0] p1_smul_76411_comb;
  wire [20:0] p1_smul_76412_comb;
  wire [20:0] p1_smul_76413_comb;
  wire [20:0] p1_smul_76414_comb;
  wire [20:0] p1_smul_76415_comb;
  wire [20:0] p1_smul_76416_comb;
  wire [20:0] p1_smul_76417_comb;
  wire [20:0] p1_smul_76418_comb;
  wire [20:0] p1_smul_76419_comb;
  wire [20:0] p1_smul_76420_comb;
  wire [20:0] p1_smul_76421_comb;
  wire [20:0] p1_smul_76422_comb;
  wire [20:0] p1_smul_76423_comb;
  wire [20:0] p1_smul_76424_comb;
  wire [20:0] p1_smul_76425_comb;
  wire [20:0] p1_smul_76426_comb;
  wire [20:0] p1_smul_76427_comb;
  wire [20:0] p1_smul_76428_comb;
  wire [20:0] p1_smul_76429_comb;
  wire [20:0] p1_smul_76430_comb;
  wire [20:0] p1_smul_76431_comb;
  wire [19:0] p1_add_76432_comb;
  wire [19:0] p1_add_76434_comb;
  wire [19:0] p1_add_76436_comb;
  wire [19:0] p1_add_76438_comb;
  wire [19:0] p1_add_76440_comb;
  wire [19:0] p1_add_76442_comb;
  wire [19:0] p1_add_76444_comb;
  wire [19:0] p1_add_76446_comb;
  wire [19:0] p1_add_76448_comb;
  wire [19:0] p1_add_76450_comb;
  wire [19:0] p1_add_76452_comb;
  wire [19:0] p1_add_76454_comb;
  wire [19:0] p1_add_76456_comb;
  wire [19:0] p1_add_76458_comb;
  wire [19:0] p1_add_76460_comb;
  wire [19:0] p1_add_76462_comb;
  wire [18:0] p1_smul_76465_comb;
  wire [18:0] p1_smul_76467_comb;
  wire [18:0] p1_smul_76468_comb;
  wire [18:0] p1_smul_76470_comb;
  wire [18:0] p1_smul_76473_comb;
  wire [18:0] p1_smul_76475_comb;
  wire [18:0] p1_smul_76476_comb;
  wire [18:0] p1_smul_76478_comb;
  wire [18:0] p1_smul_76481_comb;
  wire [18:0] p1_smul_76483_comb;
  wire [18:0] p1_smul_76484_comb;
  wire [18:0] p1_smul_76486_comb;
  wire [18:0] p1_smul_76489_comb;
  wire [18:0] p1_smul_76491_comb;
  wire [18:0] p1_smul_76492_comb;
  wire [18:0] p1_smul_76494_comb;
  wire [19:0] p1_add_76496_comb;
  wire [19:0] p1_bit_slice_76497_comb;
  wire [19:0] p1_bit_slice_76498_comb;
  wire [19:0] p1_add_76499_comb;
  wire [19:0] p1_add_76500_comb;
  wire [19:0] p1_bit_slice_76501_comb;
  wire [19:0] p1_bit_slice_76502_comb;
  wire [19:0] p1_add_76503_comb;
  wire [19:0] p1_add_76504_comb;
  wire [19:0] p1_bit_slice_76505_comb;
  wire [19:0] p1_bit_slice_76506_comb;
  wire [19:0] p1_add_76507_comb;
  wire [19:0] p1_add_76508_comb;
  wire [19:0] p1_bit_slice_76509_comb;
  wire [19:0] p1_bit_slice_76510_comb;
  wire [19:0] p1_add_76511_comb;
  wire [19:0] p1_bit_slice_76528_comb;
  wire [19:0] p1_add_76529_comb;
  wire [19:0] p1_add_76530_comb;
  wire [19:0] p1_bit_slice_76531_comb;
  wire [19:0] p1_bit_slice_76532_comb;
  wire [19:0] p1_add_76533_comb;
  wire [19:0] p1_add_76534_comb;
  wire [19:0] p1_bit_slice_76535_comb;
  wire [18:0] p1_smul_76536_comb;
  wire [18:0] p1_smul_76539_comb;
  wire [18:0] p1_smul_76540_comb;
  wire [18:0] p1_smul_76543_comb;
  wire [18:0] p1_smul_76544_comb;
  wire [18:0] p1_smul_76547_comb;
  wire [18:0] p1_smul_76548_comb;
  wire [18:0] p1_smul_76551_comb;
  wire [19:0] p1_add_76552_comb;
  wire [19:0] p1_add_76554_comb;
  wire [19:0] p1_add_76556_comb;
  wire [19:0] p1_add_76558_comb;
  wire [19:0] p1_add_76560_comb;
  wire [19:0] p1_add_76562_comb;
  wire [19:0] p1_add_76564_comb;
  wire [19:0] p1_add_76566_comb;
  wire [20:0] p1_smul_76568_comb;
  wire [20:0] p1_smul_76569_comb;
  wire [20:0] p1_smul_76570_comb;
  wire [20:0] p1_smul_76571_comb;
  wire [20:0] p1_smul_76572_comb;
  wire [20:0] p1_smul_76573_comb;
  wire [20:0] p1_smul_76574_comb;
  wire [20:0] p1_smul_76575_comb;
  wire [20:0] p1_smul_76576_comb;
  wire [20:0] p1_smul_76577_comb;
  wire [20:0] p1_smul_76578_comb;
  wire [20:0] p1_smul_76579_comb;
  wire [20:0] p1_smul_76580_comb;
  wire [20:0] p1_smul_76581_comb;
  wire [20:0] p1_smul_76582_comb;
  wire [20:0] p1_smul_76583_comb;
  wire [19:0] p1_add_76584_comb;
  wire [19:0] p1_add_76586_comb;
  wire [19:0] p1_add_76588_comb;
  wire [19:0] p1_add_76590_comb;
  wire [19:0] p1_add_76592_comb;
  wire [19:0] p1_add_76594_comb;
  wire [19:0] p1_add_76596_comb;
  wire [19:0] p1_add_76598_comb;
  wire [18:0] p1_smul_76601_comb;
  wire [18:0] p1_smul_76603_comb;
  wire [18:0] p1_smul_76604_comb;
  wire [18:0] p1_smul_76606_comb;
  wire [18:0] p1_smul_76609_comb;
  wire [18:0] p1_smul_76611_comb;
  wire [18:0] p1_smul_76612_comb;
  wire [18:0] p1_smul_76614_comb;
  wire [19:0] p1_add_76616_comb;
  wire [19:0] p1_bit_slice_76617_comb;
  wire [19:0] p1_bit_slice_76618_comb;
  wire [19:0] p1_add_76619_comb;
  wire [19:0] p1_add_76620_comb;
  wire [19:0] p1_bit_slice_76621_comb;
  wire [19:0] p1_bit_slice_76622_comb;
  wire [19:0] p1_add_76623_comb;
  wire [19:0] p1_bit_slice_76640_comb;
  wire [19:0] p1_add_76641_comb;
  wire [19:0] p1_add_76642_comb;
  wire [19:0] p1_bit_slice_76643_comb;
  wire [19:0] p1_bit_slice_76644_comb;
  wire [19:0] p1_add_76645_comb;
  wire [19:0] p1_add_76646_comb;
  wire [19:0] p1_bit_slice_76647_comb;
  wire [18:0] p1_smul_76648_comb;
  wire [18:0] p1_smul_76651_comb;
  wire [18:0] p1_smul_76652_comb;
  wire [18:0] p1_smul_76655_comb;
  wire [18:0] p1_smul_76656_comb;
  wire [18:0] p1_smul_76659_comb;
  wire [18:0] p1_smul_76660_comb;
  wire [18:0] p1_smul_76663_comb;
  wire [19:0] p1_add_76664_comb;
  wire [19:0] p1_add_76666_comb;
  wire [19:0] p1_add_76668_comb;
  wire [19:0] p1_add_76670_comb;
  wire [19:0] p1_add_76672_comb;
  wire [19:0] p1_add_76674_comb;
  wire [19:0] p1_add_76676_comb;
  wire [19:0] p1_add_76678_comb;
  wire [20:0] p1_smul_76680_comb;
  wire [20:0] p1_smul_76681_comb;
  wire [20:0] p1_smul_76682_comb;
  wire [20:0] p1_smul_76683_comb;
  wire [20:0] p1_smul_76684_comb;
  wire [20:0] p1_smul_76685_comb;
  wire [20:0] p1_smul_76686_comb;
  wire [20:0] p1_smul_76687_comb;
  wire [20:0] p1_smul_76688_comb;
  wire [20:0] p1_smul_76689_comb;
  wire [20:0] p1_smul_76690_comb;
  wire [20:0] p1_smul_76691_comb;
  wire [20:0] p1_smul_76692_comb;
  wire [20:0] p1_smul_76693_comb;
  wire [20:0] p1_smul_76694_comb;
  wire [20:0] p1_smul_76695_comb;
  wire [19:0] p1_add_76696_comb;
  wire [19:0] p1_add_76698_comb;
  wire [19:0] p1_add_76700_comb;
  wire [19:0] p1_add_76702_comb;
  wire [19:0] p1_add_76704_comb;
  wire [19:0] p1_add_76706_comb;
  wire [19:0] p1_add_76708_comb;
  wire [19:0] p1_add_76710_comb;
  wire [18:0] p1_smul_76713_comb;
  wire [18:0] p1_smul_76715_comb;
  wire [18:0] p1_smul_76716_comb;
  wire [18:0] p1_smul_76718_comb;
  wire [18:0] p1_smul_76721_comb;
  wire [18:0] p1_smul_76723_comb;
  wire [18:0] p1_smul_76724_comb;
  wire [18:0] p1_smul_76726_comb;
  wire [19:0] p1_add_76728_comb;
  wire [19:0] p1_bit_slice_76729_comb;
  wire [19:0] p1_bit_slice_76730_comb;
  wire [19:0] p1_add_76731_comb;
  wire [19:0] p1_add_76732_comb;
  wire [19:0] p1_bit_slice_76733_comb;
  wire [19:0] p1_bit_slice_76734_comb;
  wire [19:0] p1_add_76735_comb;
  wire [12:0] p1_add_76736_comb;
  wire [12:0] p1_add_76737_comb;
  wire [12:0] p1_add_76738_comb;
  wire [12:0] p1_add_76739_comb;
  wire [12:0] p1_add_76740_comb;
  wire [12:0] p1_add_76741_comb;
  wire [12:0] p1_add_76742_comb;
  wire [12:0] p1_add_76743_comb;
  wire [12:0] p1_add_76744_comb;
  wire [12:0] p1_add_76745_comb;
  wire [12:0] p1_add_76746_comb;
  wire [12:0] p1_add_76747_comb;
  wire [12:0] p1_add_76748_comb;
  wire [12:0] p1_add_76749_comb;
  wire [12:0] p1_add_76750_comb;
  wire [12:0] p1_add_76751_comb;
  wire [18:0] p1_add_76768_comb;
  wire [18:0] p1_add_76770_comb;
  wire [18:0] p1_add_76772_comb;
  wire [18:0] p1_add_76774_comb;
  wire [18:0] p1_add_76776_comb;
  wire [18:0] p1_add_76778_comb;
  wire [18:0] p1_add_76780_comb;
  wire [18:0] p1_add_76782_comb;
  wire [18:0] p1_add_76784_comb;
  wire [18:0] p1_add_76786_comb;
  wire [18:0] p1_add_76788_comb;
  wire [18:0] p1_add_76790_comb;
  wire [18:0] p1_add_76792_comb;
  wire [18:0] p1_add_76794_comb;
  wire [18:0] p1_add_76796_comb;
  wire [18:0] p1_add_76798_comb;
  wire [20:0] p1_concat_76800_comb;
  wire [20:0] p1_concat_76801_comb;
  wire [20:0] p1_concat_76802_comb;
  wire [20:0] p1_concat_76803_comb;
  wire [20:0] p1_concat_76804_comb;
  wire [20:0] p1_concat_76805_comb;
  wire [20:0] p1_concat_76806_comb;
  wire [20:0] p1_concat_76807_comb;
  wire [20:0] p1_concat_76808_comb;
  wire [20:0] p1_concat_76809_comb;
  wire [20:0] p1_concat_76810_comb;
  wire [20:0] p1_concat_76811_comb;
  wire [20:0] p1_concat_76812_comb;
  wire [20:0] p1_concat_76813_comb;
  wire [20:0] p1_concat_76814_comb;
  wire [20:0] p1_concat_76815_comb;
  wire [20:0] p1_add_76816_comb;
  wire [20:0] p1_add_76817_comb;
  wire [20:0] p1_add_76818_comb;
  wire [20:0] p1_add_76819_comb;
  wire [20:0] p1_add_76820_comb;
  wire [20:0] p1_add_76821_comb;
  wire [20:0] p1_add_76822_comb;
  wire [20:0] p1_add_76823_comb;
  wire [20:0] p1_add_76824_comb;
  wire [20:0] p1_add_76825_comb;
  wire [20:0] p1_add_76826_comb;
  wire [20:0] p1_add_76827_comb;
  wire [20:0] p1_add_76828_comb;
  wire [20:0] p1_add_76829_comb;
  wire [20:0] p1_add_76830_comb;
  wire [20:0] p1_add_76831_comb;
  wire [20:0] p1_concat_76832_comb;
  wire [20:0] p1_concat_76833_comb;
  wire [20:0] p1_concat_76834_comb;
  wire [20:0] p1_concat_76835_comb;
  wire [20:0] p1_concat_76836_comb;
  wire [20:0] p1_concat_76837_comb;
  wire [20:0] p1_concat_76838_comb;
  wire [20:0] p1_concat_76839_comb;
  wire [20:0] p1_concat_76840_comb;
  wire [20:0] p1_concat_76841_comb;
  wire [20:0] p1_concat_76842_comb;
  wire [20:0] p1_concat_76843_comb;
  wire [20:0] p1_concat_76844_comb;
  wire [20:0] p1_concat_76845_comb;
  wire [20:0] p1_concat_76846_comb;
  wire [20:0] p1_concat_76847_comb;
  wire [18:0] p1_add_76848_comb;
  wire [18:0] p1_add_76850_comb;
  wire [18:0] p1_add_76852_comb;
  wire [18:0] p1_add_76854_comb;
  wire [18:0] p1_add_76856_comb;
  wire [18:0] p1_add_76858_comb;
  wire [18:0] p1_add_76860_comb;
  wire [18:0] p1_add_76862_comb;
  wire [18:0] p1_add_76864_comb;
  wire [18:0] p1_add_76866_comb;
  wire [18:0] p1_add_76868_comb;
  wire [18:0] p1_add_76870_comb;
  wire [18:0] p1_add_76872_comb;
  wire [18:0] p1_add_76874_comb;
  wire [18:0] p1_add_76876_comb;
  wire [18:0] p1_add_76878_comb;
  wire [12:0] p1_add_76896_comb;
  wire [12:0] p1_add_76897_comb;
  wire [12:0] p1_add_76898_comb;
  wire [12:0] p1_add_76899_comb;
  wire [12:0] p1_add_76900_comb;
  wire [12:0] p1_add_76901_comb;
  wire [12:0] p1_add_76902_comb;
  wire [12:0] p1_add_76903_comb;
  wire [18:0] p1_add_76912_comb;
  wire [18:0] p1_add_76914_comb;
  wire [18:0] p1_add_76916_comb;
  wire [18:0] p1_add_76918_comb;
  wire [18:0] p1_add_76920_comb;
  wire [18:0] p1_add_76922_comb;
  wire [18:0] p1_add_76924_comb;
  wire [18:0] p1_add_76926_comb;
  wire [20:0] p1_concat_76928_comb;
  wire [20:0] p1_concat_76929_comb;
  wire [20:0] p1_concat_76930_comb;
  wire [20:0] p1_concat_76931_comb;
  wire [20:0] p1_concat_76932_comb;
  wire [20:0] p1_concat_76933_comb;
  wire [20:0] p1_concat_76934_comb;
  wire [20:0] p1_concat_76935_comb;
  wire [20:0] p1_add_76936_comb;
  wire [20:0] p1_add_76937_comb;
  wire [20:0] p1_add_76938_comb;
  wire [20:0] p1_add_76939_comb;
  wire [20:0] p1_add_76940_comb;
  wire [20:0] p1_add_76941_comb;
  wire [20:0] p1_add_76942_comb;
  wire [20:0] p1_add_76943_comb;
  wire [20:0] p1_concat_76944_comb;
  wire [20:0] p1_concat_76945_comb;
  wire [20:0] p1_concat_76946_comb;
  wire [20:0] p1_concat_76947_comb;
  wire [20:0] p1_concat_76948_comb;
  wire [20:0] p1_concat_76949_comb;
  wire [20:0] p1_concat_76950_comb;
  wire [20:0] p1_concat_76951_comb;
  wire [18:0] p1_add_76952_comb;
  wire [18:0] p1_add_76954_comb;
  wire [18:0] p1_add_76956_comb;
  wire [18:0] p1_add_76958_comb;
  wire [18:0] p1_add_76960_comb;
  wire [18:0] p1_add_76962_comb;
  wire [18:0] p1_add_76964_comb;
  wire [18:0] p1_add_76966_comb;
  wire [12:0] p1_add_76976_comb;
  wire [12:0] p1_add_76977_comb;
  wire [12:0] p1_add_76978_comb;
  wire [12:0] p1_add_76979_comb;
  wire [12:0] p1_add_76980_comb;
  wire [12:0] p1_add_76981_comb;
  wire [12:0] p1_add_76982_comb;
  wire [12:0] p1_add_76983_comb;
  wire [18:0] p1_add_76992_comb;
  wire [18:0] p1_add_76994_comb;
  wire [18:0] p1_add_76996_comb;
  wire [18:0] p1_add_76998_comb;
  wire [18:0] p1_add_77000_comb;
  wire [18:0] p1_add_77002_comb;
  wire [18:0] p1_add_77004_comb;
  wire [18:0] p1_add_77006_comb;
  wire [20:0] p1_concat_77008_comb;
  wire [20:0] p1_concat_77009_comb;
  wire [20:0] p1_concat_77010_comb;
  wire [20:0] p1_concat_77011_comb;
  wire [20:0] p1_concat_77012_comb;
  wire [20:0] p1_concat_77013_comb;
  wire [20:0] p1_concat_77014_comb;
  wire [20:0] p1_concat_77015_comb;
  wire [20:0] p1_add_77016_comb;
  wire [20:0] p1_add_77017_comb;
  wire [20:0] p1_add_77018_comb;
  wire [20:0] p1_add_77019_comb;
  wire [20:0] p1_add_77020_comb;
  wire [20:0] p1_add_77021_comb;
  wire [20:0] p1_add_77022_comb;
  wire [20:0] p1_add_77023_comb;
  wire [20:0] p1_concat_77024_comb;
  wire [20:0] p1_concat_77025_comb;
  wire [20:0] p1_concat_77026_comb;
  wire [20:0] p1_concat_77027_comb;
  wire [20:0] p1_concat_77028_comb;
  wire [20:0] p1_concat_77029_comb;
  wire [20:0] p1_concat_77030_comb;
  wire [20:0] p1_concat_77031_comb;
  wire [18:0] p1_add_77032_comb;
  wire [18:0] p1_add_77034_comb;
  wire [18:0] p1_add_77036_comb;
  wire [18:0] p1_add_77038_comb;
  wire [18:0] p1_add_77040_comb;
  wire [18:0] p1_add_77042_comb;
  wire [18:0] p1_add_77044_comb;
  wire [18:0] p1_add_77046_comb;
  wire [23:0] p1_add_77072_comb;
  wire [23:0] p1_add_77074_comb;
  wire [23:0] p1_add_77076_comb;
  wire [23:0] p1_add_77078_comb;
  wire [23:0] p1_add_77080_comb;
  wire [23:0] p1_add_77082_comb;
  wire [23:0] p1_add_77084_comb;
  wire [23:0] p1_add_77086_comb;
  wire [19:0] p1_concat_77088_comb;
  wire [19:0] p1_concat_77089_comb;
  wire [19:0] p1_concat_77090_comb;
  wire [19:0] p1_concat_77091_comb;
  wire [19:0] p1_concat_77092_comb;
  wire [19:0] p1_concat_77093_comb;
  wire [19:0] p1_concat_77094_comb;
  wire [19:0] p1_concat_77095_comb;
  wire [19:0] p1_concat_77096_comb;
  wire [19:0] p1_concat_77097_comb;
  wire [19:0] p1_concat_77098_comb;
  wire [19:0] p1_concat_77099_comb;
  wire [19:0] p1_concat_77100_comb;
  wire [19:0] p1_concat_77101_comb;
  wire [19:0] p1_concat_77102_comb;
  wire [19:0] p1_concat_77103_comb;
  wire [24:0] p1_sum__1756_comb;
  wire [24:0] p1_sum__1757_comb;
  wire [24:0] p1_sum__1758_comb;
  wire [24:0] p1_sum__1759_comb;
  wire [24:0] p1_sum__1732_comb;
  wire [24:0] p1_sum__1733_comb;
  wire [24:0] p1_sum__1734_comb;
  wire [24:0] p1_sum__1735_comb;
  wire [24:0] p1_sum__1704_comb;
  wire [24:0] p1_sum__1705_comb;
  wire [24:0] p1_sum__1706_comb;
  wire [24:0] p1_sum__1707_comb;
  wire [24:0] p1_sum__1676_comb;
  wire [24:0] p1_sum__1677_comb;
  wire [24:0] p1_sum__1678_comb;
  wire [24:0] p1_sum__1679_comb;
  wire [24:0] p1_sum__1736_comb;
  wire [24:0] p1_sum__1737_comb;
  wire [24:0] p1_sum__1738_comb;
  wire [24:0] p1_sum__1739_comb;
  wire [24:0] p1_sum__1708_comb;
  wire [24:0] p1_sum__1709_comb;
  wire [24:0] p1_sum__1710_comb;
  wire [24:0] p1_sum__1711_comb;
  wire [24:0] p1_sum__1680_comb;
  wire [24:0] p1_sum__1681_comb;
  wire [24:0] p1_sum__1682_comb;
  wire [24:0] p1_sum__1683_comb;
  wire [24:0] p1_sum__1652_comb;
  wire [24:0] p1_sum__1653_comb;
  wire [24:0] p1_sum__1654_comb;
  wire [24:0] p1_sum__1655_comb;
  wire [24:0] p1_sum__1712_comb;
  wire [24:0] p1_sum__1713_comb;
  wire [24:0] p1_sum__1714_comb;
  wire [24:0] p1_sum__1715_comb;
  wire [24:0] p1_sum__1684_comb;
  wire [24:0] p1_sum__1685_comb;
  wire [24:0] p1_sum__1686_comb;
  wire [24:0] p1_sum__1687_comb;
  wire [24:0] p1_sum__1656_comb;
  wire [24:0] p1_sum__1657_comb;
  wire [24:0] p1_sum__1658_comb;
  wire [24:0] p1_sum__1659_comb;
  wire [24:0] p1_sum__1632_comb;
  wire [24:0] p1_sum__1633_comb;
  wire [24:0] p1_sum__1634_comb;
  wire [24:0] p1_sum__1635_comb;
  wire [19:0] p1_concat_77152_comb;
  wire [19:0] p1_concat_77153_comb;
  wire [19:0] p1_concat_77154_comb;
  wire [19:0] p1_concat_77155_comb;
  wire [19:0] p1_concat_77156_comb;
  wire [19:0] p1_concat_77157_comb;
  wire [19:0] p1_concat_77158_comb;
  wire [19:0] p1_concat_77159_comb;
  wire [19:0] p1_concat_77160_comb;
  wire [19:0] p1_concat_77161_comb;
  wire [19:0] p1_concat_77162_comb;
  wire [19:0] p1_concat_77163_comb;
  wire [19:0] p1_concat_77164_comb;
  wire [19:0] p1_concat_77165_comb;
  wire [19:0] p1_concat_77166_comb;
  wire [19:0] p1_concat_77167_comb;
  wire [23:0] p1_add_77168_comb;
  wire [23:0] p1_add_77170_comb;
  wire [23:0] p1_add_77172_comb;
  wire [23:0] p1_add_77174_comb;
  wire [23:0] p1_add_77176_comb;
  wire [23:0] p1_add_77178_comb;
  wire [23:0] p1_add_77180_comb;
  wire [23:0] p1_add_77182_comb;
  wire [23:0] p1_add_77192_comb;
  wire [23:0] p1_add_77194_comb;
  wire [23:0] p1_add_77196_comb;
  wire [23:0] p1_add_77198_comb;
  wire [19:0] p1_concat_77200_comb;
  wire [19:0] p1_concat_77201_comb;
  wire [19:0] p1_concat_77202_comb;
  wire [19:0] p1_concat_77203_comb;
  wire [19:0] p1_concat_77204_comb;
  wire [19:0] p1_concat_77205_comb;
  wire [19:0] p1_concat_77206_comb;
  wire [19:0] p1_concat_77207_comb;
  wire [24:0] p1_sum__1776_comb;
  wire [24:0] p1_sum__1777_comb;
  wire [24:0] p1_sum__1778_comb;
  wire [24:0] p1_sum__1779_comb;
  wire [24:0] p1_sum__1648_comb;
  wire [24:0] p1_sum__1649_comb;
  wire [24:0] p1_sum__1650_comb;
  wire [24:0] p1_sum__1651_comb;
  wire [24:0] p1_sum__1760_comb;
  wire [24:0] p1_sum__1761_comb;
  wire [24:0] p1_sum__1762_comb;
  wire [24:0] p1_sum__1763_comb;
  wire [24:0] p1_sum__1628_comb;
  wire [24:0] p1_sum__1629_comb;
  wire [24:0] p1_sum__1630_comb;
  wire [24:0] p1_sum__1631_comb;
  wire [24:0] p1_sum__1740_comb;
  wire [24:0] p1_sum__1741_comb;
  wire [24:0] p1_sum__1742_comb;
  wire [24:0] p1_sum__1743_comb;
  wire [24:0] p1_sum__1612_comb;
  wire [24:0] p1_sum__1613_comb;
  wire [24:0] p1_sum__1614_comb;
  wire [24:0] p1_sum__1615_comb;
  wire [19:0] p1_concat_77232_comb;
  wire [19:0] p1_concat_77233_comb;
  wire [19:0] p1_concat_77234_comb;
  wire [19:0] p1_concat_77235_comb;
  wire [19:0] p1_concat_77236_comb;
  wire [19:0] p1_concat_77237_comb;
  wire [19:0] p1_concat_77238_comb;
  wire [19:0] p1_concat_77239_comb;
  wire [23:0] p1_add_77240_comb;
  wire [23:0] p1_add_77242_comb;
  wire [23:0] p1_add_77244_comb;
  wire [23:0] p1_add_77246_comb;
  wire [23:0] p1_add_77256_comb;
  wire [23:0] p1_add_77258_comb;
  wire [23:0] p1_add_77260_comb;
  wire [23:0] p1_add_77262_comb;
  wire [19:0] p1_concat_77264_comb;
  wire [19:0] p1_concat_77265_comb;
  wire [19:0] p1_concat_77266_comb;
  wire [19:0] p1_concat_77267_comb;
  wire [19:0] p1_concat_77268_comb;
  wire [19:0] p1_concat_77269_comb;
  wire [19:0] p1_concat_77270_comb;
  wire [19:0] p1_concat_77271_comb;
  wire [24:0] p1_sum__1792_comb;
  wire [24:0] p1_sum__1793_comb;
  wire [24:0] p1_sum__1794_comb;
  wire [24:0] p1_sum__1795_comb;
  wire [24:0] p1_sum__1624_comb;
  wire [24:0] p1_sum__1625_comb;
  wire [24:0] p1_sum__1626_comb;
  wire [24:0] p1_sum__1627_comb;
  wire [24:0] p1_sum__1780_comb;
  wire [24:0] p1_sum__1781_comb;
  wire [24:0] p1_sum__1782_comb;
  wire [24:0] p1_sum__1783_comb;
  wire [24:0] p1_sum__1608_comb;
  wire [24:0] p1_sum__1609_comb;
  wire [24:0] p1_sum__1610_comb;
  wire [24:0] p1_sum__1611_comb;
  wire [24:0] p1_sum__1764_comb;
  wire [24:0] p1_sum__1765_comb;
  wire [24:0] p1_sum__1766_comb;
  wire [24:0] p1_sum__1767_comb;
  wire [24:0] p1_sum__1596_comb;
  wire [24:0] p1_sum__1597_comb;
  wire [24:0] p1_sum__1598_comb;
  wire [24:0] p1_sum__1599_comb;
  wire [19:0] p1_concat_77296_comb;
  wire [19:0] p1_concat_77297_comb;
  wire [19:0] p1_concat_77298_comb;
  wire [19:0] p1_concat_77299_comb;
  wire [19:0] p1_concat_77300_comb;
  wire [19:0] p1_concat_77301_comb;
  wire [19:0] p1_concat_77302_comb;
  wire [19:0] p1_concat_77303_comb;
  wire [23:0] p1_add_77304_comb;
  wire [23:0] p1_add_77306_comb;
  wire [23:0] p1_add_77308_comb;
  wire [23:0] p1_add_77310_comb;
  wire [23:0] p1_add_77312_comb;
  wire [23:0] p1_add_77313_comb;
  wire [23:0] p1_add_77314_comb;
  wire [23:0] p1_add_77315_comb;
  wire [23:0] p1_add_77316_comb;
  wire [23:0] p1_add_77317_comb;
  wire [23:0] p1_add_77318_comb;
  wire [23:0] p1_add_77319_comb;
  wire [24:0] p1_sum__1348_comb;
  wire [24:0] p1_sum__1349_comb;
  wire [24:0] p1_sum__1340_comb;
  wire [24:0] p1_sum__1341_comb;
  wire [24:0] p1_sum__1330_comb;
  wire [24:0] p1_sum__1331_comb;
  wire [24:0] p1_sum__1318_comb;
  wire [24:0] p1_sum__1319_comb;
  wire [24:0] p1_sum__1334_comb;
  wire [24:0] p1_sum__1335_comb;
  wire [24:0] p1_sum__1322_comb;
  wire [24:0] p1_sum__1323_comb;
  wire [24:0] p1_sum__1308_comb;
  wire [24:0] p1_sum__1309_comb;
  wire [24:0] p1_sum__1294_comb;
  wire [24:0] p1_sum__1295_comb;
  wire [24:0] p1_sum__1324_comb;
  wire [24:0] p1_sum__1325_comb;
  wire [24:0] p1_sum__1310_comb;
  wire [24:0] p1_sum__1311_comb;
  wire [24:0] p1_sum__1296_comb;
  wire [24:0] p1_sum__1297_comb;
  wire [24:0] p1_sum__1282_comb;
  wire [24:0] p1_sum__1283_comb;
  wire [24:0] p1_sum__1312_comb;
  wire [24:0] p1_sum__1313_comb;
  wire [24:0] p1_sum__1298_comb;
  wire [24:0] p1_sum__1299_comb;
  wire [24:0] p1_sum__1284_comb;
  wire [24:0] p1_sum__1285_comb;
  wire [24:0] p1_sum__1272_comb;
  wire [24:0] p1_sum__1273_comb;
  wire [24:0] p1_sum__1288_comb;
  wire [24:0] p1_sum__1289_comb;
  wire [24:0] p1_sum__1276_comb;
  wire [24:0] p1_sum__1277_comb;
  wire [24:0] p1_sum__1266_comb;
  wire [24:0] p1_sum__1267_comb;
  wire [24:0] p1_sum__1258_comb;
  wire [24:0] p1_sum__1259_comb;
  wire [23:0] p1_add_77392_comb;
  wire [23:0] p1_add_77393_comb;
  wire [23:0] p1_add_77394_comb;
  wire [23:0] p1_add_77395_comb;
  wire [24:0] p1_sum__1354_comb;
  wire [24:0] p1_sum__1355_comb;
  wire [24:0] p1_sum__1304_comb;
  wire [24:0] p1_sum__1305_comb;
  wire [24:0] p1_sum__1344_comb;
  wire [24:0] p1_sum__1345_comb;
  wire [24:0] p1_sum__1280_comb;
  wire [24:0] p1_sum__1281_comb;
  wire [24:0] p1_sum__1336_comb;
  wire [24:0] p1_sum__1337_comb;
  wire [24:0] p1_sum__1270_comb;
  wire [24:0] p1_sum__1271_comb;
  wire [24:0] p1_sum__1326_comb;
  wire [24:0] p1_sum__1327_comb;
  wire [24:0] p1_sum__1262_comb;
  wire [24:0] p1_sum__1263_comb;
  wire [24:0] p1_sum__1302_comb;
  wire [24:0] p1_sum__1303_comb;
  wire [24:0] p1_sum__1252_comb;
  wire [24:0] p1_sum__1253_comb;
  wire [23:0] p1_add_77432_comb;
  wire [23:0] p1_add_77433_comb;
  wire [23:0] p1_add_77434_comb;
  wire [23:0] p1_add_77435_comb;
  wire [24:0] p1_sum__1358_comb;
  wire [24:0] p1_sum__1359_comb;
  wire [24:0] p1_sum__1290_comb;
  wire [24:0] p1_sum__1291_comb;
  wire [24:0] p1_sum__1352_comb;
  wire [24:0] p1_sum__1353_comb;
  wire [24:0] p1_sum__1268_comb;
  wire [24:0] p1_sum__1269_comb;
  wire [24:0] p1_sum__1346_comb;
  wire [24:0] p1_sum__1347_comb;
  wire [24:0] p1_sum__1260_comb;
  wire [24:0] p1_sum__1261_comb;
  wire [24:0] p1_sum__1338_comb;
  wire [24:0] p1_sum__1339_comb;
  wire [24:0] p1_sum__1254_comb;
  wire [24:0] p1_sum__1255_comb;
  wire [24:0] p1_sum__1316_comb;
  wire [24:0] p1_sum__1317_comb;
  wire [24:0] p1_sum__1248_comb;
  wire [24:0] p1_sum__1249_comb;
  wire [23:0] p1_add_77472_comb;
  wire [23:0] p1_add_77474_comb;
  wire [23:0] p1_add_77476_comb;
  wire [23:0] p1_add_77478_comb;
  wire [24:0] p1_sum__1130_comb;
  wire [24:0] p1_sum__1126_comb;
  wire [24:0] p1_sum__1121_comb;
  wire [24:0] p1_sum__1115_comb;
  wire [23:0] p1_add_77488_comb;
  wire [23:0] p1_add_77489_comb;
  wire [23:0] p1_add_77490_comb;
  wire [23:0] p1_add_77491_comb;
  wire [23:0] p1_add_77492_comb;
  wire [23:0] p1_add_77493_comb;
  wire [23:0] p1_add_77494_comb;
  wire [23:0] p1_add_77495_comb;
  wire [24:0] p1_sum__1123_comb;
  wire [24:0] p1_sum__1117_comb;
  wire [24:0] p1_sum__1110_comb;
  wire [24:0] p1_sum__1103_comb;
  wire [24:0] p1_sum__1118_comb;
  wire [24:0] p1_sum__1111_comb;
  wire [24:0] p1_sum__1104_comb;
  wire [24:0] p1_sum__1097_comb;
  wire [24:0] p1_sum__1112_comb;
  wire [24:0] p1_sum__1105_comb;
  wire [24:0] p1_sum__1098_comb;
  wire [24:0] p1_sum__1092_comb;
  wire [23:0] p1_add_77520_comb;
  wire [23:0] p1_add_77521_comb;
  wire [23:0] p1_add_77522_comb;
  wire [23:0] p1_add_77523_comb;
  wire [23:0] p1_add_77524_comb;
  wire [23:0] p1_add_77525_comb;
  wire [23:0] p1_add_77526_comb;
  wire [23:0] p1_add_77527_comb;
  wire [24:0] p1_sum__1100_comb;
  wire [24:0] p1_sum__1094_comb;
  wire [24:0] p1_sum__1089_comb;
  wire [24:0] p1_sum__1085_comb;
  wire [23:0] p1_add_77536_comb;
  wire [23:0] p1_add_77538_comb;
  wire [24:0] p1_sum__1133_comb;
  wire [24:0] p1_sum__1108_comb;
  wire [23:0] p1_add_77544_comb;
  wire [23:0] p1_add_77545_comb;
  wire [23:0] p1_add_77546_comb;
  wire [23:0] p1_add_77547_comb;
  wire [24:0] p1_sum__1128_comb;
  wire [24:0] p1_sum__1096_comb;
  wire [24:0] p1_sum__1124_comb;
  wire [24:0] p1_sum__1091_comb;
  wire [24:0] p1_sum__1119_comb;
  wire [24:0] p1_sum__1087_comb;
  wire [23:0] p1_add_77560_comb;
  wire [23:0] p1_add_77561_comb;
  wire [23:0] p1_add_77562_comb;
  wire [23:0] p1_add_77563_comb;
  wire [24:0] p1_sum__1107_comb;
  wire [24:0] p1_sum__1082_comb;
  wire [23:0] p1_add_77568_comb;
  wire [23:0] p1_add_77570_comb;
  wire [24:0] p1_sum__1135_comb;
  wire [24:0] p1_sum__1101_comb;
  wire [23:0] p1_add_77576_comb;
  wire [23:0] p1_add_77577_comb;
  wire [23:0] p1_add_77578_comb;
  wire [23:0] p1_add_77579_comb;
  wire [24:0] p1_sum__1132_comb;
  wire [24:0] p1_sum__1090_comb;
  wire [24:0] p1_sum__1129_comb;
  wire [24:0] p1_sum__1086_comb;
  wire [24:0] p1_sum__1125_comb;
  wire [24:0] p1_sum__1083_comb;
  wire [23:0] p1_add_77592_comb;
  wire [23:0] p1_add_77593_comb;
  wire [23:0] p1_add_77594_comb;
  wire [23:0] p1_add_77595_comb;
  wire [24:0] p1_sum__1114_comb;
  wire [24:0] p1_sum__1080_comb;
  wire [23:0] p1_umul_27340_NarrowedMult__comb;
  wire [23:0] p1_umul_27342_NarrowedMult__comb;
  wire [23:0] p1_umul_27344_NarrowedMult__comb;
  wire [23:0] p1_umul_27346_NarrowedMult__comb;
  wire [24:0] p1_add_77604_comb;
  wire [24:0] p1_add_77605_comb;
  wire [24:0] p1_add_77606_comb;
  wire [24:0] p1_add_77607_comb;
  wire [23:0] p1_add_77608_comb;
  wire [23:0] p1_add_77609_comb;
  wire [23:0] p1_add_77610_comb;
  wire [23:0] p1_add_77611_comb;
  wire [24:0] p1_add_77612_comb;
  wire [24:0] p1_add_77613_comb;
  wire [24:0] p1_add_77614_comb;
  wire [24:0] p1_add_77615_comb;
  wire [24:0] p1_add_77616_comb;
  wire [24:0] p1_add_77617_comb;
  wire [24:0] p1_add_77618_comb;
  wire [24:0] p1_add_77619_comb;
  wire [24:0] p1_add_77620_comb;
  wire [24:0] p1_add_77621_comb;
  wire [24:0] p1_add_77622_comb;
  wire [24:0] p1_add_77623_comb;
  wire [23:0] p1_add_77624_comb;
  wire [23:0] p1_add_77625_comb;
  wire [23:0] p1_add_77626_comb;
  wire [23:0] p1_add_77627_comb;
  wire [24:0] p1_add_77628_comb;
  wire [24:0] p1_add_77629_comb;
  wire [24:0] p1_add_77630_comb;
  wire [24:0] p1_add_77631_comb;
  wire [23:0] p1_umul_27338_NarrowedMult__comb;
  wire [23:0] p1_umul_27348_NarrowedMult__comb;
  wire [24:0] p1_add_77634_comb;
  wire [24:0] p1_add_77635_comb;
  wire [23:0] p1_add_77636_comb;
  wire [23:0] p1_add_77637_comb;
  wire [24:0] p1_add_77638_comb;
  wire [24:0] p1_add_77639_comb;
  wire [24:0] p1_add_77640_comb;
  wire [24:0] p1_add_77641_comb;
  wire [24:0] p1_add_77642_comb;
  wire [24:0] p1_add_77643_comb;
  wire [23:0] p1_add_77644_comb;
  wire [23:0] p1_add_77645_comb;
  wire [24:0] p1_add_77646_comb;
  wire [24:0] p1_add_77647_comb;
  wire [23:0] p1_umul_27336_NarrowedMult__comb;
  wire [23:0] p1_umul_27350_NarrowedMult__comb;
  wire [24:0] p1_add_77650_comb;
  wire [24:0] p1_add_77651_comb;
  wire [23:0] p1_add_77652_comb;
  wire [23:0] p1_add_77653_comb;
  wire [24:0] p1_add_77654_comb;
  wire [24:0] p1_add_77655_comb;
  wire [24:0] p1_add_77656_comb;
  wire [24:0] p1_add_77657_comb;
  wire [24:0] p1_add_77658_comb;
  wire [24:0] p1_add_77659_comb;
  wire [23:0] p1_add_77660_comb;
  wire [23:0] p1_add_77661_comb;
  wire [24:0] p1_add_77662_comb;
  wire [24:0] p1_add_77663_comb;
  wire [16:0] p1_bit_slice_77664_comb;
  wire [16:0] p1_bit_slice_77665_comb;
  wire [16:0] p1_bit_slice_77666_comb;
  wire [16:0] p1_bit_slice_77667_comb;
  wire [16:0] p1_bit_slice_77668_comb;
  wire [16:0] p1_bit_slice_77669_comb;
  wire [16:0] p1_bit_slice_77670_comb;
  wire [16:0] p1_bit_slice_77671_comb;
  wire [16:0] p1_bit_slice_77672_comb;
  wire [16:0] p1_bit_slice_77673_comb;
  wire [16:0] p1_bit_slice_77674_comb;
  wire [16:0] p1_bit_slice_77675_comb;
  wire [16:0] p1_bit_slice_77676_comb;
  wire [16:0] p1_bit_slice_77677_comb;
  wire [16:0] p1_bit_slice_77678_comb;
  wire [16:0] p1_bit_slice_77679_comb;
  wire [16:0] p1_bit_slice_77680_comb;
  wire [16:0] p1_bit_slice_77681_comb;
  wire [16:0] p1_bit_slice_77682_comb;
  wire [16:0] p1_bit_slice_77683_comb;
  wire [16:0] p1_bit_slice_77684_comb;
  wire [16:0] p1_bit_slice_77685_comb;
  wire [16:0] p1_bit_slice_77686_comb;
  wire [16:0] p1_bit_slice_77687_comb;
  wire [16:0] p1_bit_slice_77688_comb;
  wire [16:0] p1_bit_slice_77689_comb;
  wire [16:0] p1_bit_slice_77690_comb;
  wire [16:0] p1_bit_slice_77691_comb;
  wire [16:0] p1_bit_slice_77692_comb;
  wire [16:0] p1_bit_slice_77693_comb;
  wire [16:0] p1_bit_slice_77694_comb;
  wire [16:0] p1_bit_slice_77695_comb;
  wire [16:0] p1_bit_slice_77696_comb;
  wire [16:0] p1_bit_slice_77697_comb;
  wire [16:0] p1_bit_slice_77698_comb;
  wire [16:0] p1_bit_slice_77699_comb;
  wire [16:0] p1_bit_slice_77700_comb;
  wire [16:0] p1_bit_slice_77701_comb;
  wire [16:0] p1_bit_slice_77702_comb;
  wire [16:0] p1_bit_slice_77703_comb;
  wire [16:0] p1_bit_slice_77704_comb;
  wire [16:0] p1_bit_slice_77705_comb;
  wire [16:0] p1_bit_slice_77706_comb;
  wire [16:0] p1_bit_slice_77707_comb;
  wire [16:0] p1_bit_slice_77708_comb;
  wire [16:0] p1_bit_slice_77709_comb;
  wire [16:0] p1_bit_slice_77710_comb;
  wire [16:0] p1_bit_slice_77711_comb;
  wire [16:0] p1_bit_slice_77712_comb;
  wire [16:0] p1_bit_slice_77713_comb;
  wire [16:0] p1_bit_slice_77714_comb;
  wire [16:0] p1_bit_slice_77715_comb;
  wire [16:0] p1_bit_slice_77716_comb;
  wire [16:0] p1_bit_slice_77717_comb;
  wire [16:0] p1_bit_slice_77718_comb;
  wire [16:0] p1_bit_slice_77719_comb;
  wire [16:0] p1_bit_slice_77720_comb;
  wire [16:0] p1_bit_slice_77721_comb;
  wire [16:0] p1_bit_slice_77722_comb;
  wire [16:0] p1_bit_slice_77723_comb;
  wire [16:0] p1_bit_slice_77724_comb;
  wire [16:0] p1_bit_slice_77725_comb;
  wire [16:0] p1_bit_slice_77726_comb;
  wire [16:0] p1_bit_slice_77727_comb;
  wire [17:0] p1_add_77856_comb;
  wire [17:0] p1_add_77857_comb;
  wire [17:0] p1_add_77858_comb;
  wire [17:0] p1_add_77859_comb;
  wire [17:0] p1_add_77860_comb;
  wire [17:0] p1_add_77861_comb;
  wire [17:0] p1_add_77862_comb;
  wire [17:0] p1_add_77863_comb;
  wire [17:0] p1_add_77864_comb;
  wire [17:0] p1_add_77865_comb;
  wire [17:0] p1_add_77866_comb;
  wire [17:0] p1_add_77867_comb;
  wire [17:0] p1_add_77868_comb;
  wire [17:0] p1_add_77869_comb;
  wire [17:0] p1_add_77870_comb;
  wire [17:0] p1_add_77871_comb;
  wire [17:0] p1_add_77872_comb;
  wire [17:0] p1_add_77873_comb;
  wire [17:0] p1_add_77874_comb;
  wire [17:0] p1_add_77875_comb;
  wire [17:0] p1_add_77876_comb;
  wire [17:0] p1_add_77877_comb;
  wire [17:0] p1_add_77878_comb;
  wire [17:0] p1_add_77879_comb;
  wire [17:0] p1_add_77880_comb;
  wire [17:0] p1_add_77881_comb;
  wire [17:0] p1_add_77882_comb;
  wire [17:0] p1_add_77883_comb;
  wire [17:0] p1_add_77884_comb;
  wire [17:0] p1_add_77885_comb;
  wire [17:0] p1_add_77886_comb;
  wire [17:0] p1_add_77887_comb;
  wire [17:0] p1_add_77888_comb;
  wire [17:0] p1_add_77889_comb;
  wire [17:0] p1_add_77890_comb;
  wire [17:0] p1_add_77891_comb;
  wire [17:0] p1_add_77892_comb;
  wire [17:0] p1_add_77893_comb;
  wire [17:0] p1_add_77894_comb;
  wire [17:0] p1_add_77895_comb;
  wire [17:0] p1_add_77896_comb;
  wire [17:0] p1_add_77897_comb;
  wire [17:0] p1_add_77898_comb;
  wire [17:0] p1_add_77899_comb;
  wire [17:0] p1_add_77900_comb;
  wire [17:0] p1_add_77901_comb;
  wire [17:0] p1_add_77902_comb;
  wire [17:0] p1_add_77903_comb;
  wire [17:0] p1_add_77904_comb;
  wire [17:0] p1_add_77905_comb;
  wire [17:0] p1_add_77906_comb;
  wire [17:0] p1_add_77907_comb;
  wire [17:0] p1_add_77908_comb;
  wire [17:0] p1_add_77909_comb;
  wire [17:0] p1_add_77910_comb;
  wire [17:0] p1_add_77911_comb;
  wire [17:0] p1_add_77912_comb;
  wire [17:0] p1_add_77913_comb;
  wire [17:0] p1_add_77914_comb;
  wire [17:0] p1_add_77915_comb;
  wire [17:0] p1_add_77916_comb;
  wire [17:0] p1_add_77917_comb;
  wire [17:0] p1_add_77918_comb;
  wire [17:0] p1_add_77919_comb;
  wire [11:0] p1_clipped__40_comb;
  wire [11:0] p1_clipped__56_comb;
  wire [11:0] p1_clipped__72_comb;
  wire [11:0] p1_clipped__88_comb;
  wire [11:0] p1_clipped__41_comb;
  wire [11:0] p1_clipped__57_comb;
  wire [11:0] p1_clipped__73_comb;
  wire [11:0] p1_clipped__89_comb;
  wire [11:0] p1_clipped__42_comb;
  wire [11:0] p1_clipped__58_comb;
  wire [11:0] p1_clipped__74_comb;
  wire [11:0] p1_clipped__90_comb;
  wire [11:0] p1_clipped__43_comb;
  wire [11:0] p1_clipped__59_comb;
  wire [11:0] p1_clipped__75_comb;
  wire [11:0] p1_clipped__91_comb;
  wire [11:0] p1_clipped__44_comb;
  wire [11:0] p1_clipped__60_comb;
  wire [11:0] p1_clipped__76_comb;
  wire [11:0] p1_clipped__92_comb;
  wire [11:0] p1_clipped__45_comb;
  wire [11:0] p1_clipped__61_comb;
  wire [11:0] p1_clipped__77_comb;
  wire [11:0] p1_clipped__93_comb;
  wire [11:0] p1_clipped__46_comb;
  wire [11:0] p1_clipped__62_comb;
  wire [11:0] p1_clipped__78_comb;
  wire [11:0] p1_clipped__94_comb;
  wire [11:0] p1_clipped__47_comb;
  wire [11:0] p1_clipped__63_comb;
  wire [11:0] p1_clipped__79_comb;
  wire [11:0] p1_clipped__95_comb;
  wire [11:0] p1_clipped__24_comb;
  wire [11:0] p1_clipped__104_comb;
  wire [11:0] p1_clipped__25_comb;
  wire [11:0] p1_clipped__105_comb;
  wire [11:0] p1_clipped__26_comb;
  wire [11:0] p1_clipped__106_comb;
  wire [11:0] p1_clipped__27_comb;
  wire [11:0] p1_clipped__107_comb;
  wire [11:0] p1_clipped__28_comb;
  wire [11:0] p1_clipped__108_comb;
  wire [11:0] p1_clipped__29_comb;
  wire [11:0] p1_clipped__109_comb;
  wire [11:0] p1_clipped__30_comb;
  wire [11:0] p1_clipped__110_comb;
  wire [11:0] p1_clipped__31_comb;
  wire [11:0] p1_clipped__111_comb;
  wire [11:0] p1_clipped__8_comb;
  wire [11:0] p1_clipped__120_comb;
  wire [11:0] p1_clipped__9_comb;
  wire [11:0] p1_clipped__121_comb;
  wire [11:0] p1_clipped__10_comb;
  wire [11:0] p1_clipped__122_comb;
  wire [11:0] p1_clipped__11_comb;
  wire [11:0] p1_clipped__123_comb;
  wire [11:0] p1_clipped__12_comb;
  wire [11:0] p1_clipped__124_comb;
  wire [11:0] p1_clipped__13_comb;
  wire [11:0] p1_clipped__125_comb;
  wire [11:0] p1_clipped__14_comb;
  wire [11:0] p1_clipped__126_comb;
  wire [11:0] p1_clipped__15_comb;
  wire [11:0] p1_clipped__127_comb;
  wire [23:0] p1_sign_ext_78562_comb;
  wire [23:0] p1_sign_ext_78563_comb;
  wire [23:0] p1_sign_ext_78564_comb;
  wire [23:0] p1_sign_ext_78565_comb;
  wire [23:0] p1_sign_ext_78570_comb;
  wire [23:0] p1_sign_ext_78571_comb;
  wire [23:0] p1_sign_ext_78572_comb;
  wire [23:0] p1_sign_ext_78573_comb;
  wire [23:0] p1_sign_ext_78578_comb;
  wire [23:0] p1_sign_ext_78579_comb;
  wire [23:0] p1_sign_ext_78580_comb;
  wire [23:0] p1_sign_ext_78581_comb;
  wire [23:0] p1_sign_ext_78586_comb;
  wire [23:0] p1_sign_ext_78587_comb;
  wire [23:0] p1_sign_ext_78588_comb;
  wire [23:0] p1_sign_ext_78589_comb;
  wire [23:0] p1_sign_ext_78594_comb;
  wire [23:0] p1_sign_ext_78595_comb;
  wire [23:0] p1_sign_ext_78596_comb;
  wire [23:0] p1_sign_ext_78597_comb;
  wire [23:0] p1_sign_ext_78602_comb;
  wire [23:0] p1_sign_ext_78603_comb;
  wire [23:0] p1_sign_ext_78604_comb;
  wire [23:0] p1_sign_ext_78605_comb;
  wire [23:0] p1_sign_ext_78610_comb;
  wire [23:0] p1_sign_ext_78611_comb;
  wire [23:0] p1_sign_ext_78612_comb;
  wire [23:0] p1_sign_ext_78613_comb;
  wire [23:0] p1_sign_ext_78618_comb;
  wire [23:0] p1_sign_ext_78619_comb;
  wire [23:0] p1_sign_ext_78620_comb;
  wire [23:0] p1_sign_ext_78621_comb;
  wire [23:0] p1_sign_ext_78624_comb;
  wire [23:0] p1_sign_ext_78625_comb;
  wire [23:0] p1_sign_ext_78626_comb;
  wire [23:0] p1_sign_ext_78627_comb;
  wire [23:0] p1_sign_ext_78628_comb;
  wire [23:0] p1_sign_ext_78629_comb;
  wire [23:0] p1_sign_ext_78630_comb;
  wire [23:0] p1_sign_ext_78631_comb;
  wire [23:0] p1_sign_ext_78632_comb;
  wire [23:0] p1_sign_ext_78633_comb;
  wire [23:0] p1_sign_ext_78634_comb;
  wire [23:0] p1_sign_ext_78635_comb;
  wire [23:0] p1_sign_ext_78636_comb;
  wire [23:0] p1_sign_ext_78637_comb;
  wire [23:0] p1_sign_ext_78638_comb;
  wire [23:0] p1_sign_ext_78639_comb;
  wire [23:0] p1_sign_ext_78672_comb;
  wire [23:0] p1_sign_ext_78677_comb;
  wire [23:0] p1_sign_ext_78678_comb;
  wire [23:0] p1_sign_ext_78683_comb;
  wire [23:0] p1_sign_ext_78684_comb;
  wire [23:0] p1_sign_ext_78689_comb;
  wire [23:0] p1_sign_ext_78690_comb;
  wire [23:0] p1_sign_ext_78695_comb;
  wire [23:0] p1_sign_ext_78696_comb;
  wire [23:0] p1_sign_ext_78701_comb;
  wire [23:0] p1_sign_ext_78702_comb;
  wire [23:0] p1_sign_ext_78707_comb;
  wire [23:0] p1_sign_ext_78708_comb;
  wire [23:0] p1_sign_ext_78713_comb;
  wire [23:0] p1_sign_ext_78714_comb;
  wire [23:0] p1_sign_ext_78719_comb;
  wire [20:0] p1_smul_78752_comb;
  wire [20:0] p1_smul_78753_comb;
  wire [20:0] p1_smul_78762_comb;
  wire [20:0] p1_smul_78763_comb;
  wire [20:0] p1_smul_78764_comb;
  wire [20:0] p1_smul_78765_comb;
  wire [20:0] p1_smul_78774_comb;
  wire [20:0] p1_smul_78775_comb;
  wire [20:0] p1_smul_78776_comb;
  wire [20:0] p1_smul_78777_comb;
  wire [20:0] p1_smul_78786_comb;
  wire [20:0] p1_smul_78787_comb;
  wire [20:0] p1_smul_78788_comb;
  wire [20:0] p1_smul_78789_comb;
  wire [20:0] p1_smul_78798_comb;
  wire [20:0] p1_smul_78799_comb;
  wire [20:0] p1_smul_78800_comb;
  wire [20:0] p1_smul_78801_comb;
  wire [20:0] p1_smul_78810_comb;
  wire [20:0] p1_smul_78811_comb;
  wire [20:0] p1_smul_78812_comb;
  wire [20:0] p1_smul_78813_comb;
  wire [20:0] p1_smul_78822_comb;
  wire [20:0] p1_smul_78823_comb;
  wire [20:0] p1_smul_78824_comb;
  wire [20:0] p1_smul_78825_comb;
  wire [20:0] p1_smul_78834_comb;
  wire [20:0] p1_smul_78835_comb;
  wire [20:0] p1_smul_78836_comb;
  wire [20:0] p1_smul_78837_comb;
  wire [20:0] p1_smul_78846_comb;
  wire [20:0] p1_smul_78847_comb;
  wire [20:0] p1_smul_78896_comb;
  wire [20:0] p1_smul_78898_comb;
  wire [20:0] p1_smul_78901_comb;
  wire [20:0] p1_smul_78903_comb;
  wire [20:0] p1_smul_78904_comb;
  wire [20:0] p1_smul_78906_comb;
  wire [20:0] p1_smul_78909_comb;
  wire [20:0] p1_smul_78911_comb;
  wire [20:0] p1_smul_78912_comb;
  wire [20:0] p1_smul_78914_comb;
  wire [20:0] p1_smul_78917_comb;
  wire [20:0] p1_smul_78919_comb;
  wire [20:0] p1_smul_78920_comb;
  wire [20:0] p1_smul_78922_comb;
  wire [20:0] p1_smul_78925_comb;
  wire [20:0] p1_smul_78927_comb;
  wire [20:0] p1_smul_78928_comb;
  wire [20:0] p1_smul_78930_comb;
  wire [20:0] p1_smul_78933_comb;
  wire [20:0] p1_smul_78935_comb;
  wire [20:0] p1_smul_78936_comb;
  wire [20:0] p1_smul_78938_comb;
  wire [20:0] p1_smul_78941_comb;
  wire [20:0] p1_smul_78943_comb;
  wire [20:0] p1_smul_78944_comb;
  wire [20:0] p1_smul_78946_comb;
  wire [20:0] p1_smul_78949_comb;
  wire [20:0] p1_smul_78951_comb;
  wire [20:0] p1_smul_78952_comb;
  wire [20:0] p1_smul_78954_comb;
  wire [20:0] p1_smul_78957_comb;
  wire [20:0] p1_smul_78959_comb;
  wire [20:0] p1_smul_78962_comb;
  wire [20:0] p1_smul_78964_comb;
  wire [20:0] p1_smul_78965_comb;
  wire [20:0] p1_smul_78967_comb;
  wire [20:0] p1_smul_78972_comb;
  wire [20:0] p1_smul_78974_comb;
  wire [20:0] p1_smul_78975_comb;
  wire [20:0] p1_smul_78977_comb;
  wire [20:0] p1_smul_78982_comb;
  wire [20:0] p1_smul_78984_comb;
  wire [20:0] p1_smul_78985_comb;
  wire [20:0] p1_smul_78987_comb;
  wire [20:0] p1_smul_78992_comb;
  wire [20:0] p1_smul_78994_comb;
  wire [20:0] p1_smul_78995_comb;
  wire [20:0] p1_smul_78997_comb;
  wire [20:0] p1_smul_79002_comb;
  wire [20:0] p1_smul_79004_comb;
  wire [20:0] p1_smul_79005_comb;
  wire [20:0] p1_smul_79007_comb;
  wire [20:0] p1_smul_79012_comb;
  wire [20:0] p1_smul_79014_comb;
  wire [20:0] p1_smul_79015_comb;
  wire [20:0] p1_smul_79017_comb;
  wire [20:0] p1_smul_79022_comb;
  wire [20:0] p1_smul_79024_comb;
  wire [20:0] p1_smul_79025_comb;
  wire [20:0] p1_smul_79027_comb;
  wire [20:0] p1_smul_79032_comb;
  wire [20:0] p1_smul_79034_comb;
  wire [20:0] p1_smul_79035_comb;
  wire [20:0] p1_smul_79037_comb;
  wire [20:0] p1_smul_79074_comb;
  wire [20:0] p1_smul_79075_comb;
  wire [20:0] p1_smul_79076_comb;
  wire [20:0] p1_smul_79077_comb;
  wire [20:0] p1_smul_79082_comb;
  wire [20:0] p1_smul_79083_comb;
  wire [20:0] p1_smul_79084_comb;
  wire [20:0] p1_smul_79085_comb;
  wire [20:0] p1_smul_79090_comb;
  wire [20:0] p1_smul_79091_comb;
  wire [20:0] p1_smul_79092_comb;
  wire [20:0] p1_smul_79093_comb;
  wire [20:0] p1_smul_79098_comb;
  wire [20:0] p1_smul_79099_comb;
  wire [20:0] p1_smul_79100_comb;
  wire [20:0] p1_smul_79101_comb;
  wire [20:0] p1_smul_79106_comb;
  wire [20:0] p1_smul_79107_comb;
  wire [20:0] p1_smul_79108_comb;
  wire [20:0] p1_smul_79109_comb;
  wire [20:0] p1_smul_79114_comb;
  wire [20:0] p1_smul_79115_comb;
  wire [20:0] p1_smul_79116_comb;
  wire [20:0] p1_smul_79117_comb;
  wire [20:0] p1_smul_79122_comb;
  wire [20:0] p1_smul_79123_comb;
  wire [20:0] p1_smul_79124_comb;
  wire [20:0] p1_smul_79125_comb;
  wire [20:0] p1_smul_79130_comb;
  wire [20:0] p1_smul_79131_comb;
  wire [20:0] p1_smul_79132_comb;
  wire [20:0] p1_smul_79133_comb;
  wire [20:0] p1_add_79136_comb;
  wire [19:0] p1_smul_79137_comb;
  wire [19:0] p1_smul_79138_comb;
  wire [19:0] p1_smul_79139_comb;
  wire [19:0] p1_smul_79140_comb;
  wire [20:0] p1_add_79141_comb;
  wire [20:0] p1_add_79142_comb;
  wire [19:0] p1_smul_79143_comb;
  wire [19:0] p1_smul_79144_comb;
  wire [19:0] p1_smul_79145_comb;
  wire [19:0] p1_smul_79146_comb;
  wire [20:0] p1_add_79147_comb;
  wire [20:0] p1_add_79148_comb;
  wire [19:0] p1_smul_79149_comb;
  wire [19:0] p1_smul_79150_comb;
  wire [19:0] p1_smul_79151_comb;
  wire [19:0] p1_smul_79152_comb;
  wire [20:0] p1_add_79153_comb;
  wire [20:0] p1_add_79154_comb;
  wire [19:0] p1_smul_79155_comb;
  wire [19:0] p1_smul_79156_comb;
  wire [19:0] p1_smul_79157_comb;
  wire [19:0] p1_smul_79158_comb;
  wire [20:0] p1_add_79159_comb;
  wire [20:0] p1_add_79160_comb;
  wire [19:0] p1_smul_79161_comb;
  wire [19:0] p1_smul_79162_comb;
  wire [19:0] p1_smul_79163_comb;
  wire [19:0] p1_smul_79164_comb;
  wire [20:0] p1_add_79165_comb;
  wire [20:0] p1_add_79166_comb;
  wire [19:0] p1_smul_79167_comb;
  wire [19:0] p1_smul_79168_comb;
  wire [19:0] p1_smul_79169_comb;
  wire [19:0] p1_smul_79170_comb;
  wire [20:0] p1_add_79171_comb;
  wire [20:0] p1_add_79172_comb;
  wire [19:0] p1_smul_79173_comb;
  wire [19:0] p1_smul_79174_comb;
  wire [19:0] p1_smul_79175_comb;
  wire [19:0] p1_smul_79176_comb;
  wire [20:0] p1_add_79177_comb;
  wire [20:0] p1_add_79178_comb;
  wire [19:0] p1_smul_79179_comb;
  wire [19:0] p1_smul_79180_comb;
  wire [19:0] p1_smul_79181_comb;
  wire [19:0] p1_smul_79182_comb;
  wire [20:0] p1_add_79183_comb;
  wire [19:0] p1_smul_79186_comb;
  wire [19:0] p1_smul_79187_comb;
  wire [19:0] p1_smul_79192_comb;
  wire [19:0] p1_smul_79193_comb;
  wire [19:0] p1_smul_79198_comb;
  wire [19:0] p1_smul_79199_comb;
  wire [19:0] p1_smul_79204_comb;
  wire [19:0] p1_smul_79205_comb;
  wire [19:0] p1_smul_79210_comb;
  wire [19:0] p1_smul_79211_comb;
  wire [19:0] p1_smul_79216_comb;
  wire [19:0] p1_smul_79217_comb;
  wire [19:0] p1_smul_79222_comb;
  wire [19:0] p1_smul_79223_comb;
  wire [19:0] p1_smul_79228_comb;
  wire [19:0] p1_smul_79229_comb;
  wire [19:0] p1_smul_79234_comb;
  wire [19:0] p1_smul_79235_comb;
  wire [19:0] p1_smul_79240_comb;
  wire [19:0] p1_smul_79241_comb;
  wire [19:0] p1_smul_79246_comb;
  wire [19:0] p1_smul_79247_comb;
  wire [19:0] p1_smul_79252_comb;
  wire [19:0] p1_smul_79253_comb;
  wire [19:0] p1_smul_79258_comb;
  wire [19:0] p1_smul_79259_comb;
  wire [19:0] p1_smul_79264_comb;
  wire [19:0] p1_smul_79265_comb;
  wire [19:0] p1_smul_79270_comb;
  wire [19:0] p1_smul_79271_comb;
  wire [19:0] p1_smul_79276_comb;
  wire [19:0] p1_smul_79277_comb;
  wire [19:0] p1_smul_79281_comb;
  wire [19:0] p1_smul_79283_comb;
  wire [19:0] p1_smul_79284_comb;
  wire [19:0] p1_smul_79286_comb;
  wire [19:0] p1_smul_79289_comb;
  wire [19:0] p1_smul_79291_comb;
  wire [19:0] p1_smul_79292_comb;
  wire [19:0] p1_smul_79294_comb;
  wire [19:0] p1_smul_79297_comb;
  wire [19:0] p1_smul_79299_comb;
  wire [19:0] p1_smul_79300_comb;
  wire [19:0] p1_smul_79302_comb;
  wire [19:0] p1_smul_79305_comb;
  wire [19:0] p1_smul_79307_comb;
  wire [19:0] p1_smul_79308_comb;
  wire [19:0] p1_smul_79310_comb;
  wire [19:0] p1_smul_79313_comb;
  wire [19:0] p1_smul_79315_comb;
  wire [19:0] p1_smul_79316_comb;
  wire [19:0] p1_smul_79318_comb;
  wire [19:0] p1_smul_79321_comb;
  wire [19:0] p1_smul_79323_comb;
  wire [19:0] p1_smul_79324_comb;
  wire [19:0] p1_smul_79326_comb;
  wire [19:0] p1_smul_79329_comb;
  wire [19:0] p1_smul_79331_comb;
  wire [19:0] p1_smul_79332_comb;
  wire [19:0] p1_smul_79334_comb;
  wire [19:0] p1_smul_79337_comb;
  wire [19:0] p1_smul_79339_comb;
  wire [19:0] p1_smul_79340_comb;
  wire [19:0] p1_smul_79342_comb;
  wire [19:0] p1_smul_79408_comb;
  wire [19:0] p1_smul_79410_comb;
  wire [19:0] p1_smul_79413_comb;
  wire [19:0] p1_smul_79415_comb;
  wire [19:0] p1_smul_79416_comb;
  wire [19:0] p1_smul_79418_comb;
  wire [19:0] p1_smul_79421_comb;
  wire [19:0] p1_smul_79423_comb;
  wire [19:0] p1_smul_79424_comb;
  wire [19:0] p1_smul_79426_comb;
  wire [19:0] p1_smul_79429_comb;
  wire [19:0] p1_smul_79431_comb;
  wire [19:0] p1_smul_79432_comb;
  wire [19:0] p1_smul_79434_comb;
  wire [19:0] p1_smul_79437_comb;
  wire [19:0] p1_smul_79439_comb;
  wire [19:0] p1_smul_79440_comb;
  wire [19:0] p1_smul_79442_comb;
  wire [19:0] p1_smul_79445_comb;
  wire [19:0] p1_smul_79447_comb;
  wire [19:0] p1_smul_79448_comb;
  wire [19:0] p1_smul_79450_comb;
  wire [19:0] p1_smul_79453_comb;
  wire [19:0] p1_smul_79455_comb;
  wire [19:0] p1_smul_79456_comb;
  wire [19:0] p1_smul_79458_comb;
  wire [19:0] p1_smul_79461_comb;
  wire [19:0] p1_smul_79463_comb;
  wire [19:0] p1_smul_79464_comb;
  wire [19:0] p1_smul_79466_comb;
  wire [19:0] p1_smul_79469_comb;
  wire [19:0] p1_smul_79471_comb;
  wire [19:0] p1_smul_79472_comb;
  wire [19:0] p1_smul_79475_comb;
  wire [19:0] p1_smul_79478_comb;
  wire [19:0] p1_smul_79481_comb;
  wire [19:0] p1_smul_79482_comb;
  wire [19:0] p1_smul_79485_comb;
  wire [19:0] p1_smul_79488_comb;
  wire [19:0] p1_smul_79491_comb;
  wire [19:0] p1_smul_79492_comb;
  wire [19:0] p1_smul_79495_comb;
  wire [19:0] p1_smul_79498_comb;
  wire [19:0] p1_smul_79501_comb;
  wire [19:0] p1_smul_79502_comb;
  wire [19:0] p1_smul_79505_comb;
  wire [19:0] p1_smul_79508_comb;
  wire [19:0] p1_smul_79511_comb;
  wire [19:0] p1_smul_79512_comb;
  wire [19:0] p1_smul_79515_comb;
  wire [19:0] p1_smul_79518_comb;
  wire [19:0] p1_smul_79521_comb;
  wire [19:0] p1_smul_79522_comb;
  wire [19:0] p1_smul_79525_comb;
  wire [19:0] p1_smul_79528_comb;
  wire [19:0] p1_smul_79531_comb;
  wire [19:0] p1_smul_79532_comb;
  wire [19:0] p1_smul_79535_comb;
  wire [19:0] p1_smul_79538_comb;
  wire [19:0] p1_smul_79541_comb;
  wire [19:0] p1_smul_79542_comb;
  wire [19:0] p1_smul_79545_comb;
  wire [19:0] p1_smul_79548_comb;
  wire [19:0] p1_smul_79551_comb;
  wire [19:0] p1_smul_79552_comb;
  wire [19:0] p1_smul_79553_comb;
  wire [20:0] p1_add_79554_comb;
  wire [20:0] p1_add_79555_comb;
  wire [19:0] p1_smul_79556_comb;
  wire [19:0] p1_smul_79557_comb;
  wire [19:0] p1_smul_79558_comb;
  wire [19:0] p1_smul_79559_comb;
  wire [20:0] p1_add_79560_comb;
  wire [20:0] p1_add_79561_comb;
  wire [19:0] p1_smul_79562_comb;
  wire [19:0] p1_smul_79563_comb;
  wire [19:0] p1_smul_79564_comb;
  wire [19:0] p1_smul_79565_comb;
  wire [20:0] p1_add_79566_comb;
  wire [20:0] p1_add_79567_comb;
  wire [19:0] p1_smul_79568_comb;
  wire [19:0] p1_smul_79569_comb;
  wire [19:0] p1_smul_79570_comb;
  wire [19:0] p1_smul_79571_comb;
  wire [20:0] p1_add_79572_comb;
  wire [20:0] p1_add_79573_comb;
  wire [19:0] p1_smul_79574_comb;
  wire [19:0] p1_smul_79575_comb;
  wire [19:0] p1_smul_79576_comb;
  wire [19:0] p1_smul_79577_comb;
  wire [20:0] p1_add_79578_comb;
  wire [20:0] p1_add_79579_comb;
  wire [19:0] p1_smul_79580_comb;
  wire [19:0] p1_smul_79581_comb;
  wire [19:0] p1_smul_79582_comb;
  wire [19:0] p1_smul_79583_comb;
  wire [20:0] p1_add_79584_comb;
  wire [20:0] p1_add_79585_comb;
  wire [19:0] p1_smul_79586_comb;
  wire [19:0] p1_smul_79587_comb;
  wire [19:0] p1_smul_79588_comb;
  wire [19:0] p1_smul_79589_comb;
  wire [20:0] p1_add_79590_comb;
  wire [20:0] p1_add_79591_comb;
  wire [19:0] p1_smul_79592_comb;
  wire [19:0] p1_smul_79593_comb;
  wire [19:0] p1_smul_79594_comb;
  wire [19:0] p1_smul_79595_comb;
  wire [20:0] p1_add_79596_comb;
  wire [20:0] p1_add_79597_comb;
  wire [19:0] p1_smul_79598_comb;
  wire [19:0] p1_smul_79599_comb;
  wire [19:0] p1_bit_slice_79664_comb;
  wire [19:0] p1_add_79665_comb;
  wire [19:0] p1_add_79666_comb;
  wire [19:0] p1_bit_slice_79667_comb;
  wire [19:0] p1_bit_slice_79668_comb;
  wire [19:0] p1_add_79669_comb;
  wire [19:0] p1_add_79670_comb;
  wire [19:0] p1_bit_slice_79671_comb;
  wire [19:0] p1_bit_slice_79672_comb;
  wire [19:0] p1_add_79673_comb;
  wire [19:0] p1_add_79674_comb;
  wire [19:0] p1_bit_slice_79675_comb;
  wire [19:0] p1_bit_slice_79676_comb;
  wire [19:0] p1_add_79677_comb;
  wire [19:0] p1_add_79678_comb;
  wire [19:0] p1_bit_slice_79679_comb;
  wire [19:0] p1_bit_slice_79680_comb;
  wire [19:0] p1_add_79681_comb;
  wire [19:0] p1_add_79682_comb;
  wire [19:0] p1_bit_slice_79683_comb;
  wire [19:0] p1_bit_slice_79684_comb;
  wire [19:0] p1_add_79685_comb;
  wire [19:0] p1_add_79686_comb;
  wire [19:0] p1_bit_slice_79687_comb;
  wire [19:0] p1_bit_slice_79688_comb;
  wire [19:0] p1_add_79689_comb;
  wire [19:0] p1_add_79690_comb;
  wire [19:0] p1_bit_slice_79691_comb;
  wire [19:0] p1_bit_slice_79692_comb;
  wire [19:0] p1_add_79693_comb;
  wire [19:0] p1_add_79694_comb;
  wire [19:0] p1_bit_slice_79695_comb;
  wire [18:0] p1_smul_79696_comb;
  wire [18:0] p1_smul_79699_comb;
  wire [18:0] p1_smul_79700_comb;
  wire [18:0] p1_smul_79703_comb;
  wire [18:0] p1_smul_79704_comb;
  wire [18:0] p1_smul_79707_comb;
  wire [18:0] p1_smul_79708_comb;
  wire [18:0] p1_smul_79711_comb;
  wire [18:0] p1_smul_79712_comb;
  wire [18:0] p1_smul_79715_comb;
  wire [18:0] p1_smul_79716_comb;
  wire [18:0] p1_smul_79719_comb;
  wire [18:0] p1_smul_79720_comb;
  wire [18:0] p1_smul_79723_comb;
  wire [18:0] p1_smul_79724_comb;
  wire [18:0] p1_smul_79727_comb;
  wire [18:0] p1_smul_79728_comb;
  wire [18:0] p1_smul_79731_comb;
  wire [18:0] p1_smul_79732_comb;
  wire [18:0] p1_smul_79735_comb;
  wire [18:0] p1_smul_79736_comb;
  wire [18:0] p1_smul_79739_comb;
  wire [18:0] p1_smul_79740_comb;
  wire [18:0] p1_smul_79743_comb;
  wire [18:0] p1_smul_79744_comb;
  wire [18:0] p1_smul_79747_comb;
  wire [18:0] p1_smul_79748_comb;
  wire [18:0] p1_smul_79751_comb;
  wire [18:0] p1_smul_79752_comb;
  wire [18:0] p1_smul_79755_comb;
  wire [18:0] p1_smul_79756_comb;
  wire [18:0] p1_smul_79759_comb;
  wire [19:0] p1_add_79760_comb;
  wire [19:0] p1_add_79762_comb;
  wire [19:0] p1_add_79764_comb;
  wire [19:0] p1_add_79766_comb;
  wire [19:0] p1_add_79768_comb;
  wire [19:0] p1_add_79770_comb;
  wire [19:0] p1_add_79772_comb;
  wire [19:0] p1_add_79774_comb;
  wire [19:0] p1_add_79776_comb;
  wire [19:0] p1_add_79778_comb;
  wire [19:0] p1_add_79780_comb;
  wire [19:0] p1_add_79782_comb;
  wire [19:0] p1_add_79784_comb;
  wire [19:0] p1_add_79786_comb;
  wire [19:0] p1_add_79788_comb;
  wire [19:0] p1_add_79790_comb;
  wire [19:0] p1_add_79792_comb;
  wire [19:0] p1_add_79794_comb;
  wire [19:0] p1_add_79796_comb;
  wire [19:0] p1_add_79798_comb;
  wire [19:0] p1_add_79800_comb;
  wire [19:0] p1_add_79802_comb;
  wire [19:0] p1_add_79804_comb;
  wire [19:0] p1_add_79806_comb;
  wire [19:0] p1_add_79808_comb;
  wire [19:0] p1_add_79810_comb;
  wire [19:0] p1_add_79812_comb;
  wire [19:0] p1_add_79814_comb;
  wire [19:0] p1_add_79816_comb;
  wire [19:0] p1_add_79818_comb;
  wire [19:0] p1_add_79820_comb;
  wire [19:0] p1_add_79822_comb;
  wire [20:0] p1_smul_79824_comb;
  wire [20:0] p1_smul_79825_comb;
  wire [20:0] p1_smul_79826_comb;
  wire [20:0] p1_smul_79827_comb;
  wire [20:0] p1_smul_79828_comb;
  wire [20:0] p1_smul_79829_comb;
  wire [20:0] p1_smul_79830_comb;
  wire [20:0] p1_smul_79831_comb;
  wire [20:0] p1_smul_79832_comb;
  wire [20:0] p1_smul_79833_comb;
  wire [20:0] p1_smul_79834_comb;
  wire [20:0] p1_smul_79835_comb;
  wire [20:0] p1_smul_79836_comb;
  wire [20:0] p1_smul_79837_comb;
  wire [20:0] p1_smul_79838_comb;
  wire [20:0] p1_smul_79839_comb;
  wire [20:0] p1_smul_79840_comb;
  wire [20:0] p1_smul_79841_comb;
  wire [20:0] p1_smul_79842_comb;
  wire [20:0] p1_smul_79843_comb;
  wire [20:0] p1_smul_79844_comb;
  wire [20:0] p1_smul_79845_comb;
  wire [20:0] p1_smul_79846_comb;
  wire [20:0] p1_smul_79847_comb;
  wire [20:0] p1_smul_79848_comb;
  wire [20:0] p1_smul_79849_comb;
  wire [20:0] p1_smul_79850_comb;
  wire [20:0] p1_smul_79851_comb;
  wire [20:0] p1_smul_79852_comb;
  wire [20:0] p1_smul_79853_comb;
  wire [20:0] p1_smul_79854_comb;
  wire [20:0] p1_smul_79855_comb;
  wire [20:0] p1_smul_79856_comb;
  wire [20:0] p1_smul_79857_comb;
  wire [20:0] p1_smul_79858_comb;
  wire [20:0] p1_smul_79859_comb;
  wire [20:0] p1_smul_79860_comb;
  wire [20:0] p1_smul_79861_comb;
  wire [20:0] p1_smul_79862_comb;
  wire [20:0] p1_smul_79863_comb;
  wire [20:0] p1_smul_79864_comb;
  wire [20:0] p1_smul_79865_comb;
  wire [20:0] p1_smul_79866_comb;
  wire [20:0] p1_smul_79867_comb;
  wire [20:0] p1_smul_79868_comb;
  wire [20:0] p1_smul_79869_comb;
  wire [20:0] p1_smul_79870_comb;
  wire [20:0] p1_smul_79871_comb;
  wire [20:0] p1_smul_79872_comb;
  wire [20:0] p1_smul_79873_comb;
  wire [20:0] p1_smul_79874_comb;
  wire [20:0] p1_smul_79875_comb;
  wire [20:0] p1_smul_79876_comb;
  wire [20:0] p1_smul_79877_comb;
  wire [20:0] p1_smul_79878_comb;
  wire [20:0] p1_smul_79879_comb;
  wire [20:0] p1_smul_79880_comb;
  wire [20:0] p1_smul_79881_comb;
  wire [20:0] p1_smul_79882_comb;
  wire [20:0] p1_smul_79883_comb;
  wire [20:0] p1_smul_79884_comb;
  wire [20:0] p1_smul_79885_comb;
  wire [20:0] p1_smul_79886_comb;
  wire [20:0] p1_smul_79887_comb;
  wire [19:0] p1_add_79888_comb;
  wire [19:0] p1_add_79890_comb;
  wire [19:0] p1_add_79892_comb;
  wire [19:0] p1_add_79894_comb;
  wire [19:0] p1_add_79896_comb;
  wire [19:0] p1_add_79898_comb;
  wire [19:0] p1_add_79900_comb;
  wire [19:0] p1_add_79902_comb;
  wire [19:0] p1_add_79904_comb;
  wire [19:0] p1_add_79906_comb;
  wire [19:0] p1_add_79908_comb;
  wire [19:0] p1_add_79910_comb;
  wire [19:0] p1_add_79912_comb;
  wire [19:0] p1_add_79914_comb;
  wire [19:0] p1_add_79916_comb;
  wire [19:0] p1_add_79918_comb;
  wire [19:0] p1_add_79920_comb;
  wire [19:0] p1_add_79922_comb;
  wire [19:0] p1_add_79924_comb;
  wire [19:0] p1_add_79926_comb;
  wire [19:0] p1_add_79928_comb;
  wire [19:0] p1_add_79930_comb;
  wire [19:0] p1_add_79932_comb;
  wire [19:0] p1_add_79934_comb;
  wire [19:0] p1_add_79936_comb;
  wire [19:0] p1_add_79938_comb;
  wire [19:0] p1_add_79940_comb;
  wire [19:0] p1_add_79942_comb;
  wire [19:0] p1_add_79944_comb;
  wire [19:0] p1_add_79946_comb;
  wire [19:0] p1_add_79948_comb;
  wire [19:0] p1_add_79950_comb;
  wire [18:0] p1_smul_79953_comb;
  wire [18:0] p1_smul_79955_comb;
  wire [18:0] p1_smul_79956_comb;
  wire [18:0] p1_smul_79958_comb;
  wire [18:0] p1_smul_79961_comb;
  wire [18:0] p1_smul_79963_comb;
  wire [18:0] p1_smul_79964_comb;
  wire [18:0] p1_smul_79966_comb;
  wire [18:0] p1_smul_79969_comb;
  wire [18:0] p1_smul_79971_comb;
  wire [18:0] p1_smul_79972_comb;
  wire [18:0] p1_smul_79974_comb;
  wire [18:0] p1_smul_79977_comb;
  wire [18:0] p1_smul_79979_comb;
  wire [18:0] p1_smul_79980_comb;
  wire [18:0] p1_smul_79982_comb;
  wire [18:0] p1_smul_79985_comb;
  wire [18:0] p1_smul_79987_comb;
  wire [18:0] p1_smul_79988_comb;
  wire [18:0] p1_smul_79990_comb;
  wire [18:0] p1_smul_79993_comb;
  wire [18:0] p1_smul_79995_comb;
  wire [18:0] p1_smul_79996_comb;
  wire [18:0] p1_smul_79998_comb;
  wire [18:0] p1_smul_80001_comb;
  wire [18:0] p1_smul_80003_comb;
  wire [18:0] p1_smul_80004_comb;
  wire [18:0] p1_smul_80006_comb;
  wire [18:0] p1_smul_80009_comb;
  wire [18:0] p1_smul_80011_comb;
  wire [18:0] p1_smul_80012_comb;
  wire [18:0] p1_smul_80014_comb;
  wire [19:0] p1_add_80016_comb;
  wire [19:0] p1_bit_slice_80017_comb;
  wire [19:0] p1_bit_slice_80018_comb;
  wire [19:0] p1_add_80019_comb;
  wire [19:0] p1_add_80020_comb;
  wire [19:0] p1_bit_slice_80021_comb;
  wire [19:0] p1_bit_slice_80022_comb;
  wire [19:0] p1_add_80023_comb;
  wire [19:0] p1_add_80024_comb;
  wire [19:0] p1_bit_slice_80025_comb;
  wire [19:0] p1_bit_slice_80026_comb;
  wire [19:0] p1_add_80027_comb;
  wire [19:0] p1_add_80028_comb;
  wire [19:0] p1_bit_slice_80029_comb;
  wire [19:0] p1_bit_slice_80030_comb;
  wire [19:0] p1_add_80031_comb;
  wire [19:0] p1_add_80032_comb;
  wire [19:0] p1_bit_slice_80033_comb;
  wire [19:0] p1_bit_slice_80034_comb;
  wire [19:0] p1_add_80035_comb;
  wire [19:0] p1_add_80036_comb;
  wire [19:0] p1_bit_slice_80037_comb;
  wire [19:0] p1_bit_slice_80038_comb;
  wire [19:0] p1_add_80039_comb;
  wire [19:0] p1_add_80040_comb;
  wire [19:0] p1_bit_slice_80041_comb;
  wire [19:0] p1_bit_slice_80042_comb;
  wire [19:0] p1_add_80043_comb;
  wire [19:0] p1_add_80044_comb;
  wire [19:0] p1_bit_slice_80045_comb;
  wire [19:0] p1_bit_slice_80046_comb;
  wire [19:0] p1_add_80047_comb;
  wire [12:0] p1_add_80048_comb;
  wire [12:0] p1_add_80049_comb;
  wire [12:0] p1_add_80050_comb;
  wire [12:0] p1_add_80051_comb;
  wire [12:0] p1_add_80052_comb;
  wire [12:0] p1_add_80053_comb;
  wire [12:0] p1_add_80054_comb;
  wire [12:0] p1_add_80055_comb;
  wire [12:0] p1_add_80056_comb;
  wire [12:0] p1_add_80057_comb;
  wire [12:0] p1_add_80058_comb;
  wire [12:0] p1_add_80059_comb;
  wire [12:0] p1_add_80060_comb;
  wire [12:0] p1_add_80061_comb;
  wire [12:0] p1_add_80062_comb;
  wire [12:0] p1_add_80063_comb;
  wire [12:0] p1_add_80064_comb;
  wire [12:0] p1_add_80065_comb;
  wire [12:0] p1_add_80066_comb;
  wire [12:0] p1_add_80067_comb;
  wire [12:0] p1_add_80068_comb;
  wire [12:0] p1_add_80069_comb;
  wire [12:0] p1_add_80070_comb;
  wire [12:0] p1_add_80071_comb;
  wire [12:0] p1_add_80072_comb;
  wire [12:0] p1_add_80073_comb;
  wire [12:0] p1_add_80074_comb;
  wire [12:0] p1_add_80075_comb;
  wire [12:0] p1_add_80076_comb;
  wire [12:0] p1_add_80077_comb;
  wire [12:0] p1_add_80078_comb;
  wire [12:0] p1_add_80079_comb;
  wire [18:0] p1_add_80112_comb;
  wire [18:0] p1_add_80114_comb;
  wire [18:0] p1_add_80116_comb;
  wire [18:0] p1_add_80118_comb;
  wire [18:0] p1_add_80120_comb;
  wire [18:0] p1_add_80122_comb;
  wire [18:0] p1_add_80124_comb;
  wire [18:0] p1_add_80126_comb;
  wire [18:0] p1_add_80128_comb;
  wire [18:0] p1_add_80130_comb;
  wire [18:0] p1_add_80132_comb;
  wire [18:0] p1_add_80134_comb;
  wire [18:0] p1_add_80136_comb;
  wire [18:0] p1_add_80138_comb;
  wire [18:0] p1_add_80140_comb;
  wire [18:0] p1_add_80142_comb;
  wire [18:0] p1_add_80144_comb;
  wire [18:0] p1_add_80146_comb;
  wire [18:0] p1_add_80148_comb;
  wire [18:0] p1_add_80150_comb;
  wire [18:0] p1_add_80152_comb;
  wire [18:0] p1_add_80154_comb;
  wire [18:0] p1_add_80156_comb;
  wire [18:0] p1_add_80158_comb;
  wire [18:0] p1_add_80160_comb;
  wire [18:0] p1_add_80162_comb;
  wire [18:0] p1_add_80164_comb;
  wire [18:0] p1_add_80166_comb;
  wire [18:0] p1_add_80168_comb;
  wire [18:0] p1_add_80170_comb;
  wire [18:0] p1_add_80172_comb;
  wire [18:0] p1_add_80174_comb;
  wire [20:0] p1_concat_80176_comb;
  wire [20:0] p1_concat_80177_comb;
  wire [20:0] p1_concat_80178_comb;
  wire [20:0] p1_concat_80179_comb;
  wire [20:0] p1_concat_80180_comb;
  wire [20:0] p1_concat_80181_comb;
  wire [20:0] p1_concat_80182_comb;
  wire [20:0] p1_concat_80183_comb;
  wire [20:0] p1_concat_80184_comb;
  wire [20:0] p1_concat_80185_comb;
  wire [20:0] p1_concat_80186_comb;
  wire [20:0] p1_concat_80187_comb;
  wire [20:0] p1_concat_80188_comb;
  wire [20:0] p1_concat_80189_comb;
  wire [20:0] p1_concat_80190_comb;
  wire [20:0] p1_concat_80191_comb;
  wire [20:0] p1_concat_80192_comb;
  wire [20:0] p1_concat_80193_comb;
  wire [20:0] p1_concat_80194_comb;
  wire [20:0] p1_concat_80195_comb;
  wire [20:0] p1_concat_80196_comb;
  wire [20:0] p1_concat_80197_comb;
  wire [20:0] p1_concat_80198_comb;
  wire [20:0] p1_concat_80199_comb;
  wire [20:0] p1_concat_80200_comb;
  wire [20:0] p1_concat_80201_comb;
  wire [20:0] p1_concat_80202_comb;
  wire [20:0] p1_concat_80203_comb;
  wire [20:0] p1_concat_80204_comb;
  wire [20:0] p1_concat_80205_comb;
  wire [20:0] p1_concat_80206_comb;
  wire [20:0] p1_concat_80207_comb;
  wire [20:0] p1_add_80208_comb;
  wire [20:0] p1_add_80209_comb;
  wire [20:0] p1_add_80210_comb;
  wire [20:0] p1_add_80211_comb;
  wire [20:0] p1_add_80212_comb;
  wire [20:0] p1_add_80213_comb;
  wire [20:0] p1_add_80214_comb;
  wire [20:0] p1_add_80215_comb;
  wire [20:0] p1_add_80216_comb;
  wire [20:0] p1_add_80217_comb;
  wire [20:0] p1_add_80218_comb;
  wire [20:0] p1_add_80219_comb;
  wire [20:0] p1_add_80220_comb;
  wire [20:0] p1_add_80221_comb;
  wire [20:0] p1_add_80222_comb;
  wire [20:0] p1_add_80223_comb;
  wire [20:0] p1_add_80224_comb;
  wire [20:0] p1_add_80225_comb;
  wire [20:0] p1_add_80226_comb;
  wire [20:0] p1_add_80227_comb;
  wire [20:0] p1_add_80228_comb;
  wire [20:0] p1_add_80229_comb;
  wire [20:0] p1_add_80230_comb;
  wire [20:0] p1_add_80231_comb;
  wire [20:0] p1_add_80232_comb;
  wire [20:0] p1_add_80233_comb;
  wire [20:0] p1_add_80234_comb;
  wire [20:0] p1_add_80235_comb;
  wire [20:0] p1_add_80236_comb;
  wire [20:0] p1_add_80237_comb;
  wire [20:0] p1_add_80238_comb;
  wire [20:0] p1_add_80239_comb;
  wire [20:0] p1_concat_80240_comb;
  wire [20:0] p1_concat_80241_comb;
  wire [20:0] p1_concat_80242_comb;
  wire [20:0] p1_concat_80243_comb;
  wire [20:0] p1_concat_80244_comb;
  wire [20:0] p1_concat_80245_comb;
  wire [20:0] p1_concat_80246_comb;
  wire [20:0] p1_concat_80247_comb;
  wire [20:0] p1_concat_80248_comb;
  wire [20:0] p1_concat_80249_comb;
  wire [20:0] p1_concat_80250_comb;
  wire [20:0] p1_concat_80251_comb;
  wire [20:0] p1_concat_80252_comb;
  wire [20:0] p1_concat_80253_comb;
  wire [20:0] p1_concat_80254_comb;
  wire [20:0] p1_concat_80255_comb;
  wire [20:0] p1_concat_80256_comb;
  wire [20:0] p1_concat_80257_comb;
  wire [20:0] p1_concat_80258_comb;
  wire [20:0] p1_concat_80259_comb;
  wire [20:0] p1_concat_80260_comb;
  wire [20:0] p1_concat_80261_comb;
  wire [20:0] p1_concat_80262_comb;
  wire [20:0] p1_concat_80263_comb;
  wire [20:0] p1_concat_80264_comb;
  wire [20:0] p1_concat_80265_comb;
  wire [20:0] p1_concat_80266_comb;
  wire [20:0] p1_concat_80267_comb;
  wire [20:0] p1_concat_80268_comb;
  wire [20:0] p1_concat_80269_comb;
  wire [20:0] p1_concat_80270_comb;
  wire [20:0] p1_concat_80271_comb;
  wire [18:0] p1_add_80272_comb;
  wire [18:0] p1_add_80274_comb;
  wire [18:0] p1_add_80276_comb;
  wire [18:0] p1_add_80278_comb;
  wire [18:0] p1_add_80280_comb;
  wire [18:0] p1_add_80282_comb;
  wire [18:0] p1_add_80284_comb;
  wire [18:0] p1_add_80286_comb;
  wire [18:0] p1_add_80288_comb;
  wire [18:0] p1_add_80290_comb;
  wire [18:0] p1_add_80292_comb;
  wire [18:0] p1_add_80294_comb;
  wire [18:0] p1_add_80296_comb;
  wire [18:0] p1_add_80298_comb;
  wire [18:0] p1_add_80300_comb;
  wire [18:0] p1_add_80302_comb;
  wire [18:0] p1_add_80304_comb;
  wire [18:0] p1_add_80306_comb;
  wire [18:0] p1_add_80308_comb;
  wire [18:0] p1_add_80310_comb;
  wire [18:0] p1_add_80312_comb;
  wire [18:0] p1_add_80314_comb;
  wire [18:0] p1_add_80316_comb;
  wire [18:0] p1_add_80318_comb;
  wire [18:0] p1_add_80320_comb;
  wire [18:0] p1_add_80322_comb;
  wire [18:0] p1_add_80324_comb;
  wire [18:0] p1_add_80326_comb;
  wire [18:0] p1_add_80328_comb;
  wire [18:0] p1_add_80330_comb;
  wire [18:0] p1_add_80332_comb;
  wire [18:0] p1_add_80334_comb;
  wire [23:0] p1_add_80400_comb;
  wire [23:0] p1_add_80402_comb;
  wire [23:0] p1_add_80404_comb;
  wire [23:0] p1_add_80406_comb;
  wire [23:0] p1_add_80408_comb;
  wire [23:0] p1_add_80410_comb;
  wire [23:0] p1_add_80412_comb;
  wire [23:0] p1_add_80414_comb;
  wire [23:0] p1_add_80416_comb;
  wire [23:0] p1_add_80418_comb;
  wire [23:0] p1_add_80420_comb;
  wire [23:0] p1_add_80422_comb;
  wire [23:0] p1_add_80424_comb;
  wire [23:0] p1_add_80426_comb;
  wire [23:0] p1_add_80428_comb;
  wire [23:0] p1_add_80430_comb;
  wire [19:0] p1_concat_80432_comb;
  wire [19:0] p1_concat_80433_comb;
  wire [19:0] p1_concat_80434_comb;
  wire [19:0] p1_concat_80435_comb;
  wire [19:0] p1_concat_80436_comb;
  wire [19:0] p1_concat_80437_comb;
  wire [19:0] p1_concat_80438_comb;
  wire [19:0] p1_concat_80439_comb;
  wire [19:0] p1_concat_80440_comb;
  wire [19:0] p1_concat_80441_comb;
  wire [19:0] p1_concat_80442_comb;
  wire [19:0] p1_concat_80443_comb;
  wire [19:0] p1_concat_80444_comb;
  wire [19:0] p1_concat_80445_comb;
  wire [19:0] p1_concat_80446_comb;
  wire [19:0] p1_concat_80447_comb;
  wire [19:0] p1_concat_80448_comb;
  wire [19:0] p1_concat_80449_comb;
  wire [19:0] p1_concat_80450_comb;
  wire [19:0] p1_concat_80451_comb;
  wire [19:0] p1_concat_80452_comb;
  wire [19:0] p1_concat_80453_comb;
  wire [19:0] p1_concat_80454_comb;
  wire [19:0] p1_concat_80455_comb;
  wire [19:0] p1_concat_80456_comb;
  wire [19:0] p1_concat_80457_comb;
  wire [19:0] p1_concat_80458_comb;
  wire [19:0] p1_concat_80459_comb;
  wire [19:0] p1_concat_80460_comb;
  wire [19:0] p1_concat_80461_comb;
  wire [19:0] p1_concat_80462_comb;
  wire [19:0] p1_concat_80463_comb;
  wire [24:0] p1_sum__1572_comb;
  wire [24:0] p1_sum__1573_comb;
  wire [24:0] p1_sum__1574_comb;
  wire [24:0] p1_sum__1575_comb;
  wire [24:0] p1_sum__1544_comb;
  wire [24:0] p1_sum__1545_comb;
  wire [24:0] p1_sum__1546_comb;
  wire [24:0] p1_sum__1547_comb;
  wire [24:0] p1_sum__1516_comb;
  wire [24:0] p1_sum__1517_comb;
  wire [24:0] p1_sum__1518_comb;
  wire [24:0] p1_sum__1519_comb;
  wire [24:0] p1_sum__1488_comb;
  wire [24:0] p1_sum__1489_comb;
  wire [24:0] p1_sum__1490_comb;
  wire [24:0] p1_sum__1491_comb;
  wire [24:0] p1_sum__1460_comb;
  wire [24:0] p1_sum__1461_comb;
  wire [24:0] p1_sum__1462_comb;
  wire [24:0] p1_sum__1463_comb;
  wire [24:0] p1_sum__1432_comb;
  wire [24:0] p1_sum__1433_comb;
  wire [24:0] p1_sum__1434_comb;
  wire [24:0] p1_sum__1435_comb;
  wire [24:0] p1_sum__1404_comb;
  wire [24:0] p1_sum__1405_comb;
  wire [24:0] p1_sum__1406_comb;
  wire [24:0] p1_sum__1407_comb;
  wire [24:0] p1_sum__1376_comb;
  wire [24:0] p1_sum__1377_comb;
  wire [24:0] p1_sum__1378_comb;
  wire [24:0] p1_sum__1379_comb;
  wire [24:0] p1_sum__1568_comb;
  wire [24:0] p1_sum__1569_comb;
  wire [24:0] p1_sum__1570_comb;
  wire [24:0] p1_sum__1571_comb;
  wire [24:0] p1_sum__1540_comb;
  wire [24:0] p1_sum__1541_comb;
  wire [24:0] p1_sum__1542_comb;
  wire [24:0] p1_sum__1543_comb;
  wire [24:0] p1_sum__1512_comb;
  wire [24:0] p1_sum__1513_comb;
  wire [24:0] p1_sum__1514_comb;
  wire [24:0] p1_sum__1515_comb;
  wire [24:0] p1_sum__1484_comb;
  wire [24:0] p1_sum__1485_comb;
  wire [24:0] p1_sum__1486_comb;
  wire [24:0] p1_sum__1487_comb;
  wire [24:0] p1_sum__1456_comb;
  wire [24:0] p1_sum__1457_comb;
  wire [24:0] p1_sum__1458_comb;
  wire [24:0] p1_sum__1459_comb;
  wire [24:0] p1_sum__1428_comb;
  wire [24:0] p1_sum__1429_comb;
  wire [24:0] p1_sum__1430_comb;
  wire [24:0] p1_sum__1431_comb;
  wire [24:0] p1_sum__1400_comb;
  wire [24:0] p1_sum__1401_comb;
  wire [24:0] p1_sum__1402_comb;
  wire [24:0] p1_sum__1403_comb;
  wire [24:0] p1_sum__1372_comb;
  wire [24:0] p1_sum__1373_comb;
  wire [24:0] p1_sum__1374_comb;
  wire [24:0] p1_sum__1375_comb;
  wire [24:0] p1_sum__1564_comb;
  wire [24:0] p1_sum__1565_comb;
  wire [24:0] p1_sum__1566_comb;
  wire [24:0] p1_sum__1567_comb;
  wire [24:0] p1_sum__1536_comb;
  wire [24:0] p1_sum__1537_comb;
  wire [24:0] p1_sum__1538_comb;
  wire [24:0] p1_sum__1539_comb;
  wire [24:0] p1_sum__1508_comb;
  wire [24:0] p1_sum__1509_comb;
  wire [24:0] p1_sum__1510_comb;
  wire [24:0] p1_sum__1511_comb;
  wire [24:0] p1_sum__1480_comb;
  wire [24:0] p1_sum__1481_comb;
  wire [24:0] p1_sum__1482_comb;
  wire [24:0] p1_sum__1483_comb;
  wire [24:0] p1_sum__1452_comb;
  wire [24:0] p1_sum__1453_comb;
  wire [24:0] p1_sum__1454_comb;
  wire [24:0] p1_sum__1455_comb;
  wire [24:0] p1_sum__1424_comb;
  wire [24:0] p1_sum__1425_comb;
  wire [24:0] p1_sum__1426_comb;
  wire [24:0] p1_sum__1427_comb;
  wire [24:0] p1_sum__1396_comb;
  wire [24:0] p1_sum__1397_comb;
  wire [24:0] p1_sum__1398_comb;
  wire [24:0] p1_sum__1399_comb;
  wire [24:0] p1_sum__1368_comb;
  wire [24:0] p1_sum__1369_comb;
  wire [24:0] p1_sum__1370_comb;
  wire [24:0] p1_sum__1371_comb;
  wire [19:0] p1_concat_80560_comb;
  wire [19:0] p1_concat_80561_comb;
  wire [19:0] p1_concat_80562_comb;
  wire [19:0] p1_concat_80563_comb;
  wire [19:0] p1_concat_80564_comb;
  wire [19:0] p1_concat_80565_comb;
  wire [19:0] p1_concat_80566_comb;
  wire [19:0] p1_concat_80567_comb;
  wire [19:0] p1_concat_80568_comb;
  wire [19:0] p1_concat_80569_comb;
  wire [19:0] p1_concat_80570_comb;
  wire [19:0] p1_concat_80571_comb;
  wire [19:0] p1_concat_80572_comb;
  wire [19:0] p1_concat_80573_comb;
  wire [19:0] p1_concat_80574_comb;
  wire [19:0] p1_concat_80575_comb;
  wire [19:0] p1_concat_80576_comb;
  wire [19:0] p1_concat_80577_comb;
  wire [19:0] p1_concat_80578_comb;
  wire [19:0] p1_concat_80579_comb;
  wire [19:0] p1_concat_80580_comb;
  wire [19:0] p1_concat_80581_comb;
  wire [19:0] p1_concat_80582_comb;
  wire [19:0] p1_concat_80583_comb;
  wire [19:0] p1_concat_80584_comb;
  wire [19:0] p1_concat_80585_comb;
  wire [19:0] p1_concat_80586_comb;
  wire [19:0] p1_concat_80587_comb;
  wire [19:0] p1_concat_80588_comb;
  wire [19:0] p1_concat_80589_comb;
  wire [19:0] p1_concat_80590_comb;
  wire [19:0] p1_concat_80591_comb;
  wire [23:0] p1_add_80592_comb;
  wire [23:0] p1_add_80594_comb;
  wire [23:0] p1_add_80596_comb;
  wire [23:0] p1_add_80598_comb;
  wire [23:0] p1_add_80600_comb;
  wire [23:0] p1_add_80602_comb;
  wire [23:0] p1_add_80604_comb;
  wire [23:0] p1_add_80606_comb;
  wire [23:0] p1_add_80608_comb;
  wire [23:0] p1_add_80610_comb;
  wire [23:0] p1_add_80612_comb;
  wire [23:0] p1_add_80614_comb;
  wire [23:0] p1_add_80616_comb;
  wire [23:0] p1_add_80618_comb;
  wire [23:0] p1_add_80620_comb;
  wire [23:0] p1_add_80622_comb;
  wire [23:0] p1_add_80624_comb;
  wire [23:0] p1_add_80625_comb;
  wire [23:0] p1_add_80626_comb;
  wire [23:0] p1_add_80627_comb;
  wire [23:0] p1_add_80628_comb;
  wire [23:0] p1_add_80629_comb;
  wire [23:0] p1_add_80630_comb;
  wire [23:0] p1_add_80631_comb;
  wire [23:0] p1_add_80632_comb;
  wire [23:0] p1_add_80633_comb;
  wire [23:0] p1_add_80634_comb;
  wire [23:0] p1_add_80635_comb;
  wire [23:0] p1_add_80636_comb;
  wire [23:0] p1_add_80637_comb;
  wire [23:0] p1_add_80638_comb;
  wire [23:0] p1_add_80639_comb;
  wire [24:0] p1_sum__1246_comb;
  wire [24:0] p1_sum__1247_comb;
  wire [24:0] p1_sum__1232_comb;
  wire [24:0] p1_sum__1233_comb;
  wire [24:0] p1_sum__1218_comb;
  wire [24:0] p1_sum__1219_comb;
  wire [24:0] p1_sum__1204_comb;
  wire [24:0] p1_sum__1205_comb;
  wire [24:0] p1_sum__1190_comb;
  wire [24:0] p1_sum__1191_comb;
  wire [24:0] p1_sum__1176_comb;
  wire [24:0] p1_sum__1177_comb;
  wire [24:0] p1_sum__1162_comb;
  wire [24:0] p1_sum__1163_comb;
  wire [24:0] p1_sum__1148_comb;
  wire [24:0] p1_sum__1149_comb;
  wire [24:0] p1_sum__1242_comb;
  wire [24:0] p1_sum__1243_comb;
  wire [24:0] p1_sum__1228_comb;
  wire [24:0] p1_sum__1229_comb;
  wire [24:0] p1_sum__1214_comb;
  wire [24:0] p1_sum__1215_comb;
  wire [24:0] p1_sum__1200_comb;
  wire [24:0] p1_sum__1201_comb;
  wire [24:0] p1_sum__1186_comb;
  wire [24:0] p1_sum__1187_comb;
  wire [24:0] p1_sum__1172_comb;
  wire [24:0] p1_sum__1173_comb;
  wire [24:0] p1_sum__1158_comb;
  wire [24:0] p1_sum__1159_comb;
  wire [24:0] p1_sum__1144_comb;
  wire [24:0] p1_sum__1145_comb;
  wire [24:0] p1_sum__1240_comb;
  wire [24:0] p1_sum__1241_comb;
  wire [24:0] p1_sum__1226_comb;
  wire [24:0] p1_sum__1227_comb;
  wire [24:0] p1_sum__1212_comb;
  wire [24:0] p1_sum__1213_comb;
  wire [24:0] p1_sum__1198_comb;
  wire [24:0] p1_sum__1199_comb;
  wire [24:0] p1_sum__1184_comb;
  wire [24:0] p1_sum__1185_comb;
  wire [24:0] p1_sum__1170_comb;
  wire [24:0] p1_sum__1171_comb;
  wire [24:0] p1_sum__1156_comb;
  wire [24:0] p1_sum__1157_comb;
  wire [24:0] p1_sum__1142_comb;
  wire [24:0] p1_sum__1143_comb;
  wire [24:0] p1_sum__1238_comb;
  wire [24:0] p1_sum__1239_comb;
  wire [24:0] p1_sum__1224_comb;
  wire [24:0] p1_sum__1225_comb;
  wire [24:0] p1_sum__1210_comb;
  wire [24:0] p1_sum__1211_comb;
  wire [24:0] p1_sum__1196_comb;
  wire [24:0] p1_sum__1197_comb;
  wire [24:0] p1_sum__1182_comb;
  wire [24:0] p1_sum__1183_comb;
  wire [24:0] p1_sum__1168_comb;
  wire [24:0] p1_sum__1169_comb;
  wire [24:0] p1_sum__1154_comb;
  wire [24:0] p1_sum__1155_comb;
  wire [24:0] p1_sum__1140_comb;
  wire [24:0] p1_sum__1141_comb;
  wire [24:0] p1_sum__1234_comb;
  wire [24:0] p1_sum__1235_comb;
  wire [24:0] p1_sum__1220_comb;
  wire [24:0] p1_sum__1221_comb;
  wire [24:0] p1_sum__1206_comb;
  wire [24:0] p1_sum__1207_comb;
  wire [24:0] p1_sum__1192_comb;
  wire [24:0] p1_sum__1193_comb;
  wire [24:0] p1_sum__1178_comb;
  wire [24:0] p1_sum__1179_comb;
  wire [24:0] p1_sum__1164_comb;
  wire [24:0] p1_sum__1165_comb;
  wire [24:0] p1_sum__1150_comb;
  wire [24:0] p1_sum__1151_comb;
  wire [24:0] p1_sum__1136_comb;
  wire [24:0] p1_sum__1137_comb;
  wire [23:0] p1_add_80784_comb;
  wire [23:0] p1_add_80786_comb;
  wire [23:0] p1_add_80788_comb;
  wire [23:0] p1_add_80790_comb;
  wire [23:0] p1_add_80792_comb;
  wire [23:0] p1_add_80794_comb;
  wire [23:0] p1_add_80796_comb;
  wire [23:0] p1_add_80798_comb;
  wire [24:0] p1_sum__1079_comb;
  wire [24:0] p1_sum__1072_comb;
  wire [24:0] p1_sum__1065_comb;
  wire [24:0] p1_sum__1058_comb;
  wire [24:0] p1_sum__1051_comb;
  wire [24:0] p1_sum__1044_comb;
  wire [24:0] p1_sum__1037_comb;
  wire [24:0] p1_sum__1030_comb;
  wire [23:0] p1_add_80816_comb;
  wire [23:0] p1_add_80817_comb;
  wire [23:0] p1_add_80818_comb;
  wire [23:0] p1_add_80819_comb;
  wire [23:0] p1_add_80820_comb;
  wire [23:0] p1_add_80821_comb;
  wire [23:0] p1_add_80822_comb;
  wire [23:0] p1_add_80823_comb;
  wire [23:0] p1_add_80824_comb;
  wire [23:0] p1_add_80825_comb;
  wire [23:0] p1_add_80826_comb;
  wire [23:0] p1_add_80827_comb;
  wire [23:0] p1_add_80828_comb;
  wire [23:0] p1_add_80829_comb;
  wire [23:0] p1_add_80830_comb;
  wire [23:0] p1_add_80831_comb;
  wire [24:0] p1_sum__1077_comb;
  wire [24:0] p1_sum__1070_comb;
  wire [24:0] p1_sum__1063_comb;
  wire [24:0] p1_sum__1056_comb;
  wire [24:0] p1_sum__1049_comb;
  wire [24:0] p1_sum__1042_comb;
  wire [24:0] p1_sum__1035_comb;
  wire [24:0] p1_sum__1028_comb;
  wire [24:0] p1_sum__1076_comb;
  wire [24:0] p1_sum__1069_comb;
  wire [24:0] p1_sum__1062_comb;
  wire [24:0] p1_sum__1055_comb;
  wire [24:0] p1_sum__1048_comb;
  wire [24:0] p1_sum__1041_comb;
  wire [24:0] p1_sum__1034_comb;
  wire [24:0] p1_sum__1027_comb;
  wire [24:0] p1_sum__1075_comb;
  wire [24:0] p1_sum__1068_comb;
  wire [24:0] p1_sum__1061_comb;
  wire [24:0] p1_sum__1054_comb;
  wire [24:0] p1_sum__1047_comb;
  wire [24:0] p1_sum__1040_comb;
  wire [24:0] p1_sum__1033_comb;
  wire [24:0] p1_sum__1026_comb;
  wire [23:0] p1_add_80880_comb;
  wire [23:0] p1_add_80881_comb;
  wire [23:0] p1_add_80882_comb;
  wire [23:0] p1_add_80883_comb;
  wire [23:0] p1_add_80884_comb;
  wire [23:0] p1_add_80885_comb;
  wire [23:0] p1_add_80886_comb;
  wire [23:0] p1_add_80887_comb;
  wire [23:0] p1_add_80888_comb;
  wire [23:0] p1_add_80889_comb;
  wire [23:0] p1_add_80890_comb;
  wire [23:0] p1_add_80891_comb;
  wire [23:0] p1_add_80892_comb;
  wire [23:0] p1_add_80893_comb;
  wire [23:0] p1_add_80894_comb;
  wire [23:0] p1_add_80895_comb;
  wire [24:0] p1_sum__1073_comb;
  wire [24:0] p1_sum__1066_comb;
  wire [24:0] p1_sum__1059_comb;
  wire [24:0] p1_sum__1052_comb;
  wire [24:0] p1_sum__1045_comb;
  wire [24:0] p1_sum__1038_comb;
  wire [24:0] p1_sum__1031_comb;
  wire [24:0] p1_sum__1024_comb;
  wire [23:0] p1_umul_28632_NarrowedMult__comb;
  wire [23:0] p1_umul_28634_NarrowedMult__comb;
  wire [23:0] p1_umul_28636_NarrowedMult__comb;
  wire [23:0] p1_umul_28638_NarrowedMult__comb;
  wire [23:0] p1_umul_28640_NarrowedMult__comb;
  wire [23:0] p1_umul_28642_NarrowedMult__comb;
  wire [23:0] p1_umul_28644_NarrowedMult__comb;
  wire [23:0] p1_umul_28646_NarrowedMult__comb;
  wire [24:0] p1_add_80920_comb;
  wire [24:0] p1_add_80921_comb;
  wire [24:0] p1_add_80922_comb;
  wire [24:0] p1_add_80923_comb;
  wire [24:0] p1_add_80924_comb;
  wire [24:0] p1_add_80925_comb;
  wire [24:0] p1_add_80926_comb;
  wire [24:0] p1_add_80927_comb;
  wire [23:0] p1_add_80928_comb;
  wire [23:0] p1_add_80929_comb;
  wire [23:0] p1_add_80930_comb;
  wire [23:0] p1_add_80931_comb;
  wire [23:0] p1_add_80932_comb;
  wire [23:0] p1_add_80933_comb;
  wire [23:0] p1_add_80934_comb;
  wire [23:0] p1_add_80935_comb;
  wire [24:0] p1_add_80936_comb;
  wire [24:0] p1_add_80937_comb;
  wire [24:0] p1_add_80938_comb;
  wire [24:0] p1_add_80939_comb;
  wire [24:0] p1_add_80940_comb;
  wire [24:0] p1_add_80941_comb;
  wire [24:0] p1_add_80942_comb;
  wire [24:0] p1_add_80943_comb;
  wire [24:0] p1_add_80944_comb;
  wire [24:0] p1_add_80945_comb;
  wire [24:0] p1_add_80946_comb;
  wire [24:0] p1_add_80947_comb;
  wire [24:0] p1_add_80948_comb;
  wire [24:0] p1_add_80949_comb;
  wire [24:0] p1_add_80950_comb;
  wire [24:0] p1_add_80951_comb;
  wire [24:0] p1_add_80952_comb;
  wire [24:0] p1_add_80953_comb;
  wire [24:0] p1_add_80954_comb;
  wire [24:0] p1_add_80955_comb;
  wire [24:0] p1_add_80956_comb;
  wire [24:0] p1_add_80957_comb;
  wire [24:0] p1_add_80958_comb;
  wire [24:0] p1_add_80959_comb;
  wire [23:0] p1_add_80960_comb;
  wire [23:0] p1_add_80961_comb;
  wire [23:0] p1_add_80962_comb;
  wire [23:0] p1_add_80963_comb;
  wire [23:0] p1_add_80964_comb;
  wire [23:0] p1_add_80965_comb;
  wire [23:0] p1_add_80966_comb;
  wire [23:0] p1_add_80967_comb;
  wire [24:0] p1_add_80968_comb;
  wire [24:0] p1_add_80969_comb;
  wire [24:0] p1_add_80970_comb;
  wire [24:0] p1_add_80971_comb;
  wire [24:0] p1_add_80972_comb;
  wire [24:0] p1_add_80973_comb;
  wire [24:0] p1_add_80974_comb;
  wire [24:0] p1_add_80975_comb;
  wire [16:0] p1_bit_slice_80976_comb;
  wire [16:0] p1_bit_slice_80977_comb;
  wire [16:0] p1_bit_slice_80978_comb;
  wire [16:0] p1_bit_slice_80979_comb;
  wire [16:0] p1_bit_slice_80980_comb;
  wire [16:0] p1_bit_slice_80981_comb;
  wire [16:0] p1_bit_slice_80982_comb;
  wire [16:0] p1_bit_slice_80983_comb;
  wire [16:0] p1_bit_slice_80984_comb;
  wire [16:0] p1_bit_slice_80985_comb;
  wire [16:0] p1_bit_slice_80986_comb;
  wire [16:0] p1_bit_slice_80987_comb;
  wire [16:0] p1_bit_slice_80988_comb;
  wire [16:0] p1_bit_slice_80989_comb;
  wire [16:0] p1_bit_slice_80990_comb;
  wire [16:0] p1_bit_slice_80991_comb;
  wire [16:0] p1_bit_slice_80992_comb;
  wire [16:0] p1_bit_slice_80993_comb;
  wire [16:0] p1_bit_slice_80994_comb;
  wire [16:0] p1_bit_slice_80995_comb;
  wire [16:0] p1_bit_slice_80996_comb;
  wire [16:0] p1_bit_slice_80997_comb;
  wire [16:0] p1_bit_slice_80998_comb;
  wire [16:0] p1_bit_slice_80999_comb;
  wire [16:0] p1_bit_slice_81000_comb;
  wire [16:0] p1_bit_slice_81001_comb;
  wire [16:0] p1_bit_slice_81002_comb;
  wire [16:0] p1_bit_slice_81003_comb;
  wire [16:0] p1_bit_slice_81004_comb;
  wire [16:0] p1_bit_slice_81005_comb;
  wire [16:0] p1_bit_slice_81006_comb;
  wire [16:0] p1_bit_slice_81007_comb;
  wire [16:0] p1_bit_slice_81008_comb;
  wire [16:0] p1_bit_slice_81009_comb;
  wire [16:0] p1_bit_slice_81010_comb;
  wire [16:0] p1_bit_slice_81011_comb;
  wire [16:0] p1_bit_slice_81012_comb;
  wire [16:0] p1_bit_slice_81013_comb;
  wire [16:0] p1_bit_slice_81014_comb;
  wire [16:0] p1_bit_slice_81015_comb;
  wire [16:0] p1_bit_slice_81016_comb;
  wire [16:0] p1_bit_slice_81017_comb;
  wire [16:0] p1_bit_slice_81018_comb;
  wire [16:0] p1_bit_slice_81019_comb;
  wire [16:0] p1_bit_slice_81020_comb;
  wire [16:0] p1_bit_slice_81021_comb;
  wire [16:0] p1_bit_slice_81022_comb;
  wire [16:0] p1_bit_slice_81023_comb;
  wire [16:0] p1_bit_slice_81024_comb;
  wire [16:0] p1_bit_slice_81025_comb;
  wire [16:0] p1_bit_slice_81026_comb;
  wire [16:0] p1_bit_slice_81027_comb;
  wire [16:0] p1_bit_slice_81028_comb;
  wire [16:0] p1_bit_slice_81029_comb;
  wire [16:0] p1_bit_slice_81030_comb;
  wire [16:0] p1_bit_slice_81031_comb;
  wire [16:0] p1_bit_slice_81032_comb;
  wire [16:0] p1_bit_slice_81033_comb;
  wire [16:0] p1_bit_slice_81034_comb;
  wire [16:0] p1_bit_slice_81035_comb;
  wire [16:0] p1_bit_slice_81036_comb;
  wire [16:0] p1_bit_slice_81037_comb;
  wire [16:0] p1_bit_slice_81038_comb;
  wire [16:0] p1_bit_slice_81039_comb;
  wire [17:0] p1_add_81168_comb;
  wire [17:0] p1_add_81169_comb;
  wire [17:0] p1_add_81170_comb;
  wire [17:0] p1_add_81171_comb;
  wire [17:0] p1_add_81172_comb;
  wire [17:0] p1_add_81173_comb;
  wire [17:0] p1_add_81174_comb;
  wire [17:0] p1_add_81175_comb;
  wire [17:0] p1_add_81176_comb;
  wire [17:0] p1_add_81177_comb;
  wire [17:0] p1_add_81178_comb;
  wire [17:0] p1_add_81179_comb;
  wire [17:0] p1_add_81180_comb;
  wire [17:0] p1_add_81181_comb;
  wire [17:0] p1_add_81182_comb;
  wire [17:0] p1_add_81183_comb;
  wire [17:0] p1_add_81184_comb;
  wire [17:0] p1_add_81185_comb;
  wire [17:0] p1_add_81186_comb;
  wire [17:0] p1_add_81187_comb;
  wire [17:0] p1_add_81188_comb;
  wire [17:0] p1_add_81189_comb;
  wire [17:0] p1_add_81190_comb;
  wire [17:0] p1_add_81191_comb;
  wire [17:0] p1_add_81192_comb;
  wire [17:0] p1_add_81193_comb;
  wire [17:0] p1_add_81194_comb;
  wire [17:0] p1_add_81195_comb;
  wire [17:0] p1_add_81196_comb;
  wire [17:0] p1_add_81197_comb;
  wire [17:0] p1_add_81198_comb;
  wire [17:0] p1_add_81199_comb;
  wire [17:0] p1_add_81200_comb;
  wire [17:0] p1_add_81201_comb;
  wire [17:0] p1_add_81202_comb;
  wire [17:0] p1_add_81203_comb;
  wire [17:0] p1_add_81204_comb;
  wire [17:0] p1_add_81205_comb;
  wire [17:0] p1_add_81206_comb;
  wire [17:0] p1_add_81207_comb;
  wire [17:0] p1_add_81208_comb;
  wire [17:0] p1_add_81209_comb;
  wire [17:0] p1_add_81210_comb;
  wire [17:0] p1_add_81211_comb;
  wire [17:0] p1_add_81212_comb;
  wire [17:0] p1_add_81213_comb;
  wire [17:0] p1_add_81214_comb;
  wire [17:0] p1_add_81215_comb;
  wire [17:0] p1_add_81216_comb;
  wire [17:0] p1_add_81217_comb;
  wire [17:0] p1_add_81218_comb;
  wire [17:0] p1_add_81219_comb;
  wire [17:0] p1_add_81220_comb;
  wire [17:0] p1_add_81221_comb;
  wire [17:0] p1_add_81222_comb;
  wire [17:0] p1_add_81223_comb;
  wire [17:0] p1_add_81224_comb;
  wire [17:0] p1_add_81225_comb;
  wire [17:0] p1_add_81226_comb;
  wire [17:0] p1_add_81227_comb;
  wire [17:0] p1_add_81228_comb;
  wire [17:0] p1_add_81229_comb;
  wire [17:0] p1_add_81230_comb;
  wire [17:0] p1_add_81231_comb;
  wire [11:0] p1_clipped__136_comb;
  wire [11:0] p1_clipped__152_comb;
  wire [11:0] p1_clipped__168_comb;
  wire [11:0] p1_clipped__184_comb;
  wire [11:0] p1_clipped__200_comb;
  wire [11:0] p1_clipped__216_comb;
  wire [11:0] p1_clipped__232_comb;
  wire [11:0] p1_clipped__248_comb;
  wire [11:0] p1_clipped__137_comb;
  wire [11:0] p1_clipped__153_comb;
  wire [11:0] p1_clipped__169_comb;
  wire [11:0] p1_clipped__185_comb;
  wire [11:0] p1_clipped__201_comb;
  wire [11:0] p1_clipped__217_comb;
  wire [11:0] p1_clipped__233_comb;
  wire [11:0] p1_clipped__249_comb;
  wire [11:0] p1_clipped__138_comb;
  wire [11:0] p1_clipped__154_comb;
  wire [11:0] p1_clipped__170_comb;
  wire [11:0] p1_clipped__186_comb;
  wire [11:0] p1_clipped__202_comb;
  wire [11:0] p1_clipped__218_comb;
  wire [11:0] p1_clipped__234_comb;
  wire [11:0] p1_clipped__250_comb;
  wire [11:0] p1_clipped__139_comb;
  wire [11:0] p1_clipped__155_comb;
  wire [11:0] p1_clipped__171_comb;
  wire [11:0] p1_clipped__187_comb;
  wire [11:0] p1_clipped__203_comb;
  wire [11:0] p1_clipped__219_comb;
  wire [11:0] p1_clipped__235_comb;
  wire [11:0] p1_clipped__251_comb;
  wire [11:0] p1_clipped__140_comb;
  wire [11:0] p1_clipped__156_comb;
  wire [11:0] p1_clipped__172_comb;
  wire [11:0] p1_clipped__188_comb;
  wire [11:0] p1_clipped__204_comb;
  wire [11:0] p1_clipped__220_comb;
  wire [11:0] p1_clipped__236_comb;
  wire [11:0] p1_clipped__252_comb;
  wire [11:0] p1_clipped__141_comb;
  wire [11:0] p1_clipped__157_comb;
  wire [11:0] p1_clipped__173_comb;
  wire [11:0] p1_clipped__189_comb;
  wire [11:0] p1_clipped__205_comb;
  wire [11:0] p1_clipped__221_comb;
  wire [11:0] p1_clipped__237_comb;
  wire [11:0] p1_clipped__253_comb;
  wire [11:0] p1_clipped__142_comb;
  wire [11:0] p1_clipped__158_comb;
  wire [11:0] p1_clipped__174_comb;
  wire [11:0] p1_clipped__190_comb;
  wire [11:0] p1_clipped__206_comb;
  wire [11:0] p1_clipped__222_comb;
  wire [11:0] p1_clipped__238_comb;
  wire [11:0] p1_clipped__254_comb;
  wire [11:0] p1_clipped__143_comb;
  wire [11:0] p1_clipped__159_comb;
  wire [11:0] p1_clipped__175_comb;
  wire [11:0] p1_clipped__191_comb;
  wire [11:0] p1_clipped__207_comb;
  wire [11:0] p1_clipped__223_comb;
  wire [11:0] p1_clipped__239_comb;
  wire [11:0] p1_clipped__255_comb;
  wire [11:0] p1_array_81872_comb[0:7];
  wire [11:0] p1_array_81873_comb[0:7];
  wire [11:0] p1_array_81874_comb[0:7];
  wire [11:0] p1_array_81875_comb[0:7];
  wire [11:0] p1_array_81876_comb[0:7];
  wire [11:0] p1_array_81877_comb[0:7];
  wire [11:0] p1_array_81878_comb[0:7];
  wire [11:0] p1_array_81879_comb[0:7];
  wire [11:0] p1_col_transformed_comb[0:7][0:7];
  assign p1_array_index_75184_comb = p0_x[3'h2][3'h2];
  assign p1_array_index_75185_comb = p0_x[3'h2][3'h3];
  assign p1_array_index_75186_comb = p0_x[3'h2][3'h4];
  assign p1_array_index_75187_comb = p0_x[3'h2][3'h5];
  assign p1_array_index_75188_comb = p0_x[3'h3][3'h2];
  assign p1_array_index_75189_comb = p0_x[3'h3][3'h3];
  assign p1_array_index_75190_comb = p0_x[3'h3][3'h4];
  assign p1_array_index_75191_comb = p0_x[3'h3][3'h5];
  assign p1_array_index_75192_comb = p0_x[3'h4][3'h2];
  assign p1_array_index_75193_comb = p0_x[3'h4][3'h3];
  assign p1_array_index_75194_comb = p0_x[3'h4][3'h4];
  assign p1_array_index_75195_comb = p0_x[3'h4][3'h5];
  assign p1_array_index_75196_comb = p0_x[3'h5][3'h2];
  assign p1_array_index_75197_comb = p0_x[3'h5][3'h3];
  assign p1_array_index_75198_comb = p0_x[3'h5][3'h4];
  assign p1_array_index_75199_comb = p0_x[3'h5][3'h5];
  assign p1_array_index_75200_comb = p0_x[3'h2][3'h1];
  assign p1_array_index_75201_comb = p0_x[3'h2][3'h6];
  assign p1_array_index_75202_comb = p0_x[3'h3][3'h1];
  assign p1_array_index_75203_comb = p0_x[3'h3][3'h6];
  assign p1_array_index_75204_comb = p0_x[3'h4][3'h1];
  assign p1_array_index_75205_comb = p0_x[3'h4][3'h6];
  assign p1_array_index_75206_comb = p0_x[3'h5][3'h1];
  assign p1_array_index_75207_comb = p0_x[3'h5][3'h6];
  assign p1_array_index_75208_comb = p0_x[3'h2][3'h0];
  assign p1_array_index_75209_comb = p0_x[3'h2][3'h7];
  assign p1_array_index_75210_comb = p0_x[3'h3][3'h0];
  assign p1_array_index_75211_comb = p0_x[3'h3][3'h7];
  assign p1_array_index_75212_comb = p0_x[3'h4][3'h0];
  assign p1_array_index_75213_comb = p0_x[3'h4][3'h7];
  assign p1_array_index_75214_comb = p0_x[3'h5][3'h0];
  assign p1_array_index_75215_comb = p0_x[3'h5][3'h7];
  assign p1_array_index_75216_comb = p0_x[3'h1][3'h2];
  assign p1_array_index_75217_comb = p0_x[3'h1][3'h3];
  assign p1_array_index_75218_comb = p0_x[3'h1][3'h4];
  assign p1_array_index_75219_comb = p0_x[3'h1][3'h5];
  assign p1_array_index_75220_comb = p0_x[3'h6][3'h2];
  assign p1_array_index_75221_comb = p0_x[3'h6][3'h3];
  assign p1_array_index_75222_comb = p0_x[3'h6][3'h4];
  assign p1_array_index_75223_comb = p0_x[3'h6][3'h5];
  assign p1_array_index_75224_comb = p0_x[3'h1][3'h1];
  assign p1_array_index_75225_comb = p0_x[3'h1][3'h6];
  assign p1_array_index_75226_comb = p0_x[3'h6][3'h1];
  assign p1_array_index_75227_comb = p0_x[3'h6][3'h6];
  assign p1_array_index_75228_comb = p0_x[3'h1][3'h0];
  assign p1_array_index_75229_comb = p0_x[3'h1][3'h7];
  assign p1_array_index_75230_comb = p0_x[3'h6][3'h0];
  assign p1_array_index_75231_comb = p0_x[3'h6][3'h7];
  assign p1_array_index_75232_comb = p0_x[3'h0][3'h2];
  assign p1_array_index_75233_comb = p0_x[3'h0][3'h3];
  assign p1_array_index_75234_comb = p0_x[3'h0][3'h4];
  assign p1_array_index_75235_comb = p0_x[3'h0][3'h5];
  assign p1_array_index_75236_comb = p0_x[3'h7][3'h2];
  assign p1_array_index_75237_comb = p0_x[3'h7][3'h3];
  assign p1_array_index_75238_comb = p0_x[3'h7][3'h4];
  assign p1_array_index_75239_comb = p0_x[3'h7][3'h5];
  assign p1_array_index_75240_comb = p0_x[3'h0][3'h1];
  assign p1_array_index_75241_comb = p0_x[3'h0][3'h6];
  assign p1_array_index_75242_comb = p0_x[3'h7][3'h1];
  assign p1_array_index_75243_comb = p0_x[3'h7][3'h6];
  assign p1_array_index_75244_comb = p0_x[3'h0][3'h0];
  assign p1_array_index_75245_comb = p0_x[3'h0][3'h7];
  assign p1_array_index_75246_comb = p0_x[3'h7][3'h0];
  assign p1_array_index_75247_comb = p0_x[3'h7][3'h7];
  assign p1_sign_ext_75250_comb = {{12{p1_array_index_75184_comb[11]}}, p1_array_index_75184_comb};
  assign p1_sign_ext_75251_comb = {{12{p1_array_index_75185_comb[11]}}, p1_array_index_75185_comb};
  assign p1_sign_ext_75252_comb = {{12{p1_array_index_75186_comb[11]}}, p1_array_index_75186_comb};
  assign p1_sign_ext_75253_comb = {{12{p1_array_index_75187_comb[11]}}, p1_array_index_75187_comb};
  assign p1_sign_ext_75258_comb = {{12{p1_array_index_75188_comb[11]}}, p1_array_index_75188_comb};
  assign p1_sign_ext_75259_comb = {{12{p1_array_index_75189_comb[11]}}, p1_array_index_75189_comb};
  assign p1_sign_ext_75260_comb = {{12{p1_array_index_75190_comb[11]}}, p1_array_index_75190_comb};
  assign p1_sign_ext_75261_comb = {{12{p1_array_index_75191_comb[11]}}, p1_array_index_75191_comb};
  assign p1_sign_ext_75266_comb = {{12{p1_array_index_75192_comb[11]}}, p1_array_index_75192_comb};
  assign p1_sign_ext_75267_comb = {{12{p1_array_index_75193_comb[11]}}, p1_array_index_75193_comb};
  assign p1_sign_ext_75268_comb = {{12{p1_array_index_75194_comb[11]}}, p1_array_index_75194_comb};
  assign p1_sign_ext_75269_comb = {{12{p1_array_index_75195_comb[11]}}, p1_array_index_75195_comb};
  assign p1_sign_ext_75274_comb = {{12{p1_array_index_75196_comb[11]}}, p1_array_index_75196_comb};
  assign p1_sign_ext_75275_comb = {{12{p1_array_index_75197_comb[11]}}, p1_array_index_75197_comb};
  assign p1_sign_ext_75276_comb = {{12{p1_array_index_75198_comb[11]}}, p1_array_index_75198_comb};
  assign p1_sign_ext_75277_comb = {{12{p1_array_index_75199_comb[11]}}, p1_array_index_75199_comb};
  assign p1_sign_ext_75280_comb = {{12{p1_array_index_75200_comb[11]}}, p1_array_index_75200_comb};
  assign p1_sign_ext_75281_comb = {{12{p1_array_index_75201_comb[11]}}, p1_array_index_75201_comb};
  assign p1_sign_ext_75282_comb = {{12{p1_array_index_75202_comb[11]}}, p1_array_index_75202_comb};
  assign p1_sign_ext_75283_comb = {{12{p1_array_index_75203_comb[11]}}, p1_array_index_75203_comb};
  assign p1_sign_ext_75284_comb = {{12{p1_array_index_75204_comb[11]}}, p1_array_index_75204_comb};
  assign p1_sign_ext_75285_comb = {{12{p1_array_index_75205_comb[11]}}, p1_array_index_75205_comb};
  assign p1_sign_ext_75286_comb = {{12{p1_array_index_75206_comb[11]}}, p1_array_index_75206_comb};
  assign p1_sign_ext_75287_comb = {{12{p1_array_index_75207_comb[11]}}, p1_array_index_75207_comb};
  assign p1_sign_ext_75304_comb = {{12{p1_array_index_75208_comb[11]}}, p1_array_index_75208_comb};
  assign p1_sign_ext_75309_comb = {{12{p1_array_index_75209_comb[11]}}, p1_array_index_75209_comb};
  assign p1_sign_ext_75310_comb = {{12{p1_array_index_75210_comb[11]}}, p1_array_index_75210_comb};
  assign p1_sign_ext_75315_comb = {{12{p1_array_index_75211_comb[11]}}, p1_array_index_75211_comb};
  assign p1_sign_ext_75316_comb = {{12{p1_array_index_75212_comb[11]}}, p1_array_index_75212_comb};
  assign p1_sign_ext_75321_comb = {{12{p1_array_index_75213_comb[11]}}, p1_array_index_75213_comb};
  assign p1_sign_ext_75322_comb = {{12{p1_array_index_75214_comb[11]}}, p1_array_index_75214_comb};
  assign p1_sign_ext_75327_comb = {{12{p1_array_index_75215_comb[11]}}, p1_array_index_75215_comb};
  assign p1_sign_ext_75346_comb = {{12{p1_array_index_75216_comb[11]}}, p1_array_index_75216_comb};
  assign p1_sign_ext_75347_comb = {{12{p1_array_index_75217_comb[11]}}, p1_array_index_75217_comb};
  assign p1_sign_ext_75348_comb = {{12{p1_array_index_75218_comb[11]}}, p1_array_index_75218_comb};
  assign p1_sign_ext_75349_comb = {{12{p1_array_index_75219_comb[11]}}, p1_array_index_75219_comb};
  assign p1_sign_ext_75354_comb = {{12{p1_array_index_75220_comb[11]}}, p1_array_index_75220_comb};
  assign p1_sign_ext_75355_comb = {{12{p1_array_index_75221_comb[11]}}, p1_array_index_75221_comb};
  assign p1_sign_ext_75356_comb = {{12{p1_array_index_75222_comb[11]}}, p1_array_index_75222_comb};
  assign p1_sign_ext_75357_comb = {{12{p1_array_index_75223_comb[11]}}, p1_array_index_75223_comb};
  assign p1_sign_ext_75360_comb = {{12{p1_array_index_75224_comb[11]}}, p1_array_index_75224_comb};
  assign p1_sign_ext_75361_comb = {{12{p1_array_index_75225_comb[11]}}, p1_array_index_75225_comb};
  assign p1_sign_ext_75362_comb = {{12{p1_array_index_75226_comb[11]}}, p1_array_index_75226_comb};
  assign p1_sign_ext_75363_comb = {{12{p1_array_index_75227_comb[11]}}, p1_array_index_75227_comb};
  assign p1_sign_ext_75372_comb = {{12{p1_array_index_75228_comb[11]}}, p1_array_index_75228_comb};
  assign p1_sign_ext_75377_comb = {{12{p1_array_index_75229_comb[11]}}, p1_array_index_75229_comb};
  assign p1_sign_ext_75378_comb = {{12{p1_array_index_75230_comb[11]}}, p1_array_index_75230_comb};
  assign p1_sign_ext_75383_comb = {{12{p1_array_index_75231_comb[11]}}, p1_array_index_75231_comb};
  assign p1_sign_ext_75394_comb = {{12{p1_array_index_75232_comb[11]}}, p1_array_index_75232_comb};
  assign p1_sign_ext_75395_comb = {{12{p1_array_index_75233_comb[11]}}, p1_array_index_75233_comb};
  assign p1_sign_ext_75396_comb = {{12{p1_array_index_75234_comb[11]}}, p1_array_index_75234_comb};
  assign p1_sign_ext_75397_comb = {{12{p1_array_index_75235_comb[11]}}, p1_array_index_75235_comb};
  assign p1_sign_ext_75402_comb = {{12{p1_array_index_75236_comb[11]}}, p1_array_index_75236_comb};
  assign p1_sign_ext_75403_comb = {{12{p1_array_index_75237_comb[11]}}, p1_array_index_75237_comb};
  assign p1_sign_ext_75404_comb = {{12{p1_array_index_75238_comb[11]}}, p1_array_index_75238_comb};
  assign p1_sign_ext_75405_comb = {{12{p1_array_index_75239_comb[11]}}, p1_array_index_75239_comb};
  assign p1_sign_ext_75408_comb = {{12{p1_array_index_75240_comb[11]}}, p1_array_index_75240_comb};
  assign p1_sign_ext_75409_comb = {{12{p1_array_index_75241_comb[11]}}, p1_array_index_75241_comb};
  assign p1_sign_ext_75410_comb = {{12{p1_array_index_75242_comb[11]}}, p1_array_index_75242_comb};
  assign p1_sign_ext_75411_comb = {{12{p1_array_index_75243_comb[11]}}, p1_array_index_75243_comb};
  assign p1_sign_ext_75420_comb = {{12{p1_array_index_75244_comb[11]}}, p1_array_index_75244_comb};
  assign p1_sign_ext_75425_comb = {{12{p1_array_index_75245_comb[11]}}, p1_array_index_75245_comb};
  assign p1_sign_ext_75426_comb = {{12{p1_array_index_75246_comb[11]}}, p1_array_index_75246_comb};
  assign p1_sign_ext_75431_comb = {{12{p1_array_index_75247_comb[11]}}, p1_array_index_75247_comb};
  assign p1_smul_75440_comb = smul21b_12b_x_9b(p1_array_index_75208_comb, 9'h0fb);
  assign p1_smul_75441_comb = smul21b_12b_x_9b(p1_array_index_75200_comb, 9'h0d5);
  assign p1_smul_75450_comb = smul21b_12b_x_9b(p1_array_index_75201_comb, 9'h12b);
  assign p1_smul_75451_comb = smul21b_12b_x_9b(p1_array_index_75209_comb, 9'h105);
  assign p1_smul_75452_comb = smul21b_12b_x_9b(p1_array_index_75210_comb, 9'h0fb);
  assign p1_smul_75453_comb = smul21b_12b_x_9b(p1_array_index_75202_comb, 9'h0d5);
  assign p1_smul_75462_comb = smul21b_12b_x_9b(p1_array_index_75203_comb, 9'h12b);
  assign p1_smul_75463_comb = smul21b_12b_x_9b(p1_array_index_75211_comb, 9'h105);
  assign p1_smul_75464_comb = smul21b_12b_x_9b(p1_array_index_75212_comb, 9'h0fb);
  assign p1_smul_75465_comb = smul21b_12b_x_9b(p1_array_index_75204_comb, 9'h0d5);
  assign p1_smul_75474_comb = smul21b_12b_x_9b(p1_array_index_75205_comb, 9'h12b);
  assign p1_smul_75475_comb = smul21b_12b_x_9b(p1_array_index_75213_comb, 9'h105);
  assign p1_smul_75476_comb = smul21b_12b_x_9b(p1_array_index_75214_comb, 9'h0fb);
  assign p1_smul_75477_comb = smul21b_12b_x_9b(p1_array_index_75206_comb, 9'h0d5);
  assign p1_smul_75486_comb = smul21b_12b_x_9b(p1_array_index_75207_comb, 9'h12b);
  assign p1_smul_75487_comb = smul21b_12b_x_9b(p1_array_index_75215_comb, 9'h105);
  assign p1_smul_75512_comb = smul21b_12b_x_9b(p1_array_index_75208_comb, 9'h0d5);
  assign p1_smul_75514_comb = smul21b_12b_x_9b(p1_array_index_75184_comb, 9'h105);
  assign p1_smul_75517_comb = smul21b_12b_x_9b(p1_array_index_75187_comb, 9'h0fb);
  assign p1_smul_75519_comb = smul21b_12b_x_9b(p1_array_index_75209_comb, 9'h12b);
  assign p1_smul_75520_comb = smul21b_12b_x_9b(p1_array_index_75210_comb, 9'h0d5);
  assign p1_smul_75522_comb = smul21b_12b_x_9b(p1_array_index_75188_comb, 9'h105);
  assign p1_smul_75525_comb = smul21b_12b_x_9b(p1_array_index_75191_comb, 9'h0fb);
  assign p1_smul_75527_comb = smul21b_12b_x_9b(p1_array_index_75211_comb, 9'h12b);
  assign p1_smul_75528_comb = smul21b_12b_x_9b(p1_array_index_75212_comb, 9'h0d5);
  assign p1_smul_75530_comb = smul21b_12b_x_9b(p1_array_index_75192_comb, 9'h105);
  assign p1_smul_75533_comb = smul21b_12b_x_9b(p1_array_index_75195_comb, 9'h0fb);
  assign p1_smul_75535_comb = smul21b_12b_x_9b(p1_array_index_75213_comb, 9'h12b);
  assign p1_smul_75536_comb = smul21b_12b_x_9b(p1_array_index_75214_comb, 9'h0d5);
  assign p1_smul_75538_comb = smul21b_12b_x_9b(p1_array_index_75196_comb, 9'h105);
  assign p1_smul_75541_comb = smul21b_12b_x_9b(p1_array_index_75199_comb, 9'h0fb);
  assign p1_smul_75543_comb = smul21b_12b_x_9b(p1_array_index_75215_comb, 9'h12b);
  assign p1_smul_75546_comb = smul21b_12b_x_9b(p1_array_index_75200_comb, 9'h105);
  assign p1_smul_75548_comb = smul21b_12b_x_9b(p1_array_index_75185_comb, 9'h0d5);
  assign p1_smul_75549_comb = smul21b_12b_x_9b(p1_array_index_75186_comb, 9'h0d5);
  assign p1_smul_75551_comb = smul21b_12b_x_9b(p1_array_index_75201_comb, 9'h105);
  assign p1_smul_75556_comb = smul21b_12b_x_9b(p1_array_index_75202_comb, 9'h105);
  assign p1_smul_75558_comb = smul21b_12b_x_9b(p1_array_index_75189_comb, 9'h0d5);
  assign p1_smul_75559_comb = smul21b_12b_x_9b(p1_array_index_75190_comb, 9'h0d5);
  assign p1_smul_75561_comb = smul21b_12b_x_9b(p1_array_index_75203_comb, 9'h105);
  assign p1_smul_75566_comb = smul21b_12b_x_9b(p1_array_index_75204_comb, 9'h105);
  assign p1_smul_75568_comb = smul21b_12b_x_9b(p1_array_index_75193_comb, 9'h0d5);
  assign p1_smul_75569_comb = smul21b_12b_x_9b(p1_array_index_75194_comb, 9'h0d5);
  assign p1_smul_75571_comb = smul21b_12b_x_9b(p1_array_index_75205_comb, 9'h105);
  assign p1_smul_75576_comb = smul21b_12b_x_9b(p1_array_index_75206_comb, 9'h105);
  assign p1_smul_75578_comb = smul21b_12b_x_9b(p1_array_index_75197_comb, 9'h0d5);
  assign p1_smul_75579_comb = smul21b_12b_x_9b(p1_array_index_75198_comb, 9'h0d5);
  assign p1_smul_75581_comb = smul21b_12b_x_9b(p1_array_index_75207_comb, 9'h105);
  assign p1_smul_75602_comb = smul21b_12b_x_9b(p1_array_index_75184_comb, 9'h0d5);
  assign p1_smul_75603_comb = smul21b_12b_x_9b(p1_array_index_75185_comb, 9'h105);
  assign p1_smul_75604_comb = smul21b_12b_x_9b(p1_array_index_75186_comb, 9'h105);
  assign p1_smul_75605_comb = smul21b_12b_x_9b(p1_array_index_75187_comb, 9'h0d5);
  assign p1_smul_75610_comb = smul21b_12b_x_9b(p1_array_index_75188_comb, 9'h0d5);
  assign p1_smul_75611_comb = smul21b_12b_x_9b(p1_array_index_75189_comb, 9'h105);
  assign p1_smul_75612_comb = smul21b_12b_x_9b(p1_array_index_75190_comb, 9'h105);
  assign p1_smul_75613_comb = smul21b_12b_x_9b(p1_array_index_75191_comb, 9'h0d5);
  assign p1_smul_75618_comb = smul21b_12b_x_9b(p1_array_index_75192_comb, 9'h0d5);
  assign p1_smul_75619_comb = smul21b_12b_x_9b(p1_array_index_75193_comb, 9'h105);
  assign p1_smul_75620_comb = smul21b_12b_x_9b(p1_array_index_75194_comb, 9'h105);
  assign p1_smul_75621_comb = smul21b_12b_x_9b(p1_array_index_75195_comb, 9'h0d5);
  assign p1_smul_75626_comb = smul21b_12b_x_9b(p1_array_index_75196_comb, 9'h0d5);
  assign p1_smul_75627_comb = smul21b_12b_x_9b(p1_array_index_75197_comb, 9'h105);
  assign p1_smul_75628_comb = smul21b_12b_x_9b(p1_array_index_75198_comb, 9'h105);
  assign p1_smul_75629_comb = smul21b_12b_x_9b(p1_array_index_75199_comb, 9'h0d5);
  assign p1_smul_75632_comb = smul21b_12b_x_9b(p1_array_index_75228_comb, 9'h0fb);
  assign p1_smul_75633_comb = smul21b_12b_x_9b(p1_array_index_75224_comb, 9'h0d5);
  assign p1_smul_75642_comb = smul21b_12b_x_9b(p1_array_index_75225_comb, 9'h12b);
  assign p1_smul_75643_comb = smul21b_12b_x_9b(p1_array_index_75229_comb, 9'h105);
  assign p1_smul_75644_comb = smul21b_12b_x_9b(p1_array_index_75230_comb, 9'h0fb);
  assign p1_smul_75645_comb = smul21b_12b_x_9b(p1_array_index_75226_comb, 9'h0d5);
  assign p1_smul_75654_comb = smul21b_12b_x_9b(p1_array_index_75227_comb, 9'h12b);
  assign p1_smul_75655_comb = smul21b_12b_x_9b(p1_array_index_75231_comb, 9'h105);
  assign p1_smul_75668_comb = smul21b_12b_x_9b(p1_array_index_75228_comb, 9'h0d5);
  assign p1_smul_75670_comb = smul21b_12b_x_9b(p1_array_index_75216_comb, 9'h105);
  assign p1_smul_75673_comb = smul21b_12b_x_9b(p1_array_index_75219_comb, 9'h0fb);
  assign p1_smul_75675_comb = smul21b_12b_x_9b(p1_array_index_75229_comb, 9'h12b);
  assign p1_smul_75676_comb = smul21b_12b_x_9b(p1_array_index_75230_comb, 9'h0d5);
  assign p1_smul_75678_comb = smul21b_12b_x_9b(p1_array_index_75220_comb, 9'h105);
  assign p1_smul_75681_comb = smul21b_12b_x_9b(p1_array_index_75223_comb, 9'h0fb);
  assign p1_smul_75683_comb = smul21b_12b_x_9b(p1_array_index_75231_comb, 9'h12b);
  assign p1_smul_75686_comb = smul21b_12b_x_9b(p1_array_index_75224_comb, 9'h105);
  assign p1_smul_75688_comb = smul21b_12b_x_9b(p1_array_index_75217_comb, 9'h0d5);
  assign p1_smul_75689_comb = smul21b_12b_x_9b(p1_array_index_75218_comb, 9'h0d5);
  assign p1_smul_75691_comb = smul21b_12b_x_9b(p1_array_index_75225_comb, 9'h105);
  assign p1_smul_75696_comb = smul21b_12b_x_9b(p1_array_index_75226_comb, 9'h105);
  assign p1_smul_75698_comb = smul21b_12b_x_9b(p1_array_index_75221_comb, 9'h0d5);
  assign p1_smul_75699_comb = smul21b_12b_x_9b(p1_array_index_75222_comb, 9'h0d5);
  assign p1_smul_75701_comb = smul21b_12b_x_9b(p1_array_index_75227_comb, 9'h105);
  assign p1_smul_75714_comb = smul21b_12b_x_9b(p1_array_index_75216_comb, 9'h0d5);
  assign p1_smul_75715_comb = smul21b_12b_x_9b(p1_array_index_75217_comb, 9'h105);
  assign p1_smul_75716_comb = smul21b_12b_x_9b(p1_array_index_75218_comb, 9'h105);
  assign p1_smul_75717_comb = smul21b_12b_x_9b(p1_array_index_75219_comb, 9'h0d5);
  assign p1_smul_75722_comb = smul21b_12b_x_9b(p1_array_index_75220_comb, 9'h0d5);
  assign p1_smul_75723_comb = smul21b_12b_x_9b(p1_array_index_75221_comb, 9'h105);
  assign p1_smul_75724_comb = smul21b_12b_x_9b(p1_array_index_75222_comb, 9'h105);
  assign p1_smul_75725_comb = smul21b_12b_x_9b(p1_array_index_75223_comb, 9'h0d5);
  assign p1_smul_75728_comb = smul21b_12b_x_9b(p1_array_index_75244_comb, 9'h0fb);
  assign p1_smul_75729_comb = smul21b_12b_x_9b(p1_array_index_75240_comb, 9'h0d5);
  assign p1_smul_75738_comb = smul21b_12b_x_9b(p1_array_index_75241_comb, 9'h12b);
  assign p1_smul_75739_comb = smul21b_12b_x_9b(p1_array_index_75245_comb, 9'h105);
  assign p1_smul_75740_comb = smul21b_12b_x_9b(p1_array_index_75246_comb, 9'h0fb);
  assign p1_smul_75741_comb = smul21b_12b_x_9b(p1_array_index_75242_comb, 9'h0d5);
  assign p1_smul_75750_comb = smul21b_12b_x_9b(p1_array_index_75243_comb, 9'h12b);
  assign p1_smul_75751_comb = smul21b_12b_x_9b(p1_array_index_75247_comb, 9'h105);
  assign p1_smul_75764_comb = smul21b_12b_x_9b(p1_array_index_75244_comb, 9'h0d5);
  assign p1_smul_75766_comb = smul21b_12b_x_9b(p1_array_index_75232_comb, 9'h105);
  assign p1_smul_75769_comb = smul21b_12b_x_9b(p1_array_index_75235_comb, 9'h0fb);
  assign p1_smul_75771_comb = smul21b_12b_x_9b(p1_array_index_75245_comb, 9'h12b);
  assign p1_smul_75772_comb = smul21b_12b_x_9b(p1_array_index_75246_comb, 9'h0d5);
  assign p1_smul_75774_comb = smul21b_12b_x_9b(p1_array_index_75236_comb, 9'h105);
  assign p1_smul_75777_comb = smul21b_12b_x_9b(p1_array_index_75239_comb, 9'h0fb);
  assign p1_smul_75779_comb = smul21b_12b_x_9b(p1_array_index_75247_comb, 9'h12b);
  assign p1_smul_75782_comb = smul21b_12b_x_9b(p1_array_index_75240_comb, 9'h105);
  assign p1_smul_75784_comb = smul21b_12b_x_9b(p1_array_index_75233_comb, 9'h0d5);
  assign p1_smul_75785_comb = smul21b_12b_x_9b(p1_array_index_75234_comb, 9'h0d5);
  assign p1_smul_75787_comb = smul21b_12b_x_9b(p1_array_index_75241_comb, 9'h105);
  assign p1_smul_75792_comb = smul21b_12b_x_9b(p1_array_index_75242_comb, 9'h105);
  assign p1_smul_75794_comb = smul21b_12b_x_9b(p1_array_index_75237_comb, 9'h0d5);
  assign p1_smul_75795_comb = smul21b_12b_x_9b(p1_array_index_75238_comb, 9'h0d5);
  assign p1_smul_75797_comb = smul21b_12b_x_9b(p1_array_index_75243_comb, 9'h105);
  assign p1_smul_75810_comb = smul21b_12b_x_9b(p1_array_index_75232_comb, 9'h0d5);
  assign p1_smul_75811_comb = smul21b_12b_x_9b(p1_array_index_75233_comb, 9'h105);
  assign p1_smul_75812_comb = smul21b_12b_x_9b(p1_array_index_75234_comb, 9'h105);
  assign p1_smul_75813_comb = smul21b_12b_x_9b(p1_array_index_75235_comb, 9'h0d5);
  assign p1_smul_75818_comb = smul21b_12b_x_9b(p1_array_index_75236_comb, 9'h0d5);
  assign p1_smul_75819_comb = smul21b_12b_x_9b(p1_array_index_75237_comb, 9'h105);
  assign p1_smul_75820_comb = smul21b_12b_x_9b(p1_array_index_75238_comb, 9'h105);
  assign p1_smul_75821_comb = smul21b_12b_x_9b(p1_array_index_75239_comb, 9'h0d5);
  assign p1_add_75824_comb = p1_smul_75440_comb + p1_smul_75441_comb;
  assign p1_smul_75825_comb = smul20b_20b_x_8b(p1_sign_ext_75250_comb[19:0], 8'h47);
  assign p1_smul_75826_comb = smul20b_20b_x_6b(p1_sign_ext_75251_comb[19:0], 6'h19);
  assign p1_smul_75827_comb = smul20b_20b_x_6b(p1_sign_ext_75252_comb[19:0], 6'h27);
  assign p1_smul_75828_comb = smul20b_20b_x_8b(p1_sign_ext_75253_comb[19:0], 8'hb9);
  assign p1_add_75829_comb = p1_smul_75450_comb + p1_smul_75451_comb;
  assign p1_add_75830_comb = p1_smul_75452_comb + p1_smul_75453_comb;
  assign p1_smul_75831_comb = smul20b_20b_x_8b(p1_sign_ext_75258_comb[19:0], 8'h47);
  assign p1_smul_75832_comb = smul20b_20b_x_6b(p1_sign_ext_75259_comb[19:0], 6'h19);
  assign p1_smul_75833_comb = smul20b_20b_x_6b(p1_sign_ext_75260_comb[19:0], 6'h27);
  assign p1_smul_75834_comb = smul20b_20b_x_8b(p1_sign_ext_75261_comb[19:0], 8'hb9);
  assign p1_add_75835_comb = p1_smul_75462_comb + p1_smul_75463_comb;
  assign p1_add_75836_comb = p1_smul_75464_comb + p1_smul_75465_comb;
  assign p1_smul_75837_comb = smul20b_20b_x_8b(p1_sign_ext_75266_comb[19:0], 8'h47);
  assign p1_smul_75838_comb = smul20b_20b_x_6b(p1_sign_ext_75267_comb[19:0], 6'h19);
  assign p1_smul_75839_comb = smul20b_20b_x_6b(p1_sign_ext_75268_comb[19:0], 6'h27);
  assign p1_smul_75840_comb = smul20b_20b_x_8b(p1_sign_ext_75269_comb[19:0], 8'hb9);
  assign p1_add_75841_comb = p1_smul_75474_comb + p1_smul_75475_comb;
  assign p1_add_75842_comb = p1_smul_75476_comb + p1_smul_75477_comb;
  assign p1_smul_75843_comb = smul20b_20b_x_8b(p1_sign_ext_75274_comb[19:0], 8'h47);
  assign p1_smul_75844_comb = smul20b_20b_x_6b(p1_sign_ext_75275_comb[19:0], 6'h19);
  assign p1_smul_75845_comb = smul20b_20b_x_6b(p1_sign_ext_75276_comb[19:0], 6'h27);
  assign p1_smul_75846_comb = smul20b_20b_x_8b(p1_sign_ext_75277_comb[19:0], 8'hb9);
  assign p1_add_75847_comb = p1_smul_75486_comb + p1_smul_75487_comb;
  assign p1_smul_75850_comb = smul20b_20b_x_7b(p1_sign_ext_75280_comb[19:0], 7'h31);
  assign p1_smul_75851_comb = smul20b_20b_x_7b(p1_sign_ext_75250_comb[19:0], 7'h4f);
  assign p1_smul_75856_comb = smul20b_20b_x_7b(p1_sign_ext_75253_comb[19:0], 7'h4f);
  assign p1_smul_75857_comb = smul20b_20b_x_7b(p1_sign_ext_75281_comb[19:0], 7'h31);
  assign p1_smul_75862_comb = smul20b_20b_x_7b(p1_sign_ext_75282_comb[19:0], 7'h31);
  assign p1_smul_75863_comb = smul20b_20b_x_7b(p1_sign_ext_75258_comb[19:0], 7'h4f);
  assign p1_smul_75868_comb = smul20b_20b_x_7b(p1_sign_ext_75261_comb[19:0], 7'h4f);
  assign p1_smul_75869_comb = smul20b_20b_x_7b(p1_sign_ext_75283_comb[19:0], 7'h31);
  assign p1_smul_75874_comb = smul20b_20b_x_7b(p1_sign_ext_75284_comb[19:0], 7'h31);
  assign p1_smul_75875_comb = smul20b_20b_x_7b(p1_sign_ext_75266_comb[19:0], 7'h4f);
  assign p1_smul_75880_comb = smul20b_20b_x_7b(p1_sign_ext_75269_comb[19:0], 7'h4f);
  assign p1_smul_75881_comb = smul20b_20b_x_7b(p1_sign_ext_75285_comb[19:0], 7'h31);
  assign p1_smul_75886_comb = smul20b_20b_x_7b(p1_sign_ext_75286_comb[19:0], 7'h31);
  assign p1_smul_75887_comb = smul20b_20b_x_7b(p1_sign_ext_75274_comb[19:0], 7'h4f);
  assign p1_smul_75892_comb = smul20b_20b_x_7b(p1_sign_ext_75277_comb[19:0], 7'h4f);
  assign p1_smul_75893_comb = smul20b_20b_x_7b(p1_sign_ext_75287_comb[19:0], 7'h31);
  assign p1_smul_75897_comb = smul20b_20b_x_6b(p1_sign_ext_75280_comb[19:0], 6'h27);
  assign p1_smul_75899_comb = smul20b_20b_x_8b(p1_sign_ext_75251_comb[19:0], 8'hb9);
  assign p1_smul_75900_comb = smul20b_20b_x_8b(p1_sign_ext_75252_comb[19:0], 8'h47);
  assign p1_smul_75902_comb = smul20b_20b_x_6b(p1_sign_ext_75281_comb[19:0], 6'h19);
  assign p1_smul_75905_comb = smul20b_20b_x_6b(p1_sign_ext_75282_comb[19:0], 6'h27);
  assign p1_smul_75907_comb = smul20b_20b_x_8b(p1_sign_ext_75259_comb[19:0], 8'hb9);
  assign p1_smul_75908_comb = smul20b_20b_x_8b(p1_sign_ext_75260_comb[19:0], 8'h47);
  assign p1_smul_75910_comb = smul20b_20b_x_6b(p1_sign_ext_75283_comb[19:0], 6'h19);
  assign p1_smul_75913_comb = smul20b_20b_x_6b(p1_sign_ext_75284_comb[19:0], 6'h27);
  assign p1_smul_75915_comb = smul20b_20b_x_8b(p1_sign_ext_75267_comb[19:0], 8'hb9);
  assign p1_smul_75916_comb = smul20b_20b_x_8b(p1_sign_ext_75268_comb[19:0], 8'h47);
  assign p1_smul_75918_comb = smul20b_20b_x_6b(p1_sign_ext_75285_comb[19:0], 6'h19);
  assign p1_smul_75921_comb = smul20b_20b_x_6b(p1_sign_ext_75286_comb[19:0], 6'h27);
  assign p1_smul_75923_comb = smul20b_20b_x_8b(p1_sign_ext_75275_comb[19:0], 8'hb9);
  assign p1_smul_75924_comb = smul20b_20b_x_8b(p1_sign_ext_75276_comb[19:0], 8'h47);
  assign p1_smul_75926_comb = smul20b_20b_x_6b(p1_sign_ext_75287_comb[19:0], 6'h19);
  assign p1_smul_75960_comb = smul20b_20b_x_8b(p1_sign_ext_75304_comb[19:0], 8'h47);
  assign p1_smul_75962_comb = smul20b_20b_x_6b(p1_sign_ext_75250_comb[19:0], 6'h27);
  assign p1_smul_75965_comb = smul20b_20b_x_6b(p1_sign_ext_75253_comb[19:0], 6'h27);
  assign p1_smul_75967_comb = smul20b_20b_x_8b(p1_sign_ext_75309_comb[19:0], 8'h47);
  assign p1_smul_75968_comb = smul20b_20b_x_8b(p1_sign_ext_75310_comb[19:0], 8'h47);
  assign p1_smul_75970_comb = smul20b_20b_x_6b(p1_sign_ext_75258_comb[19:0], 6'h27);
  assign p1_smul_75973_comb = smul20b_20b_x_6b(p1_sign_ext_75261_comb[19:0], 6'h27);
  assign p1_smul_75975_comb = smul20b_20b_x_8b(p1_sign_ext_75315_comb[19:0], 8'h47);
  assign p1_smul_75976_comb = smul20b_20b_x_8b(p1_sign_ext_75316_comb[19:0], 8'h47);
  assign p1_smul_75978_comb = smul20b_20b_x_6b(p1_sign_ext_75266_comb[19:0], 6'h27);
  assign p1_smul_75981_comb = smul20b_20b_x_6b(p1_sign_ext_75269_comb[19:0], 6'h27);
  assign p1_smul_75983_comb = smul20b_20b_x_8b(p1_sign_ext_75321_comb[19:0], 8'h47);
  assign p1_smul_75984_comb = smul20b_20b_x_8b(p1_sign_ext_75322_comb[19:0], 8'h47);
  assign p1_smul_75986_comb = smul20b_20b_x_6b(p1_sign_ext_75274_comb[19:0], 6'h27);
  assign p1_smul_75989_comb = smul20b_20b_x_6b(p1_sign_ext_75277_comb[19:0], 6'h27);
  assign p1_smul_75991_comb = smul20b_20b_x_8b(p1_sign_ext_75327_comb[19:0], 8'h47);
  assign p1_smul_75992_comb = smul20b_20b_x_7b(p1_sign_ext_75304_comb[19:0], 7'h31);
  assign p1_smul_75995_comb = smul20b_20b_x_7b(p1_sign_ext_75250_comb[19:0], 7'h31);
  assign p1_smul_75998_comb = smul20b_20b_x_7b(p1_sign_ext_75253_comb[19:0], 7'h31);
  assign p1_smul_76001_comb = smul20b_20b_x_7b(p1_sign_ext_75309_comb[19:0], 7'h31);
  assign p1_smul_76002_comb = smul20b_20b_x_7b(p1_sign_ext_75310_comb[19:0], 7'h31);
  assign p1_smul_76005_comb = smul20b_20b_x_7b(p1_sign_ext_75258_comb[19:0], 7'h31);
  assign p1_smul_76008_comb = smul20b_20b_x_7b(p1_sign_ext_75261_comb[19:0], 7'h31);
  assign p1_smul_76011_comb = smul20b_20b_x_7b(p1_sign_ext_75315_comb[19:0], 7'h31);
  assign p1_smul_76012_comb = smul20b_20b_x_7b(p1_sign_ext_75316_comb[19:0], 7'h31);
  assign p1_smul_76015_comb = smul20b_20b_x_7b(p1_sign_ext_75266_comb[19:0], 7'h31);
  assign p1_smul_76018_comb = smul20b_20b_x_7b(p1_sign_ext_75269_comb[19:0], 7'h31);
  assign p1_smul_76021_comb = smul20b_20b_x_7b(p1_sign_ext_75321_comb[19:0], 7'h31);
  assign p1_smul_76022_comb = smul20b_20b_x_7b(p1_sign_ext_75322_comb[19:0], 7'h31);
  assign p1_smul_76025_comb = smul20b_20b_x_7b(p1_sign_ext_75274_comb[19:0], 7'h31);
  assign p1_smul_76028_comb = smul20b_20b_x_7b(p1_sign_ext_75277_comb[19:0], 7'h31);
  assign p1_smul_76031_comb = smul20b_20b_x_7b(p1_sign_ext_75327_comb[19:0], 7'h31);
  assign p1_smul_76032_comb = smul20b_20b_x_6b(p1_sign_ext_75304_comb[19:0], 6'h19);
  assign p1_smul_76033_comb = smul20b_20b_x_8b(p1_sign_ext_75280_comb[19:0], 8'hb9);
  assign p1_add_76034_comb = p1_smul_75602_comb + p1_smul_75603_comb;
  assign p1_add_76035_comb = p1_smul_75604_comb + p1_smul_75605_comb;
  assign p1_smul_76036_comb = smul20b_20b_x_8b(p1_sign_ext_75281_comb[19:0], 8'hb9);
  assign p1_smul_76037_comb = smul20b_20b_x_6b(p1_sign_ext_75309_comb[19:0], 6'h19);
  assign p1_smul_76038_comb = smul20b_20b_x_6b(p1_sign_ext_75310_comb[19:0], 6'h19);
  assign p1_smul_76039_comb = smul20b_20b_x_8b(p1_sign_ext_75282_comb[19:0], 8'hb9);
  assign p1_add_76040_comb = p1_smul_75610_comb + p1_smul_75611_comb;
  assign p1_add_76041_comb = p1_smul_75612_comb + p1_smul_75613_comb;
  assign p1_smul_76042_comb = smul20b_20b_x_8b(p1_sign_ext_75283_comb[19:0], 8'hb9);
  assign p1_smul_76043_comb = smul20b_20b_x_6b(p1_sign_ext_75315_comb[19:0], 6'h19);
  assign p1_smul_76044_comb = smul20b_20b_x_6b(p1_sign_ext_75316_comb[19:0], 6'h19);
  assign p1_smul_76045_comb = smul20b_20b_x_8b(p1_sign_ext_75284_comb[19:0], 8'hb9);
  assign p1_add_76046_comb = p1_smul_75618_comb + p1_smul_75619_comb;
  assign p1_add_76047_comb = p1_smul_75620_comb + p1_smul_75621_comb;
  assign p1_smul_76048_comb = smul20b_20b_x_8b(p1_sign_ext_75285_comb[19:0], 8'hb9);
  assign p1_smul_76049_comb = smul20b_20b_x_6b(p1_sign_ext_75321_comb[19:0], 6'h19);
  assign p1_smul_76050_comb = smul20b_20b_x_6b(p1_sign_ext_75322_comb[19:0], 6'h19);
  assign p1_smul_76051_comb = smul20b_20b_x_8b(p1_sign_ext_75286_comb[19:0], 8'hb9);
  assign p1_add_76052_comb = p1_smul_75626_comb + p1_smul_75627_comb;
  assign p1_add_76053_comb = p1_smul_75628_comb + p1_smul_75629_comb;
  assign p1_smul_76054_comb = smul20b_20b_x_8b(p1_sign_ext_75287_comb[19:0], 8'hb9);
  assign p1_smul_76055_comb = smul20b_20b_x_6b(p1_sign_ext_75327_comb[19:0], 6'h19);
  assign p1_add_76056_comb = p1_smul_75632_comb + p1_smul_75633_comb;
  assign p1_smul_76057_comb = smul20b_20b_x_8b(p1_sign_ext_75346_comb[19:0], 8'h47);
  assign p1_smul_76058_comb = smul20b_20b_x_6b(p1_sign_ext_75347_comb[19:0], 6'h19);
  assign p1_smul_76059_comb = smul20b_20b_x_6b(p1_sign_ext_75348_comb[19:0], 6'h27);
  assign p1_smul_76060_comb = smul20b_20b_x_8b(p1_sign_ext_75349_comb[19:0], 8'hb9);
  assign p1_add_76061_comb = p1_smul_75642_comb + p1_smul_75643_comb;
  assign p1_add_76062_comb = p1_smul_75644_comb + p1_smul_75645_comb;
  assign p1_smul_76063_comb = smul20b_20b_x_8b(p1_sign_ext_75354_comb[19:0], 8'h47);
  assign p1_smul_76064_comb = smul20b_20b_x_6b(p1_sign_ext_75355_comb[19:0], 6'h19);
  assign p1_smul_76065_comb = smul20b_20b_x_6b(p1_sign_ext_75356_comb[19:0], 6'h27);
  assign p1_smul_76066_comb = smul20b_20b_x_8b(p1_sign_ext_75357_comb[19:0], 8'hb9);
  assign p1_add_76067_comb = p1_smul_75654_comb + p1_smul_75655_comb;
  assign p1_smul_76070_comb = smul20b_20b_x_7b(p1_sign_ext_75360_comb[19:0], 7'h31);
  assign p1_smul_76071_comb = smul20b_20b_x_7b(p1_sign_ext_75346_comb[19:0], 7'h4f);
  assign p1_smul_76076_comb = smul20b_20b_x_7b(p1_sign_ext_75349_comb[19:0], 7'h4f);
  assign p1_smul_76077_comb = smul20b_20b_x_7b(p1_sign_ext_75361_comb[19:0], 7'h31);
  assign p1_smul_76082_comb = smul20b_20b_x_7b(p1_sign_ext_75362_comb[19:0], 7'h31);
  assign p1_smul_76083_comb = smul20b_20b_x_7b(p1_sign_ext_75354_comb[19:0], 7'h4f);
  assign p1_smul_76088_comb = smul20b_20b_x_7b(p1_sign_ext_75357_comb[19:0], 7'h4f);
  assign p1_smul_76089_comb = smul20b_20b_x_7b(p1_sign_ext_75363_comb[19:0], 7'h31);
  assign p1_smul_76093_comb = smul20b_20b_x_6b(p1_sign_ext_75360_comb[19:0], 6'h27);
  assign p1_smul_76095_comb = smul20b_20b_x_8b(p1_sign_ext_75347_comb[19:0], 8'hb9);
  assign p1_smul_76096_comb = smul20b_20b_x_8b(p1_sign_ext_75348_comb[19:0], 8'h47);
  assign p1_smul_76098_comb = smul20b_20b_x_6b(p1_sign_ext_75361_comb[19:0], 6'h19);
  assign p1_smul_76101_comb = smul20b_20b_x_6b(p1_sign_ext_75362_comb[19:0], 6'h27);
  assign p1_smul_76103_comb = smul20b_20b_x_8b(p1_sign_ext_75355_comb[19:0], 8'hb9);
  assign p1_smul_76104_comb = smul20b_20b_x_8b(p1_sign_ext_75356_comb[19:0], 8'h47);
  assign p1_smul_76106_comb = smul20b_20b_x_6b(p1_sign_ext_75363_comb[19:0], 6'h19);
  assign p1_smul_76124_comb = smul20b_20b_x_8b(p1_sign_ext_75372_comb[19:0], 8'h47);
  assign p1_smul_76126_comb = smul20b_20b_x_6b(p1_sign_ext_75346_comb[19:0], 6'h27);
  assign p1_smul_76129_comb = smul20b_20b_x_6b(p1_sign_ext_75349_comb[19:0], 6'h27);
  assign p1_smul_76131_comb = smul20b_20b_x_8b(p1_sign_ext_75377_comb[19:0], 8'h47);
  assign p1_smul_76132_comb = smul20b_20b_x_8b(p1_sign_ext_75378_comb[19:0], 8'h47);
  assign p1_smul_76134_comb = smul20b_20b_x_6b(p1_sign_ext_75354_comb[19:0], 6'h27);
  assign p1_smul_76137_comb = smul20b_20b_x_6b(p1_sign_ext_75357_comb[19:0], 6'h27);
  assign p1_smul_76139_comb = smul20b_20b_x_8b(p1_sign_ext_75383_comb[19:0], 8'h47);
  assign p1_smul_76140_comb = smul20b_20b_x_7b(p1_sign_ext_75372_comb[19:0], 7'h31);
  assign p1_smul_76143_comb = smul20b_20b_x_7b(p1_sign_ext_75346_comb[19:0], 7'h31);
  assign p1_smul_76146_comb = smul20b_20b_x_7b(p1_sign_ext_75349_comb[19:0], 7'h31);
  assign p1_smul_76149_comb = smul20b_20b_x_7b(p1_sign_ext_75377_comb[19:0], 7'h31);
  assign p1_smul_76150_comb = smul20b_20b_x_7b(p1_sign_ext_75378_comb[19:0], 7'h31);
  assign p1_smul_76153_comb = smul20b_20b_x_7b(p1_sign_ext_75354_comb[19:0], 7'h31);
  assign p1_smul_76156_comb = smul20b_20b_x_7b(p1_sign_ext_75357_comb[19:0], 7'h31);
  assign p1_smul_76159_comb = smul20b_20b_x_7b(p1_sign_ext_75383_comb[19:0], 7'h31);
  assign p1_smul_76160_comb = smul20b_20b_x_6b(p1_sign_ext_75372_comb[19:0], 6'h19);
  assign p1_smul_76161_comb = smul20b_20b_x_8b(p1_sign_ext_75360_comb[19:0], 8'hb9);
  assign p1_add_76162_comb = p1_smul_75714_comb + p1_smul_75715_comb;
  assign p1_add_76163_comb = p1_smul_75716_comb + p1_smul_75717_comb;
  assign p1_smul_76164_comb = smul20b_20b_x_8b(p1_sign_ext_75361_comb[19:0], 8'hb9);
  assign p1_smul_76165_comb = smul20b_20b_x_6b(p1_sign_ext_75377_comb[19:0], 6'h19);
  assign p1_smul_76166_comb = smul20b_20b_x_6b(p1_sign_ext_75378_comb[19:0], 6'h19);
  assign p1_smul_76167_comb = smul20b_20b_x_8b(p1_sign_ext_75362_comb[19:0], 8'hb9);
  assign p1_add_76168_comb = p1_smul_75722_comb + p1_smul_75723_comb;
  assign p1_add_76169_comb = p1_smul_75724_comb + p1_smul_75725_comb;
  assign p1_smul_76170_comb = smul20b_20b_x_8b(p1_sign_ext_75363_comb[19:0], 8'hb9);
  assign p1_smul_76171_comb = smul20b_20b_x_6b(p1_sign_ext_75383_comb[19:0], 6'h19);
  assign p1_add_76172_comb = p1_smul_75728_comb + p1_smul_75729_comb;
  assign p1_smul_76173_comb = smul20b_20b_x_8b(p1_sign_ext_75394_comb[19:0], 8'h47);
  assign p1_smul_76174_comb = smul20b_20b_x_6b(p1_sign_ext_75395_comb[19:0], 6'h19);
  assign p1_smul_76175_comb = smul20b_20b_x_6b(p1_sign_ext_75396_comb[19:0], 6'h27);
  assign p1_smul_76176_comb = smul20b_20b_x_8b(p1_sign_ext_75397_comb[19:0], 8'hb9);
  assign p1_add_76177_comb = p1_smul_75738_comb + p1_smul_75739_comb;
  assign p1_add_76178_comb = p1_smul_75740_comb + p1_smul_75741_comb;
  assign p1_smul_76179_comb = smul20b_20b_x_8b(p1_sign_ext_75402_comb[19:0], 8'h47);
  assign p1_smul_76180_comb = smul20b_20b_x_6b(p1_sign_ext_75403_comb[19:0], 6'h19);
  assign p1_smul_76181_comb = smul20b_20b_x_6b(p1_sign_ext_75404_comb[19:0], 6'h27);
  assign p1_smul_76182_comb = smul20b_20b_x_8b(p1_sign_ext_75405_comb[19:0], 8'hb9);
  assign p1_add_76183_comb = p1_smul_75750_comb + p1_smul_75751_comb;
  assign p1_smul_76186_comb = smul20b_20b_x_7b(p1_sign_ext_75408_comb[19:0], 7'h31);
  assign p1_smul_76187_comb = smul20b_20b_x_7b(p1_sign_ext_75394_comb[19:0], 7'h4f);
  assign p1_smul_76192_comb = smul20b_20b_x_7b(p1_sign_ext_75397_comb[19:0], 7'h4f);
  assign p1_smul_76193_comb = smul20b_20b_x_7b(p1_sign_ext_75409_comb[19:0], 7'h31);
  assign p1_smul_76198_comb = smul20b_20b_x_7b(p1_sign_ext_75410_comb[19:0], 7'h31);
  assign p1_smul_76199_comb = smul20b_20b_x_7b(p1_sign_ext_75402_comb[19:0], 7'h4f);
  assign p1_smul_76204_comb = smul20b_20b_x_7b(p1_sign_ext_75405_comb[19:0], 7'h4f);
  assign p1_smul_76205_comb = smul20b_20b_x_7b(p1_sign_ext_75411_comb[19:0], 7'h31);
  assign p1_smul_76209_comb = smul20b_20b_x_6b(p1_sign_ext_75408_comb[19:0], 6'h27);
  assign p1_smul_76211_comb = smul20b_20b_x_8b(p1_sign_ext_75395_comb[19:0], 8'hb9);
  assign p1_smul_76212_comb = smul20b_20b_x_8b(p1_sign_ext_75396_comb[19:0], 8'h47);
  assign p1_smul_76214_comb = smul20b_20b_x_6b(p1_sign_ext_75409_comb[19:0], 6'h19);
  assign p1_smul_76217_comb = smul20b_20b_x_6b(p1_sign_ext_75410_comb[19:0], 6'h27);
  assign p1_smul_76219_comb = smul20b_20b_x_8b(p1_sign_ext_75403_comb[19:0], 8'hb9);
  assign p1_smul_76220_comb = smul20b_20b_x_8b(p1_sign_ext_75404_comb[19:0], 8'h47);
  assign p1_smul_76222_comb = smul20b_20b_x_6b(p1_sign_ext_75411_comb[19:0], 6'h19);
  assign p1_smul_76240_comb = smul20b_20b_x_8b(p1_sign_ext_75420_comb[19:0], 8'h47);
  assign p1_smul_76242_comb = smul20b_20b_x_6b(p1_sign_ext_75394_comb[19:0], 6'h27);
  assign p1_smul_76245_comb = smul20b_20b_x_6b(p1_sign_ext_75397_comb[19:0], 6'h27);
  assign p1_smul_76247_comb = smul20b_20b_x_8b(p1_sign_ext_75425_comb[19:0], 8'h47);
  assign p1_smul_76248_comb = smul20b_20b_x_8b(p1_sign_ext_75426_comb[19:0], 8'h47);
  assign p1_smul_76250_comb = smul20b_20b_x_6b(p1_sign_ext_75402_comb[19:0], 6'h27);
  assign p1_smul_76253_comb = smul20b_20b_x_6b(p1_sign_ext_75405_comb[19:0], 6'h27);
  assign p1_smul_76255_comb = smul20b_20b_x_8b(p1_sign_ext_75431_comb[19:0], 8'h47);
  assign p1_smul_76256_comb = smul20b_20b_x_7b(p1_sign_ext_75420_comb[19:0], 7'h31);
  assign p1_smul_76259_comb = smul20b_20b_x_7b(p1_sign_ext_75394_comb[19:0], 7'h31);
  assign p1_smul_76262_comb = smul20b_20b_x_7b(p1_sign_ext_75397_comb[19:0], 7'h31);
  assign p1_smul_76265_comb = smul20b_20b_x_7b(p1_sign_ext_75425_comb[19:0], 7'h31);
  assign p1_smul_76266_comb = smul20b_20b_x_7b(p1_sign_ext_75426_comb[19:0], 7'h31);
  assign p1_smul_76269_comb = smul20b_20b_x_7b(p1_sign_ext_75402_comb[19:0], 7'h31);
  assign p1_smul_76272_comb = smul20b_20b_x_7b(p1_sign_ext_75405_comb[19:0], 7'h31);
  assign p1_smul_76275_comb = smul20b_20b_x_7b(p1_sign_ext_75431_comb[19:0], 7'h31);
  assign p1_smul_76276_comb = smul20b_20b_x_6b(p1_sign_ext_75420_comb[19:0], 6'h19);
  assign p1_smul_76277_comb = smul20b_20b_x_8b(p1_sign_ext_75408_comb[19:0], 8'hb9);
  assign p1_add_76278_comb = p1_smul_75810_comb + p1_smul_75811_comb;
  assign p1_add_76279_comb = p1_smul_75812_comb + p1_smul_75813_comb;
  assign p1_smul_76280_comb = smul20b_20b_x_8b(p1_sign_ext_75409_comb[19:0], 8'hb9);
  assign p1_smul_76281_comb = smul20b_20b_x_6b(p1_sign_ext_75425_comb[19:0], 6'h19);
  assign p1_smul_76282_comb = smul20b_20b_x_6b(p1_sign_ext_75426_comb[19:0], 6'h19);
  assign p1_smul_76283_comb = smul20b_20b_x_8b(p1_sign_ext_75410_comb[19:0], 8'hb9);
  assign p1_add_76284_comb = p1_smul_75818_comb + p1_smul_75819_comb;
  assign p1_add_76285_comb = p1_smul_75820_comb + p1_smul_75821_comb;
  assign p1_smul_76286_comb = smul20b_20b_x_8b(p1_sign_ext_75411_comb[19:0], 8'hb9);
  assign p1_smul_76287_comb = smul20b_20b_x_6b(p1_sign_ext_75431_comb[19:0], 6'h19);
  assign p1_bit_slice_76320_comb = p1_add_75824_comb[20:1];
  assign p1_add_76321_comb = p1_smul_75825_comb + p1_smul_75826_comb;
  assign p1_add_76322_comb = p1_smul_75827_comb + p1_smul_75828_comb;
  assign p1_bit_slice_76323_comb = p1_add_75829_comb[20:1];
  assign p1_bit_slice_76324_comb = p1_add_75830_comb[20:1];
  assign p1_add_76325_comb = p1_smul_75831_comb + p1_smul_75832_comb;
  assign p1_add_76326_comb = p1_smul_75833_comb + p1_smul_75834_comb;
  assign p1_bit_slice_76327_comb = p1_add_75835_comb[20:1];
  assign p1_bit_slice_76328_comb = p1_add_75836_comb[20:1];
  assign p1_add_76329_comb = p1_smul_75837_comb + p1_smul_75838_comb;
  assign p1_add_76330_comb = p1_smul_75839_comb + p1_smul_75840_comb;
  assign p1_bit_slice_76331_comb = p1_add_75841_comb[20:1];
  assign p1_bit_slice_76332_comb = p1_add_75842_comb[20:1];
  assign p1_add_76333_comb = p1_smul_75843_comb + p1_smul_75844_comb;
  assign p1_add_76334_comb = p1_smul_75845_comb + p1_smul_75846_comb;
  assign p1_bit_slice_76335_comb = p1_add_75847_comb[20:1];
  assign p1_smul_76336_comb = smul19b_19b_x_7b(p1_sign_ext_75304_comb[18:0], 7'h3b);
  assign p1_smul_76339_comb = smul19b_19b_x_7b(p1_sign_ext_75251_comb[18:0], 7'h45);
  assign p1_smul_76340_comb = smul19b_19b_x_7b(p1_sign_ext_75252_comb[18:0], 7'h45);
  assign p1_smul_76343_comb = smul19b_19b_x_7b(p1_sign_ext_75309_comb[18:0], 7'h3b);
  assign p1_smul_76344_comb = smul19b_19b_x_7b(p1_sign_ext_75310_comb[18:0], 7'h3b);
  assign p1_smul_76347_comb = smul19b_19b_x_7b(p1_sign_ext_75259_comb[18:0], 7'h45);
  assign p1_smul_76348_comb = smul19b_19b_x_7b(p1_sign_ext_75260_comb[18:0], 7'h45);
  assign p1_smul_76351_comb = smul19b_19b_x_7b(p1_sign_ext_75315_comb[18:0], 7'h3b);
  assign p1_smul_76352_comb = smul19b_19b_x_7b(p1_sign_ext_75316_comb[18:0], 7'h3b);
  assign p1_smul_76355_comb = smul19b_19b_x_7b(p1_sign_ext_75267_comb[18:0], 7'h45);
  assign p1_smul_76356_comb = smul19b_19b_x_7b(p1_sign_ext_75268_comb[18:0], 7'h45);
  assign p1_smul_76359_comb = smul19b_19b_x_7b(p1_sign_ext_75321_comb[18:0], 7'h3b);
  assign p1_smul_76360_comb = smul19b_19b_x_7b(p1_sign_ext_75322_comb[18:0], 7'h3b);
  assign p1_smul_76363_comb = smul19b_19b_x_7b(p1_sign_ext_75275_comb[18:0], 7'h45);
  assign p1_smul_76364_comb = smul19b_19b_x_7b(p1_sign_ext_75276_comb[18:0], 7'h45);
  assign p1_smul_76367_comb = smul19b_19b_x_7b(p1_sign_ext_75327_comb[18:0], 7'h3b);
  assign p1_add_76368_comb = p1_smul_75512_comb[20:1] + p1_smul_75897_comb;
  assign p1_add_76370_comb = p1_smul_75514_comb[20:1] + p1_smul_75899_comb;
  assign p1_add_76372_comb = p1_smul_75900_comb + p1_smul_75517_comb[20:1];
  assign p1_add_76374_comb = p1_smul_75902_comb + p1_smul_75519_comb[20:1];
  assign p1_add_76376_comb = p1_smul_75520_comb[20:1] + p1_smul_75905_comb;
  assign p1_add_76378_comb = p1_smul_75522_comb[20:1] + p1_smul_75907_comb;
  assign p1_add_76380_comb = p1_smul_75908_comb + p1_smul_75525_comb[20:1];
  assign p1_add_76382_comb = p1_smul_75910_comb + p1_smul_75527_comb[20:1];
  assign p1_add_76384_comb = p1_smul_75528_comb[20:1] + p1_smul_75913_comb;
  assign p1_add_76386_comb = p1_smul_75530_comb[20:1] + p1_smul_75915_comb;
  assign p1_add_76388_comb = p1_smul_75916_comb + p1_smul_75533_comb[20:1];
  assign p1_add_76390_comb = p1_smul_75918_comb + p1_smul_75535_comb[20:1];
  assign p1_add_76392_comb = p1_smul_75536_comb[20:1] + p1_smul_75921_comb;
  assign p1_add_76394_comb = p1_smul_75538_comb[20:1] + p1_smul_75923_comb;
  assign p1_add_76396_comb = p1_smul_75924_comb + p1_smul_75541_comb[20:1];
  assign p1_add_76398_comb = p1_smul_75926_comb + p1_smul_75543_comb[20:1];
  assign p1_smul_76400_comb = smul21b_12b_x_9b(p1_array_index_75208_comb, 9'h0b5);
  assign p1_smul_76401_comb = smul21b_12b_x_9b(p1_array_index_75200_comb, 9'h14b);
  assign p1_smul_76402_comb = smul21b_12b_x_9b(p1_array_index_75184_comb, 9'h14b);
  assign p1_smul_76403_comb = smul21b_12b_x_9b(p1_array_index_75185_comb, 9'h0b5);
  assign p1_smul_76404_comb = smul21b_12b_x_9b(p1_array_index_75186_comb, 9'h0b5);
  assign p1_smul_76405_comb = smul21b_12b_x_9b(p1_array_index_75187_comb, 9'h14b);
  assign p1_smul_76406_comb = smul21b_12b_x_9b(p1_array_index_75201_comb, 9'h14b);
  assign p1_smul_76407_comb = smul21b_12b_x_9b(p1_array_index_75209_comb, 9'h0b5);
  assign p1_smul_76408_comb = smul21b_12b_x_9b(p1_array_index_75210_comb, 9'h0b5);
  assign p1_smul_76409_comb = smul21b_12b_x_9b(p1_array_index_75202_comb, 9'h14b);
  assign p1_smul_76410_comb = smul21b_12b_x_9b(p1_array_index_75188_comb, 9'h14b);
  assign p1_smul_76411_comb = smul21b_12b_x_9b(p1_array_index_75189_comb, 9'h0b5);
  assign p1_smul_76412_comb = smul21b_12b_x_9b(p1_array_index_75190_comb, 9'h0b5);
  assign p1_smul_76413_comb = smul21b_12b_x_9b(p1_array_index_75191_comb, 9'h14b);
  assign p1_smul_76414_comb = smul21b_12b_x_9b(p1_array_index_75203_comb, 9'h14b);
  assign p1_smul_76415_comb = smul21b_12b_x_9b(p1_array_index_75211_comb, 9'h0b5);
  assign p1_smul_76416_comb = smul21b_12b_x_9b(p1_array_index_75212_comb, 9'h0b5);
  assign p1_smul_76417_comb = smul21b_12b_x_9b(p1_array_index_75204_comb, 9'h14b);
  assign p1_smul_76418_comb = smul21b_12b_x_9b(p1_array_index_75192_comb, 9'h14b);
  assign p1_smul_76419_comb = smul21b_12b_x_9b(p1_array_index_75193_comb, 9'h0b5);
  assign p1_smul_76420_comb = smul21b_12b_x_9b(p1_array_index_75194_comb, 9'h0b5);
  assign p1_smul_76421_comb = smul21b_12b_x_9b(p1_array_index_75195_comb, 9'h14b);
  assign p1_smul_76422_comb = smul21b_12b_x_9b(p1_array_index_75205_comb, 9'h14b);
  assign p1_smul_76423_comb = smul21b_12b_x_9b(p1_array_index_75213_comb, 9'h0b5);
  assign p1_smul_76424_comb = smul21b_12b_x_9b(p1_array_index_75214_comb, 9'h0b5);
  assign p1_smul_76425_comb = smul21b_12b_x_9b(p1_array_index_75206_comb, 9'h14b);
  assign p1_smul_76426_comb = smul21b_12b_x_9b(p1_array_index_75196_comb, 9'h14b);
  assign p1_smul_76427_comb = smul21b_12b_x_9b(p1_array_index_75197_comb, 9'h0b5);
  assign p1_smul_76428_comb = smul21b_12b_x_9b(p1_array_index_75198_comb, 9'h0b5);
  assign p1_smul_76429_comb = smul21b_12b_x_9b(p1_array_index_75199_comb, 9'h14b);
  assign p1_smul_76430_comb = smul21b_12b_x_9b(p1_array_index_75207_comb, 9'h14b);
  assign p1_smul_76431_comb = smul21b_12b_x_9b(p1_array_index_75215_comb, 9'h0b5);
  assign p1_add_76432_comb = p1_smul_75960_comb + p1_smul_75546_comb[20:1];
  assign p1_add_76434_comb = p1_smul_75962_comb + p1_smul_75548_comb[20:1];
  assign p1_add_76436_comb = p1_smul_75549_comb[20:1] + p1_smul_75965_comb;
  assign p1_add_76438_comb = p1_smul_75551_comb[20:1] + p1_smul_75967_comb;
  assign p1_add_76440_comb = p1_smul_75968_comb + p1_smul_75556_comb[20:1];
  assign p1_add_76442_comb = p1_smul_75970_comb + p1_smul_75558_comb[20:1];
  assign p1_add_76444_comb = p1_smul_75559_comb[20:1] + p1_smul_75973_comb;
  assign p1_add_76446_comb = p1_smul_75561_comb[20:1] + p1_smul_75975_comb;
  assign p1_add_76448_comb = p1_smul_75976_comb + p1_smul_75566_comb[20:1];
  assign p1_add_76450_comb = p1_smul_75978_comb + p1_smul_75568_comb[20:1];
  assign p1_add_76452_comb = p1_smul_75569_comb[20:1] + p1_smul_75981_comb;
  assign p1_add_76454_comb = p1_smul_75571_comb[20:1] + p1_smul_75983_comb;
  assign p1_add_76456_comb = p1_smul_75984_comb + p1_smul_75576_comb[20:1];
  assign p1_add_76458_comb = p1_smul_75986_comb + p1_smul_75578_comb[20:1];
  assign p1_add_76460_comb = p1_smul_75579_comb[20:1] + p1_smul_75989_comb;
  assign p1_add_76462_comb = p1_smul_75581_comb[20:1] + p1_smul_75991_comb;
  assign p1_smul_76465_comb = smul19b_19b_x_7b(p1_sign_ext_75280_comb[18:0], 7'h45);
  assign p1_smul_76467_comb = smul19b_19b_x_7b(p1_sign_ext_75251_comb[18:0], 7'h3b);
  assign p1_smul_76468_comb = smul19b_19b_x_7b(p1_sign_ext_75252_comb[18:0], 7'h3b);
  assign p1_smul_76470_comb = smul19b_19b_x_7b(p1_sign_ext_75281_comb[18:0], 7'h45);
  assign p1_smul_76473_comb = smul19b_19b_x_7b(p1_sign_ext_75282_comb[18:0], 7'h45);
  assign p1_smul_76475_comb = smul19b_19b_x_7b(p1_sign_ext_75259_comb[18:0], 7'h3b);
  assign p1_smul_76476_comb = smul19b_19b_x_7b(p1_sign_ext_75260_comb[18:0], 7'h3b);
  assign p1_smul_76478_comb = smul19b_19b_x_7b(p1_sign_ext_75283_comb[18:0], 7'h45);
  assign p1_smul_76481_comb = smul19b_19b_x_7b(p1_sign_ext_75284_comb[18:0], 7'h45);
  assign p1_smul_76483_comb = smul19b_19b_x_7b(p1_sign_ext_75267_comb[18:0], 7'h3b);
  assign p1_smul_76484_comb = smul19b_19b_x_7b(p1_sign_ext_75268_comb[18:0], 7'h3b);
  assign p1_smul_76486_comb = smul19b_19b_x_7b(p1_sign_ext_75285_comb[18:0], 7'h45);
  assign p1_smul_76489_comb = smul19b_19b_x_7b(p1_sign_ext_75286_comb[18:0], 7'h45);
  assign p1_smul_76491_comb = smul19b_19b_x_7b(p1_sign_ext_75275_comb[18:0], 7'h3b);
  assign p1_smul_76492_comb = smul19b_19b_x_7b(p1_sign_ext_75276_comb[18:0], 7'h3b);
  assign p1_smul_76494_comb = smul19b_19b_x_7b(p1_sign_ext_75287_comb[18:0], 7'h45);
  assign p1_add_76496_comb = p1_smul_76032_comb + p1_smul_76033_comb;
  assign p1_bit_slice_76497_comb = p1_add_76034_comb[20:1];
  assign p1_bit_slice_76498_comb = p1_add_76035_comb[20:1];
  assign p1_add_76499_comb = p1_smul_76036_comb + p1_smul_76037_comb;
  assign p1_add_76500_comb = p1_smul_76038_comb + p1_smul_76039_comb;
  assign p1_bit_slice_76501_comb = p1_add_76040_comb[20:1];
  assign p1_bit_slice_76502_comb = p1_add_76041_comb[20:1];
  assign p1_add_76503_comb = p1_smul_76042_comb + p1_smul_76043_comb;
  assign p1_add_76504_comb = p1_smul_76044_comb + p1_smul_76045_comb;
  assign p1_bit_slice_76505_comb = p1_add_76046_comb[20:1];
  assign p1_bit_slice_76506_comb = p1_add_76047_comb[20:1];
  assign p1_add_76507_comb = p1_smul_76048_comb + p1_smul_76049_comb;
  assign p1_add_76508_comb = p1_smul_76050_comb + p1_smul_76051_comb;
  assign p1_bit_slice_76509_comb = p1_add_76052_comb[20:1];
  assign p1_bit_slice_76510_comb = p1_add_76053_comb[20:1];
  assign p1_add_76511_comb = p1_smul_76054_comb + p1_smul_76055_comb;
  assign p1_bit_slice_76528_comb = p1_add_76056_comb[20:1];
  assign p1_add_76529_comb = p1_smul_76057_comb + p1_smul_76058_comb;
  assign p1_add_76530_comb = p1_smul_76059_comb + p1_smul_76060_comb;
  assign p1_bit_slice_76531_comb = p1_add_76061_comb[20:1];
  assign p1_bit_slice_76532_comb = p1_add_76062_comb[20:1];
  assign p1_add_76533_comb = p1_smul_76063_comb + p1_smul_76064_comb;
  assign p1_add_76534_comb = p1_smul_76065_comb + p1_smul_76066_comb;
  assign p1_bit_slice_76535_comb = p1_add_76067_comb[20:1];
  assign p1_smul_76536_comb = smul19b_19b_x_7b(p1_sign_ext_75372_comb[18:0], 7'h3b);
  assign p1_smul_76539_comb = smul19b_19b_x_7b(p1_sign_ext_75347_comb[18:0], 7'h45);
  assign p1_smul_76540_comb = smul19b_19b_x_7b(p1_sign_ext_75348_comb[18:0], 7'h45);
  assign p1_smul_76543_comb = smul19b_19b_x_7b(p1_sign_ext_75377_comb[18:0], 7'h3b);
  assign p1_smul_76544_comb = smul19b_19b_x_7b(p1_sign_ext_75378_comb[18:0], 7'h3b);
  assign p1_smul_76547_comb = smul19b_19b_x_7b(p1_sign_ext_75355_comb[18:0], 7'h45);
  assign p1_smul_76548_comb = smul19b_19b_x_7b(p1_sign_ext_75356_comb[18:0], 7'h45);
  assign p1_smul_76551_comb = smul19b_19b_x_7b(p1_sign_ext_75383_comb[18:0], 7'h3b);
  assign p1_add_76552_comb = p1_smul_75668_comb[20:1] + p1_smul_76093_comb;
  assign p1_add_76554_comb = p1_smul_75670_comb[20:1] + p1_smul_76095_comb;
  assign p1_add_76556_comb = p1_smul_76096_comb + p1_smul_75673_comb[20:1];
  assign p1_add_76558_comb = p1_smul_76098_comb + p1_smul_75675_comb[20:1];
  assign p1_add_76560_comb = p1_smul_75676_comb[20:1] + p1_smul_76101_comb;
  assign p1_add_76562_comb = p1_smul_75678_comb[20:1] + p1_smul_76103_comb;
  assign p1_add_76564_comb = p1_smul_76104_comb + p1_smul_75681_comb[20:1];
  assign p1_add_76566_comb = p1_smul_76106_comb + p1_smul_75683_comb[20:1];
  assign p1_smul_76568_comb = smul21b_12b_x_9b(p1_array_index_75228_comb, 9'h0b5);
  assign p1_smul_76569_comb = smul21b_12b_x_9b(p1_array_index_75224_comb, 9'h14b);
  assign p1_smul_76570_comb = smul21b_12b_x_9b(p1_array_index_75216_comb, 9'h14b);
  assign p1_smul_76571_comb = smul21b_12b_x_9b(p1_array_index_75217_comb, 9'h0b5);
  assign p1_smul_76572_comb = smul21b_12b_x_9b(p1_array_index_75218_comb, 9'h0b5);
  assign p1_smul_76573_comb = smul21b_12b_x_9b(p1_array_index_75219_comb, 9'h14b);
  assign p1_smul_76574_comb = smul21b_12b_x_9b(p1_array_index_75225_comb, 9'h14b);
  assign p1_smul_76575_comb = smul21b_12b_x_9b(p1_array_index_75229_comb, 9'h0b5);
  assign p1_smul_76576_comb = smul21b_12b_x_9b(p1_array_index_75230_comb, 9'h0b5);
  assign p1_smul_76577_comb = smul21b_12b_x_9b(p1_array_index_75226_comb, 9'h14b);
  assign p1_smul_76578_comb = smul21b_12b_x_9b(p1_array_index_75220_comb, 9'h14b);
  assign p1_smul_76579_comb = smul21b_12b_x_9b(p1_array_index_75221_comb, 9'h0b5);
  assign p1_smul_76580_comb = smul21b_12b_x_9b(p1_array_index_75222_comb, 9'h0b5);
  assign p1_smul_76581_comb = smul21b_12b_x_9b(p1_array_index_75223_comb, 9'h14b);
  assign p1_smul_76582_comb = smul21b_12b_x_9b(p1_array_index_75227_comb, 9'h14b);
  assign p1_smul_76583_comb = smul21b_12b_x_9b(p1_array_index_75231_comb, 9'h0b5);
  assign p1_add_76584_comb = p1_smul_76124_comb + p1_smul_75686_comb[20:1];
  assign p1_add_76586_comb = p1_smul_76126_comb + p1_smul_75688_comb[20:1];
  assign p1_add_76588_comb = p1_smul_75689_comb[20:1] + p1_smul_76129_comb;
  assign p1_add_76590_comb = p1_smul_75691_comb[20:1] + p1_smul_76131_comb;
  assign p1_add_76592_comb = p1_smul_76132_comb + p1_smul_75696_comb[20:1];
  assign p1_add_76594_comb = p1_smul_76134_comb + p1_smul_75698_comb[20:1];
  assign p1_add_76596_comb = p1_smul_75699_comb[20:1] + p1_smul_76137_comb;
  assign p1_add_76598_comb = p1_smul_75701_comb[20:1] + p1_smul_76139_comb;
  assign p1_smul_76601_comb = smul19b_19b_x_7b(p1_sign_ext_75360_comb[18:0], 7'h45);
  assign p1_smul_76603_comb = smul19b_19b_x_7b(p1_sign_ext_75347_comb[18:0], 7'h3b);
  assign p1_smul_76604_comb = smul19b_19b_x_7b(p1_sign_ext_75348_comb[18:0], 7'h3b);
  assign p1_smul_76606_comb = smul19b_19b_x_7b(p1_sign_ext_75361_comb[18:0], 7'h45);
  assign p1_smul_76609_comb = smul19b_19b_x_7b(p1_sign_ext_75362_comb[18:0], 7'h45);
  assign p1_smul_76611_comb = smul19b_19b_x_7b(p1_sign_ext_75355_comb[18:0], 7'h3b);
  assign p1_smul_76612_comb = smul19b_19b_x_7b(p1_sign_ext_75356_comb[18:0], 7'h3b);
  assign p1_smul_76614_comb = smul19b_19b_x_7b(p1_sign_ext_75363_comb[18:0], 7'h45);
  assign p1_add_76616_comb = p1_smul_76160_comb + p1_smul_76161_comb;
  assign p1_bit_slice_76617_comb = p1_add_76162_comb[20:1];
  assign p1_bit_slice_76618_comb = p1_add_76163_comb[20:1];
  assign p1_add_76619_comb = p1_smul_76164_comb + p1_smul_76165_comb;
  assign p1_add_76620_comb = p1_smul_76166_comb + p1_smul_76167_comb;
  assign p1_bit_slice_76621_comb = p1_add_76168_comb[20:1];
  assign p1_bit_slice_76622_comb = p1_add_76169_comb[20:1];
  assign p1_add_76623_comb = p1_smul_76170_comb + p1_smul_76171_comb;
  assign p1_bit_slice_76640_comb = p1_add_76172_comb[20:1];
  assign p1_add_76641_comb = p1_smul_76173_comb + p1_smul_76174_comb;
  assign p1_add_76642_comb = p1_smul_76175_comb + p1_smul_76176_comb;
  assign p1_bit_slice_76643_comb = p1_add_76177_comb[20:1];
  assign p1_bit_slice_76644_comb = p1_add_76178_comb[20:1];
  assign p1_add_76645_comb = p1_smul_76179_comb + p1_smul_76180_comb;
  assign p1_add_76646_comb = p1_smul_76181_comb + p1_smul_76182_comb;
  assign p1_bit_slice_76647_comb = p1_add_76183_comb[20:1];
  assign p1_smul_76648_comb = smul19b_19b_x_7b(p1_sign_ext_75420_comb[18:0], 7'h3b);
  assign p1_smul_76651_comb = smul19b_19b_x_7b(p1_sign_ext_75395_comb[18:0], 7'h45);
  assign p1_smul_76652_comb = smul19b_19b_x_7b(p1_sign_ext_75396_comb[18:0], 7'h45);
  assign p1_smul_76655_comb = smul19b_19b_x_7b(p1_sign_ext_75425_comb[18:0], 7'h3b);
  assign p1_smul_76656_comb = smul19b_19b_x_7b(p1_sign_ext_75426_comb[18:0], 7'h3b);
  assign p1_smul_76659_comb = smul19b_19b_x_7b(p1_sign_ext_75403_comb[18:0], 7'h45);
  assign p1_smul_76660_comb = smul19b_19b_x_7b(p1_sign_ext_75404_comb[18:0], 7'h45);
  assign p1_smul_76663_comb = smul19b_19b_x_7b(p1_sign_ext_75431_comb[18:0], 7'h3b);
  assign p1_add_76664_comb = p1_smul_75764_comb[20:1] + p1_smul_76209_comb;
  assign p1_add_76666_comb = p1_smul_75766_comb[20:1] + p1_smul_76211_comb;
  assign p1_add_76668_comb = p1_smul_76212_comb + p1_smul_75769_comb[20:1];
  assign p1_add_76670_comb = p1_smul_76214_comb + p1_smul_75771_comb[20:1];
  assign p1_add_76672_comb = p1_smul_75772_comb[20:1] + p1_smul_76217_comb;
  assign p1_add_76674_comb = p1_smul_75774_comb[20:1] + p1_smul_76219_comb;
  assign p1_add_76676_comb = p1_smul_76220_comb + p1_smul_75777_comb[20:1];
  assign p1_add_76678_comb = p1_smul_76222_comb + p1_smul_75779_comb[20:1];
  assign p1_smul_76680_comb = smul21b_12b_x_9b(p1_array_index_75244_comb, 9'h0b5);
  assign p1_smul_76681_comb = smul21b_12b_x_9b(p1_array_index_75240_comb, 9'h14b);
  assign p1_smul_76682_comb = smul21b_12b_x_9b(p1_array_index_75232_comb, 9'h14b);
  assign p1_smul_76683_comb = smul21b_12b_x_9b(p1_array_index_75233_comb, 9'h0b5);
  assign p1_smul_76684_comb = smul21b_12b_x_9b(p1_array_index_75234_comb, 9'h0b5);
  assign p1_smul_76685_comb = smul21b_12b_x_9b(p1_array_index_75235_comb, 9'h14b);
  assign p1_smul_76686_comb = smul21b_12b_x_9b(p1_array_index_75241_comb, 9'h14b);
  assign p1_smul_76687_comb = smul21b_12b_x_9b(p1_array_index_75245_comb, 9'h0b5);
  assign p1_smul_76688_comb = smul21b_12b_x_9b(p1_array_index_75246_comb, 9'h0b5);
  assign p1_smul_76689_comb = smul21b_12b_x_9b(p1_array_index_75242_comb, 9'h14b);
  assign p1_smul_76690_comb = smul21b_12b_x_9b(p1_array_index_75236_comb, 9'h14b);
  assign p1_smul_76691_comb = smul21b_12b_x_9b(p1_array_index_75237_comb, 9'h0b5);
  assign p1_smul_76692_comb = smul21b_12b_x_9b(p1_array_index_75238_comb, 9'h0b5);
  assign p1_smul_76693_comb = smul21b_12b_x_9b(p1_array_index_75239_comb, 9'h14b);
  assign p1_smul_76694_comb = smul21b_12b_x_9b(p1_array_index_75243_comb, 9'h14b);
  assign p1_smul_76695_comb = smul21b_12b_x_9b(p1_array_index_75247_comb, 9'h0b5);
  assign p1_add_76696_comb = p1_smul_76240_comb + p1_smul_75782_comb[20:1];
  assign p1_add_76698_comb = p1_smul_76242_comb + p1_smul_75784_comb[20:1];
  assign p1_add_76700_comb = p1_smul_75785_comb[20:1] + p1_smul_76245_comb;
  assign p1_add_76702_comb = p1_smul_75787_comb[20:1] + p1_smul_76247_comb;
  assign p1_add_76704_comb = p1_smul_76248_comb + p1_smul_75792_comb[20:1];
  assign p1_add_76706_comb = p1_smul_76250_comb + p1_smul_75794_comb[20:1];
  assign p1_add_76708_comb = p1_smul_75795_comb[20:1] + p1_smul_76253_comb;
  assign p1_add_76710_comb = p1_smul_75797_comb[20:1] + p1_smul_76255_comb;
  assign p1_smul_76713_comb = smul19b_19b_x_7b(p1_sign_ext_75408_comb[18:0], 7'h45);
  assign p1_smul_76715_comb = smul19b_19b_x_7b(p1_sign_ext_75395_comb[18:0], 7'h3b);
  assign p1_smul_76716_comb = smul19b_19b_x_7b(p1_sign_ext_75396_comb[18:0], 7'h3b);
  assign p1_smul_76718_comb = smul19b_19b_x_7b(p1_sign_ext_75409_comb[18:0], 7'h45);
  assign p1_smul_76721_comb = smul19b_19b_x_7b(p1_sign_ext_75410_comb[18:0], 7'h45);
  assign p1_smul_76723_comb = smul19b_19b_x_7b(p1_sign_ext_75403_comb[18:0], 7'h3b);
  assign p1_smul_76724_comb = smul19b_19b_x_7b(p1_sign_ext_75404_comb[18:0], 7'h3b);
  assign p1_smul_76726_comb = smul19b_19b_x_7b(p1_sign_ext_75411_comb[18:0], 7'h45);
  assign p1_add_76728_comb = p1_smul_76276_comb + p1_smul_76277_comb;
  assign p1_bit_slice_76729_comb = p1_add_76278_comb[20:1];
  assign p1_bit_slice_76730_comb = p1_add_76279_comb[20:1];
  assign p1_add_76731_comb = p1_smul_76280_comb + p1_smul_76281_comb;
  assign p1_add_76732_comb = p1_smul_76282_comb + p1_smul_76283_comb;
  assign p1_bit_slice_76733_comb = p1_add_76284_comb[20:1];
  assign p1_bit_slice_76734_comb = p1_add_76285_comb[20:1];
  assign p1_add_76735_comb = p1_smul_76286_comb + p1_smul_76287_comb;
  assign p1_add_76736_comb = p1_sign_ext_75304_comb[12:0] + p1_sign_ext_75280_comb[12:0];
  assign p1_add_76737_comb = p1_sign_ext_75250_comb[12:0] + p1_sign_ext_75251_comb[12:0];
  assign p1_add_76738_comb = p1_sign_ext_75252_comb[12:0] + p1_sign_ext_75253_comb[12:0];
  assign p1_add_76739_comb = p1_sign_ext_75281_comb[12:0] + p1_sign_ext_75309_comb[12:0];
  assign p1_add_76740_comb = p1_sign_ext_75310_comb[12:0] + p1_sign_ext_75282_comb[12:0];
  assign p1_add_76741_comb = p1_sign_ext_75258_comb[12:0] + p1_sign_ext_75259_comb[12:0];
  assign p1_add_76742_comb = p1_sign_ext_75260_comb[12:0] + p1_sign_ext_75261_comb[12:0];
  assign p1_add_76743_comb = p1_sign_ext_75283_comb[12:0] + p1_sign_ext_75315_comb[12:0];
  assign p1_add_76744_comb = p1_sign_ext_75316_comb[12:0] + p1_sign_ext_75284_comb[12:0];
  assign p1_add_76745_comb = p1_sign_ext_75266_comb[12:0] + p1_sign_ext_75267_comb[12:0];
  assign p1_add_76746_comb = p1_sign_ext_75268_comb[12:0] + p1_sign_ext_75269_comb[12:0];
  assign p1_add_76747_comb = p1_sign_ext_75285_comb[12:0] + p1_sign_ext_75321_comb[12:0];
  assign p1_add_76748_comb = p1_sign_ext_75322_comb[12:0] + p1_sign_ext_75286_comb[12:0];
  assign p1_add_76749_comb = p1_sign_ext_75274_comb[12:0] + p1_sign_ext_75275_comb[12:0];
  assign p1_add_76750_comb = p1_sign_ext_75276_comb[12:0] + p1_sign_ext_75277_comb[12:0];
  assign p1_add_76751_comb = p1_sign_ext_75287_comb[12:0] + p1_sign_ext_75327_comb[12:0];
  assign p1_add_76768_comb = p1_smul_76336_comb + p1_smul_75850_comb[19:1];
  assign p1_add_76770_comb = p1_smul_75851_comb[19:1] + p1_smul_76339_comb;
  assign p1_add_76772_comb = p1_smul_76340_comb + p1_smul_75856_comb[19:1];
  assign p1_add_76774_comb = p1_smul_75857_comb[19:1] + p1_smul_76343_comb;
  assign p1_add_76776_comb = p1_smul_76344_comb + p1_smul_75862_comb[19:1];
  assign p1_add_76778_comb = p1_smul_75863_comb[19:1] + p1_smul_76347_comb;
  assign p1_add_76780_comb = p1_smul_76348_comb + p1_smul_75868_comb[19:1];
  assign p1_add_76782_comb = p1_smul_75869_comb[19:1] + p1_smul_76351_comb;
  assign p1_add_76784_comb = p1_smul_76352_comb + p1_smul_75874_comb[19:1];
  assign p1_add_76786_comb = p1_smul_75875_comb[19:1] + p1_smul_76355_comb;
  assign p1_add_76788_comb = p1_smul_76356_comb + p1_smul_75880_comb[19:1];
  assign p1_add_76790_comb = p1_smul_75881_comb[19:1] + p1_smul_76359_comb;
  assign p1_add_76792_comb = p1_smul_76360_comb + p1_smul_75886_comb[19:1];
  assign p1_add_76794_comb = p1_smul_75887_comb[19:1] + p1_smul_76363_comb;
  assign p1_add_76796_comb = p1_smul_76364_comb + p1_smul_75892_comb[19:1];
  assign p1_add_76798_comb = p1_smul_75893_comb[19:1] + p1_smul_76367_comb;
  assign p1_concat_76800_comb = {p1_add_76368_comb, p1_smul_75512_comb[0]};
  assign p1_concat_76801_comb = {p1_add_76370_comb, p1_smul_75514_comb[0]};
  assign p1_concat_76802_comb = {p1_add_76372_comb, p1_smul_75517_comb[0]};
  assign p1_concat_76803_comb = {p1_add_76374_comb, p1_smul_75519_comb[0]};
  assign p1_concat_76804_comb = {p1_add_76376_comb, p1_smul_75520_comb[0]};
  assign p1_concat_76805_comb = {p1_add_76378_comb, p1_smul_75522_comb[0]};
  assign p1_concat_76806_comb = {p1_add_76380_comb, p1_smul_75525_comb[0]};
  assign p1_concat_76807_comb = {p1_add_76382_comb, p1_smul_75527_comb[0]};
  assign p1_concat_76808_comb = {p1_add_76384_comb, p1_smul_75528_comb[0]};
  assign p1_concat_76809_comb = {p1_add_76386_comb, p1_smul_75530_comb[0]};
  assign p1_concat_76810_comb = {p1_add_76388_comb, p1_smul_75533_comb[0]};
  assign p1_concat_76811_comb = {p1_add_76390_comb, p1_smul_75535_comb[0]};
  assign p1_concat_76812_comb = {p1_add_76392_comb, p1_smul_75536_comb[0]};
  assign p1_concat_76813_comb = {p1_add_76394_comb, p1_smul_75538_comb[0]};
  assign p1_concat_76814_comb = {p1_add_76396_comb, p1_smul_75541_comb[0]};
  assign p1_concat_76815_comb = {p1_add_76398_comb, p1_smul_75543_comb[0]};
  assign p1_add_76816_comb = p1_smul_76400_comb + p1_smul_76401_comb;
  assign p1_add_76817_comb = p1_smul_76402_comb + p1_smul_76403_comb;
  assign p1_add_76818_comb = p1_smul_76404_comb + p1_smul_76405_comb;
  assign p1_add_76819_comb = p1_smul_76406_comb + p1_smul_76407_comb;
  assign p1_add_76820_comb = p1_smul_76408_comb + p1_smul_76409_comb;
  assign p1_add_76821_comb = p1_smul_76410_comb + p1_smul_76411_comb;
  assign p1_add_76822_comb = p1_smul_76412_comb + p1_smul_76413_comb;
  assign p1_add_76823_comb = p1_smul_76414_comb + p1_smul_76415_comb;
  assign p1_add_76824_comb = p1_smul_76416_comb + p1_smul_76417_comb;
  assign p1_add_76825_comb = p1_smul_76418_comb + p1_smul_76419_comb;
  assign p1_add_76826_comb = p1_smul_76420_comb + p1_smul_76421_comb;
  assign p1_add_76827_comb = p1_smul_76422_comb + p1_smul_76423_comb;
  assign p1_add_76828_comb = p1_smul_76424_comb + p1_smul_76425_comb;
  assign p1_add_76829_comb = p1_smul_76426_comb + p1_smul_76427_comb;
  assign p1_add_76830_comb = p1_smul_76428_comb + p1_smul_76429_comb;
  assign p1_add_76831_comb = p1_smul_76430_comb + p1_smul_76431_comb;
  assign p1_concat_76832_comb = {p1_add_76432_comb, p1_smul_75546_comb[0]};
  assign p1_concat_76833_comb = {p1_add_76434_comb, p1_smul_75548_comb[0]};
  assign p1_concat_76834_comb = {p1_add_76436_comb, p1_smul_75549_comb[0]};
  assign p1_concat_76835_comb = {p1_add_76438_comb, p1_smul_75551_comb[0]};
  assign p1_concat_76836_comb = {p1_add_76440_comb, p1_smul_75556_comb[0]};
  assign p1_concat_76837_comb = {p1_add_76442_comb, p1_smul_75558_comb[0]};
  assign p1_concat_76838_comb = {p1_add_76444_comb, p1_smul_75559_comb[0]};
  assign p1_concat_76839_comb = {p1_add_76446_comb, p1_smul_75561_comb[0]};
  assign p1_concat_76840_comb = {p1_add_76448_comb, p1_smul_75566_comb[0]};
  assign p1_concat_76841_comb = {p1_add_76450_comb, p1_smul_75568_comb[0]};
  assign p1_concat_76842_comb = {p1_add_76452_comb, p1_smul_75569_comb[0]};
  assign p1_concat_76843_comb = {p1_add_76454_comb, p1_smul_75571_comb[0]};
  assign p1_concat_76844_comb = {p1_add_76456_comb, p1_smul_75576_comb[0]};
  assign p1_concat_76845_comb = {p1_add_76458_comb, p1_smul_75578_comb[0]};
  assign p1_concat_76846_comb = {p1_add_76460_comb, p1_smul_75579_comb[0]};
  assign p1_concat_76847_comb = {p1_add_76462_comb, p1_smul_75581_comb[0]};
  assign p1_add_76848_comb = p1_smul_75992_comb[19:1] + p1_smul_76465_comb;
  assign p1_add_76850_comb = p1_smul_75995_comb[19:1] + p1_smul_76467_comb;
  assign p1_add_76852_comb = p1_smul_76468_comb + p1_smul_75998_comb[19:1];
  assign p1_add_76854_comb = p1_smul_76470_comb + p1_smul_76001_comb[19:1];
  assign p1_add_76856_comb = p1_smul_76002_comb[19:1] + p1_smul_76473_comb;
  assign p1_add_76858_comb = p1_smul_76005_comb[19:1] + p1_smul_76475_comb;
  assign p1_add_76860_comb = p1_smul_76476_comb + p1_smul_76008_comb[19:1];
  assign p1_add_76862_comb = p1_smul_76478_comb + p1_smul_76011_comb[19:1];
  assign p1_add_76864_comb = p1_smul_76012_comb[19:1] + p1_smul_76481_comb;
  assign p1_add_76866_comb = p1_smul_76015_comb[19:1] + p1_smul_76483_comb;
  assign p1_add_76868_comb = p1_smul_76484_comb + p1_smul_76018_comb[19:1];
  assign p1_add_76870_comb = p1_smul_76486_comb + p1_smul_76021_comb[19:1];
  assign p1_add_76872_comb = p1_smul_76022_comb[19:1] + p1_smul_76489_comb;
  assign p1_add_76874_comb = p1_smul_76025_comb[19:1] + p1_smul_76491_comb;
  assign p1_add_76876_comb = p1_smul_76492_comb + p1_smul_76028_comb[19:1];
  assign p1_add_76878_comb = p1_smul_76494_comb + p1_smul_76031_comb[19:1];
  assign p1_add_76896_comb = p1_sign_ext_75372_comb[12:0] + p1_sign_ext_75360_comb[12:0];
  assign p1_add_76897_comb = p1_sign_ext_75346_comb[12:0] + p1_sign_ext_75347_comb[12:0];
  assign p1_add_76898_comb = p1_sign_ext_75348_comb[12:0] + p1_sign_ext_75349_comb[12:0];
  assign p1_add_76899_comb = p1_sign_ext_75361_comb[12:0] + p1_sign_ext_75377_comb[12:0];
  assign p1_add_76900_comb = p1_sign_ext_75378_comb[12:0] + p1_sign_ext_75362_comb[12:0];
  assign p1_add_76901_comb = p1_sign_ext_75354_comb[12:0] + p1_sign_ext_75355_comb[12:0];
  assign p1_add_76902_comb = p1_sign_ext_75356_comb[12:0] + p1_sign_ext_75357_comb[12:0];
  assign p1_add_76903_comb = p1_sign_ext_75363_comb[12:0] + p1_sign_ext_75383_comb[12:0];
  assign p1_add_76912_comb = p1_smul_76536_comb + p1_smul_76070_comb[19:1];
  assign p1_add_76914_comb = p1_smul_76071_comb[19:1] + p1_smul_76539_comb;
  assign p1_add_76916_comb = p1_smul_76540_comb + p1_smul_76076_comb[19:1];
  assign p1_add_76918_comb = p1_smul_76077_comb[19:1] + p1_smul_76543_comb;
  assign p1_add_76920_comb = p1_smul_76544_comb + p1_smul_76082_comb[19:1];
  assign p1_add_76922_comb = p1_smul_76083_comb[19:1] + p1_smul_76547_comb;
  assign p1_add_76924_comb = p1_smul_76548_comb + p1_smul_76088_comb[19:1];
  assign p1_add_76926_comb = p1_smul_76089_comb[19:1] + p1_smul_76551_comb;
  assign p1_concat_76928_comb = {p1_add_76552_comb, p1_smul_75668_comb[0]};
  assign p1_concat_76929_comb = {p1_add_76554_comb, p1_smul_75670_comb[0]};
  assign p1_concat_76930_comb = {p1_add_76556_comb, p1_smul_75673_comb[0]};
  assign p1_concat_76931_comb = {p1_add_76558_comb, p1_smul_75675_comb[0]};
  assign p1_concat_76932_comb = {p1_add_76560_comb, p1_smul_75676_comb[0]};
  assign p1_concat_76933_comb = {p1_add_76562_comb, p1_smul_75678_comb[0]};
  assign p1_concat_76934_comb = {p1_add_76564_comb, p1_smul_75681_comb[0]};
  assign p1_concat_76935_comb = {p1_add_76566_comb, p1_smul_75683_comb[0]};
  assign p1_add_76936_comb = p1_smul_76568_comb + p1_smul_76569_comb;
  assign p1_add_76937_comb = p1_smul_76570_comb + p1_smul_76571_comb;
  assign p1_add_76938_comb = p1_smul_76572_comb + p1_smul_76573_comb;
  assign p1_add_76939_comb = p1_smul_76574_comb + p1_smul_76575_comb;
  assign p1_add_76940_comb = p1_smul_76576_comb + p1_smul_76577_comb;
  assign p1_add_76941_comb = p1_smul_76578_comb + p1_smul_76579_comb;
  assign p1_add_76942_comb = p1_smul_76580_comb + p1_smul_76581_comb;
  assign p1_add_76943_comb = p1_smul_76582_comb + p1_smul_76583_comb;
  assign p1_concat_76944_comb = {p1_add_76584_comb, p1_smul_75686_comb[0]};
  assign p1_concat_76945_comb = {p1_add_76586_comb, p1_smul_75688_comb[0]};
  assign p1_concat_76946_comb = {p1_add_76588_comb, p1_smul_75689_comb[0]};
  assign p1_concat_76947_comb = {p1_add_76590_comb, p1_smul_75691_comb[0]};
  assign p1_concat_76948_comb = {p1_add_76592_comb, p1_smul_75696_comb[0]};
  assign p1_concat_76949_comb = {p1_add_76594_comb, p1_smul_75698_comb[0]};
  assign p1_concat_76950_comb = {p1_add_76596_comb, p1_smul_75699_comb[0]};
  assign p1_concat_76951_comb = {p1_add_76598_comb, p1_smul_75701_comb[0]};
  assign p1_add_76952_comb = p1_smul_76140_comb[19:1] + p1_smul_76601_comb;
  assign p1_add_76954_comb = p1_smul_76143_comb[19:1] + p1_smul_76603_comb;
  assign p1_add_76956_comb = p1_smul_76604_comb + p1_smul_76146_comb[19:1];
  assign p1_add_76958_comb = p1_smul_76606_comb + p1_smul_76149_comb[19:1];
  assign p1_add_76960_comb = p1_smul_76150_comb[19:1] + p1_smul_76609_comb;
  assign p1_add_76962_comb = p1_smul_76153_comb[19:1] + p1_smul_76611_comb;
  assign p1_add_76964_comb = p1_smul_76612_comb + p1_smul_76156_comb[19:1];
  assign p1_add_76966_comb = p1_smul_76614_comb + p1_smul_76159_comb[19:1];
  assign p1_add_76976_comb = p1_sign_ext_75420_comb[12:0] + p1_sign_ext_75408_comb[12:0];
  assign p1_add_76977_comb = p1_sign_ext_75394_comb[12:0] + p1_sign_ext_75395_comb[12:0];
  assign p1_add_76978_comb = p1_sign_ext_75396_comb[12:0] + p1_sign_ext_75397_comb[12:0];
  assign p1_add_76979_comb = p1_sign_ext_75409_comb[12:0] + p1_sign_ext_75425_comb[12:0];
  assign p1_add_76980_comb = p1_sign_ext_75426_comb[12:0] + p1_sign_ext_75410_comb[12:0];
  assign p1_add_76981_comb = p1_sign_ext_75402_comb[12:0] + p1_sign_ext_75403_comb[12:0];
  assign p1_add_76982_comb = p1_sign_ext_75404_comb[12:0] + p1_sign_ext_75405_comb[12:0];
  assign p1_add_76983_comb = p1_sign_ext_75411_comb[12:0] + p1_sign_ext_75431_comb[12:0];
  assign p1_add_76992_comb = p1_smul_76648_comb + p1_smul_76186_comb[19:1];
  assign p1_add_76994_comb = p1_smul_76187_comb[19:1] + p1_smul_76651_comb;
  assign p1_add_76996_comb = p1_smul_76652_comb + p1_smul_76192_comb[19:1];
  assign p1_add_76998_comb = p1_smul_76193_comb[19:1] + p1_smul_76655_comb;
  assign p1_add_77000_comb = p1_smul_76656_comb + p1_smul_76198_comb[19:1];
  assign p1_add_77002_comb = p1_smul_76199_comb[19:1] + p1_smul_76659_comb;
  assign p1_add_77004_comb = p1_smul_76660_comb + p1_smul_76204_comb[19:1];
  assign p1_add_77006_comb = p1_smul_76205_comb[19:1] + p1_smul_76663_comb;
  assign p1_concat_77008_comb = {p1_add_76664_comb, p1_smul_75764_comb[0]};
  assign p1_concat_77009_comb = {p1_add_76666_comb, p1_smul_75766_comb[0]};
  assign p1_concat_77010_comb = {p1_add_76668_comb, p1_smul_75769_comb[0]};
  assign p1_concat_77011_comb = {p1_add_76670_comb, p1_smul_75771_comb[0]};
  assign p1_concat_77012_comb = {p1_add_76672_comb, p1_smul_75772_comb[0]};
  assign p1_concat_77013_comb = {p1_add_76674_comb, p1_smul_75774_comb[0]};
  assign p1_concat_77014_comb = {p1_add_76676_comb, p1_smul_75777_comb[0]};
  assign p1_concat_77015_comb = {p1_add_76678_comb, p1_smul_75779_comb[0]};
  assign p1_add_77016_comb = p1_smul_76680_comb + p1_smul_76681_comb;
  assign p1_add_77017_comb = p1_smul_76682_comb + p1_smul_76683_comb;
  assign p1_add_77018_comb = p1_smul_76684_comb + p1_smul_76685_comb;
  assign p1_add_77019_comb = p1_smul_76686_comb + p1_smul_76687_comb;
  assign p1_add_77020_comb = p1_smul_76688_comb + p1_smul_76689_comb;
  assign p1_add_77021_comb = p1_smul_76690_comb + p1_smul_76691_comb;
  assign p1_add_77022_comb = p1_smul_76692_comb + p1_smul_76693_comb;
  assign p1_add_77023_comb = p1_smul_76694_comb + p1_smul_76695_comb;
  assign p1_concat_77024_comb = {p1_add_76696_comb, p1_smul_75782_comb[0]};
  assign p1_concat_77025_comb = {p1_add_76698_comb, p1_smul_75784_comb[0]};
  assign p1_concat_77026_comb = {p1_add_76700_comb, p1_smul_75785_comb[0]};
  assign p1_concat_77027_comb = {p1_add_76702_comb, p1_smul_75787_comb[0]};
  assign p1_concat_77028_comb = {p1_add_76704_comb, p1_smul_75792_comb[0]};
  assign p1_concat_77029_comb = {p1_add_76706_comb, p1_smul_75794_comb[0]};
  assign p1_concat_77030_comb = {p1_add_76708_comb, p1_smul_75795_comb[0]};
  assign p1_concat_77031_comb = {p1_add_76710_comb, p1_smul_75797_comb[0]};
  assign p1_add_77032_comb = p1_smul_76256_comb[19:1] + p1_smul_76713_comb;
  assign p1_add_77034_comb = p1_smul_76259_comb[19:1] + p1_smul_76715_comb;
  assign p1_add_77036_comb = p1_smul_76716_comb + p1_smul_76262_comb[19:1];
  assign p1_add_77038_comb = p1_smul_76718_comb + p1_smul_76265_comb[19:1];
  assign p1_add_77040_comb = p1_smul_76266_comb[19:1] + p1_smul_76721_comb;
  assign p1_add_77042_comb = p1_smul_76269_comb[19:1] + p1_smul_76723_comb;
  assign p1_add_77044_comb = p1_smul_76724_comb + p1_smul_76272_comb[19:1];
  assign p1_add_77046_comb = p1_smul_76726_comb + p1_smul_76275_comb[19:1];
  assign p1_add_77072_comb = {{4{p1_bit_slice_76320_comb[19]}}, p1_bit_slice_76320_comb} + {{4{p1_add_76321_comb[19]}}, p1_add_76321_comb};
  assign p1_add_77074_comb = {{4{p1_add_76322_comb[19]}}, p1_add_76322_comb} + {{4{p1_bit_slice_76323_comb[19]}}, p1_bit_slice_76323_comb};
  assign p1_add_77076_comb = {{4{p1_bit_slice_76324_comb[19]}}, p1_bit_slice_76324_comb} + {{4{p1_add_76325_comb[19]}}, p1_add_76325_comb};
  assign p1_add_77078_comb = {{4{p1_add_76326_comb[19]}}, p1_add_76326_comb} + {{4{p1_bit_slice_76327_comb[19]}}, p1_bit_slice_76327_comb};
  assign p1_add_77080_comb = {{4{p1_bit_slice_76328_comb[19]}}, p1_bit_slice_76328_comb} + {{4{p1_add_76329_comb[19]}}, p1_add_76329_comb};
  assign p1_add_77082_comb = {{4{p1_add_76330_comb[19]}}, p1_add_76330_comb} + {{4{p1_bit_slice_76331_comb[19]}}, p1_bit_slice_76331_comb};
  assign p1_add_77084_comb = {{4{p1_bit_slice_76332_comb[19]}}, p1_bit_slice_76332_comb} + {{4{p1_add_76333_comb[19]}}, p1_add_76333_comb};
  assign p1_add_77086_comb = {{4{p1_add_76334_comb[19]}}, p1_add_76334_comb} + {{4{p1_bit_slice_76335_comb[19]}}, p1_bit_slice_76335_comb};
  assign p1_concat_77088_comb = {p1_add_76768_comb, p1_smul_75850_comb[0]};
  assign p1_concat_77089_comb = {p1_add_76770_comb, p1_smul_75851_comb[0]};
  assign p1_concat_77090_comb = {p1_add_76772_comb, p1_smul_75856_comb[0]};
  assign p1_concat_77091_comb = {p1_add_76774_comb, p1_smul_75857_comb[0]};
  assign p1_concat_77092_comb = {p1_add_76776_comb, p1_smul_75862_comb[0]};
  assign p1_concat_77093_comb = {p1_add_76778_comb, p1_smul_75863_comb[0]};
  assign p1_concat_77094_comb = {p1_add_76780_comb, p1_smul_75868_comb[0]};
  assign p1_concat_77095_comb = {p1_add_76782_comb, p1_smul_75869_comb[0]};
  assign p1_concat_77096_comb = {p1_add_76784_comb, p1_smul_75874_comb[0]};
  assign p1_concat_77097_comb = {p1_add_76786_comb, p1_smul_75875_comb[0]};
  assign p1_concat_77098_comb = {p1_add_76788_comb, p1_smul_75880_comb[0]};
  assign p1_concat_77099_comb = {p1_add_76790_comb, p1_smul_75881_comb[0]};
  assign p1_concat_77100_comb = {p1_add_76792_comb, p1_smul_75886_comb[0]};
  assign p1_concat_77101_comb = {p1_add_76794_comb, p1_smul_75887_comb[0]};
  assign p1_concat_77102_comb = {p1_add_76796_comb, p1_smul_75892_comb[0]};
  assign p1_concat_77103_comb = {p1_add_76798_comb, p1_smul_75893_comb[0]};
  assign p1_sum__1756_comb = {{4{p1_concat_76800_comb[20]}}, p1_concat_76800_comb};
  assign p1_sum__1757_comb = {{4{p1_concat_76801_comb[20]}}, p1_concat_76801_comb};
  assign p1_sum__1758_comb = {{4{p1_concat_76802_comb[20]}}, p1_concat_76802_comb};
  assign p1_sum__1759_comb = {{4{p1_concat_76803_comb[20]}}, p1_concat_76803_comb};
  assign p1_sum__1732_comb = {{4{p1_concat_76804_comb[20]}}, p1_concat_76804_comb};
  assign p1_sum__1733_comb = {{4{p1_concat_76805_comb[20]}}, p1_concat_76805_comb};
  assign p1_sum__1734_comb = {{4{p1_concat_76806_comb[20]}}, p1_concat_76806_comb};
  assign p1_sum__1735_comb = {{4{p1_concat_76807_comb[20]}}, p1_concat_76807_comb};
  assign p1_sum__1704_comb = {{4{p1_concat_76808_comb[20]}}, p1_concat_76808_comb};
  assign p1_sum__1705_comb = {{4{p1_concat_76809_comb[20]}}, p1_concat_76809_comb};
  assign p1_sum__1706_comb = {{4{p1_concat_76810_comb[20]}}, p1_concat_76810_comb};
  assign p1_sum__1707_comb = {{4{p1_concat_76811_comb[20]}}, p1_concat_76811_comb};
  assign p1_sum__1676_comb = {{4{p1_concat_76812_comb[20]}}, p1_concat_76812_comb};
  assign p1_sum__1677_comb = {{4{p1_concat_76813_comb[20]}}, p1_concat_76813_comb};
  assign p1_sum__1678_comb = {{4{p1_concat_76814_comb[20]}}, p1_concat_76814_comb};
  assign p1_sum__1679_comb = {{4{p1_concat_76815_comb[20]}}, p1_concat_76815_comb};
  assign p1_sum__1736_comb = {{4{p1_add_76816_comb[20]}}, p1_add_76816_comb};
  assign p1_sum__1737_comb = {{4{p1_add_76817_comb[20]}}, p1_add_76817_comb};
  assign p1_sum__1738_comb = {{4{p1_add_76818_comb[20]}}, p1_add_76818_comb};
  assign p1_sum__1739_comb = {{4{p1_add_76819_comb[20]}}, p1_add_76819_comb};
  assign p1_sum__1708_comb = {{4{p1_add_76820_comb[20]}}, p1_add_76820_comb};
  assign p1_sum__1709_comb = {{4{p1_add_76821_comb[20]}}, p1_add_76821_comb};
  assign p1_sum__1710_comb = {{4{p1_add_76822_comb[20]}}, p1_add_76822_comb};
  assign p1_sum__1711_comb = {{4{p1_add_76823_comb[20]}}, p1_add_76823_comb};
  assign p1_sum__1680_comb = {{4{p1_add_76824_comb[20]}}, p1_add_76824_comb};
  assign p1_sum__1681_comb = {{4{p1_add_76825_comb[20]}}, p1_add_76825_comb};
  assign p1_sum__1682_comb = {{4{p1_add_76826_comb[20]}}, p1_add_76826_comb};
  assign p1_sum__1683_comb = {{4{p1_add_76827_comb[20]}}, p1_add_76827_comb};
  assign p1_sum__1652_comb = {{4{p1_add_76828_comb[20]}}, p1_add_76828_comb};
  assign p1_sum__1653_comb = {{4{p1_add_76829_comb[20]}}, p1_add_76829_comb};
  assign p1_sum__1654_comb = {{4{p1_add_76830_comb[20]}}, p1_add_76830_comb};
  assign p1_sum__1655_comb = {{4{p1_add_76831_comb[20]}}, p1_add_76831_comb};
  assign p1_sum__1712_comb = {{4{p1_concat_76832_comb[20]}}, p1_concat_76832_comb};
  assign p1_sum__1713_comb = {{4{p1_concat_76833_comb[20]}}, p1_concat_76833_comb};
  assign p1_sum__1714_comb = {{4{p1_concat_76834_comb[20]}}, p1_concat_76834_comb};
  assign p1_sum__1715_comb = {{4{p1_concat_76835_comb[20]}}, p1_concat_76835_comb};
  assign p1_sum__1684_comb = {{4{p1_concat_76836_comb[20]}}, p1_concat_76836_comb};
  assign p1_sum__1685_comb = {{4{p1_concat_76837_comb[20]}}, p1_concat_76837_comb};
  assign p1_sum__1686_comb = {{4{p1_concat_76838_comb[20]}}, p1_concat_76838_comb};
  assign p1_sum__1687_comb = {{4{p1_concat_76839_comb[20]}}, p1_concat_76839_comb};
  assign p1_sum__1656_comb = {{4{p1_concat_76840_comb[20]}}, p1_concat_76840_comb};
  assign p1_sum__1657_comb = {{4{p1_concat_76841_comb[20]}}, p1_concat_76841_comb};
  assign p1_sum__1658_comb = {{4{p1_concat_76842_comb[20]}}, p1_concat_76842_comb};
  assign p1_sum__1659_comb = {{4{p1_concat_76843_comb[20]}}, p1_concat_76843_comb};
  assign p1_sum__1632_comb = {{4{p1_concat_76844_comb[20]}}, p1_concat_76844_comb};
  assign p1_sum__1633_comb = {{4{p1_concat_76845_comb[20]}}, p1_concat_76845_comb};
  assign p1_sum__1634_comb = {{4{p1_concat_76846_comb[20]}}, p1_concat_76846_comb};
  assign p1_sum__1635_comb = {{4{p1_concat_76847_comb[20]}}, p1_concat_76847_comb};
  assign p1_concat_77152_comb = {p1_add_76848_comb, p1_smul_75992_comb[0]};
  assign p1_concat_77153_comb = {p1_add_76850_comb, p1_smul_75995_comb[0]};
  assign p1_concat_77154_comb = {p1_add_76852_comb, p1_smul_75998_comb[0]};
  assign p1_concat_77155_comb = {p1_add_76854_comb, p1_smul_76001_comb[0]};
  assign p1_concat_77156_comb = {p1_add_76856_comb, p1_smul_76002_comb[0]};
  assign p1_concat_77157_comb = {p1_add_76858_comb, p1_smul_76005_comb[0]};
  assign p1_concat_77158_comb = {p1_add_76860_comb, p1_smul_76008_comb[0]};
  assign p1_concat_77159_comb = {p1_add_76862_comb, p1_smul_76011_comb[0]};
  assign p1_concat_77160_comb = {p1_add_76864_comb, p1_smul_76012_comb[0]};
  assign p1_concat_77161_comb = {p1_add_76866_comb, p1_smul_76015_comb[0]};
  assign p1_concat_77162_comb = {p1_add_76868_comb, p1_smul_76018_comb[0]};
  assign p1_concat_77163_comb = {p1_add_76870_comb, p1_smul_76021_comb[0]};
  assign p1_concat_77164_comb = {p1_add_76872_comb, p1_smul_76022_comb[0]};
  assign p1_concat_77165_comb = {p1_add_76874_comb, p1_smul_76025_comb[0]};
  assign p1_concat_77166_comb = {p1_add_76876_comb, p1_smul_76028_comb[0]};
  assign p1_concat_77167_comb = {p1_add_76878_comb, p1_smul_76031_comb[0]};
  assign p1_add_77168_comb = {{4{p1_add_76496_comb[19]}}, p1_add_76496_comb} + {{4{p1_bit_slice_76497_comb[19]}}, p1_bit_slice_76497_comb};
  assign p1_add_77170_comb = {{4{p1_bit_slice_76498_comb[19]}}, p1_bit_slice_76498_comb} + {{4{p1_add_76499_comb[19]}}, p1_add_76499_comb};
  assign p1_add_77172_comb = {{4{p1_add_76500_comb[19]}}, p1_add_76500_comb} + {{4{p1_bit_slice_76501_comb[19]}}, p1_bit_slice_76501_comb};
  assign p1_add_77174_comb = {{4{p1_bit_slice_76502_comb[19]}}, p1_bit_slice_76502_comb} + {{4{p1_add_76503_comb[19]}}, p1_add_76503_comb};
  assign p1_add_77176_comb = {{4{p1_add_76504_comb[19]}}, p1_add_76504_comb} + {{4{p1_bit_slice_76505_comb[19]}}, p1_bit_slice_76505_comb};
  assign p1_add_77178_comb = {{4{p1_bit_slice_76506_comb[19]}}, p1_bit_slice_76506_comb} + {{4{p1_add_76507_comb[19]}}, p1_add_76507_comb};
  assign p1_add_77180_comb = {{4{p1_add_76508_comb[19]}}, p1_add_76508_comb} + {{4{p1_bit_slice_76509_comb[19]}}, p1_bit_slice_76509_comb};
  assign p1_add_77182_comb = {{4{p1_bit_slice_76510_comb[19]}}, p1_bit_slice_76510_comb} + {{4{p1_add_76511_comb[19]}}, p1_add_76511_comb};
  assign p1_add_77192_comb = {{4{p1_bit_slice_76528_comb[19]}}, p1_bit_slice_76528_comb} + {{4{p1_add_76529_comb[19]}}, p1_add_76529_comb};
  assign p1_add_77194_comb = {{4{p1_add_76530_comb[19]}}, p1_add_76530_comb} + {{4{p1_bit_slice_76531_comb[19]}}, p1_bit_slice_76531_comb};
  assign p1_add_77196_comb = {{4{p1_bit_slice_76532_comb[19]}}, p1_bit_slice_76532_comb} + {{4{p1_add_76533_comb[19]}}, p1_add_76533_comb};
  assign p1_add_77198_comb = {{4{p1_add_76534_comb[19]}}, p1_add_76534_comb} + {{4{p1_bit_slice_76535_comb[19]}}, p1_bit_slice_76535_comb};
  assign p1_concat_77200_comb = {p1_add_76912_comb, p1_smul_76070_comb[0]};
  assign p1_concat_77201_comb = {p1_add_76914_comb, p1_smul_76071_comb[0]};
  assign p1_concat_77202_comb = {p1_add_76916_comb, p1_smul_76076_comb[0]};
  assign p1_concat_77203_comb = {p1_add_76918_comb, p1_smul_76077_comb[0]};
  assign p1_concat_77204_comb = {p1_add_76920_comb, p1_smul_76082_comb[0]};
  assign p1_concat_77205_comb = {p1_add_76922_comb, p1_smul_76083_comb[0]};
  assign p1_concat_77206_comb = {p1_add_76924_comb, p1_smul_76088_comb[0]};
  assign p1_concat_77207_comb = {p1_add_76926_comb, p1_smul_76089_comb[0]};
  assign p1_sum__1776_comb = {{4{p1_concat_76928_comb[20]}}, p1_concat_76928_comb};
  assign p1_sum__1777_comb = {{4{p1_concat_76929_comb[20]}}, p1_concat_76929_comb};
  assign p1_sum__1778_comb = {{4{p1_concat_76930_comb[20]}}, p1_concat_76930_comb};
  assign p1_sum__1779_comb = {{4{p1_concat_76931_comb[20]}}, p1_concat_76931_comb};
  assign p1_sum__1648_comb = {{4{p1_concat_76932_comb[20]}}, p1_concat_76932_comb};
  assign p1_sum__1649_comb = {{4{p1_concat_76933_comb[20]}}, p1_concat_76933_comb};
  assign p1_sum__1650_comb = {{4{p1_concat_76934_comb[20]}}, p1_concat_76934_comb};
  assign p1_sum__1651_comb = {{4{p1_concat_76935_comb[20]}}, p1_concat_76935_comb};
  assign p1_sum__1760_comb = {{4{p1_add_76936_comb[20]}}, p1_add_76936_comb};
  assign p1_sum__1761_comb = {{4{p1_add_76937_comb[20]}}, p1_add_76937_comb};
  assign p1_sum__1762_comb = {{4{p1_add_76938_comb[20]}}, p1_add_76938_comb};
  assign p1_sum__1763_comb = {{4{p1_add_76939_comb[20]}}, p1_add_76939_comb};
  assign p1_sum__1628_comb = {{4{p1_add_76940_comb[20]}}, p1_add_76940_comb};
  assign p1_sum__1629_comb = {{4{p1_add_76941_comb[20]}}, p1_add_76941_comb};
  assign p1_sum__1630_comb = {{4{p1_add_76942_comb[20]}}, p1_add_76942_comb};
  assign p1_sum__1631_comb = {{4{p1_add_76943_comb[20]}}, p1_add_76943_comb};
  assign p1_sum__1740_comb = {{4{p1_concat_76944_comb[20]}}, p1_concat_76944_comb};
  assign p1_sum__1741_comb = {{4{p1_concat_76945_comb[20]}}, p1_concat_76945_comb};
  assign p1_sum__1742_comb = {{4{p1_concat_76946_comb[20]}}, p1_concat_76946_comb};
  assign p1_sum__1743_comb = {{4{p1_concat_76947_comb[20]}}, p1_concat_76947_comb};
  assign p1_sum__1612_comb = {{4{p1_concat_76948_comb[20]}}, p1_concat_76948_comb};
  assign p1_sum__1613_comb = {{4{p1_concat_76949_comb[20]}}, p1_concat_76949_comb};
  assign p1_sum__1614_comb = {{4{p1_concat_76950_comb[20]}}, p1_concat_76950_comb};
  assign p1_sum__1615_comb = {{4{p1_concat_76951_comb[20]}}, p1_concat_76951_comb};
  assign p1_concat_77232_comb = {p1_add_76952_comb, p1_smul_76140_comb[0]};
  assign p1_concat_77233_comb = {p1_add_76954_comb, p1_smul_76143_comb[0]};
  assign p1_concat_77234_comb = {p1_add_76956_comb, p1_smul_76146_comb[0]};
  assign p1_concat_77235_comb = {p1_add_76958_comb, p1_smul_76149_comb[0]};
  assign p1_concat_77236_comb = {p1_add_76960_comb, p1_smul_76150_comb[0]};
  assign p1_concat_77237_comb = {p1_add_76962_comb, p1_smul_76153_comb[0]};
  assign p1_concat_77238_comb = {p1_add_76964_comb, p1_smul_76156_comb[0]};
  assign p1_concat_77239_comb = {p1_add_76966_comb, p1_smul_76159_comb[0]};
  assign p1_add_77240_comb = {{4{p1_add_76616_comb[19]}}, p1_add_76616_comb} + {{4{p1_bit_slice_76617_comb[19]}}, p1_bit_slice_76617_comb};
  assign p1_add_77242_comb = {{4{p1_bit_slice_76618_comb[19]}}, p1_bit_slice_76618_comb} + {{4{p1_add_76619_comb[19]}}, p1_add_76619_comb};
  assign p1_add_77244_comb = {{4{p1_add_76620_comb[19]}}, p1_add_76620_comb} + {{4{p1_bit_slice_76621_comb[19]}}, p1_bit_slice_76621_comb};
  assign p1_add_77246_comb = {{4{p1_bit_slice_76622_comb[19]}}, p1_bit_slice_76622_comb} + {{4{p1_add_76623_comb[19]}}, p1_add_76623_comb};
  assign p1_add_77256_comb = {{4{p1_bit_slice_76640_comb[19]}}, p1_bit_slice_76640_comb} + {{4{p1_add_76641_comb[19]}}, p1_add_76641_comb};
  assign p1_add_77258_comb = {{4{p1_add_76642_comb[19]}}, p1_add_76642_comb} + {{4{p1_bit_slice_76643_comb[19]}}, p1_bit_slice_76643_comb};
  assign p1_add_77260_comb = {{4{p1_bit_slice_76644_comb[19]}}, p1_bit_slice_76644_comb} + {{4{p1_add_76645_comb[19]}}, p1_add_76645_comb};
  assign p1_add_77262_comb = {{4{p1_add_76646_comb[19]}}, p1_add_76646_comb} + {{4{p1_bit_slice_76647_comb[19]}}, p1_bit_slice_76647_comb};
  assign p1_concat_77264_comb = {p1_add_76992_comb, p1_smul_76186_comb[0]};
  assign p1_concat_77265_comb = {p1_add_76994_comb, p1_smul_76187_comb[0]};
  assign p1_concat_77266_comb = {p1_add_76996_comb, p1_smul_76192_comb[0]};
  assign p1_concat_77267_comb = {p1_add_76998_comb, p1_smul_76193_comb[0]};
  assign p1_concat_77268_comb = {p1_add_77000_comb, p1_smul_76198_comb[0]};
  assign p1_concat_77269_comb = {p1_add_77002_comb, p1_smul_76199_comb[0]};
  assign p1_concat_77270_comb = {p1_add_77004_comb, p1_smul_76204_comb[0]};
  assign p1_concat_77271_comb = {p1_add_77006_comb, p1_smul_76205_comb[0]};
  assign p1_sum__1792_comb = {{4{p1_concat_77008_comb[20]}}, p1_concat_77008_comb};
  assign p1_sum__1793_comb = {{4{p1_concat_77009_comb[20]}}, p1_concat_77009_comb};
  assign p1_sum__1794_comb = {{4{p1_concat_77010_comb[20]}}, p1_concat_77010_comb};
  assign p1_sum__1795_comb = {{4{p1_concat_77011_comb[20]}}, p1_concat_77011_comb};
  assign p1_sum__1624_comb = {{4{p1_concat_77012_comb[20]}}, p1_concat_77012_comb};
  assign p1_sum__1625_comb = {{4{p1_concat_77013_comb[20]}}, p1_concat_77013_comb};
  assign p1_sum__1626_comb = {{4{p1_concat_77014_comb[20]}}, p1_concat_77014_comb};
  assign p1_sum__1627_comb = {{4{p1_concat_77015_comb[20]}}, p1_concat_77015_comb};
  assign p1_sum__1780_comb = {{4{p1_add_77016_comb[20]}}, p1_add_77016_comb};
  assign p1_sum__1781_comb = {{4{p1_add_77017_comb[20]}}, p1_add_77017_comb};
  assign p1_sum__1782_comb = {{4{p1_add_77018_comb[20]}}, p1_add_77018_comb};
  assign p1_sum__1783_comb = {{4{p1_add_77019_comb[20]}}, p1_add_77019_comb};
  assign p1_sum__1608_comb = {{4{p1_add_77020_comb[20]}}, p1_add_77020_comb};
  assign p1_sum__1609_comb = {{4{p1_add_77021_comb[20]}}, p1_add_77021_comb};
  assign p1_sum__1610_comb = {{4{p1_add_77022_comb[20]}}, p1_add_77022_comb};
  assign p1_sum__1611_comb = {{4{p1_add_77023_comb[20]}}, p1_add_77023_comb};
  assign p1_sum__1764_comb = {{4{p1_concat_77024_comb[20]}}, p1_concat_77024_comb};
  assign p1_sum__1765_comb = {{4{p1_concat_77025_comb[20]}}, p1_concat_77025_comb};
  assign p1_sum__1766_comb = {{4{p1_concat_77026_comb[20]}}, p1_concat_77026_comb};
  assign p1_sum__1767_comb = {{4{p1_concat_77027_comb[20]}}, p1_concat_77027_comb};
  assign p1_sum__1596_comb = {{4{p1_concat_77028_comb[20]}}, p1_concat_77028_comb};
  assign p1_sum__1597_comb = {{4{p1_concat_77029_comb[20]}}, p1_concat_77029_comb};
  assign p1_sum__1598_comb = {{4{p1_concat_77030_comb[20]}}, p1_concat_77030_comb};
  assign p1_sum__1599_comb = {{4{p1_concat_77031_comb[20]}}, p1_concat_77031_comb};
  assign p1_concat_77296_comb = {p1_add_77032_comb, p1_smul_76256_comb[0]};
  assign p1_concat_77297_comb = {p1_add_77034_comb, p1_smul_76259_comb[0]};
  assign p1_concat_77298_comb = {p1_add_77036_comb, p1_smul_76262_comb[0]};
  assign p1_concat_77299_comb = {p1_add_77038_comb, p1_smul_76265_comb[0]};
  assign p1_concat_77300_comb = {p1_add_77040_comb, p1_smul_76266_comb[0]};
  assign p1_concat_77301_comb = {p1_add_77042_comb, p1_smul_76269_comb[0]};
  assign p1_concat_77302_comb = {p1_add_77044_comb, p1_smul_76272_comb[0]};
  assign p1_concat_77303_comb = {p1_add_77046_comb, p1_smul_76275_comb[0]};
  assign p1_add_77304_comb = {{4{p1_add_76728_comb[19]}}, p1_add_76728_comb} + {{4{p1_bit_slice_76729_comb[19]}}, p1_bit_slice_76729_comb};
  assign p1_add_77306_comb = {{4{p1_bit_slice_76730_comb[19]}}, p1_bit_slice_76730_comb} + {{4{p1_add_76731_comb[19]}}, p1_add_76731_comb};
  assign p1_add_77308_comb = {{4{p1_add_76732_comb[19]}}, p1_add_76732_comb} + {{4{p1_bit_slice_76733_comb[19]}}, p1_bit_slice_76733_comb};
  assign p1_add_77310_comb = {{4{p1_bit_slice_76734_comb[19]}}, p1_bit_slice_76734_comb} + {{4{p1_add_76735_comb[19]}}, p1_add_76735_comb};
  assign p1_add_77312_comb = {{11{p1_add_76736_comb[12]}}, p1_add_76736_comb} + {{11{p1_add_76737_comb[12]}}, p1_add_76737_comb};
  assign p1_add_77313_comb = {{11{p1_add_76738_comb[12]}}, p1_add_76738_comb} + {{11{p1_add_76739_comb[12]}}, p1_add_76739_comb};
  assign p1_add_77314_comb = {{11{p1_add_76740_comb[12]}}, p1_add_76740_comb} + {{11{p1_add_76741_comb[12]}}, p1_add_76741_comb};
  assign p1_add_77315_comb = {{11{p1_add_76742_comb[12]}}, p1_add_76742_comb} + {{11{p1_add_76743_comb[12]}}, p1_add_76743_comb};
  assign p1_add_77316_comb = {{11{p1_add_76744_comb[12]}}, p1_add_76744_comb} + {{11{p1_add_76745_comb[12]}}, p1_add_76745_comb};
  assign p1_add_77317_comb = {{11{p1_add_76746_comb[12]}}, p1_add_76746_comb} + {{11{p1_add_76747_comb[12]}}, p1_add_76747_comb};
  assign p1_add_77318_comb = {{11{p1_add_76748_comb[12]}}, p1_add_76748_comb} + {{11{p1_add_76749_comb[12]}}, p1_add_76749_comb};
  assign p1_add_77319_comb = {{11{p1_add_76750_comb[12]}}, p1_add_76750_comb} + {{11{p1_add_76751_comb[12]}}, p1_add_76751_comb};
  assign p1_sum__1348_comb = {p1_add_77072_comb, p1_add_75824_comb[0]};
  assign p1_sum__1349_comb = {p1_add_77074_comb, p1_add_75829_comb[0]};
  assign p1_sum__1340_comb = {p1_add_77076_comb, p1_add_75830_comb[0]};
  assign p1_sum__1341_comb = {p1_add_77078_comb, p1_add_75835_comb[0]};
  assign p1_sum__1330_comb = {p1_add_77080_comb, p1_add_75836_comb[0]};
  assign p1_sum__1331_comb = {p1_add_77082_comb, p1_add_75841_comb[0]};
  assign p1_sum__1318_comb = {p1_add_77084_comb, p1_add_75842_comb[0]};
  assign p1_sum__1319_comb = {p1_add_77086_comb, p1_add_75847_comb[0]};
  assign p1_sum__1334_comb = p1_sum__1756_comb + p1_sum__1757_comb;
  assign p1_sum__1335_comb = p1_sum__1758_comb + p1_sum__1759_comb;
  assign p1_sum__1322_comb = p1_sum__1732_comb + p1_sum__1733_comb;
  assign p1_sum__1323_comb = p1_sum__1734_comb + p1_sum__1735_comb;
  assign p1_sum__1308_comb = p1_sum__1704_comb + p1_sum__1705_comb;
  assign p1_sum__1309_comb = p1_sum__1706_comb + p1_sum__1707_comb;
  assign p1_sum__1294_comb = p1_sum__1676_comb + p1_sum__1677_comb;
  assign p1_sum__1295_comb = p1_sum__1678_comb + p1_sum__1679_comb;
  assign p1_sum__1324_comb = p1_sum__1736_comb + p1_sum__1737_comb;
  assign p1_sum__1325_comb = p1_sum__1738_comb + p1_sum__1739_comb;
  assign p1_sum__1310_comb = p1_sum__1708_comb + p1_sum__1709_comb;
  assign p1_sum__1311_comb = p1_sum__1710_comb + p1_sum__1711_comb;
  assign p1_sum__1296_comb = p1_sum__1680_comb + p1_sum__1681_comb;
  assign p1_sum__1297_comb = p1_sum__1682_comb + p1_sum__1683_comb;
  assign p1_sum__1282_comb = p1_sum__1652_comb + p1_sum__1653_comb;
  assign p1_sum__1283_comb = p1_sum__1654_comb + p1_sum__1655_comb;
  assign p1_sum__1312_comb = p1_sum__1712_comb + p1_sum__1713_comb;
  assign p1_sum__1313_comb = p1_sum__1714_comb + p1_sum__1715_comb;
  assign p1_sum__1298_comb = p1_sum__1684_comb + p1_sum__1685_comb;
  assign p1_sum__1299_comb = p1_sum__1686_comb + p1_sum__1687_comb;
  assign p1_sum__1284_comb = p1_sum__1656_comb + p1_sum__1657_comb;
  assign p1_sum__1285_comb = p1_sum__1658_comb + p1_sum__1659_comb;
  assign p1_sum__1272_comb = p1_sum__1632_comb + p1_sum__1633_comb;
  assign p1_sum__1273_comb = p1_sum__1634_comb + p1_sum__1635_comb;
  assign p1_sum__1288_comb = {p1_add_77168_comb, p1_add_76034_comb[0]};
  assign p1_sum__1289_comb = {p1_add_77170_comb, p1_add_76035_comb[0]};
  assign p1_sum__1276_comb = {p1_add_77172_comb, p1_add_76040_comb[0]};
  assign p1_sum__1277_comb = {p1_add_77174_comb, p1_add_76041_comb[0]};
  assign p1_sum__1266_comb = {p1_add_77176_comb, p1_add_76046_comb[0]};
  assign p1_sum__1267_comb = {p1_add_77178_comb, p1_add_76047_comb[0]};
  assign p1_sum__1258_comb = {p1_add_77180_comb, p1_add_76052_comb[0]};
  assign p1_sum__1259_comb = {p1_add_77182_comb, p1_add_76053_comb[0]};
  assign p1_add_77392_comb = {{11{p1_add_76896_comb[12]}}, p1_add_76896_comb} + {{11{p1_add_76897_comb[12]}}, p1_add_76897_comb};
  assign p1_add_77393_comb = {{11{p1_add_76898_comb[12]}}, p1_add_76898_comb} + {{11{p1_add_76899_comb[12]}}, p1_add_76899_comb};
  assign p1_add_77394_comb = {{11{p1_add_76900_comb[12]}}, p1_add_76900_comb} + {{11{p1_add_76901_comb[12]}}, p1_add_76901_comb};
  assign p1_add_77395_comb = {{11{p1_add_76902_comb[12]}}, p1_add_76902_comb} + {{11{p1_add_76903_comb[12]}}, p1_add_76903_comb};
  assign p1_sum__1354_comb = {p1_add_77192_comb, p1_add_76056_comb[0]};
  assign p1_sum__1355_comb = {p1_add_77194_comb, p1_add_76061_comb[0]};
  assign p1_sum__1304_comb = {p1_add_77196_comb, p1_add_76062_comb[0]};
  assign p1_sum__1305_comb = {p1_add_77198_comb, p1_add_76067_comb[0]};
  assign p1_sum__1344_comb = p1_sum__1776_comb + p1_sum__1777_comb;
  assign p1_sum__1345_comb = p1_sum__1778_comb + p1_sum__1779_comb;
  assign p1_sum__1280_comb = p1_sum__1648_comb + p1_sum__1649_comb;
  assign p1_sum__1281_comb = p1_sum__1650_comb + p1_sum__1651_comb;
  assign p1_sum__1336_comb = p1_sum__1760_comb + p1_sum__1761_comb;
  assign p1_sum__1337_comb = p1_sum__1762_comb + p1_sum__1763_comb;
  assign p1_sum__1270_comb = p1_sum__1628_comb + p1_sum__1629_comb;
  assign p1_sum__1271_comb = p1_sum__1630_comb + p1_sum__1631_comb;
  assign p1_sum__1326_comb = p1_sum__1740_comb + p1_sum__1741_comb;
  assign p1_sum__1327_comb = p1_sum__1742_comb + p1_sum__1743_comb;
  assign p1_sum__1262_comb = p1_sum__1612_comb + p1_sum__1613_comb;
  assign p1_sum__1263_comb = p1_sum__1614_comb + p1_sum__1615_comb;
  assign p1_sum__1302_comb = {p1_add_77240_comb, p1_add_76162_comb[0]};
  assign p1_sum__1303_comb = {p1_add_77242_comb, p1_add_76163_comb[0]};
  assign p1_sum__1252_comb = {p1_add_77244_comb, p1_add_76168_comb[0]};
  assign p1_sum__1253_comb = {p1_add_77246_comb, p1_add_76169_comb[0]};
  assign p1_add_77432_comb = {{11{p1_add_76976_comb[12]}}, p1_add_76976_comb} + {{11{p1_add_76977_comb[12]}}, p1_add_76977_comb};
  assign p1_add_77433_comb = {{11{p1_add_76978_comb[12]}}, p1_add_76978_comb} + {{11{p1_add_76979_comb[12]}}, p1_add_76979_comb};
  assign p1_add_77434_comb = {{11{p1_add_76980_comb[12]}}, p1_add_76980_comb} + {{11{p1_add_76981_comb[12]}}, p1_add_76981_comb};
  assign p1_add_77435_comb = {{11{p1_add_76982_comb[12]}}, p1_add_76982_comb} + {{11{p1_add_76983_comb[12]}}, p1_add_76983_comb};
  assign p1_sum__1358_comb = {p1_add_77256_comb, p1_add_76172_comb[0]};
  assign p1_sum__1359_comb = {p1_add_77258_comb, p1_add_76177_comb[0]};
  assign p1_sum__1290_comb = {p1_add_77260_comb, p1_add_76178_comb[0]};
  assign p1_sum__1291_comb = {p1_add_77262_comb, p1_add_76183_comb[0]};
  assign p1_sum__1352_comb = p1_sum__1792_comb + p1_sum__1793_comb;
  assign p1_sum__1353_comb = p1_sum__1794_comb + p1_sum__1795_comb;
  assign p1_sum__1268_comb = p1_sum__1624_comb + p1_sum__1625_comb;
  assign p1_sum__1269_comb = p1_sum__1626_comb + p1_sum__1627_comb;
  assign p1_sum__1346_comb = p1_sum__1780_comb + p1_sum__1781_comb;
  assign p1_sum__1347_comb = p1_sum__1782_comb + p1_sum__1783_comb;
  assign p1_sum__1260_comb = p1_sum__1608_comb + p1_sum__1609_comb;
  assign p1_sum__1261_comb = p1_sum__1610_comb + p1_sum__1611_comb;
  assign p1_sum__1338_comb = p1_sum__1764_comb + p1_sum__1765_comb;
  assign p1_sum__1339_comb = p1_sum__1766_comb + p1_sum__1767_comb;
  assign p1_sum__1254_comb = p1_sum__1596_comb + p1_sum__1597_comb;
  assign p1_sum__1255_comb = p1_sum__1598_comb + p1_sum__1599_comb;
  assign p1_sum__1316_comb = {p1_add_77304_comb, p1_add_76278_comb[0]};
  assign p1_sum__1317_comb = {p1_add_77306_comb, p1_add_76279_comb[0]};
  assign p1_sum__1248_comb = {p1_add_77308_comb, p1_add_76284_comb[0]};
  assign p1_sum__1249_comb = {p1_add_77310_comb, p1_add_76285_comb[0]};
  assign p1_add_77472_comb = p1_add_77312_comb + p1_add_77313_comb;
  assign p1_add_77474_comb = p1_add_77314_comb + p1_add_77315_comb;
  assign p1_add_77476_comb = p1_add_77316_comb + p1_add_77317_comb;
  assign p1_add_77478_comb = p1_add_77318_comb + p1_add_77319_comb;
  assign p1_sum__1130_comb = p1_sum__1348_comb + p1_sum__1349_comb;
  assign p1_sum__1126_comb = p1_sum__1340_comb + p1_sum__1341_comb;
  assign p1_sum__1121_comb = p1_sum__1330_comb + p1_sum__1331_comb;
  assign p1_sum__1115_comb = p1_sum__1318_comb + p1_sum__1319_comb;
  assign p1_add_77488_comb = {{4{p1_concat_77088_comb[19]}}, p1_concat_77088_comb} + {{4{p1_concat_77089_comb[19]}}, p1_concat_77089_comb};
  assign p1_add_77489_comb = {{4{p1_concat_77090_comb[19]}}, p1_concat_77090_comb} + {{4{p1_concat_77091_comb[19]}}, p1_concat_77091_comb};
  assign p1_add_77490_comb = {{4{p1_concat_77092_comb[19]}}, p1_concat_77092_comb} + {{4{p1_concat_77093_comb[19]}}, p1_concat_77093_comb};
  assign p1_add_77491_comb = {{4{p1_concat_77094_comb[19]}}, p1_concat_77094_comb} + {{4{p1_concat_77095_comb[19]}}, p1_concat_77095_comb};
  assign p1_add_77492_comb = {{4{p1_concat_77096_comb[19]}}, p1_concat_77096_comb} + {{4{p1_concat_77097_comb[19]}}, p1_concat_77097_comb};
  assign p1_add_77493_comb = {{4{p1_concat_77098_comb[19]}}, p1_concat_77098_comb} + {{4{p1_concat_77099_comb[19]}}, p1_concat_77099_comb};
  assign p1_add_77494_comb = {{4{p1_concat_77100_comb[19]}}, p1_concat_77100_comb} + {{4{p1_concat_77101_comb[19]}}, p1_concat_77101_comb};
  assign p1_add_77495_comb = {{4{p1_concat_77102_comb[19]}}, p1_concat_77102_comb} + {{4{p1_concat_77103_comb[19]}}, p1_concat_77103_comb};
  assign p1_sum__1123_comb = p1_sum__1334_comb + p1_sum__1335_comb;
  assign p1_sum__1117_comb = p1_sum__1322_comb + p1_sum__1323_comb;
  assign p1_sum__1110_comb = p1_sum__1308_comb + p1_sum__1309_comb;
  assign p1_sum__1103_comb = p1_sum__1294_comb + p1_sum__1295_comb;
  assign p1_sum__1118_comb = p1_sum__1324_comb + p1_sum__1325_comb;
  assign p1_sum__1111_comb = p1_sum__1310_comb + p1_sum__1311_comb;
  assign p1_sum__1104_comb = p1_sum__1296_comb + p1_sum__1297_comb;
  assign p1_sum__1097_comb = p1_sum__1282_comb + p1_sum__1283_comb;
  assign p1_sum__1112_comb = p1_sum__1312_comb + p1_sum__1313_comb;
  assign p1_sum__1105_comb = p1_sum__1298_comb + p1_sum__1299_comb;
  assign p1_sum__1098_comb = p1_sum__1284_comb + p1_sum__1285_comb;
  assign p1_sum__1092_comb = p1_sum__1272_comb + p1_sum__1273_comb;
  assign p1_add_77520_comb = {{4{p1_concat_77152_comb[19]}}, p1_concat_77152_comb} + {{4{p1_concat_77153_comb[19]}}, p1_concat_77153_comb};
  assign p1_add_77521_comb = {{4{p1_concat_77154_comb[19]}}, p1_concat_77154_comb} + {{4{p1_concat_77155_comb[19]}}, p1_concat_77155_comb};
  assign p1_add_77522_comb = {{4{p1_concat_77156_comb[19]}}, p1_concat_77156_comb} + {{4{p1_concat_77157_comb[19]}}, p1_concat_77157_comb};
  assign p1_add_77523_comb = {{4{p1_concat_77158_comb[19]}}, p1_concat_77158_comb} + {{4{p1_concat_77159_comb[19]}}, p1_concat_77159_comb};
  assign p1_add_77524_comb = {{4{p1_concat_77160_comb[19]}}, p1_concat_77160_comb} + {{4{p1_concat_77161_comb[19]}}, p1_concat_77161_comb};
  assign p1_add_77525_comb = {{4{p1_concat_77162_comb[19]}}, p1_concat_77162_comb} + {{4{p1_concat_77163_comb[19]}}, p1_concat_77163_comb};
  assign p1_add_77526_comb = {{4{p1_concat_77164_comb[19]}}, p1_concat_77164_comb} + {{4{p1_concat_77165_comb[19]}}, p1_concat_77165_comb};
  assign p1_add_77527_comb = {{4{p1_concat_77166_comb[19]}}, p1_concat_77166_comb} + {{4{p1_concat_77167_comb[19]}}, p1_concat_77167_comb};
  assign p1_sum__1100_comb = p1_sum__1288_comb + p1_sum__1289_comb;
  assign p1_sum__1094_comb = p1_sum__1276_comb + p1_sum__1277_comb;
  assign p1_sum__1089_comb = p1_sum__1266_comb + p1_sum__1267_comb;
  assign p1_sum__1085_comb = p1_sum__1258_comb + p1_sum__1259_comb;
  assign p1_add_77536_comb = p1_add_77392_comb + p1_add_77393_comb;
  assign p1_add_77538_comb = p1_add_77394_comb + p1_add_77395_comb;
  assign p1_sum__1133_comb = p1_sum__1354_comb + p1_sum__1355_comb;
  assign p1_sum__1108_comb = p1_sum__1304_comb + p1_sum__1305_comb;
  assign p1_add_77544_comb = {{4{p1_concat_77200_comb[19]}}, p1_concat_77200_comb} + {{4{p1_concat_77201_comb[19]}}, p1_concat_77201_comb};
  assign p1_add_77545_comb = {{4{p1_concat_77202_comb[19]}}, p1_concat_77202_comb} + {{4{p1_concat_77203_comb[19]}}, p1_concat_77203_comb};
  assign p1_add_77546_comb = {{4{p1_concat_77204_comb[19]}}, p1_concat_77204_comb} + {{4{p1_concat_77205_comb[19]}}, p1_concat_77205_comb};
  assign p1_add_77547_comb = {{4{p1_concat_77206_comb[19]}}, p1_concat_77206_comb} + {{4{p1_concat_77207_comb[19]}}, p1_concat_77207_comb};
  assign p1_sum__1128_comb = p1_sum__1344_comb + p1_sum__1345_comb;
  assign p1_sum__1096_comb = p1_sum__1280_comb + p1_sum__1281_comb;
  assign p1_sum__1124_comb = p1_sum__1336_comb + p1_sum__1337_comb;
  assign p1_sum__1091_comb = p1_sum__1270_comb + p1_sum__1271_comb;
  assign p1_sum__1119_comb = p1_sum__1326_comb + p1_sum__1327_comb;
  assign p1_sum__1087_comb = p1_sum__1262_comb + p1_sum__1263_comb;
  assign p1_add_77560_comb = {{4{p1_concat_77232_comb[19]}}, p1_concat_77232_comb} + {{4{p1_concat_77233_comb[19]}}, p1_concat_77233_comb};
  assign p1_add_77561_comb = {{4{p1_concat_77234_comb[19]}}, p1_concat_77234_comb} + {{4{p1_concat_77235_comb[19]}}, p1_concat_77235_comb};
  assign p1_add_77562_comb = {{4{p1_concat_77236_comb[19]}}, p1_concat_77236_comb} + {{4{p1_concat_77237_comb[19]}}, p1_concat_77237_comb};
  assign p1_add_77563_comb = {{4{p1_concat_77238_comb[19]}}, p1_concat_77238_comb} + {{4{p1_concat_77239_comb[19]}}, p1_concat_77239_comb};
  assign p1_sum__1107_comb = p1_sum__1302_comb + p1_sum__1303_comb;
  assign p1_sum__1082_comb = p1_sum__1252_comb + p1_sum__1253_comb;
  assign p1_add_77568_comb = p1_add_77432_comb + p1_add_77433_comb;
  assign p1_add_77570_comb = p1_add_77434_comb + p1_add_77435_comb;
  assign p1_sum__1135_comb = p1_sum__1358_comb + p1_sum__1359_comb;
  assign p1_sum__1101_comb = p1_sum__1290_comb + p1_sum__1291_comb;
  assign p1_add_77576_comb = {{4{p1_concat_77264_comb[19]}}, p1_concat_77264_comb} + {{4{p1_concat_77265_comb[19]}}, p1_concat_77265_comb};
  assign p1_add_77577_comb = {{4{p1_concat_77266_comb[19]}}, p1_concat_77266_comb} + {{4{p1_concat_77267_comb[19]}}, p1_concat_77267_comb};
  assign p1_add_77578_comb = {{4{p1_concat_77268_comb[19]}}, p1_concat_77268_comb} + {{4{p1_concat_77269_comb[19]}}, p1_concat_77269_comb};
  assign p1_add_77579_comb = {{4{p1_concat_77270_comb[19]}}, p1_concat_77270_comb} + {{4{p1_concat_77271_comb[19]}}, p1_concat_77271_comb};
  assign p1_sum__1132_comb = p1_sum__1352_comb + p1_sum__1353_comb;
  assign p1_sum__1090_comb = p1_sum__1268_comb + p1_sum__1269_comb;
  assign p1_sum__1129_comb = p1_sum__1346_comb + p1_sum__1347_comb;
  assign p1_sum__1086_comb = p1_sum__1260_comb + p1_sum__1261_comb;
  assign p1_sum__1125_comb = p1_sum__1338_comb + p1_sum__1339_comb;
  assign p1_sum__1083_comb = p1_sum__1254_comb + p1_sum__1255_comb;
  assign p1_add_77592_comb = {{4{p1_concat_77296_comb[19]}}, p1_concat_77296_comb} + {{4{p1_concat_77297_comb[19]}}, p1_concat_77297_comb};
  assign p1_add_77593_comb = {{4{p1_concat_77298_comb[19]}}, p1_concat_77298_comb} + {{4{p1_concat_77299_comb[19]}}, p1_concat_77299_comb};
  assign p1_add_77594_comb = {{4{p1_concat_77300_comb[19]}}, p1_concat_77300_comb} + {{4{p1_concat_77301_comb[19]}}, p1_concat_77301_comb};
  assign p1_add_77595_comb = {{4{p1_concat_77302_comb[19]}}, p1_concat_77302_comb} + {{4{p1_concat_77303_comb[19]}}, p1_concat_77303_comb};
  assign p1_sum__1114_comb = p1_sum__1316_comb + p1_sum__1317_comb;
  assign p1_sum__1080_comb = p1_sum__1248_comb + p1_sum__1249_comb;
  assign p1_umul_27340_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_77472_comb, 7'h5b);
  assign p1_umul_27342_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_77474_comb, 7'h5b);
  assign p1_umul_27344_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_77476_comb, 7'h5b);
  assign p1_umul_27346_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_77478_comb, 7'h5b);
  assign p1_add_77604_comb = p1_sum__1130_comb + 25'h000_0001;
  assign p1_add_77605_comb = p1_sum__1126_comb + 25'h000_0001;
  assign p1_add_77606_comb = p1_sum__1121_comb + 25'h000_0001;
  assign p1_add_77607_comb = p1_sum__1115_comb + 25'h000_0001;
  assign p1_add_77608_comb = p1_add_77488_comb + p1_add_77489_comb;
  assign p1_add_77609_comb = p1_add_77490_comb + p1_add_77491_comb;
  assign p1_add_77610_comb = p1_add_77492_comb + p1_add_77493_comb;
  assign p1_add_77611_comb = p1_add_77494_comb + p1_add_77495_comb;
  assign p1_add_77612_comb = p1_sum__1123_comb + 25'h000_0001;
  assign p1_add_77613_comb = p1_sum__1117_comb + 25'h000_0001;
  assign p1_add_77614_comb = p1_sum__1110_comb + 25'h000_0001;
  assign p1_add_77615_comb = p1_sum__1103_comb + 25'h000_0001;
  assign p1_add_77616_comb = p1_sum__1118_comb + 25'h000_0001;
  assign p1_add_77617_comb = p1_sum__1111_comb + 25'h000_0001;
  assign p1_add_77618_comb = p1_sum__1104_comb + 25'h000_0001;
  assign p1_add_77619_comb = p1_sum__1097_comb + 25'h000_0001;
  assign p1_add_77620_comb = p1_sum__1112_comb + 25'h000_0001;
  assign p1_add_77621_comb = p1_sum__1105_comb + 25'h000_0001;
  assign p1_add_77622_comb = p1_sum__1098_comb + 25'h000_0001;
  assign p1_add_77623_comb = p1_sum__1092_comb + 25'h000_0001;
  assign p1_add_77624_comb = p1_add_77520_comb + p1_add_77521_comb;
  assign p1_add_77625_comb = p1_add_77522_comb + p1_add_77523_comb;
  assign p1_add_77626_comb = p1_add_77524_comb + p1_add_77525_comb;
  assign p1_add_77627_comb = p1_add_77526_comb + p1_add_77527_comb;
  assign p1_add_77628_comb = p1_sum__1100_comb + 25'h000_0001;
  assign p1_add_77629_comb = p1_sum__1094_comb + 25'h000_0001;
  assign p1_add_77630_comb = p1_sum__1089_comb + 25'h000_0001;
  assign p1_add_77631_comb = p1_sum__1085_comb + 25'h000_0001;
  assign p1_umul_27338_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_77536_comb, 7'h5b);
  assign p1_umul_27348_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_77538_comb, 7'h5b);
  assign p1_add_77634_comb = p1_sum__1133_comb + 25'h000_0001;
  assign p1_add_77635_comb = p1_sum__1108_comb + 25'h000_0001;
  assign p1_add_77636_comb = p1_add_77544_comb + p1_add_77545_comb;
  assign p1_add_77637_comb = p1_add_77546_comb + p1_add_77547_comb;
  assign p1_add_77638_comb = p1_sum__1128_comb + 25'h000_0001;
  assign p1_add_77639_comb = p1_sum__1096_comb + 25'h000_0001;
  assign p1_add_77640_comb = p1_sum__1124_comb + 25'h000_0001;
  assign p1_add_77641_comb = p1_sum__1091_comb + 25'h000_0001;
  assign p1_add_77642_comb = p1_sum__1119_comb + 25'h000_0001;
  assign p1_add_77643_comb = p1_sum__1087_comb + 25'h000_0001;
  assign p1_add_77644_comb = p1_add_77560_comb + p1_add_77561_comb;
  assign p1_add_77645_comb = p1_add_77562_comb + p1_add_77563_comb;
  assign p1_add_77646_comb = p1_sum__1107_comb + 25'h000_0001;
  assign p1_add_77647_comb = p1_sum__1082_comb + 25'h000_0001;
  assign p1_umul_27336_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_77568_comb, 7'h5b);
  assign p1_umul_27350_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_77570_comb, 7'h5b);
  assign p1_add_77650_comb = p1_sum__1135_comb + 25'h000_0001;
  assign p1_add_77651_comb = p1_sum__1101_comb + 25'h000_0001;
  assign p1_add_77652_comb = p1_add_77576_comb + p1_add_77577_comb;
  assign p1_add_77653_comb = p1_add_77578_comb + p1_add_77579_comb;
  assign p1_add_77654_comb = p1_sum__1132_comb + 25'h000_0001;
  assign p1_add_77655_comb = p1_sum__1090_comb + 25'h000_0001;
  assign p1_add_77656_comb = p1_sum__1129_comb + 25'h000_0001;
  assign p1_add_77657_comb = p1_sum__1086_comb + 25'h000_0001;
  assign p1_add_77658_comb = p1_sum__1125_comb + 25'h000_0001;
  assign p1_add_77659_comb = p1_sum__1083_comb + 25'h000_0001;
  assign p1_add_77660_comb = p1_add_77592_comb + p1_add_77593_comb;
  assign p1_add_77661_comb = p1_add_77594_comb + p1_add_77595_comb;
  assign p1_add_77662_comb = p1_sum__1114_comb + 25'h000_0001;
  assign p1_add_77663_comb = p1_sum__1080_comb + 25'h000_0001;
  assign p1_bit_slice_77664_comb = p1_umul_27340_NarrowedMult__comb[23:7];
  assign p1_bit_slice_77665_comb = p1_umul_27342_NarrowedMult__comb[23:7];
  assign p1_bit_slice_77666_comb = p1_umul_27344_NarrowedMult__comb[23:7];
  assign p1_bit_slice_77667_comb = p1_umul_27346_NarrowedMult__comb[23:7];
  assign p1_bit_slice_77668_comb = p1_add_77604_comb[24:8];
  assign p1_bit_slice_77669_comb = p1_add_77605_comb[24:8];
  assign p1_bit_slice_77670_comb = p1_add_77606_comb[24:8];
  assign p1_bit_slice_77671_comb = p1_add_77607_comb[24:8];
  assign p1_bit_slice_77672_comb = p1_add_77608_comb[23:7];
  assign p1_bit_slice_77673_comb = p1_add_77609_comb[23:7];
  assign p1_bit_slice_77674_comb = p1_add_77610_comb[23:7];
  assign p1_bit_slice_77675_comb = p1_add_77611_comb[23:7];
  assign p1_bit_slice_77676_comb = p1_add_77612_comb[24:8];
  assign p1_bit_slice_77677_comb = p1_add_77613_comb[24:8];
  assign p1_bit_slice_77678_comb = p1_add_77614_comb[24:8];
  assign p1_bit_slice_77679_comb = p1_add_77615_comb[24:8];
  assign p1_bit_slice_77680_comb = p1_add_77616_comb[24:8];
  assign p1_bit_slice_77681_comb = p1_add_77617_comb[24:8];
  assign p1_bit_slice_77682_comb = p1_add_77618_comb[24:8];
  assign p1_bit_slice_77683_comb = p1_add_77619_comb[24:8];
  assign p1_bit_slice_77684_comb = p1_add_77620_comb[24:8];
  assign p1_bit_slice_77685_comb = p1_add_77621_comb[24:8];
  assign p1_bit_slice_77686_comb = p1_add_77622_comb[24:8];
  assign p1_bit_slice_77687_comb = p1_add_77623_comb[24:8];
  assign p1_bit_slice_77688_comb = p1_add_77624_comb[23:7];
  assign p1_bit_slice_77689_comb = p1_add_77625_comb[23:7];
  assign p1_bit_slice_77690_comb = p1_add_77626_comb[23:7];
  assign p1_bit_slice_77691_comb = p1_add_77627_comb[23:7];
  assign p1_bit_slice_77692_comb = p1_add_77628_comb[24:8];
  assign p1_bit_slice_77693_comb = p1_add_77629_comb[24:8];
  assign p1_bit_slice_77694_comb = p1_add_77630_comb[24:8];
  assign p1_bit_slice_77695_comb = p1_add_77631_comb[24:8];
  assign p1_bit_slice_77696_comb = p1_umul_27338_NarrowedMult__comb[23:7];
  assign p1_bit_slice_77697_comb = p1_umul_27348_NarrowedMult__comb[23:7];
  assign p1_bit_slice_77698_comb = p1_add_77634_comb[24:8];
  assign p1_bit_slice_77699_comb = p1_add_77635_comb[24:8];
  assign p1_bit_slice_77700_comb = p1_add_77636_comb[23:7];
  assign p1_bit_slice_77701_comb = p1_add_77637_comb[23:7];
  assign p1_bit_slice_77702_comb = p1_add_77638_comb[24:8];
  assign p1_bit_slice_77703_comb = p1_add_77639_comb[24:8];
  assign p1_bit_slice_77704_comb = p1_add_77640_comb[24:8];
  assign p1_bit_slice_77705_comb = p1_add_77641_comb[24:8];
  assign p1_bit_slice_77706_comb = p1_add_77642_comb[24:8];
  assign p1_bit_slice_77707_comb = p1_add_77643_comb[24:8];
  assign p1_bit_slice_77708_comb = p1_add_77644_comb[23:7];
  assign p1_bit_slice_77709_comb = p1_add_77645_comb[23:7];
  assign p1_bit_slice_77710_comb = p1_add_77646_comb[24:8];
  assign p1_bit_slice_77711_comb = p1_add_77647_comb[24:8];
  assign p1_bit_slice_77712_comb = p1_umul_27336_NarrowedMult__comb[23:7];
  assign p1_bit_slice_77713_comb = p1_umul_27350_NarrowedMult__comb[23:7];
  assign p1_bit_slice_77714_comb = p1_add_77650_comb[24:8];
  assign p1_bit_slice_77715_comb = p1_add_77651_comb[24:8];
  assign p1_bit_slice_77716_comb = p1_add_77652_comb[23:7];
  assign p1_bit_slice_77717_comb = p1_add_77653_comb[23:7];
  assign p1_bit_slice_77718_comb = p1_add_77654_comb[24:8];
  assign p1_bit_slice_77719_comb = p1_add_77655_comb[24:8];
  assign p1_bit_slice_77720_comb = p1_add_77656_comb[24:8];
  assign p1_bit_slice_77721_comb = p1_add_77657_comb[24:8];
  assign p1_bit_slice_77722_comb = p1_add_77658_comb[24:8];
  assign p1_bit_slice_77723_comb = p1_add_77659_comb[24:8];
  assign p1_bit_slice_77724_comb = p1_add_77660_comb[23:7];
  assign p1_bit_slice_77725_comb = p1_add_77661_comb[23:7];
  assign p1_bit_slice_77726_comb = p1_add_77662_comb[24:8];
  assign p1_bit_slice_77727_comb = p1_add_77663_comb[24:8];
  assign p1_add_77856_comb = {{1{p1_bit_slice_77664_comb[16]}}, p1_bit_slice_77664_comb} + 18'h0_0001;
  assign p1_add_77857_comb = {{1{p1_bit_slice_77665_comb[16]}}, p1_bit_slice_77665_comb} + 18'h0_0001;
  assign p1_add_77858_comb = {{1{p1_bit_slice_77666_comb[16]}}, p1_bit_slice_77666_comb} + 18'h0_0001;
  assign p1_add_77859_comb = {{1{p1_bit_slice_77667_comb[16]}}, p1_bit_slice_77667_comb} + 18'h0_0001;
  assign p1_add_77860_comb = {{1{p1_bit_slice_77668_comb[16]}}, p1_bit_slice_77668_comb} + 18'h0_0001;
  assign p1_add_77861_comb = {{1{p1_bit_slice_77669_comb[16]}}, p1_bit_slice_77669_comb} + 18'h0_0001;
  assign p1_add_77862_comb = {{1{p1_bit_slice_77670_comb[16]}}, p1_bit_slice_77670_comb} + 18'h0_0001;
  assign p1_add_77863_comb = {{1{p1_bit_slice_77671_comb[16]}}, p1_bit_slice_77671_comb} + 18'h0_0001;
  assign p1_add_77864_comb = {{1{p1_bit_slice_77672_comb[16]}}, p1_bit_slice_77672_comb} + 18'h0_0001;
  assign p1_add_77865_comb = {{1{p1_bit_slice_77673_comb[16]}}, p1_bit_slice_77673_comb} + 18'h0_0001;
  assign p1_add_77866_comb = {{1{p1_bit_slice_77674_comb[16]}}, p1_bit_slice_77674_comb} + 18'h0_0001;
  assign p1_add_77867_comb = {{1{p1_bit_slice_77675_comb[16]}}, p1_bit_slice_77675_comb} + 18'h0_0001;
  assign p1_add_77868_comb = {{1{p1_bit_slice_77676_comb[16]}}, p1_bit_slice_77676_comb} + 18'h0_0001;
  assign p1_add_77869_comb = {{1{p1_bit_slice_77677_comb[16]}}, p1_bit_slice_77677_comb} + 18'h0_0001;
  assign p1_add_77870_comb = {{1{p1_bit_slice_77678_comb[16]}}, p1_bit_slice_77678_comb} + 18'h0_0001;
  assign p1_add_77871_comb = {{1{p1_bit_slice_77679_comb[16]}}, p1_bit_slice_77679_comb} + 18'h0_0001;
  assign p1_add_77872_comb = {{1{p1_bit_slice_77680_comb[16]}}, p1_bit_slice_77680_comb} + 18'h0_0001;
  assign p1_add_77873_comb = {{1{p1_bit_slice_77681_comb[16]}}, p1_bit_slice_77681_comb} + 18'h0_0001;
  assign p1_add_77874_comb = {{1{p1_bit_slice_77682_comb[16]}}, p1_bit_slice_77682_comb} + 18'h0_0001;
  assign p1_add_77875_comb = {{1{p1_bit_slice_77683_comb[16]}}, p1_bit_slice_77683_comb} + 18'h0_0001;
  assign p1_add_77876_comb = {{1{p1_bit_slice_77684_comb[16]}}, p1_bit_slice_77684_comb} + 18'h0_0001;
  assign p1_add_77877_comb = {{1{p1_bit_slice_77685_comb[16]}}, p1_bit_slice_77685_comb} + 18'h0_0001;
  assign p1_add_77878_comb = {{1{p1_bit_slice_77686_comb[16]}}, p1_bit_slice_77686_comb} + 18'h0_0001;
  assign p1_add_77879_comb = {{1{p1_bit_slice_77687_comb[16]}}, p1_bit_slice_77687_comb} + 18'h0_0001;
  assign p1_add_77880_comb = {{1{p1_bit_slice_77688_comb[16]}}, p1_bit_slice_77688_comb} + 18'h0_0001;
  assign p1_add_77881_comb = {{1{p1_bit_slice_77689_comb[16]}}, p1_bit_slice_77689_comb} + 18'h0_0001;
  assign p1_add_77882_comb = {{1{p1_bit_slice_77690_comb[16]}}, p1_bit_slice_77690_comb} + 18'h0_0001;
  assign p1_add_77883_comb = {{1{p1_bit_slice_77691_comb[16]}}, p1_bit_slice_77691_comb} + 18'h0_0001;
  assign p1_add_77884_comb = {{1{p1_bit_slice_77692_comb[16]}}, p1_bit_slice_77692_comb} + 18'h0_0001;
  assign p1_add_77885_comb = {{1{p1_bit_slice_77693_comb[16]}}, p1_bit_slice_77693_comb} + 18'h0_0001;
  assign p1_add_77886_comb = {{1{p1_bit_slice_77694_comb[16]}}, p1_bit_slice_77694_comb} + 18'h0_0001;
  assign p1_add_77887_comb = {{1{p1_bit_slice_77695_comb[16]}}, p1_bit_slice_77695_comb} + 18'h0_0001;
  assign p1_add_77888_comb = {{1{p1_bit_slice_77696_comb[16]}}, p1_bit_slice_77696_comb} + 18'h0_0001;
  assign p1_add_77889_comb = {{1{p1_bit_slice_77697_comb[16]}}, p1_bit_slice_77697_comb} + 18'h0_0001;
  assign p1_add_77890_comb = {{1{p1_bit_slice_77698_comb[16]}}, p1_bit_slice_77698_comb} + 18'h0_0001;
  assign p1_add_77891_comb = {{1{p1_bit_slice_77699_comb[16]}}, p1_bit_slice_77699_comb} + 18'h0_0001;
  assign p1_add_77892_comb = {{1{p1_bit_slice_77700_comb[16]}}, p1_bit_slice_77700_comb} + 18'h0_0001;
  assign p1_add_77893_comb = {{1{p1_bit_slice_77701_comb[16]}}, p1_bit_slice_77701_comb} + 18'h0_0001;
  assign p1_add_77894_comb = {{1{p1_bit_slice_77702_comb[16]}}, p1_bit_slice_77702_comb} + 18'h0_0001;
  assign p1_add_77895_comb = {{1{p1_bit_slice_77703_comb[16]}}, p1_bit_slice_77703_comb} + 18'h0_0001;
  assign p1_add_77896_comb = {{1{p1_bit_slice_77704_comb[16]}}, p1_bit_slice_77704_comb} + 18'h0_0001;
  assign p1_add_77897_comb = {{1{p1_bit_slice_77705_comb[16]}}, p1_bit_slice_77705_comb} + 18'h0_0001;
  assign p1_add_77898_comb = {{1{p1_bit_slice_77706_comb[16]}}, p1_bit_slice_77706_comb} + 18'h0_0001;
  assign p1_add_77899_comb = {{1{p1_bit_slice_77707_comb[16]}}, p1_bit_slice_77707_comb} + 18'h0_0001;
  assign p1_add_77900_comb = {{1{p1_bit_slice_77708_comb[16]}}, p1_bit_slice_77708_comb} + 18'h0_0001;
  assign p1_add_77901_comb = {{1{p1_bit_slice_77709_comb[16]}}, p1_bit_slice_77709_comb} + 18'h0_0001;
  assign p1_add_77902_comb = {{1{p1_bit_slice_77710_comb[16]}}, p1_bit_slice_77710_comb} + 18'h0_0001;
  assign p1_add_77903_comb = {{1{p1_bit_slice_77711_comb[16]}}, p1_bit_slice_77711_comb} + 18'h0_0001;
  assign p1_add_77904_comb = {{1{p1_bit_slice_77712_comb[16]}}, p1_bit_slice_77712_comb} + 18'h0_0001;
  assign p1_add_77905_comb = {{1{p1_bit_slice_77713_comb[16]}}, p1_bit_slice_77713_comb} + 18'h0_0001;
  assign p1_add_77906_comb = {{1{p1_bit_slice_77714_comb[16]}}, p1_bit_slice_77714_comb} + 18'h0_0001;
  assign p1_add_77907_comb = {{1{p1_bit_slice_77715_comb[16]}}, p1_bit_slice_77715_comb} + 18'h0_0001;
  assign p1_add_77908_comb = {{1{p1_bit_slice_77716_comb[16]}}, p1_bit_slice_77716_comb} + 18'h0_0001;
  assign p1_add_77909_comb = {{1{p1_bit_slice_77717_comb[16]}}, p1_bit_slice_77717_comb} + 18'h0_0001;
  assign p1_add_77910_comb = {{1{p1_bit_slice_77718_comb[16]}}, p1_bit_slice_77718_comb} + 18'h0_0001;
  assign p1_add_77911_comb = {{1{p1_bit_slice_77719_comb[16]}}, p1_bit_slice_77719_comb} + 18'h0_0001;
  assign p1_add_77912_comb = {{1{p1_bit_slice_77720_comb[16]}}, p1_bit_slice_77720_comb} + 18'h0_0001;
  assign p1_add_77913_comb = {{1{p1_bit_slice_77721_comb[16]}}, p1_bit_slice_77721_comb} + 18'h0_0001;
  assign p1_add_77914_comb = {{1{p1_bit_slice_77722_comb[16]}}, p1_bit_slice_77722_comb} + 18'h0_0001;
  assign p1_add_77915_comb = {{1{p1_bit_slice_77723_comb[16]}}, p1_bit_slice_77723_comb} + 18'h0_0001;
  assign p1_add_77916_comb = {{1{p1_bit_slice_77724_comb[16]}}, p1_bit_slice_77724_comb} + 18'h0_0001;
  assign p1_add_77917_comb = {{1{p1_bit_slice_77725_comb[16]}}, p1_bit_slice_77725_comb} + 18'h0_0001;
  assign p1_add_77918_comb = {{1{p1_bit_slice_77726_comb[16]}}, p1_bit_slice_77726_comb} + 18'h0_0001;
  assign p1_add_77919_comb = {{1{p1_bit_slice_77727_comb[16]}}, p1_bit_slice_77727_comb} + 18'h0_0001;
  assign p1_clipped__40_comb = $signed(p1_add_77856_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77856_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77856_comb[12:1]);
  assign p1_clipped__56_comb = $signed(p1_add_77857_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77857_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77857_comb[12:1]);
  assign p1_clipped__72_comb = $signed(p1_add_77858_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77858_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77858_comb[12:1]);
  assign p1_clipped__88_comb = $signed(p1_add_77859_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77859_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77859_comb[12:1]);
  assign p1_clipped__41_comb = $signed(p1_add_77860_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77860_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77860_comb[12:1]);
  assign p1_clipped__57_comb = $signed(p1_add_77861_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77861_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77861_comb[12:1]);
  assign p1_clipped__73_comb = $signed(p1_add_77862_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77862_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77862_comb[12:1]);
  assign p1_clipped__89_comb = $signed(p1_add_77863_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77863_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77863_comb[12:1]);
  assign p1_clipped__42_comb = $signed(p1_add_77864_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77864_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77864_comb[12:1]);
  assign p1_clipped__58_comb = $signed(p1_add_77865_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77865_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77865_comb[12:1]);
  assign p1_clipped__74_comb = $signed(p1_add_77866_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77866_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77866_comb[12:1]);
  assign p1_clipped__90_comb = $signed(p1_add_77867_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77867_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77867_comb[12:1]);
  assign p1_clipped__43_comb = $signed(p1_add_77868_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77868_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77868_comb[12:1]);
  assign p1_clipped__59_comb = $signed(p1_add_77869_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77869_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77869_comb[12:1]);
  assign p1_clipped__75_comb = $signed(p1_add_77870_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77870_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77870_comb[12:1]);
  assign p1_clipped__91_comb = $signed(p1_add_77871_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77871_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77871_comb[12:1]);
  assign p1_clipped__44_comb = $signed(p1_add_77872_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77872_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77872_comb[12:1]);
  assign p1_clipped__60_comb = $signed(p1_add_77873_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77873_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77873_comb[12:1]);
  assign p1_clipped__76_comb = $signed(p1_add_77874_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77874_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77874_comb[12:1]);
  assign p1_clipped__92_comb = $signed(p1_add_77875_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77875_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77875_comb[12:1]);
  assign p1_clipped__45_comb = $signed(p1_add_77876_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77876_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77876_comb[12:1]);
  assign p1_clipped__61_comb = $signed(p1_add_77877_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77877_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77877_comb[12:1]);
  assign p1_clipped__77_comb = $signed(p1_add_77878_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77878_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77878_comb[12:1]);
  assign p1_clipped__93_comb = $signed(p1_add_77879_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77879_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77879_comb[12:1]);
  assign p1_clipped__46_comb = $signed(p1_add_77880_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77880_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77880_comb[12:1]);
  assign p1_clipped__62_comb = $signed(p1_add_77881_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77881_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77881_comb[12:1]);
  assign p1_clipped__78_comb = $signed(p1_add_77882_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77882_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77882_comb[12:1]);
  assign p1_clipped__94_comb = $signed(p1_add_77883_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77883_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77883_comb[12:1]);
  assign p1_clipped__47_comb = $signed(p1_add_77884_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77884_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77884_comb[12:1]);
  assign p1_clipped__63_comb = $signed(p1_add_77885_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77885_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77885_comb[12:1]);
  assign p1_clipped__79_comb = $signed(p1_add_77886_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77886_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77886_comb[12:1]);
  assign p1_clipped__95_comb = $signed(p1_add_77887_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77887_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77887_comb[12:1]);
  assign p1_clipped__24_comb = $signed(p1_add_77888_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77888_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77888_comb[12:1]);
  assign p1_clipped__104_comb = $signed(p1_add_77889_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77889_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77889_comb[12:1]);
  assign p1_clipped__25_comb = $signed(p1_add_77890_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77890_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77890_comb[12:1]);
  assign p1_clipped__105_comb = $signed(p1_add_77891_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77891_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77891_comb[12:1]);
  assign p1_clipped__26_comb = $signed(p1_add_77892_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77892_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77892_comb[12:1]);
  assign p1_clipped__106_comb = $signed(p1_add_77893_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77893_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77893_comb[12:1]);
  assign p1_clipped__27_comb = $signed(p1_add_77894_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77894_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77894_comb[12:1]);
  assign p1_clipped__107_comb = $signed(p1_add_77895_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77895_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77895_comb[12:1]);
  assign p1_clipped__28_comb = $signed(p1_add_77896_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77896_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77896_comb[12:1]);
  assign p1_clipped__108_comb = $signed(p1_add_77897_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77897_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77897_comb[12:1]);
  assign p1_clipped__29_comb = $signed(p1_add_77898_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77898_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77898_comb[12:1]);
  assign p1_clipped__109_comb = $signed(p1_add_77899_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77899_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77899_comb[12:1]);
  assign p1_clipped__30_comb = $signed(p1_add_77900_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77900_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77900_comb[12:1]);
  assign p1_clipped__110_comb = $signed(p1_add_77901_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77901_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77901_comb[12:1]);
  assign p1_clipped__31_comb = $signed(p1_add_77902_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77902_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77902_comb[12:1]);
  assign p1_clipped__111_comb = $signed(p1_add_77903_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77903_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77903_comb[12:1]);
  assign p1_clipped__8_comb = $signed(p1_add_77904_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77904_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77904_comb[12:1]);
  assign p1_clipped__120_comb = $signed(p1_add_77905_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77905_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77905_comb[12:1]);
  assign p1_clipped__9_comb = $signed(p1_add_77906_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77906_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77906_comb[12:1]);
  assign p1_clipped__121_comb = $signed(p1_add_77907_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77907_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77907_comb[12:1]);
  assign p1_clipped__10_comb = $signed(p1_add_77908_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77908_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77908_comb[12:1]);
  assign p1_clipped__122_comb = $signed(p1_add_77909_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77909_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77909_comb[12:1]);
  assign p1_clipped__11_comb = $signed(p1_add_77910_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77910_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77910_comb[12:1]);
  assign p1_clipped__123_comb = $signed(p1_add_77911_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77911_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77911_comb[12:1]);
  assign p1_clipped__12_comb = $signed(p1_add_77912_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77912_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77912_comb[12:1]);
  assign p1_clipped__124_comb = $signed(p1_add_77913_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77913_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77913_comb[12:1]);
  assign p1_clipped__13_comb = $signed(p1_add_77914_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77914_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77914_comb[12:1]);
  assign p1_clipped__125_comb = $signed(p1_add_77915_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77915_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77915_comb[12:1]);
  assign p1_clipped__14_comb = $signed(p1_add_77916_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77916_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77916_comb[12:1]);
  assign p1_clipped__126_comb = $signed(p1_add_77917_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77917_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77917_comb[12:1]);
  assign p1_clipped__15_comb = $signed(p1_add_77918_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77918_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77918_comb[12:1]);
  assign p1_clipped__127_comb = $signed(p1_add_77919_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_77919_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_77919_comb[12:1]);
  assign p1_sign_ext_78562_comb = {{12{p1_clipped__40_comb[11]}}, p1_clipped__40_comb};
  assign p1_sign_ext_78563_comb = {{12{p1_clipped__56_comb[11]}}, p1_clipped__56_comb};
  assign p1_sign_ext_78564_comb = {{12{p1_clipped__72_comb[11]}}, p1_clipped__72_comb};
  assign p1_sign_ext_78565_comb = {{12{p1_clipped__88_comb[11]}}, p1_clipped__88_comb};
  assign p1_sign_ext_78570_comb = {{12{p1_clipped__41_comb[11]}}, p1_clipped__41_comb};
  assign p1_sign_ext_78571_comb = {{12{p1_clipped__57_comb[11]}}, p1_clipped__57_comb};
  assign p1_sign_ext_78572_comb = {{12{p1_clipped__73_comb[11]}}, p1_clipped__73_comb};
  assign p1_sign_ext_78573_comb = {{12{p1_clipped__89_comb[11]}}, p1_clipped__89_comb};
  assign p1_sign_ext_78578_comb = {{12{p1_clipped__42_comb[11]}}, p1_clipped__42_comb};
  assign p1_sign_ext_78579_comb = {{12{p1_clipped__58_comb[11]}}, p1_clipped__58_comb};
  assign p1_sign_ext_78580_comb = {{12{p1_clipped__74_comb[11]}}, p1_clipped__74_comb};
  assign p1_sign_ext_78581_comb = {{12{p1_clipped__90_comb[11]}}, p1_clipped__90_comb};
  assign p1_sign_ext_78586_comb = {{12{p1_clipped__43_comb[11]}}, p1_clipped__43_comb};
  assign p1_sign_ext_78587_comb = {{12{p1_clipped__59_comb[11]}}, p1_clipped__59_comb};
  assign p1_sign_ext_78588_comb = {{12{p1_clipped__75_comb[11]}}, p1_clipped__75_comb};
  assign p1_sign_ext_78589_comb = {{12{p1_clipped__91_comb[11]}}, p1_clipped__91_comb};
  assign p1_sign_ext_78594_comb = {{12{p1_clipped__44_comb[11]}}, p1_clipped__44_comb};
  assign p1_sign_ext_78595_comb = {{12{p1_clipped__60_comb[11]}}, p1_clipped__60_comb};
  assign p1_sign_ext_78596_comb = {{12{p1_clipped__76_comb[11]}}, p1_clipped__76_comb};
  assign p1_sign_ext_78597_comb = {{12{p1_clipped__92_comb[11]}}, p1_clipped__92_comb};
  assign p1_sign_ext_78602_comb = {{12{p1_clipped__45_comb[11]}}, p1_clipped__45_comb};
  assign p1_sign_ext_78603_comb = {{12{p1_clipped__61_comb[11]}}, p1_clipped__61_comb};
  assign p1_sign_ext_78604_comb = {{12{p1_clipped__77_comb[11]}}, p1_clipped__77_comb};
  assign p1_sign_ext_78605_comb = {{12{p1_clipped__93_comb[11]}}, p1_clipped__93_comb};
  assign p1_sign_ext_78610_comb = {{12{p1_clipped__46_comb[11]}}, p1_clipped__46_comb};
  assign p1_sign_ext_78611_comb = {{12{p1_clipped__62_comb[11]}}, p1_clipped__62_comb};
  assign p1_sign_ext_78612_comb = {{12{p1_clipped__78_comb[11]}}, p1_clipped__78_comb};
  assign p1_sign_ext_78613_comb = {{12{p1_clipped__94_comb[11]}}, p1_clipped__94_comb};
  assign p1_sign_ext_78618_comb = {{12{p1_clipped__47_comb[11]}}, p1_clipped__47_comb};
  assign p1_sign_ext_78619_comb = {{12{p1_clipped__63_comb[11]}}, p1_clipped__63_comb};
  assign p1_sign_ext_78620_comb = {{12{p1_clipped__79_comb[11]}}, p1_clipped__79_comb};
  assign p1_sign_ext_78621_comb = {{12{p1_clipped__95_comb[11]}}, p1_clipped__95_comb};
  assign p1_sign_ext_78624_comb = {{12{p1_clipped__24_comb[11]}}, p1_clipped__24_comb};
  assign p1_sign_ext_78625_comb = {{12{p1_clipped__104_comb[11]}}, p1_clipped__104_comb};
  assign p1_sign_ext_78626_comb = {{12{p1_clipped__25_comb[11]}}, p1_clipped__25_comb};
  assign p1_sign_ext_78627_comb = {{12{p1_clipped__105_comb[11]}}, p1_clipped__105_comb};
  assign p1_sign_ext_78628_comb = {{12{p1_clipped__26_comb[11]}}, p1_clipped__26_comb};
  assign p1_sign_ext_78629_comb = {{12{p1_clipped__106_comb[11]}}, p1_clipped__106_comb};
  assign p1_sign_ext_78630_comb = {{12{p1_clipped__27_comb[11]}}, p1_clipped__27_comb};
  assign p1_sign_ext_78631_comb = {{12{p1_clipped__107_comb[11]}}, p1_clipped__107_comb};
  assign p1_sign_ext_78632_comb = {{12{p1_clipped__28_comb[11]}}, p1_clipped__28_comb};
  assign p1_sign_ext_78633_comb = {{12{p1_clipped__108_comb[11]}}, p1_clipped__108_comb};
  assign p1_sign_ext_78634_comb = {{12{p1_clipped__29_comb[11]}}, p1_clipped__29_comb};
  assign p1_sign_ext_78635_comb = {{12{p1_clipped__109_comb[11]}}, p1_clipped__109_comb};
  assign p1_sign_ext_78636_comb = {{12{p1_clipped__30_comb[11]}}, p1_clipped__30_comb};
  assign p1_sign_ext_78637_comb = {{12{p1_clipped__110_comb[11]}}, p1_clipped__110_comb};
  assign p1_sign_ext_78638_comb = {{12{p1_clipped__31_comb[11]}}, p1_clipped__31_comb};
  assign p1_sign_ext_78639_comb = {{12{p1_clipped__111_comb[11]}}, p1_clipped__111_comb};
  assign p1_sign_ext_78672_comb = {{12{p1_clipped__8_comb[11]}}, p1_clipped__8_comb};
  assign p1_sign_ext_78677_comb = {{12{p1_clipped__120_comb[11]}}, p1_clipped__120_comb};
  assign p1_sign_ext_78678_comb = {{12{p1_clipped__9_comb[11]}}, p1_clipped__9_comb};
  assign p1_sign_ext_78683_comb = {{12{p1_clipped__121_comb[11]}}, p1_clipped__121_comb};
  assign p1_sign_ext_78684_comb = {{12{p1_clipped__10_comb[11]}}, p1_clipped__10_comb};
  assign p1_sign_ext_78689_comb = {{12{p1_clipped__122_comb[11]}}, p1_clipped__122_comb};
  assign p1_sign_ext_78690_comb = {{12{p1_clipped__11_comb[11]}}, p1_clipped__11_comb};
  assign p1_sign_ext_78695_comb = {{12{p1_clipped__123_comb[11]}}, p1_clipped__123_comb};
  assign p1_sign_ext_78696_comb = {{12{p1_clipped__12_comb[11]}}, p1_clipped__12_comb};
  assign p1_sign_ext_78701_comb = {{12{p1_clipped__124_comb[11]}}, p1_clipped__124_comb};
  assign p1_sign_ext_78702_comb = {{12{p1_clipped__13_comb[11]}}, p1_clipped__13_comb};
  assign p1_sign_ext_78707_comb = {{12{p1_clipped__125_comb[11]}}, p1_clipped__125_comb};
  assign p1_sign_ext_78708_comb = {{12{p1_clipped__14_comb[11]}}, p1_clipped__14_comb};
  assign p1_sign_ext_78713_comb = {{12{p1_clipped__126_comb[11]}}, p1_clipped__126_comb};
  assign p1_sign_ext_78714_comb = {{12{p1_clipped__15_comb[11]}}, p1_clipped__15_comb};
  assign p1_sign_ext_78719_comb = {{12{p1_clipped__127_comb[11]}}, p1_clipped__127_comb};
  assign p1_smul_78752_comb = smul21b_12b_x_9b(p1_clipped__8_comb, 9'h0fb);
  assign p1_smul_78753_comb = smul21b_12b_x_9b(p1_clipped__24_comb, 9'h0d5);
  assign p1_smul_78762_comb = smul21b_12b_x_9b(p1_clipped__104_comb, 9'h12b);
  assign p1_smul_78763_comb = smul21b_12b_x_9b(p1_clipped__120_comb, 9'h105);
  assign p1_smul_78764_comb = smul21b_12b_x_9b(p1_clipped__9_comb, 9'h0fb);
  assign p1_smul_78765_comb = smul21b_12b_x_9b(p1_clipped__25_comb, 9'h0d5);
  assign p1_smul_78774_comb = smul21b_12b_x_9b(p1_clipped__105_comb, 9'h12b);
  assign p1_smul_78775_comb = smul21b_12b_x_9b(p1_clipped__121_comb, 9'h105);
  assign p1_smul_78776_comb = smul21b_12b_x_9b(p1_clipped__10_comb, 9'h0fb);
  assign p1_smul_78777_comb = smul21b_12b_x_9b(p1_clipped__26_comb, 9'h0d5);
  assign p1_smul_78786_comb = smul21b_12b_x_9b(p1_clipped__106_comb, 9'h12b);
  assign p1_smul_78787_comb = smul21b_12b_x_9b(p1_clipped__122_comb, 9'h105);
  assign p1_smul_78788_comb = smul21b_12b_x_9b(p1_clipped__11_comb, 9'h0fb);
  assign p1_smul_78789_comb = smul21b_12b_x_9b(p1_clipped__27_comb, 9'h0d5);
  assign p1_smul_78798_comb = smul21b_12b_x_9b(p1_clipped__107_comb, 9'h12b);
  assign p1_smul_78799_comb = smul21b_12b_x_9b(p1_clipped__123_comb, 9'h105);
  assign p1_smul_78800_comb = smul21b_12b_x_9b(p1_clipped__12_comb, 9'h0fb);
  assign p1_smul_78801_comb = smul21b_12b_x_9b(p1_clipped__28_comb, 9'h0d5);
  assign p1_smul_78810_comb = smul21b_12b_x_9b(p1_clipped__108_comb, 9'h12b);
  assign p1_smul_78811_comb = smul21b_12b_x_9b(p1_clipped__124_comb, 9'h105);
  assign p1_smul_78812_comb = smul21b_12b_x_9b(p1_clipped__13_comb, 9'h0fb);
  assign p1_smul_78813_comb = smul21b_12b_x_9b(p1_clipped__29_comb, 9'h0d5);
  assign p1_smul_78822_comb = smul21b_12b_x_9b(p1_clipped__109_comb, 9'h12b);
  assign p1_smul_78823_comb = smul21b_12b_x_9b(p1_clipped__125_comb, 9'h105);
  assign p1_smul_78824_comb = smul21b_12b_x_9b(p1_clipped__14_comb, 9'h0fb);
  assign p1_smul_78825_comb = smul21b_12b_x_9b(p1_clipped__30_comb, 9'h0d5);
  assign p1_smul_78834_comb = smul21b_12b_x_9b(p1_clipped__110_comb, 9'h12b);
  assign p1_smul_78835_comb = smul21b_12b_x_9b(p1_clipped__126_comb, 9'h105);
  assign p1_smul_78836_comb = smul21b_12b_x_9b(p1_clipped__15_comb, 9'h0fb);
  assign p1_smul_78837_comb = smul21b_12b_x_9b(p1_clipped__31_comb, 9'h0d5);
  assign p1_smul_78846_comb = smul21b_12b_x_9b(p1_clipped__111_comb, 9'h12b);
  assign p1_smul_78847_comb = smul21b_12b_x_9b(p1_clipped__127_comb, 9'h105);
  assign p1_smul_78896_comb = smul21b_12b_x_9b(p1_clipped__8_comb, 9'h0d5);
  assign p1_smul_78898_comb = smul21b_12b_x_9b(p1_clipped__40_comb, 9'h105);
  assign p1_smul_78901_comb = smul21b_12b_x_9b(p1_clipped__88_comb, 9'h0fb);
  assign p1_smul_78903_comb = smul21b_12b_x_9b(p1_clipped__120_comb, 9'h12b);
  assign p1_smul_78904_comb = smul21b_12b_x_9b(p1_clipped__9_comb, 9'h0d5);
  assign p1_smul_78906_comb = smul21b_12b_x_9b(p1_clipped__41_comb, 9'h105);
  assign p1_smul_78909_comb = smul21b_12b_x_9b(p1_clipped__89_comb, 9'h0fb);
  assign p1_smul_78911_comb = smul21b_12b_x_9b(p1_clipped__121_comb, 9'h12b);
  assign p1_smul_78912_comb = smul21b_12b_x_9b(p1_clipped__10_comb, 9'h0d5);
  assign p1_smul_78914_comb = smul21b_12b_x_9b(p1_clipped__42_comb, 9'h105);
  assign p1_smul_78917_comb = smul21b_12b_x_9b(p1_clipped__90_comb, 9'h0fb);
  assign p1_smul_78919_comb = smul21b_12b_x_9b(p1_clipped__122_comb, 9'h12b);
  assign p1_smul_78920_comb = smul21b_12b_x_9b(p1_clipped__11_comb, 9'h0d5);
  assign p1_smul_78922_comb = smul21b_12b_x_9b(p1_clipped__43_comb, 9'h105);
  assign p1_smul_78925_comb = smul21b_12b_x_9b(p1_clipped__91_comb, 9'h0fb);
  assign p1_smul_78927_comb = smul21b_12b_x_9b(p1_clipped__123_comb, 9'h12b);
  assign p1_smul_78928_comb = smul21b_12b_x_9b(p1_clipped__12_comb, 9'h0d5);
  assign p1_smul_78930_comb = smul21b_12b_x_9b(p1_clipped__44_comb, 9'h105);
  assign p1_smul_78933_comb = smul21b_12b_x_9b(p1_clipped__92_comb, 9'h0fb);
  assign p1_smul_78935_comb = smul21b_12b_x_9b(p1_clipped__124_comb, 9'h12b);
  assign p1_smul_78936_comb = smul21b_12b_x_9b(p1_clipped__13_comb, 9'h0d5);
  assign p1_smul_78938_comb = smul21b_12b_x_9b(p1_clipped__45_comb, 9'h105);
  assign p1_smul_78941_comb = smul21b_12b_x_9b(p1_clipped__93_comb, 9'h0fb);
  assign p1_smul_78943_comb = smul21b_12b_x_9b(p1_clipped__125_comb, 9'h12b);
  assign p1_smul_78944_comb = smul21b_12b_x_9b(p1_clipped__14_comb, 9'h0d5);
  assign p1_smul_78946_comb = smul21b_12b_x_9b(p1_clipped__46_comb, 9'h105);
  assign p1_smul_78949_comb = smul21b_12b_x_9b(p1_clipped__94_comb, 9'h0fb);
  assign p1_smul_78951_comb = smul21b_12b_x_9b(p1_clipped__126_comb, 9'h12b);
  assign p1_smul_78952_comb = smul21b_12b_x_9b(p1_clipped__15_comb, 9'h0d5);
  assign p1_smul_78954_comb = smul21b_12b_x_9b(p1_clipped__47_comb, 9'h105);
  assign p1_smul_78957_comb = smul21b_12b_x_9b(p1_clipped__95_comb, 9'h0fb);
  assign p1_smul_78959_comb = smul21b_12b_x_9b(p1_clipped__127_comb, 9'h12b);
  assign p1_smul_78962_comb = smul21b_12b_x_9b(p1_clipped__24_comb, 9'h105);
  assign p1_smul_78964_comb = smul21b_12b_x_9b(p1_clipped__56_comb, 9'h0d5);
  assign p1_smul_78965_comb = smul21b_12b_x_9b(p1_clipped__72_comb, 9'h0d5);
  assign p1_smul_78967_comb = smul21b_12b_x_9b(p1_clipped__104_comb, 9'h105);
  assign p1_smul_78972_comb = smul21b_12b_x_9b(p1_clipped__25_comb, 9'h105);
  assign p1_smul_78974_comb = smul21b_12b_x_9b(p1_clipped__57_comb, 9'h0d5);
  assign p1_smul_78975_comb = smul21b_12b_x_9b(p1_clipped__73_comb, 9'h0d5);
  assign p1_smul_78977_comb = smul21b_12b_x_9b(p1_clipped__105_comb, 9'h105);
  assign p1_smul_78982_comb = smul21b_12b_x_9b(p1_clipped__26_comb, 9'h105);
  assign p1_smul_78984_comb = smul21b_12b_x_9b(p1_clipped__58_comb, 9'h0d5);
  assign p1_smul_78985_comb = smul21b_12b_x_9b(p1_clipped__74_comb, 9'h0d5);
  assign p1_smul_78987_comb = smul21b_12b_x_9b(p1_clipped__106_comb, 9'h105);
  assign p1_smul_78992_comb = smul21b_12b_x_9b(p1_clipped__27_comb, 9'h105);
  assign p1_smul_78994_comb = smul21b_12b_x_9b(p1_clipped__59_comb, 9'h0d5);
  assign p1_smul_78995_comb = smul21b_12b_x_9b(p1_clipped__75_comb, 9'h0d5);
  assign p1_smul_78997_comb = smul21b_12b_x_9b(p1_clipped__107_comb, 9'h105);
  assign p1_smul_79002_comb = smul21b_12b_x_9b(p1_clipped__28_comb, 9'h105);
  assign p1_smul_79004_comb = smul21b_12b_x_9b(p1_clipped__60_comb, 9'h0d5);
  assign p1_smul_79005_comb = smul21b_12b_x_9b(p1_clipped__76_comb, 9'h0d5);
  assign p1_smul_79007_comb = smul21b_12b_x_9b(p1_clipped__108_comb, 9'h105);
  assign p1_smul_79012_comb = smul21b_12b_x_9b(p1_clipped__29_comb, 9'h105);
  assign p1_smul_79014_comb = smul21b_12b_x_9b(p1_clipped__61_comb, 9'h0d5);
  assign p1_smul_79015_comb = smul21b_12b_x_9b(p1_clipped__77_comb, 9'h0d5);
  assign p1_smul_79017_comb = smul21b_12b_x_9b(p1_clipped__109_comb, 9'h105);
  assign p1_smul_79022_comb = smul21b_12b_x_9b(p1_clipped__30_comb, 9'h105);
  assign p1_smul_79024_comb = smul21b_12b_x_9b(p1_clipped__62_comb, 9'h0d5);
  assign p1_smul_79025_comb = smul21b_12b_x_9b(p1_clipped__78_comb, 9'h0d5);
  assign p1_smul_79027_comb = smul21b_12b_x_9b(p1_clipped__110_comb, 9'h105);
  assign p1_smul_79032_comb = smul21b_12b_x_9b(p1_clipped__31_comb, 9'h105);
  assign p1_smul_79034_comb = smul21b_12b_x_9b(p1_clipped__63_comb, 9'h0d5);
  assign p1_smul_79035_comb = smul21b_12b_x_9b(p1_clipped__79_comb, 9'h0d5);
  assign p1_smul_79037_comb = smul21b_12b_x_9b(p1_clipped__111_comb, 9'h105);
  assign p1_smul_79074_comb = smul21b_12b_x_9b(p1_clipped__40_comb, 9'h0d5);
  assign p1_smul_79075_comb = smul21b_12b_x_9b(p1_clipped__56_comb, 9'h105);
  assign p1_smul_79076_comb = smul21b_12b_x_9b(p1_clipped__72_comb, 9'h105);
  assign p1_smul_79077_comb = smul21b_12b_x_9b(p1_clipped__88_comb, 9'h0d5);
  assign p1_smul_79082_comb = smul21b_12b_x_9b(p1_clipped__41_comb, 9'h0d5);
  assign p1_smul_79083_comb = smul21b_12b_x_9b(p1_clipped__57_comb, 9'h105);
  assign p1_smul_79084_comb = smul21b_12b_x_9b(p1_clipped__73_comb, 9'h105);
  assign p1_smul_79085_comb = smul21b_12b_x_9b(p1_clipped__89_comb, 9'h0d5);
  assign p1_smul_79090_comb = smul21b_12b_x_9b(p1_clipped__42_comb, 9'h0d5);
  assign p1_smul_79091_comb = smul21b_12b_x_9b(p1_clipped__58_comb, 9'h105);
  assign p1_smul_79092_comb = smul21b_12b_x_9b(p1_clipped__74_comb, 9'h105);
  assign p1_smul_79093_comb = smul21b_12b_x_9b(p1_clipped__90_comb, 9'h0d5);
  assign p1_smul_79098_comb = smul21b_12b_x_9b(p1_clipped__43_comb, 9'h0d5);
  assign p1_smul_79099_comb = smul21b_12b_x_9b(p1_clipped__59_comb, 9'h105);
  assign p1_smul_79100_comb = smul21b_12b_x_9b(p1_clipped__75_comb, 9'h105);
  assign p1_smul_79101_comb = smul21b_12b_x_9b(p1_clipped__91_comb, 9'h0d5);
  assign p1_smul_79106_comb = smul21b_12b_x_9b(p1_clipped__44_comb, 9'h0d5);
  assign p1_smul_79107_comb = smul21b_12b_x_9b(p1_clipped__60_comb, 9'h105);
  assign p1_smul_79108_comb = smul21b_12b_x_9b(p1_clipped__76_comb, 9'h105);
  assign p1_smul_79109_comb = smul21b_12b_x_9b(p1_clipped__92_comb, 9'h0d5);
  assign p1_smul_79114_comb = smul21b_12b_x_9b(p1_clipped__45_comb, 9'h0d5);
  assign p1_smul_79115_comb = smul21b_12b_x_9b(p1_clipped__61_comb, 9'h105);
  assign p1_smul_79116_comb = smul21b_12b_x_9b(p1_clipped__77_comb, 9'h105);
  assign p1_smul_79117_comb = smul21b_12b_x_9b(p1_clipped__93_comb, 9'h0d5);
  assign p1_smul_79122_comb = smul21b_12b_x_9b(p1_clipped__46_comb, 9'h0d5);
  assign p1_smul_79123_comb = smul21b_12b_x_9b(p1_clipped__62_comb, 9'h105);
  assign p1_smul_79124_comb = smul21b_12b_x_9b(p1_clipped__78_comb, 9'h105);
  assign p1_smul_79125_comb = smul21b_12b_x_9b(p1_clipped__94_comb, 9'h0d5);
  assign p1_smul_79130_comb = smul21b_12b_x_9b(p1_clipped__47_comb, 9'h0d5);
  assign p1_smul_79131_comb = smul21b_12b_x_9b(p1_clipped__63_comb, 9'h105);
  assign p1_smul_79132_comb = smul21b_12b_x_9b(p1_clipped__79_comb, 9'h105);
  assign p1_smul_79133_comb = smul21b_12b_x_9b(p1_clipped__95_comb, 9'h0d5);
  assign p1_add_79136_comb = p1_smul_78752_comb + p1_smul_78753_comb;
  assign p1_smul_79137_comb = smul20b_20b_x_8b(p1_sign_ext_78562_comb[19:0], 8'h47);
  assign p1_smul_79138_comb = smul20b_20b_x_6b(p1_sign_ext_78563_comb[19:0], 6'h19);
  assign p1_smul_79139_comb = smul20b_20b_x_6b(p1_sign_ext_78564_comb[19:0], 6'h27);
  assign p1_smul_79140_comb = smul20b_20b_x_8b(p1_sign_ext_78565_comb[19:0], 8'hb9);
  assign p1_add_79141_comb = p1_smul_78762_comb + p1_smul_78763_comb;
  assign p1_add_79142_comb = p1_smul_78764_comb + p1_smul_78765_comb;
  assign p1_smul_79143_comb = smul20b_20b_x_8b(p1_sign_ext_78570_comb[19:0], 8'h47);
  assign p1_smul_79144_comb = smul20b_20b_x_6b(p1_sign_ext_78571_comb[19:0], 6'h19);
  assign p1_smul_79145_comb = smul20b_20b_x_6b(p1_sign_ext_78572_comb[19:0], 6'h27);
  assign p1_smul_79146_comb = smul20b_20b_x_8b(p1_sign_ext_78573_comb[19:0], 8'hb9);
  assign p1_add_79147_comb = p1_smul_78774_comb + p1_smul_78775_comb;
  assign p1_add_79148_comb = p1_smul_78776_comb + p1_smul_78777_comb;
  assign p1_smul_79149_comb = smul20b_20b_x_8b(p1_sign_ext_78578_comb[19:0], 8'h47);
  assign p1_smul_79150_comb = smul20b_20b_x_6b(p1_sign_ext_78579_comb[19:0], 6'h19);
  assign p1_smul_79151_comb = smul20b_20b_x_6b(p1_sign_ext_78580_comb[19:0], 6'h27);
  assign p1_smul_79152_comb = smul20b_20b_x_8b(p1_sign_ext_78581_comb[19:0], 8'hb9);
  assign p1_add_79153_comb = p1_smul_78786_comb + p1_smul_78787_comb;
  assign p1_add_79154_comb = p1_smul_78788_comb + p1_smul_78789_comb;
  assign p1_smul_79155_comb = smul20b_20b_x_8b(p1_sign_ext_78586_comb[19:0], 8'h47);
  assign p1_smul_79156_comb = smul20b_20b_x_6b(p1_sign_ext_78587_comb[19:0], 6'h19);
  assign p1_smul_79157_comb = smul20b_20b_x_6b(p1_sign_ext_78588_comb[19:0], 6'h27);
  assign p1_smul_79158_comb = smul20b_20b_x_8b(p1_sign_ext_78589_comb[19:0], 8'hb9);
  assign p1_add_79159_comb = p1_smul_78798_comb + p1_smul_78799_comb;
  assign p1_add_79160_comb = p1_smul_78800_comb + p1_smul_78801_comb;
  assign p1_smul_79161_comb = smul20b_20b_x_8b(p1_sign_ext_78594_comb[19:0], 8'h47);
  assign p1_smul_79162_comb = smul20b_20b_x_6b(p1_sign_ext_78595_comb[19:0], 6'h19);
  assign p1_smul_79163_comb = smul20b_20b_x_6b(p1_sign_ext_78596_comb[19:0], 6'h27);
  assign p1_smul_79164_comb = smul20b_20b_x_8b(p1_sign_ext_78597_comb[19:0], 8'hb9);
  assign p1_add_79165_comb = p1_smul_78810_comb + p1_smul_78811_comb;
  assign p1_add_79166_comb = p1_smul_78812_comb + p1_smul_78813_comb;
  assign p1_smul_79167_comb = smul20b_20b_x_8b(p1_sign_ext_78602_comb[19:0], 8'h47);
  assign p1_smul_79168_comb = smul20b_20b_x_6b(p1_sign_ext_78603_comb[19:0], 6'h19);
  assign p1_smul_79169_comb = smul20b_20b_x_6b(p1_sign_ext_78604_comb[19:0], 6'h27);
  assign p1_smul_79170_comb = smul20b_20b_x_8b(p1_sign_ext_78605_comb[19:0], 8'hb9);
  assign p1_add_79171_comb = p1_smul_78822_comb + p1_smul_78823_comb;
  assign p1_add_79172_comb = p1_smul_78824_comb + p1_smul_78825_comb;
  assign p1_smul_79173_comb = smul20b_20b_x_8b(p1_sign_ext_78610_comb[19:0], 8'h47);
  assign p1_smul_79174_comb = smul20b_20b_x_6b(p1_sign_ext_78611_comb[19:0], 6'h19);
  assign p1_smul_79175_comb = smul20b_20b_x_6b(p1_sign_ext_78612_comb[19:0], 6'h27);
  assign p1_smul_79176_comb = smul20b_20b_x_8b(p1_sign_ext_78613_comb[19:0], 8'hb9);
  assign p1_add_79177_comb = p1_smul_78834_comb + p1_smul_78835_comb;
  assign p1_add_79178_comb = p1_smul_78836_comb + p1_smul_78837_comb;
  assign p1_smul_79179_comb = smul20b_20b_x_8b(p1_sign_ext_78618_comb[19:0], 8'h47);
  assign p1_smul_79180_comb = smul20b_20b_x_6b(p1_sign_ext_78619_comb[19:0], 6'h19);
  assign p1_smul_79181_comb = smul20b_20b_x_6b(p1_sign_ext_78620_comb[19:0], 6'h27);
  assign p1_smul_79182_comb = smul20b_20b_x_8b(p1_sign_ext_78621_comb[19:0], 8'hb9);
  assign p1_add_79183_comb = p1_smul_78846_comb + p1_smul_78847_comb;
  assign p1_smul_79186_comb = smul20b_20b_x_7b(p1_sign_ext_78624_comb[19:0], 7'h31);
  assign p1_smul_79187_comb = smul20b_20b_x_7b(p1_sign_ext_78562_comb[19:0], 7'h4f);
  assign p1_smul_79192_comb = smul20b_20b_x_7b(p1_sign_ext_78565_comb[19:0], 7'h4f);
  assign p1_smul_79193_comb = smul20b_20b_x_7b(p1_sign_ext_78625_comb[19:0], 7'h31);
  assign p1_smul_79198_comb = smul20b_20b_x_7b(p1_sign_ext_78626_comb[19:0], 7'h31);
  assign p1_smul_79199_comb = smul20b_20b_x_7b(p1_sign_ext_78570_comb[19:0], 7'h4f);
  assign p1_smul_79204_comb = smul20b_20b_x_7b(p1_sign_ext_78573_comb[19:0], 7'h4f);
  assign p1_smul_79205_comb = smul20b_20b_x_7b(p1_sign_ext_78627_comb[19:0], 7'h31);
  assign p1_smul_79210_comb = smul20b_20b_x_7b(p1_sign_ext_78628_comb[19:0], 7'h31);
  assign p1_smul_79211_comb = smul20b_20b_x_7b(p1_sign_ext_78578_comb[19:0], 7'h4f);
  assign p1_smul_79216_comb = smul20b_20b_x_7b(p1_sign_ext_78581_comb[19:0], 7'h4f);
  assign p1_smul_79217_comb = smul20b_20b_x_7b(p1_sign_ext_78629_comb[19:0], 7'h31);
  assign p1_smul_79222_comb = smul20b_20b_x_7b(p1_sign_ext_78630_comb[19:0], 7'h31);
  assign p1_smul_79223_comb = smul20b_20b_x_7b(p1_sign_ext_78586_comb[19:0], 7'h4f);
  assign p1_smul_79228_comb = smul20b_20b_x_7b(p1_sign_ext_78589_comb[19:0], 7'h4f);
  assign p1_smul_79229_comb = smul20b_20b_x_7b(p1_sign_ext_78631_comb[19:0], 7'h31);
  assign p1_smul_79234_comb = smul20b_20b_x_7b(p1_sign_ext_78632_comb[19:0], 7'h31);
  assign p1_smul_79235_comb = smul20b_20b_x_7b(p1_sign_ext_78594_comb[19:0], 7'h4f);
  assign p1_smul_79240_comb = smul20b_20b_x_7b(p1_sign_ext_78597_comb[19:0], 7'h4f);
  assign p1_smul_79241_comb = smul20b_20b_x_7b(p1_sign_ext_78633_comb[19:0], 7'h31);
  assign p1_smul_79246_comb = smul20b_20b_x_7b(p1_sign_ext_78634_comb[19:0], 7'h31);
  assign p1_smul_79247_comb = smul20b_20b_x_7b(p1_sign_ext_78602_comb[19:0], 7'h4f);
  assign p1_smul_79252_comb = smul20b_20b_x_7b(p1_sign_ext_78605_comb[19:0], 7'h4f);
  assign p1_smul_79253_comb = smul20b_20b_x_7b(p1_sign_ext_78635_comb[19:0], 7'h31);
  assign p1_smul_79258_comb = smul20b_20b_x_7b(p1_sign_ext_78636_comb[19:0], 7'h31);
  assign p1_smul_79259_comb = smul20b_20b_x_7b(p1_sign_ext_78610_comb[19:0], 7'h4f);
  assign p1_smul_79264_comb = smul20b_20b_x_7b(p1_sign_ext_78613_comb[19:0], 7'h4f);
  assign p1_smul_79265_comb = smul20b_20b_x_7b(p1_sign_ext_78637_comb[19:0], 7'h31);
  assign p1_smul_79270_comb = smul20b_20b_x_7b(p1_sign_ext_78638_comb[19:0], 7'h31);
  assign p1_smul_79271_comb = smul20b_20b_x_7b(p1_sign_ext_78618_comb[19:0], 7'h4f);
  assign p1_smul_79276_comb = smul20b_20b_x_7b(p1_sign_ext_78621_comb[19:0], 7'h4f);
  assign p1_smul_79277_comb = smul20b_20b_x_7b(p1_sign_ext_78639_comb[19:0], 7'h31);
  assign p1_smul_79281_comb = smul20b_20b_x_6b(p1_sign_ext_78624_comb[19:0], 6'h27);
  assign p1_smul_79283_comb = smul20b_20b_x_8b(p1_sign_ext_78563_comb[19:0], 8'hb9);
  assign p1_smul_79284_comb = smul20b_20b_x_8b(p1_sign_ext_78564_comb[19:0], 8'h47);
  assign p1_smul_79286_comb = smul20b_20b_x_6b(p1_sign_ext_78625_comb[19:0], 6'h19);
  assign p1_smul_79289_comb = smul20b_20b_x_6b(p1_sign_ext_78626_comb[19:0], 6'h27);
  assign p1_smul_79291_comb = smul20b_20b_x_8b(p1_sign_ext_78571_comb[19:0], 8'hb9);
  assign p1_smul_79292_comb = smul20b_20b_x_8b(p1_sign_ext_78572_comb[19:0], 8'h47);
  assign p1_smul_79294_comb = smul20b_20b_x_6b(p1_sign_ext_78627_comb[19:0], 6'h19);
  assign p1_smul_79297_comb = smul20b_20b_x_6b(p1_sign_ext_78628_comb[19:0], 6'h27);
  assign p1_smul_79299_comb = smul20b_20b_x_8b(p1_sign_ext_78579_comb[19:0], 8'hb9);
  assign p1_smul_79300_comb = smul20b_20b_x_8b(p1_sign_ext_78580_comb[19:0], 8'h47);
  assign p1_smul_79302_comb = smul20b_20b_x_6b(p1_sign_ext_78629_comb[19:0], 6'h19);
  assign p1_smul_79305_comb = smul20b_20b_x_6b(p1_sign_ext_78630_comb[19:0], 6'h27);
  assign p1_smul_79307_comb = smul20b_20b_x_8b(p1_sign_ext_78587_comb[19:0], 8'hb9);
  assign p1_smul_79308_comb = smul20b_20b_x_8b(p1_sign_ext_78588_comb[19:0], 8'h47);
  assign p1_smul_79310_comb = smul20b_20b_x_6b(p1_sign_ext_78631_comb[19:0], 6'h19);
  assign p1_smul_79313_comb = smul20b_20b_x_6b(p1_sign_ext_78632_comb[19:0], 6'h27);
  assign p1_smul_79315_comb = smul20b_20b_x_8b(p1_sign_ext_78595_comb[19:0], 8'hb9);
  assign p1_smul_79316_comb = smul20b_20b_x_8b(p1_sign_ext_78596_comb[19:0], 8'h47);
  assign p1_smul_79318_comb = smul20b_20b_x_6b(p1_sign_ext_78633_comb[19:0], 6'h19);
  assign p1_smul_79321_comb = smul20b_20b_x_6b(p1_sign_ext_78634_comb[19:0], 6'h27);
  assign p1_smul_79323_comb = smul20b_20b_x_8b(p1_sign_ext_78603_comb[19:0], 8'hb9);
  assign p1_smul_79324_comb = smul20b_20b_x_8b(p1_sign_ext_78604_comb[19:0], 8'h47);
  assign p1_smul_79326_comb = smul20b_20b_x_6b(p1_sign_ext_78635_comb[19:0], 6'h19);
  assign p1_smul_79329_comb = smul20b_20b_x_6b(p1_sign_ext_78636_comb[19:0], 6'h27);
  assign p1_smul_79331_comb = smul20b_20b_x_8b(p1_sign_ext_78611_comb[19:0], 8'hb9);
  assign p1_smul_79332_comb = smul20b_20b_x_8b(p1_sign_ext_78612_comb[19:0], 8'h47);
  assign p1_smul_79334_comb = smul20b_20b_x_6b(p1_sign_ext_78637_comb[19:0], 6'h19);
  assign p1_smul_79337_comb = smul20b_20b_x_6b(p1_sign_ext_78638_comb[19:0], 6'h27);
  assign p1_smul_79339_comb = smul20b_20b_x_8b(p1_sign_ext_78619_comb[19:0], 8'hb9);
  assign p1_smul_79340_comb = smul20b_20b_x_8b(p1_sign_ext_78620_comb[19:0], 8'h47);
  assign p1_smul_79342_comb = smul20b_20b_x_6b(p1_sign_ext_78639_comb[19:0], 6'h19);
  assign p1_smul_79408_comb = smul20b_20b_x_8b(p1_sign_ext_78672_comb[19:0], 8'h47);
  assign p1_smul_79410_comb = smul20b_20b_x_6b(p1_sign_ext_78562_comb[19:0], 6'h27);
  assign p1_smul_79413_comb = smul20b_20b_x_6b(p1_sign_ext_78565_comb[19:0], 6'h27);
  assign p1_smul_79415_comb = smul20b_20b_x_8b(p1_sign_ext_78677_comb[19:0], 8'h47);
  assign p1_smul_79416_comb = smul20b_20b_x_8b(p1_sign_ext_78678_comb[19:0], 8'h47);
  assign p1_smul_79418_comb = smul20b_20b_x_6b(p1_sign_ext_78570_comb[19:0], 6'h27);
  assign p1_smul_79421_comb = smul20b_20b_x_6b(p1_sign_ext_78573_comb[19:0], 6'h27);
  assign p1_smul_79423_comb = smul20b_20b_x_8b(p1_sign_ext_78683_comb[19:0], 8'h47);
  assign p1_smul_79424_comb = smul20b_20b_x_8b(p1_sign_ext_78684_comb[19:0], 8'h47);
  assign p1_smul_79426_comb = smul20b_20b_x_6b(p1_sign_ext_78578_comb[19:0], 6'h27);
  assign p1_smul_79429_comb = smul20b_20b_x_6b(p1_sign_ext_78581_comb[19:0], 6'h27);
  assign p1_smul_79431_comb = smul20b_20b_x_8b(p1_sign_ext_78689_comb[19:0], 8'h47);
  assign p1_smul_79432_comb = smul20b_20b_x_8b(p1_sign_ext_78690_comb[19:0], 8'h47);
  assign p1_smul_79434_comb = smul20b_20b_x_6b(p1_sign_ext_78586_comb[19:0], 6'h27);
  assign p1_smul_79437_comb = smul20b_20b_x_6b(p1_sign_ext_78589_comb[19:0], 6'h27);
  assign p1_smul_79439_comb = smul20b_20b_x_8b(p1_sign_ext_78695_comb[19:0], 8'h47);
  assign p1_smul_79440_comb = smul20b_20b_x_8b(p1_sign_ext_78696_comb[19:0], 8'h47);
  assign p1_smul_79442_comb = smul20b_20b_x_6b(p1_sign_ext_78594_comb[19:0], 6'h27);
  assign p1_smul_79445_comb = smul20b_20b_x_6b(p1_sign_ext_78597_comb[19:0], 6'h27);
  assign p1_smul_79447_comb = smul20b_20b_x_8b(p1_sign_ext_78701_comb[19:0], 8'h47);
  assign p1_smul_79448_comb = smul20b_20b_x_8b(p1_sign_ext_78702_comb[19:0], 8'h47);
  assign p1_smul_79450_comb = smul20b_20b_x_6b(p1_sign_ext_78602_comb[19:0], 6'h27);
  assign p1_smul_79453_comb = smul20b_20b_x_6b(p1_sign_ext_78605_comb[19:0], 6'h27);
  assign p1_smul_79455_comb = smul20b_20b_x_8b(p1_sign_ext_78707_comb[19:0], 8'h47);
  assign p1_smul_79456_comb = smul20b_20b_x_8b(p1_sign_ext_78708_comb[19:0], 8'h47);
  assign p1_smul_79458_comb = smul20b_20b_x_6b(p1_sign_ext_78610_comb[19:0], 6'h27);
  assign p1_smul_79461_comb = smul20b_20b_x_6b(p1_sign_ext_78613_comb[19:0], 6'h27);
  assign p1_smul_79463_comb = smul20b_20b_x_8b(p1_sign_ext_78713_comb[19:0], 8'h47);
  assign p1_smul_79464_comb = smul20b_20b_x_8b(p1_sign_ext_78714_comb[19:0], 8'h47);
  assign p1_smul_79466_comb = smul20b_20b_x_6b(p1_sign_ext_78618_comb[19:0], 6'h27);
  assign p1_smul_79469_comb = smul20b_20b_x_6b(p1_sign_ext_78621_comb[19:0], 6'h27);
  assign p1_smul_79471_comb = smul20b_20b_x_8b(p1_sign_ext_78719_comb[19:0], 8'h47);
  assign p1_smul_79472_comb = smul20b_20b_x_7b(p1_sign_ext_78672_comb[19:0], 7'h31);
  assign p1_smul_79475_comb = smul20b_20b_x_7b(p1_sign_ext_78562_comb[19:0], 7'h31);
  assign p1_smul_79478_comb = smul20b_20b_x_7b(p1_sign_ext_78565_comb[19:0], 7'h31);
  assign p1_smul_79481_comb = smul20b_20b_x_7b(p1_sign_ext_78677_comb[19:0], 7'h31);
  assign p1_smul_79482_comb = smul20b_20b_x_7b(p1_sign_ext_78678_comb[19:0], 7'h31);
  assign p1_smul_79485_comb = smul20b_20b_x_7b(p1_sign_ext_78570_comb[19:0], 7'h31);
  assign p1_smul_79488_comb = smul20b_20b_x_7b(p1_sign_ext_78573_comb[19:0], 7'h31);
  assign p1_smul_79491_comb = smul20b_20b_x_7b(p1_sign_ext_78683_comb[19:0], 7'h31);
  assign p1_smul_79492_comb = smul20b_20b_x_7b(p1_sign_ext_78684_comb[19:0], 7'h31);
  assign p1_smul_79495_comb = smul20b_20b_x_7b(p1_sign_ext_78578_comb[19:0], 7'h31);
  assign p1_smul_79498_comb = smul20b_20b_x_7b(p1_sign_ext_78581_comb[19:0], 7'h31);
  assign p1_smul_79501_comb = smul20b_20b_x_7b(p1_sign_ext_78689_comb[19:0], 7'h31);
  assign p1_smul_79502_comb = smul20b_20b_x_7b(p1_sign_ext_78690_comb[19:0], 7'h31);
  assign p1_smul_79505_comb = smul20b_20b_x_7b(p1_sign_ext_78586_comb[19:0], 7'h31);
  assign p1_smul_79508_comb = smul20b_20b_x_7b(p1_sign_ext_78589_comb[19:0], 7'h31);
  assign p1_smul_79511_comb = smul20b_20b_x_7b(p1_sign_ext_78695_comb[19:0], 7'h31);
  assign p1_smul_79512_comb = smul20b_20b_x_7b(p1_sign_ext_78696_comb[19:0], 7'h31);
  assign p1_smul_79515_comb = smul20b_20b_x_7b(p1_sign_ext_78594_comb[19:0], 7'h31);
  assign p1_smul_79518_comb = smul20b_20b_x_7b(p1_sign_ext_78597_comb[19:0], 7'h31);
  assign p1_smul_79521_comb = smul20b_20b_x_7b(p1_sign_ext_78701_comb[19:0], 7'h31);
  assign p1_smul_79522_comb = smul20b_20b_x_7b(p1_sign_ext_78702_comb[19:0], 7'h31);
  assign p1_smul_79525_comb = smul20b_20b_x_7b(p1_sign_ext_78602_comb[19:0], 7'h31);
  assign p1_smul_79528_comb = smul20b_20b_x_7b(p1_sign_ext_78605_comb[19:0], 7'h31);
  assign p1_smul_79531_comb = smul20b_20b_x_7b(p1_sign_ext_78707_comb[19:0], 7'h31);
  assign p1_smul_79532_comb = smul20b_20b_x_7b(p1_sign_ext_78708_comb[19:0], 7'h31);
  assign p1_smul_79535_comb = smul20b_20b_x_7b(p1_sign_ext_78610_comb[19:0], 7'h31);
  assign p1_smul_79538_comb = smul20b_20b_x_7b(p1_sign_ext_78613_comb[19:0], 7'h31);
  assign p1_smul_79541_comb = smul20b_20b_x_7b(p1_sign_ext_78713_comb[19:0], 7'h31);
  assign p1_smul_79542_comb = smul20b_20b_x_7b(p1_sign_ext_78714_comb[19:0], 7'h31);
  assign p1_smul_79545_comb = smul20b_20b_x_7b(p1_sign_ext_78618_comb[19:0], 7'h31);
  assign p1_smul_79548_comb = smul20b_20b_x_7b(p1_sign_ext_78621_comb[19:0], 7'h31);
  assign p1_smul_79551_comb = smul20b_20b_x_7b(p1_sign_ext_78719_comb[19:0], 7'h31);
  assign p1_smul_79552_comb = smul20b_20b_x_6b(p1_sign_ext_78672_comb[19:0], 6'h19);
  assign p1_smul_79553_comb = smul20b_20b_x_8b(p1_sign_ext_78624_comb[19:0], 8'hb9);
  assign p1_add_79554_comb = p1_smul_79074_comb + p1_smul_79075_comb;
  assign p1_add_79555_comb = p1_smul_79076_comb + p1_smul_79077_comb;
  assign p1_smul_79556_comb = smul20b_20b_x_8b(p1_sign_ext_78625_comb[19:0], 8'hb9);
  assign p1_smul_79557_comb = smul20b_20b_x_6b(p1_sign_ext_78677_comb[19:0], 6'h19);
  assign p1_smul_79558_comb = smul20b_20b_x_6b(p1_sign_ext_78678_comb[19:0], 6'h19);
  assign p1_smul_79559_comb = smul20b_20b_x_8b(p1_sign_ext_78626_comb[19:0], 8'hb9);
  assign p1_add_79560_comb = p1_smul_79082_comb + p1_smul_79083_comb;
  assign p1_add_79561_comb = p1_smul_79084_comb + p1_smul_79085_comb;
  assign p1_smul_79562_comb = smul20b_20b_x_8b(p1_sign_ext_78627_comb[19:0], 8'hb9);
  assign p1_smul_79563_comb = smul20b_20b_x_6b(p1_sign_ext_78683_comb[19:0], 6'h19);
  assign p1_smul_79564_comb = smul20b_20b_x_6b(p1_sign_ext_78684_comb[19:0], 6'h19);
  assign p1_smul_79565_comb = smul20b_20b_x_8b(p1_sign_ext_78628_comb[19:0], 8'hb9);
  assign p1_add_79566_comb = p1_smul_79090_comb + p1_smul_79091_comb;
  assign p1_add_79567_comb = p1_smul_79092_comb + p1_smul_79093_comb;
  assign p1_smul_79568_comb = smul20b_20b_x_8b(p1_sign_ext_78629_comb[19:0], 8'hb9);
  assign p1_smul_79569_comb = smul20b_20b_x_6b(p1_sign_ext_78689_comb[19:0], 6'h19);
  assign p1_smul_79570_comb = smul20b_20b_x_6b(p1_sign_ext_78690_comb[19:0], 6'h19);
  assign p1_smul_79571_comb = smul20b_20b_x_8b(p1_sign_ext_78630_comb[19:0], 8'hb9);
  assign p1_add_79572_comb = p1_smul_79098_comb + p1_smul_79099_comb;
  assign p1_add_79573_comb = p1_smul_79100_comb + p1_smul_79101_comb;
  assign p1_smul_79574_comb = smul20b_20b_x_8b(p1_sign_ext_78631_comb[19:0], 8'hb9);
  assign p1_smul_79575_comb = smul20b_20b_x_6b(p1_sign_ext_78695_comb[19:0], 6'h19);
  assign p1_smul_79576_comb = smul20b_20b_x_6b(p1_sign_ext_78696_comb[19:0], 6'h19);
  assign p1_smul_79577_comb = smul20b_20b_x_8b(p1_sign_ext_78632_comb[19:0], 8'hb9);
  assign p1_add_79578_comb = p1_smul_79106_comb + p1_smul_79107_comb;
  assign p1_add_79579_comb = p1_smul_79108_comb + p1_smul_79109_comb;
  assign p1_smul_79580_comb = smul20b_20b_x_8b(p1_sign_ext_78633_comb[19:0], 8'hb9);
  assign p1_smul_79581_comb = smul20b_20b_x_6b(p1_sign_ext_78701_comb[19:0], 6'h19);
  assign p1_smul_79582_comb = smul20b_20b_x_6b(p1_sign_ext_78702_comb[19:0], 6'h19);
  assign p1_smul_79583_comb = smul20b_20b_x_8b(p1_sign_ext_78634_comb[19:0], 8'hb9);
  assign p1_add_79584_comb = p1_smul_79114_comb + p1_smul_79115_comb;
  assign p1_add_79585_comb = p1_smul_79116_comb + p1_smul_79117_comb;
  assign p1_smul_79586_comb = smul20b_20b_x_8b(p1_sign_ext_78635_comb[19:0], 8'hb9);
  assign p1_smul_79587_comb = smul20b_20b_x_6b(p1_sign_ext_78707_comb[19:0], 6'h19);
  assign p1_smul_79588_comb = smul20b_20b_x_6b(p1_sign_ext_78708_comb[19:0], 6'h19);
  assign p1_smul_79589_comb = smul20b_20b_x_8b(p1_sign_ext_78636_comb[19:0], 8'hb9);
  assign p1_add_79590_comb = p1_smul_79122_comb + p1_smul_79123_comb;
  assign p1_add_79591_comb = p1_smul_79124_comb + p1_smul_79125_comb;
  assign p1_smul_79592_comb = smul20b_20b_x_8b(p1_sign_ext_78637_comb[19:0], 8'hb9);
  assign p1_smul_79593_comb = smul20b_20b_x_6b(p1_sign_ext_78713_comb[19:0], 6'h19);
  assign p1_smul_79594_comb = smul20b_20b_x_6b(p1_sign_ext_78714_comb[19:0], 6'h19);
  assign p1_smul_79595_comb = smul20b_20b_x_8b(p1_sign_ext_78638_comb[19:0], 8'hb9);
  assign p1_add_79596_comb = p1_smul_79130_comb + p1_smul_79131_comb;
  assign p1_add_79597_comb = p1_smul_79132_comb + p1_smul_79133_comb;
  assign p1_smul_79598_comb = smul20b_20b_x_8b(p1_sign_ext_78639_comb[19:0], 8'hb9);
  assign p1_smul_79599_comb = smul20b_20b_x_6b(p1_sign_ext_78719_comb[19:0], 6'h19);
  assign p1_bit_slice_79664_comb = p1_add_79136_comb[20:1];
  assign p1_add_79665_comb = p1_smul_79137_comb + p1_smul_79138_comb;
  assign p1_add_79666_comb = p1_smul_79139_comb + p1_smul_79140_comb;
  assign p1_bit_slice_79667_comb = p1_add_79141_comb[20:1];
  assign p1_bit_slice_79668_comb = p1_add_79142_comb[20:1];
  assign p1_add_79669_comb = p1_smul_79143_comb + p1_smul_79144_comb;
  assign p1_add_79670_comb = p1_smul_79145_comb + p1_smul_79146_comb;
  assign p1_bit_slice_79671_comb = p1_add_79147_comb[20:1];
  assign p1_bit_slice_79672_comb = p1_add_79148_comb[20:1];
  assign p1_add_79673_comb = p1_smul_79149_comb + p1_smul_79150_comb;
  assign p1_add_79674_comb = p1_smul_79151_comb + p1_smul_79152_comb;
  assign p1_bit_slice_79675_comb = p1_add_79153_comb[20:1];
  assign p1_bit_slice_79676_comb = p1_add_79154_comb[20:1];
  assign p1_add_79677_comb = p1_smul_79155_comb + p1_smul_79156_comb;
  assign p1_add_79678_comb = p1_smul_79157_comb + p1_smul_79158_comb;
  assign p1_bit_slice_79679_comb = p1_add_79159_comb[20:1];
  assign p1_bit_slice_79680_comb = p1_add_79160_comb[20:1];
  assign p1_add_79681_comb = p1_smul_79161_comb + p1_smul_79162_comb;
  assign p1_add_79682_comb = p1_smul_79163_comb + p1_smul_79164_comb;
  assign p1_bit_slice_79683_comb = p1_add_79165_comb[20:1];
  assign p1_bit_slice_79684_comb = p1_add_79166_comb[20:1];
  assign p1_add_79685_comb = p1_smul_79167_comb + p1_smul_79168_comb;
  assign p1_add_79686_comb = p1_smul_79169_comb + p1_smul_79170_comb;
  assign p1_bit_slice_79687_comb = p1_add_79171_comb[20:1];
  assign p1_bit_slice_79688_comb = p1_add_79172_comb[20:1];
  assign p1_add_79689_comb = p1_smul_79173_comb + p1_smul_79174_comb;
  assign p1_add_79690_comb = p1_smul_79175_comb + p1_smul_79176_comb;
  assign p1_bit_slice_79691_comb = p1_add_79177_comb[20:1];
  assign p1_bit_slice_79692_comb = p1_add_79178_comb[20:1];
  assign p1_add_79693_comb = p1_smul_79179_comb + p1_smul_79180_comb;
  assign p1_add_79694_comb = p1_smul_79181_comb + p1_smul_79182_comb;
  assign p1_bit_slice_79695_comb = p1_add_79183_comb[20:1];
  assign p1_smul_79696_comb = smul19b_19b_x_7b(p1_sign_ext_78672_comb[18:0], 7'h3b);
  assign p1_smul_79699_comb = smul19b_19b_x_7b(p1_sign_ext_78563_comb[18:0], 7'h45);
  assign p1_smul_79700_comb = smul19b_19b_x_7b(p1_sign_ext_78564_comb[18:0], 7'h45);
  assign p1_smul_79703_comb = smul19b_19b_x_7b(p1_sign_ext_78677_comb[18:0], 7'h3b);
  assign p1_smul_79704_comb = smul19b_19b_x_7b(p1_sign_ext_78678_comb[18:0], 7'h3b);
  assign p1_smul_79707_comb = smul19b_19b_x_7b(p1_sign_ext_78571_comb[18:0], 7'h45);
  assign p1_smul_79708_comb = smul19b_19b_x_7b(p1_sign_ext_78572_comb[18:0], 7'h45);
  assign p1_smul_79711_comb = smul19b_19b_x_7b(p1_sign_ext_78683_comb[18:0], 7'h3b);
  assign p1_smul_79712_comb = smul19b_19b_x_7b(p1_sign_ext_78684_comb[18:0], 7'h3b);
  assign p1_smul_79715_comb = smul19b_19b_x_7b(p1_sign_ext_78579_comb[18:0], 7'h45);
  assign p1_smul_79716_comb = smul19b_19b_x_7b(p1_sign_ext_78580_comb[18:0], 7'h45);
  assign p1_smul_79719_comb = smul19b_19b_x_7b(p1_sign_ext_78689_comb[18:0], 7'h3b);
  assign p1_smul_79720_comb = smul19b_19b_x_7b(p1_sign_ext_78690_comb[18:0], 7'h3b);
  assign p1_smul_79723_comb = smul19b_19b_x_7b(p1_sign_ext_78587_comb[18:0], 7'h45);
  assign p1_smul_79724_comb = smul19b_19b_x_7b(p1_sign_ext_78588_comb[18:0], 7'h45);
  assign p1_smul_79727_comb = smul19b_19b_x_7b(p1_sign_ext_78695_comb[18:0], 7'h3b);
  assign p1_smul_79728_comb = smul19b_19b_x_7b(p1_sign_ext_78696_comb[18:0], 7'h3b);
  assign p1_smul_79731_comb = smul19b_19b_x_7b(p1_sign_ext_78595_comb[18:0], 7'h45);
  assign p1_smul_79732_comb = smul19b_19b_x_7b(p1_sign_ext_78596_comb[18:0], 7'h45);
  assign p1_smul_79735_comb = smul19b_19b_x_7b(p1_sign_ext_78701_comb[18:0], 7'h3b);
  assign p1_smul_79736_comb = smul19b_19b_x_7b(p1_sign_ext_78702_comb[18:0], 7'h3b);
  assign p1_smul_79739_comb = smul19b_19b_x_7b(p1_sign_ext_78603_comb[18:0], 7'h45);
  assign p1_smul_79740_comb = smul19b_19b_x_7b(p1_sign_ext_78604_comb[18:0], 7'h45);
  assign p1_smul_79743_comb = smul19b_19b_x_7b(p1_sign_ext_78707_comb[18:0], 7'h3b);
  assign p1_smul_79744_comb = smul19b_19b_x_7b(p1_sign_ext_78708_comb[18:0], 7'h3b);
  assign p1_smul_79747_comb = smul19b_19b_x_7b(p1_sign_ext_78611_comb[18:0], 7'h45);
  assign p1_smul_79748_comb = smul19b_19b_x_7b(p1_sign_ext_78612_comb[18:0], 7'h45);
  assign p1_smul_79751_comb = smul19b_19b_x_7b(p1_sign_ext_78713_comb[18:0], 7'h3b);
  assign p1_smul_79752_comb = smul19b_19b_x_7b(p1_sign_ext_78714_comb[18:0], 7'h3b);
  assign p1_smul_79755_comb = smul19b_19b_x_7b(p1_sign_ext_78619_comb[18:0], 7'h45);
  assign p1_smul_79756_comb = smul19b_19b_x_7b(p1_sign_ext_78620_comb[18:0], 7'h45);
  assign p1_smul_79759_comb = smul19b_19b_x_7b(p1_sign_ext_78719_comb[18:0], 7'h3b);
  assign p1_add_79760_comb = p1_smul_78896_comb[20:1] + p1_smul_79281_comb;
  assign p1_add_79762_comb = p1_smul_78898_comb[20:1] + p1_smul_79283_comb;
  assign p1_add_79764_comb = p1_smul_79284_comb + p1_smul_78901_comb[20:1];
  assign p1_add_79766_comb = p1_smul_79286_comb + p1_smul_78903_comb[20:1];
  assign p1_add_79768_comb = p1_smul_78904_comb[20:1] + p1_smul_79289_comb;
  assign p1_add_79770_comb = p1_smul_78906_comb[20:1] + p1_smul_79291_comb;
  assign p1_add_79772_comb = p1_smul_79292_comb + p1_smul_78909_comb[20:1];
  assign p1_add_79774_comb = p1_smul_79294_comb + p1_smul_78911_comb[20:1];
  assign p1_add_79776_comb = p1_smul_78912_comb[20:1] + p1_smul_79297_comb;
  assign p1_add_79778_comb = p1_smul_78914_comb[20:1] + p1_smul_79299_comb;
  assign p1_add_79780_comb = p1_smul_79300_comb + p1_smul_78917_comb[20:1];
  assign p1_add_79782_comb = p1_smul_79302_comb + p1_smul_78919_comb[20:1];
  assign p1_add_79784_comb = p1_smul_78920_comb[20:1] + p1_smul_79305_comb;
  assign p1_add_79786_comb = p1_smul_78922_comb[20:1] + p1_smul_79307_comb;
  assign p1_add_79788_comb = p1_smul_79308_comb + p1_smul_78925_comb[20:1];
  assign p1_add_79790_comb = p1_smul_79310_comb + p1_smul_78927_comb[20:1];
  assign p1_add_79792_comb = p1_smul_78928_comb[20:1] + p1_smul_79313_comb;
  assign p1_add_79794_comb = p1_smul_78930_comb[20:1] + p1_smul_79315_comb;
  assign p1_add_79796_comb = p1_smul_79316_comb + p1_smul_78933_comb[20:1];
  assign p1_add_79798_comb = p1_smul_79318_comb + p1_smul_78935_comb[20:1];
  assign p1_add_79800_comb = p1_smul_78936_comb[20:1] + p1_smul_79321_comb;
  assign p1_add_79802_comb = p1_smul_78938_comb[20:1] + p1_smul_79323_comb;
  assign p1_add_79804_comb = p1_smul_79324_comb + p1_smul_78941_comb[20:1];
  assign p1_add_79806_comb = p1_smul_79326_comb + p1_smul_78943_comb[20:1];
  assign p1_add_79808_comb = p1_smul_78944_comb[20:1] + p1_smul_79329_comb;
  assign p1_add_79810_comb = p1_smul_78946_comb[20:1] + p1_smul_79331_comb;
  assign p1_add_79812_comb = p1_smul_79332_comb + p1_smul_78949_comb[20:1];
  assign p1_add_79814_comb = p1_smul_79334_comb + p1_smul_78951_comb[20:1];
  assign p1_add_79816_comb = p1_smul_78952_comb[20:1] + p1_smul_79337_comb;
  assign p1_add_79818_comb = p1_smul_78954_comb[20:1] + p1_smul_79339_comb;
  assign p1_add_79820_comb = p1_smul_79340_comb + p1_smul_78957_comb[20:1];
  assign p1_add_79822_comb = p1_smul_79342_comb + p1_smul_78959_comb[20:1];
  assign p1_smul_79824_comb = smul21b_12b_x_9b(p1_clipped__8_comb, 9'h0b5);
  assign p1_smul_79825_comb = smul21b_12b_x_9b(p1_clipped__24_comb, 9'h14b);
  assign p1_smul_79826_comb = smul21b_12b_x_9b(p1_clipped__40_comb, 9'h14b);
  assign p1_smul_79827_comb = smul21b_12b_x_9b(p1_clipped__56_comb, 9'h0b5);
  assign p1_smul_79828_comb = smul21b_12b_x_9b(p1_clipped__72_comb, 9'h0b5);
  assign p1_smul_79829_comb = smul21b_12b_x_9b(p1_clipped__88_comb, 9'h14b);
  assign p1_smul_79830_comb = smul21b_12b_x_9b(p1_clipped__104_comb, 9'h14b);
  assign p1_smul_79831_comb = smul21b_12b_x_9b(p1_clipped__120_comb, 9'h0b5);
  assign p1_smul_79832_comb = smul21b_12b_x_9b(p1_clipped__9_comb, 9'h0b5);
  assign p1_smul_79833_comb = smul21b_12b_x_9b(p1_clipped__25_comb, 9'h14b);
  assign p1_smul_79834_comb = smul21b_12b_x_9b(p1_clipped__41_comb, 9'h14b);
  assign p1_smul_79835_comb = smul21b_12b_x_9b(p1_clipped__57_comb, 9'h0b5);
  assign p1_smul_79836_comb = smul21b_12b_x_9b(p1_clipped__73_comb, 9'h0b5);
  assign p1_smul_79837_comb = smul21b_12b_x_9b(p1_clipped__89_comb, 9'h14b);
  assign p1_smul_79838_comb = smul21b_12b_x_9b(p1_clipped__105_comb, 9'h14b);
  assign p1_smul_79839_comb = smul21b_12b_x_9b(p1_clipped__121_comb, 9'h0b5);
  assign p1_smul_79840_comb = smul21b_12b_x_9b(p1_clipped__10_comb, 9'h0b5);
  assign p1_smul_79841_comb = smul21b_12b_x_9b(p1_clipped__26_comb, 9'h14b);
  assign p1_smul_79842_comb = smul21b_12b_x_9b(p1_clipped__42_comb, 9'h14b);
  assign p1_smul_79843_comb = smul21b_12b_x_9b(p1_clipped__58_comb, 9'h0b5);
  assign p1_smul_79844_comb = smul21b_12b_x_9b(p1_clipped__74_comb, 9'h0b5);
  assign p1_smul_79845_comb = smul21b_12b_x_9b(p1_clipped__90_comb, 9'h14b);
  assign p1_smul_79846_comb = smul21b_12b_x_9b(p1_clipped__106_comb, 9'h14b);
  assign p1_smul_79847_comb = smul21b_12b_x_9b(p1_clipped__122_comb, 9'h0b5);
  assign p1_smul_79848_comb = smul21b_12b_x_9b(p1_clipped__11_comb, 9'h0b5);
  assign p1_smul_79849_comb = smul21b_12b_x_9b(p1_clipped__27_comb, 9'h14b);
  assign p1_smul_79850_comb = smul21b_12b_x_9b(p1_clipped__43_comb, 9'h14b);
  assign p1_smul_79851_comb = smul21b_12b_x_9b(p1_clipped__59_comb, 9'h0b5);
  assign p1_smul_79852_comb = smul21b_12b_x_9b(p1_clipped__75_comb, 9'h0b5);
  assign p1_smul_79853_comb = smul21b_12b_x_9b(p1_clipped__91_comb, 9'h14b);
  assign p1_smul_79854_comb = smul21b_12b_x_9b(p1_clipped__107_comb, 9'h14b);
  assign p1_smul_79855_comb = smul21b_12b_x_9b(p1_clipped__123_comb, 9'h0b5);
  assign p1_smul_79856_comb = smul21b_12b_x_9b(p1_clipped__12_comb, 9'h0b5);
  assign p1_smul_79857_comb = smul21b_12b_x_9b(p1_clipped__28_comb, 9'h14b);
  assign p1_smul_79858_comb = smul21b_12b_x_9b(p1_clipped__44_comb, 9'h14b);
  assign p1_smul_79859_comb = smul21b_12b_x_9b(p1_clipped__60_comb, 9'h0b5);
  assign p1_smul_79860_comb = smul21b_12b_x_9b(p1_clipped__76_comb, 9'h0b5);
  assign p1_smul_79861_comb = smul21b_12b_x_9b(p1_clipped__92_comb, 9'h14b);
  assign p1_smul_79862_comb = smul21b_12b_x_9b(p1_clipped__108_comb, 9'h14b);
  assign p1_smul_79863_comb = smul21b_12b_x_9b(p1_clipped__124_comb, 9'h0b5);
  assign p1_smul_79864_comb = smul21b_12b_x_9b(p1_clipped__13_comb, 9'h0b5);
  assign p1_smul_79865_comb = smul21b_12b_x_9b(p1_clipped__29_comb, 9'h14b);
  assign p1_smul_79866_comb = smul21b_12b_x_9b(p1_clipped__45_comb, 9'h14b);
  assign p1_smul_79867_comb = smul21b_12b_x_9b(p1_clipped__61_comb, 9'h0b5);
  assign p1_smul_79868_comb = smul21b_12b_x_9b(p1_clipped__77_comb, 9'h0b5);
  assign p1_smul_79869_comb = smul21b_12b_x_9b(p1_clipped__93_comb, 9'h14b);
  assign p1_smul_79870_comb = smul21b_12b_x_9b(p1_clipped__109_comb, 9'h14b);
  assign p1_smul_79871_comb = smul21b_12b_x_9b(p1_clipped__125_comb, 9'h0b5);
  assign p1_smul_79872_comb = smul21b_12b_x_9b(p1_clipped__14_comb, 9'h0b5);
  assign p1_smul_79873_comb = smul21b_12b_x_9b(p1_clipped__30_comb, 9'h14b);
  assign p1_smul_79874_comb = smul21b_12b_x_9b(p1_clipped__46_comb, 9'h14b);
  assign p1_smul_79875_comb = smul21b_12b_x_9b(p1_clipped__62_comb, 9'h0b5);
  assign p1_smul_79876_comb = smul21b_12b_x_9b(p1_clipped__78_comb, 9'h0b5);
  assign p1_smul_79877_comb = smul21b_12b_x_9b(p1_clipped__94_comb, 9'h14b);
  assign p1_smul_79878_comb = smul21b_12b_x_9b(p1_clipped__110_comb, 9'h14b);
  assign p1_smul_79879_comb = smul21b_12b_x_9b(p1_clipped__126_comb, 9'h0b5);
  assign p1_smul_79880_comb = smul21b_12b_x_9b(p1_clipped__15_comb, 9'h0b5);
  assign p1_smul_79881_comb = smul21b_12b_x_9b(p1_clipped__31_comb, 9'h14b);
  assign p1_smul_79882_comb = smul21b_12b_x_9b(p1_clipped__47_comb, 9'h14b);
  assign p1_smul_79883_comb = smul21b_12b_x_9b(p1_clipped__63_comb, 9'h0b5);
  assign p1_smul_79884_comb = smul21b_12b_x_9b(p1_clipped__79_comb, 9'h0b5);
  assign p1_smul_79885_comb = smul21b_12b_x_9b(p1_clipped__95_comb, 9'h14b);
  assign p1_smul_79886_comb = smul21b_12b_x_9b(p1_clipped__111_comb, 9'h14b);
  assign p1_smul_79887_comb = smul21b_12b_x_9b(p1_clipped__127_comb, 9'h0b5);
  assign p1_add_79888_comb = p1_smul_79408_comb + p1_smul_78962_comb[20:1];
  assign p1_add_79890_comb = p1_smul_79410_comb + p1_smul_78964_comb[20:1];
  assign p1_add_79892_comb = p1_smul_78965_comb[20:1] + p1_smul_79413_comb;
  assign p1_add_79894_comb = p1_smul_78967_comb[20:1] + p1_smul_79415_comb;
  assign p1_add_79896_comb = p1_smul_79416_comb + p1_smul_78972_comb[20:1];
  assign p1_add_79898_comb = p1_smul_79418_comb + p1_smul_78974_comb[20:1];
  assign p1_add_79900_comb = p1_smul_78975_comb[20:1] + p1_smul_79421_comb;
  assign p1_add_79902_comb = p1_smul_78977_comb[20:1] + p1_smul_79423_comb;
  assign p1_add_79904_comb = p1_smul_79424_comb + p1_smul_78982_comb[20:1];
  assign p1_add_79906_comb = p1_smul_79426_comb + p1_smul_78984_comb[20:1];
  assign p1_add_79908_comb = p1_smul_78985_comb[20:1] + p1_smul_79429_comb;
  assign p1_add_79910_comb = p1_smul_78987_comb[20:1] + p1_smul_79431_comb;
  assign p1_add_79912_comb = p1_smul_79432_comb + p1_smul_78992_comb[20:1];
  assign p1_add_79914_comb = p1_smul_79434_comb + p1_smul_78994_comb[20:1];
  assign p1_add_79916_comb = p1_smul_78995_comb[20:1] + p1_smul_79437_comb;
  assign p1_add_79918_comb = p1_smul_78997_comb[20:1] + p1_smul_79439_comb;
  assign p1_add_79920_comb = p1_smul_79440_comb + p1_smul_79002_comb[20:1];
  assign p1_add_79922_comb = p1_smul_79442_comb + p1_smul_79004_comb[20:1];
  assign p1_add_79924_comb = p1_smul_79005_comb[20:1] + p1_smul_79445_comb;
  assign p1_add_79926_comb = p1_smul_79007_comb[20:1] + p1_smul_79447_comb;
  assign p1_add_79928_comb = p1_smul_79448_comb + p1_smul_79012_comb[20:1];
  assign p1_add_79930_comb = p1_smul_79450_comb + p1_smul_79014_comb[20:1];
  assign p1_add_79932_comb = p1_smul_79015_comb[20:1] + p1_smul_79453_comb;
  assign p1_add_79934_comb = p1_smul_79017_comb[20:1] + p1_smul_79455_comb;
  assign p1_add_79936_comb = p1_smul_79456_comb + p1_smul_79022_comb[20:1];
  assign p1_add_79938_comb = p1_smul_79458_comb + p1_smul_79024_comb[20:1];
  assign p1_add_79940_comb = p1_smul_79025_comb[20:1] + p1_smul_79461_comb;
  assign p1_add_79942_comb = p1_smul_79027_comb[20:1] + p1_smul_79463_comb;
  assign p1_add_79944_comb = p1_smul_79464_comb + p1_smul_79032_comb[20:1];
  assign p1_add_79946_comb = p1_smul_79466_comb + p1_smul_79034_comb[20:1];
  assign p1_add_79948_comb = p1_smul_79035_comb[20:1] + p1_smul_79469_comb;
  assign p1_add_79950_comb = p1_smul_79037_comb[20:1] + p1_smul_79471_comb;
  assign p1_smul_79953_comb = smul19b_19b_x_7b(p1_sign_ext_78624_comb[18:0], 7'h45);
  assign p1_smul_79955_comb = smul19b_19b_x_7b(p1_sign_ext_78563_comb[18:0], 7'h3b);
  assign p1_smul_79956_comb = smul19b_19b_x_7b(p1_sign_ext_78564_comb[18:0], 7'h3b);
  assign p1_smul_79958_comb = smul19b_19b_x_7b(p1_sign_ext_78625_comb[18:0], 7'h45);
  assign p1_smul_79961_comb = smul19b_19b_x_7b(p1_sign_ext_78626_comb[18:0], 7'h45);
  assign p1_smul_79963_comb = smul19b_19b_x_7b(p1_sign_ext_78571_comb[18:0], 7'h3b);
  assign p1_smul_79964_comb = smul19b_19b_x_7b(p1_sign_ext_78572_comb[18:0], 7'h3b);
  assign p1_smul_79966_comb = smul19b_19b_x_7b(p1_sign_ext_78627_comb[18:0], 7'h45);
  assign p1_smul_79969_comb = smul19b_19b_x_7b(p1_sign_ext_78628_comb[18:0], 7'h45);
  assign p1_smul_79971_comb = smul19b_19b_x_7b(p1_sign_ext_78579_comb[18:0], 7'h3b);
  assign p1_smul_79972_comb = smul19b_19b_x_7b(p1_sign_ext_78580_comb[18:0], 7'h3b);
  assign p1_smul_79974_comb = smul19b_19b_x_7b(p1_sign_ext_78629_comb[18:0], 7'h45);
  assign p1_smul_79977_comb = smul19b_19b_x_7b(p1_sign_ext_78630_comb[18:0], 7'h45);
  assign p1_smul_79979_comb = smul19b_19b_x_7b(p1_sign_ext_78587_comb[18:0], 7'h3b);
  assign p1_smul_79980_comb = smul19b_19b_x_7b(p1_sign_ext_78588_comb[18:0], 7'h3b);
  assign p1_smul_79982_comb = smul19b_19b_x_7b(p1_sign_ext_78631_comb[18:0], 7'h45);
  assign p1_smul_79985_comb = smul19b_19b_x_7b(p1_sign_ext_78632_comb[18:0], 7'h45);
  assign p1_smul_79987_comb = smul19b_19b_x_7b(p1_sign_ext_78595_comb[18:0], 7'h3b);
  assign p1_smul_79988_comb = smul19b_19b_x_7b(p1_sign_ext_78596_comb[18:0], 7'h3b);
  assign p1_smul_79990_comb = smul19b_19b_x_7b(p1_sign_ext_78633_comb[18:0], 7'h45);
  assign p1_smul_79993_comb = smul19b_19b_x_7b(p1_sign_ext_78634_comb[18:0], 7'h45);
  assign p1_smul_79995_comb = smul19b_19b_x_7b(p1_sign_ext_78603_comb[18:0], 7'h3b);
  assign p1_smul_79996_comb = smul19b_19b_x_7b(p1_sign_ext_78604_comb[18:0], 7'h3b);
  assign p1_smul_79998_comb = smul19b_19b_x_7b(p1_sign_ext_78635_comb[18:0], 7'h45);
  assign p1_smul_80001_comb = smul19b_19b_x_7b(p1_sign_ext_78636_comb[18:0], 7'h45);
  assign p1_smul_80003_comb = smul19b_19b_x_7b(p1_sign_ext_78611_comb[18:0], 7'h3b);
  assign p1_smul_80004_comb = smul19b_19b_x_7b(p1_sign_ext_78612_comb[18:0], 7'h3b);
  assign p1_smul_80006_comb = smul19b_19b_x_7b(p1_sign_ext_78637_comb[18:0], 7'h45);
  assign p1_smul_80009_comb = smul19b_19b_x_7b(p1_sign_ext_78638_comb[18:0], 7'h45);
  assign p1_smul_80011_comb = smul19b_19b_x_7b(p1_sign_ext_78619_comb[18:0], 7'h3b);
  assign p1_smul_80012_comb = smul19b_19b_x_7b(p1_sign_ext_78620_comb[18:0], 7'h3b);
  assign p1_smul_80014_comb = smul19b_19b_x_7b(p1_sign_ext_78639_comb[18:0], 7'h45);
  assign p1_add_80016_comb = p1_smul_79552_comb + p1_smul_79553_comb;
  assign p1_bit_slice_80017_comb = p1_add_79554_comb[20:1];
  assign p1_bit_slice_80018_comb = p1_add_79555_comb[20:1];
  assign p1_add_80019_comb = p1_smul_79556_comb + p1_smul_79557_comb;
  assign p1_add_80020_comb = p1_smul_79558_comb + p1_smul_79559_comb;
  assign p1_bit_slice_80021_comb = p1_add_79560_comb[20:1];
  assign p1_bit_slice_80022_comb = p1_add_79561_comb[20:1];
  assign p1_add_80023_comb = p1_smul_79562_comb + p1_smul_79563_comb;
  assign p1_add_80024_comb = p1_smul_79564_comb + p1_smul_79565_comb;
  assign p1_bit_slice_80025_comb = p1_add_79566_comb[20:1];
  assign p1_bit_slice_80026_comb = p1_add_79567_comb[20:1];
  assign p1_add_80027_comb = p1_smul_79568_comb + p1_smul_79569_comb;
  assign p1_add_80028_comb = p1_smul_79570_comb + p1_smul_79571_comb;
  assign p1_bit_slice_80029_comb = p1_add_79572_comb[20:1];
  assign p1_bit_slice_80030_comb = p1_add_79573_comb[20:1];
  assign p1_add_80031_comb = p1_smul_79574_comb + p1_smul_79575_comb;
  assign p1_add_80032_comb = p1_smul_79576_comb + p1_smul_79577_comb;
  assign p1_bit_slice_80033_comb = p1_add_79578_comb[20:1];
  assign p1_bit_slice_80034_comb = p1_add_79579_comb[20:1];
  assign p1_add_80035_comb = p1_smul_79580_comb + p1_smul_79581_comb;
  assign p1_add_80036_comb = p1_smul_79582_comb + p1_smul_79583_comb;
  assign p1_bit_slice_80037_comb = p1_add_79584_comb[20:1];
  assign p1_bit_slice_80038_comb = p1_add_79585_comb[20:1];
  assign p1_add_80039_comb = p1_smul_79586_comb + p1_smul_79587_comb;
  assign p1_add_80040_comb = p1_smul_79588_comb + p1_smul_79589_comb;
  assign p1_bit_slice_80041_comb = p1_add_79590_comb[20:1];
  assign p1_bit_slice_80042_comb = p1_add_79591_comb[20:1];
  assign p1_add_80043_comb = p1_smul_79592_comb + p1_smul_79593_comb;
  assign p1_add_80044_comb = p1_smul_79594_comb + p1_smul_79595_comb;
  assign p1_bit_slice_80045_comb = p1_add_79596_comb[20:1];
  assign p1_bit_slice_80046_comb = p1_add_79597_comb[20:1];
  assign p1_add_80047_comb = p1_smul_79598_comb + p1_smul_79599_comb;
  assign p1_add_80048_comb = p1_sign_ext_78672_comb[12:0] + p1_sign_ext_78624_comb[12:0];
  assign p1_add_80049_comb = p1_sign_ext_78562_comb[12:0] + p1_sign_ext_78563_comb[12:0];
  assign p1_add_80050_comb = p1_sign_ext_78564_comb[12:0] + p1_sign_ext_78565_comb[12:0];
  assign p1_add_80051_comb = p1_sign_ext_78625_comb[12:0] + p1_sign_ext_78677_comb[12:0];
  assign p1_add_80052_comb = p1_sign_ext_78678_comb[12:0] + p1_sign_ext_78626_comb[12:0];
  assign p1_add_80053_comb = p1_sign_ext_78570_comb[12:0] + p1_sign_ext_78571_comb[12:0];
  assign p1_add_80054_comb = p1_sign_ext_78572_comb[12:0] + p1_sign_ext_78573_comb[12:0];
  assign p1_add_80055_comb = p1_sign_ext_78627_comb[12:0] + p1_sign_ext_78683_comb[12:0];
  assign p1_add_80056_comb = p1_sign_ext_78684_comb[12:0] + p1_sign_ext_78628_comb[12:0];
  assign p1_add_80057_comb = p1_sign_ext_78578_comb[12:0] + p1_sign_ext_78579_comb[12:0];
  assign p1_add_80058_comb = p1_sign_ext_78580_comb[12:0] + p1_sign_ext_78581_comb[12:0];
  assign p1_add_80059_comb = p1_sign_ext_78629_comb[12:0] + p1_sign_ext_78689_comb[12:0];
  assign p1_add_80060_comb = p1_sign_ext_78690_comb[12:0] + p1_sign_ext_78630_comb[12:0];
  assign p1_add_80061_comb = p1_sign_ext_78586_comb[12:0] + p1_sign_ext_78587_comb[12:0];
  assign p1_add_80062_comb = p1_sign_ext_78588_comb[12:0] + p1_sign_ext_78589_comb[12:0];
  assign p1_add_80063_comb = p1_sign_ext_78631_comb[12:0] + p1_sign_ext_78695_comb[12:0];
  assign p1_add_80064_comb = p1_sign_ext_78696_comb[12:0] + p1_sign_ext_78632_comb[12:0];
  assign p1_add_80065_comb = p1_sign_ext_78594_comb[12:0] + p1_sign_ext_78595_comb[12:0];
  assign p1_add_80066_comb = p1_sign_ext_78596_comb[12:0] + p1_sign_ext_78597_comb[12:0];
  assign p1_add_80067_comb = p1_sign_ext_78633_comb[12:0] + p1_sign_ext_78701_comb[12:0];
  assign p1_add_80068_comb = p1_sign_ext_78702_comb[12:0] + p1_sign_ext_78634_comb[12:0];
  assign p1_add_80069_comb = p1_sign_ext_78602_comb[12:0] + p1_sign_ext_78603_comb[12:0];
  assign p1_add_80070_comb = p1_sign_ext_78604_comb[12:0] + p1_sign_ext_78605_comb[12:0];
  assign p1_add_80071_comb = p1_sign_ext_78635_comb[12:0] + p1_sign_ext_78707_comb[12:0];
  assign p1_add_80072_comb = p1_sign_ext_78708_comb[12:0] + p1_sign_ext_78636_comb[12:0];
  assign p1_add_80073_comb = p1_sign_ext_78610_comb[12:0] + p1_sign_ext_78611_comb[12:0];
  assign p1_add_80074_comb = p1_sign_ext_78612_comb[12:0] + p1_sign_ext_78613_comb[12:0];
  assign p1_add_80075_comb = p1_sign_ext_78637_comb[12:0] + p1_sign_ext_78713_comb[12:0];
  assign p1_add_80076_comb = p1_sign_ext_78714_comb[12:0] + p1_sign_ext_78638_comb[12:0];
  assign p1_add_80077_comb = p1_sign_ext_78618_comb[12:0] + p1_sign_ext_78619_comb[12:0];
  assign p1_add_80078_comb = p1_sign_ext_78620_comb[12:0] + p1_sign_ext_78621_comb[12:0];
  assign p1_add_80079_comb = p1_sign_ext_78639_comb[12:0] + p1_sign_ext_78719_comb[12:0];
  assign p1_add_80112_comb = p1_smul_79696_comb + p1_smul_79186_comb[19:1];
  assign p1_add_80114_comb = p1_smul_79187_comb[19:1] + p1_smul_79699_comb;
  assign p1_add_80116_comb = p1_smul_79700_comb + p1_smul_79192_comb[19:1];
  assign p1_add_80118_comb = p1_smul_79193_comb[19:1] + p1_smul_79703_comb;
  assign p1_add_80120_comb = p1_smul_79704_comb + p1_smul_79198_comb[19:1];
  assign p1_add_80122_comb = p1_smul_79199_comb[19:1] + p1_smul_79707_comb;
  assign p1_add_80124_comb = p1_smul_79708_comb + p1_smul_79204_comb[19:1];
  assign p1_add_80126_comb = p1_smul_79205_comb[19:1] + p1_smul_79711_comb;
  assign p1_add_80128_comb = p1_smul_79712_comb + p1_smul_79210_comb[19:1];
  assign p1_add_80130_comb = p1_smul_79211_comb[19:1] + p1_smul_79715_comb;
  assign p1_add_80132_comb = p1_smul_79716_comb + p1_smul_79216_comb[19:1];
  assign p1_add_80134_comb = p1_smul_79217_comb[19:1] + p1_smul_79719_comb;
  assign p1_add_80136_comb = p1_smul_79720_comb + p1_smul_79222_comb[19:1];
  assign p1_add_80138_comb = p1_smul_79223_comb[19:1] + p1_smul_79723_comb;
  assign p1_add_80140_comb = p1_smul_79724_comb + p1_smul_79228_comb[19:1];
  assign p1_add_80142_comb = p1_smul_79229_comb[19:1] + p1_smul_79727_comb;
  assign p1_add_80144_comb = p1_smul_79728_comb + p1_smul_79234_comb[19:1];
  assign p1_add_80146_comb = p1_smul_79235_comb[19:1] + p1_smul_79731_comb;
  assign p1_add_80148_comb = p1_smul_79732_comb + p1_smul_79240_comb[19:1];
  assign p1_add_80150_comb = p1_smul_79241_comb[19:1] + p1_smul_79735_comb;
  assign p1_add_80152_comb = p1_smul_79736_comb + p1_smul_79246_comb[19:1];
  assign p1_add_80154_comb = p1_smul_79247_comb[19:1] + p1_smul_79739_comb;
  assign p1_add_80156_comb = p1_smul_79740_comb + p1_smul_79252_comb[19:1];
  assign p1_add_80158_comb = p1_smul_79253_comb[19:1] + p1_smul_79743_comb;
  assign p1_add_80160_comb = p1_smul_79744_comb + p1_smul_79258_comb[19:1];
  assign p1_add_80162_comb = p1_smul_79259_comb[19:1] + p1_smul_79747_comb;
  assign p1_add_80164_comb = p1_smul_79748_comb + p1_smul_79264_comb[19:1];
  assign p1_add_80166_comb = p1_smul_79265_comb[19:1] + p1_smul_79751_comb;
  assign p1_add_80168_comb = p1_smul_79752_comb + p1_smul_79270_comb[19:1];
  assign p1_add_80170_comb = p1_smul_79271_comb[19:1] + p1_smul_79755_comb;
  assign p1_add_80172_comb = p1_smul_79756_comb + p1_smul_79276_comb[19:1];
  assign p1_add_80174_comb = p1_smul_79277_comb[19:1] + p1_smul_79759_comb;
  assign p1_concat_80176_comb = {p1_add_79760_comb, p1_smul_78896_comb[0]};
  assign p1_concat_80177_comb = {p1_add_79762_comb, p1_smul_78898_comb[0]};
  assign p1_concat_80178_comb = {p1_add_79764_comb, p1_smul_78901_comb[0]};
  assign p1_concat_80179_comb = {p1_add_79766_comb, p1_smul_78903_comb[0]};
  assign p1_concat_80180_comb = {p1_add_79768_comb, p1_smul_78904_comb[0]};
  assign p1_concat_80181_comb = {p1_add_79770_comb, p1_smul_78906_comb[0]};
  assign p1_concat_80182_comb = {p1_add_79772_comb, p1_smul_78909_comb[0]};
  assign p1_concat_80183_comb = {p1_add_79774_comb, p1_smul_78911_comb[0]};
  assign p1_concat_80184_comb = {p1_add_79776_comb, p1_smul_78912_comb[0]};
  assign p1_concat_80185_comb = {p1_add_79778_comb, p1_smul_78914_comb[0]};
  assign p1_concat_80186_comb = {p1_add_79780_comb, p1_smul_78917_comb[0]};
  assign p1_concat_80187_comb = {p1_add_79782_comb, p1_smul_78919_comb[0]};
  assign p1_concat_80188_comb = {p1_add_79784_comb, p1_smul_78920_comb[0]};
  assign p1_concat_80189_comb = {p1_add_79786_comb, p1_smul_78922_comb[0]};
  assign p1_concat_80190_comb = {p1_add_79788_comb, p1_smul_78925_comb[0]};
  assign p1_concat_80191_comb = {p1_add_79790_comb, p1_smul_78927_comb[0]};
  assign p1_concat_80192_comb = {p1_add_79792_comb, p1_smul_78928_comb[0]};
  assign p1_concat_80193_comb = {p1_add_79794_comb, p1_smul_78930_comb[0]};
  assign p1_concat_80194_comb = {p1_add_79796_comb, p1_smul_78933_comb[0]};
  assign p1_concat_80195_comb = {p1_add_79798_comb, p1_smul_78935_comb[0]};
  assign p1_concat_80196_comb = {p1_add_79800_comb, p1_smul_78936_comb[0]};
  assign p1_concat_80197_comb = {p1_add_79802_comb, p1_smul_78938_comb[0]};
  assign p1_concat_80198_comb = {p1_add_79804_comb, p1_smul_78941_comb[0]};
  assign p1_concat_80199_comb = {p1_add_79806_comb, p1_smul_78943_comb[0]};
  assign p1_concat_80200_comb = {p1_add_79808_comb, p1_smul_78944_comb[0]};
  assign p1_concat_80201_comb = {p1_add_79810_comb, p1_smul_78946_comb[0]};
  assign p1_concat_80202_comb = {p1_add_79812_comb, p1_smul_78949_comb[0]};
  assign p1_concat_80203_comb = {p1_add_79814_comb, p1_smul_78951_comb[0]};
  assign p1_concat_80204_comb = {p1_add_79816_comb, p1_smul_78952_comb[0]};
  assign p1_concat_80205_comb = {p1_add_79818_comb, p1_smul_78954_comb[0]};
  assign p1_concat_80206_comb = {p1_add_79820_comb, p1_smul_78957_comb[0]};
  assign p1_concat_80207_comb = {p1_add_79822_comb, p1_smul_78959_comb[0]};
  assign p1_add_80208_comb = p1_smul_79824_comb + p1_smul_79825_comb;
  assign p1_add_80209_comb = p1_smul_79826_comb + p1_smul_79827_comb;
  assign p1_add_80210_comb = p1_smul_79828_comb + p1_smul_79829_comb;
  assign p1_add_80211_comb = p1_smul_79830_comb + p1_smul_79831_comb;
  assign p1_add_80212_comb = p1_smul_79832_comb + p1_smul_79833_comb;
  assign p1_add_80213_comb = p1_smul_79834_comb + p1_smul_79835_comb;
  assign p1_add_80214_comb = p1_smul_79836_comb + p1_smul_79837_comb;
  assign p1_add_80215_comb = p1_smul_79838_comb + p1_smul_79839_comb;
  assign p1_add_80216_comb = p1_smul_79840_comb + p1_smul_79841_comb;
  assign p1_add_80217_comb = p1_smul_79842_comb + p1_smul_79843_comb;
  assign p1_add_80218_comb = p1_smul_79844_comb + p1_smul_79845_comb;
  assign p1_add_80219_comb = p1_smul_79846_comb + p1_smul_79847_comb;
  assign p1_add_80220_comb = p1_smul_79848_comb + p1_smul_79849_comb;
  assign p1_add_80221_comb = p1_smul_79850_comb + p1_smul_79851_comb;
  assign p1_add_80222_comb = p1_smul_79852_comb + p1_smul_79853_comb;
  assign p1_add_80223_comb = p1_smul_79854_comb + p1_smul_79855_comb;
  assign p1_add_80224_comb = p1_smul_79856_comb + p1_smul_79857_comb;
  assign p1_add_80225_comb = p1_smul_79858_comb + p1_smul_79859_comb;
  assign p1_add_80226_comb = p1_smul_79860_comb + p1_smul_79861_comb;
  assign p1_add_80227_comb = p1_smul_79862_comb + p1_smul_79863_comb;
  assign p1_add_80228_comb = p1_smul_79864_comb + p1_smul_79865_comb;
  assign p1_add_80229_comb = p1_smul_79866_comb + p1_smul_79867_comb;
  assign p1_add_80230_comb = p1_smul_79868_comb + p1_smul_79869_comb;
  assign p1_add_80231_comb = p1_smul_79870_comb + p1_smul_79871_comb;
  assign p1_add_80232_comb = p1_smul_79872_comb + p1_smul_79873_comb;
  assign p1_add_80233_comb = p1_smul_79874_comb + p1_smul_79875_comb;
  assign p1_add_80234_comb = p1_smul_79876_comb + p1_smul_79877_comb;
  assign p1_add_80235_comb = p1_smul_79878_comb + p1_smul_79879_comb;
  assign p1_add_80236_comb = p1_smul_79880_comb + p1_smul_79881_comb;
  assign p1_add_80237_comb = p1_smul_79882_comb + p1_smul_79883_comb;
  assign p1_add_80238_comb = p1_smul_79884_comb + p1_smul_79885_comb;
  assign p1_add_80239_comb = p1_smul_79886_comb + p1_smul_79887_comb;
  assign p1_concat_80240_comb = {p1_add_79888_comb, p1_smul_78962_comb[0]};
  assign p1_concat_80241_comb = {p1_add_79890_comb, p1_smul_78964_comb[0]};
  assign p1_concat_80242_comb = {p1_add_79892_comb, p1_smul_78965_comb[0]};
  assign p1_concat_80243_comb = {p1_add_79894_comb, p1_smul_78967_comb[0]};
  assign p1_concat_80244_comb = {p1_add_79896_comb, p1_smul_78972_comb[0]};
  assign p1_concat_80245_comb = {p1_add_79898_comb, p1_smul_78974_comb[0]};
  assign p1_concat_80246_comb = {p1_add_79900_comb, p1_smul_78975_comb[0]};
  assign p1_concat_80247_comb = {p1_add_79902_comb, p1_smul_78977_comb[0]};
  assign p1_concat_80248_comb = {p1_add_79904_comb, p1_smul_78982_comb[0]};
  assign p1_concat_80249_comb = {p1_add_79906_comb, p1_smul_78984_comb[0]};
  assign p1_concat_80250_comb = {p1_add_79908_comb, p1_smul_78985_comb[0]};
  assign p1_concat_80251_comb = {p1_add_79910_comb, p1_smul_78987_comb[0]};
  assign p1_concat_80252_comb = {p1_add_79912_comb, p1_smul_78992_comb[0]};
  assign p1_concat_80253_comb = {p1_add_79914_comb, p1_smul_78994_comb[0]};
  assign p1_concat_80254_comb = {p1_add_79916_comb, p1_smul_78995_comb[0]};
  assign p1_concat_80255_comb = {p1_add_79918_comb, p1_smul_78997_comb[0]};
  assign p1_concat_80256_comb = {p1_add_79920_comb, p1_smul_79002_comb[0]};
  assign p1_concat_80257_comb = {p1_add_79922_comb, p1_smul_79004_comb[0]};
  assign p1_concat_80258_comb = {p1_add_79924_comb, p1_smul_79005_comb[0]};
  assign p1_concat_80259_comb = {p1_add_79926_comb, p1_smul_79007_comb[0]};
  assign p1_concat_80260_comb = {p1_add_79928_comb, p1_smul_79012_comb[0]};
  assign p1_concat_80261_comb = {p1_add_79930_comb, p1_smul_79014_comb[0]};
  assign p1_concat_80262_comb = {p1_add_79932_comb, p1_smul_79015_comb[0]};
  assign p1_concat_80263_comb = {p1_add_79934_comb, p1_smul_79017_comb[0]};
  assign p1_concat_80264_comb = {p1_add_79936_comb, p1_smul_79022_comb[0]};
  assign p1_concat_80265_comb = {p1_add_79938_comb, p1_smul_79024_comb[0]};
  assign p1_concat_80266_comb = {p1_add_79940_comb, p1_smul_79025_comb[0]};
  assign p1_concat_80267_comb = {p1_add_79942_comb, p1_smul_79027_comb[0]};
  assign p1_concat_80268_comb = {p1_add_79944_comb, p1_smul_79032_comb[0]};
  assign p1_concat_80269_comb = {p1_add_79946_comb, p1_smul_79034_comb[0]};
  assign p1_concat_80270_comb = {p1_add_79948_comb, p1_smul_79035_comb[0]};
  assign p1_concat_80271_comb = {p1_add_79950_comb, p1_smul_79037_comb[0]};
  assign p1_add_80272_comb = p1_smul_79472_comb[19:1] + p1_smul_79953_comb;
  assign p1_add_80274_comb = p1_smul_79475_comb[19:1] + p1_smul_79955_comb;
  assign p1_add_80276_comb = p1_smul_79956_comb + p1_smul_79478_comb[19:1];
  assign p1_add_80278_comb = p1_smul_79958_comb + p1_smul_79481_comb[19:1];
  assign p1_add_80280_comb = p1_smul_79482_comb[19:1] + p1_smul_79961_comb;
  assign p1_add_80282_comb = p1_smul_79485_comb[19:1] + p1_smul_79963_comb;
  assign p1_add_80284_comb = p1_smul_79964_comb + p1_smul_79488_comb[19:1];
  assign p1_add_80286_comb = p1_smul_79966_comb + p1_smul_79491_comb[19:1];
  assign p1_add_80288_comb = p1_smul_79492_comb[19:1] + p1_smul_79969_comb;
  assign p1_add_80290_comb = p1_smul_79495_comb[19:1] + p1_smul_79971_comb;
  assign p1_add_80292_comb = p1_smul_79972_comb + p1_smul_79498_comb[19:1];
  assign p1_add_80294_comb = p1_smul_79974_comb + p1_smul_79501_comb[19:1];
  assign p1_add_80296_comb = p1_smul_79502_comb[19:1] + p1_smul_79977_comb;
  assign p1_add_80298_comb = p1_smul_79505_comb[19:1] + p1_smul_79979_comb;
  assign p1_add_80300_comb = p1_smul_79980_comb + p1_smul_79508_comb[19:1];
  assign p1_add_80302_comb = p1_smul_79982_comb + p1_smul_79511_comb[19:1];
  assign p1_add_80304_comb = p1_smul_79512_comb[19:1] + p1_smul_79985_comb;
  assign p1_add_80306_comb = p1_smul_79515_comb[19:1] + p1_smul_79987_comb;
  assign p1_add_80308_comb = p1_smul_79988_comb + p1_smul_79518_comb[19:1];
  assign p1_add_80310_comb = p1_smul_79990_comb + p1_smul_79521_comb[19:1];
  assign p1_add_80312_comb = p1_smul_79522_comb[19:1] + p1_smul_79993_comb;
  assign p1_add_80314_comb = p1_smul_79525_comb[19:1] + p1_smul_79995_comb;
  assign p1_add_80316_comb = p1_smul_79996_comb + p1_smul_79528_comb[19:1];
  assign p1_add_80318_comb = p1_smul_79998_comb + p1_smul_79531_comb[19:1];
  assign p1_add_80320_comb = p1_smul_79532_comb[19:1] + p1_smul_80001_comb;
  assign p1_add_80322_comb = p1_smul_79535_comb[19:1] + p1_smul_80003_comb;
  assign p1_add_80324_comb = p1_smul_80004_comb + p1_smul_79538_comb[19:1];
  assign p1_add_80326_comb = p1_smul_80006_comb + p1_smul_79541_comb[19:1];
  assign p1_add_80328_comb = p1_smul_79542_comb[19:1] + p1_smul_80009_comb;
  assign p1_add_80330_comb = p1_smul_79545_comb[19:1] + p1_smul_80011_comb;
  assign p1_add_80332_comb = p1_smul_80012_comb + p1_smul_79548_comb[19:1];
  assign p1_add_80334_comb = p1_smul_80014_comb + p1_smul_79551_comb[19:1];
  assign p1_add_80400_comb = {{4{p1_bit_slice_79664_comb[19]}}, p1_bit_slice_79664_comb} + {{4{p1_add_79665_comb[19]}}, p1_add_79665_comb};
  assign p1_add_80402_comb = {{4{p1_add_79666_comb[19]}}, p1_add_79666_comb} + {{4{p1_bit_slice_79667_comb[19]}}, p1_bit_slice_79667_comb};
  assign p1_add_80404_comb = {{4{p1_bit_slice_79668_comb[19]}}, p1_bit_slice_79668_comb} + {{4{p1_add_79669_comb[19]}}, p1_add_79669_comb};
  assign p1_add_80406_comb = {{4{p1_add_79670_comb[19]}}, p1_add_79670_comb} + {{4{p1_bit_slice_79671_comb[19]}}, p1_bit_slice_79671_comb};
  assign p1_add_80408_comb = {{4{p1_bit_slice_79672_comb[19]}}, p1_bit_slice_79672_comb} + {{4{p1_add_79673_comb[19]}}, p1_add_79673_comb};
  assign p1_add_80410_comb = {{4{p1_add_79674_comb[19]}}, p1_add_79674_comb} + {{4{p1_bit_slice_79675_comb[19]}}, p1_bit_slice_79675_comb};
  assign p1_add_80412_comb = {{4{p1_bit_slice_79676_comb[19]}}, p1_bit_slice_79676_comb} + {{4{p1_add_79677_comb[19]}}, p1_add_79677_comb};
  assign p1_add_80414_comb = {{4{p1_add_79678_comb[19]}}, p1_add_79678_comb} + {{4{p1_bit_slice_79679_comb[19]}}, p1_bit_slice_79679_comb};
  assign p1_add_80416_comb = {{4{p1_bit_slice_79680_comb[19]}}, p1_bit_slice_79680_comb} + {{4{p1_add_79681_comb[19]}}, p1_add_79681_comb};
  assign p1_add_80418_comb = {{4{p1_add_79682_comb[19]}}, p1_add_79682_comb} + {{4{p1_bit_slice_79683_comb[19]}}, p1_bit_slice_79683_comb};
  assign p1_add_80420_comb = {{4{p1_bit_slice_79684_comb[19]}}, p1_bit_slice_79684_comb} + {{4{p1_add_79685_comb[19]}}, p1_add_79685_comb};
  assign p1_add_80422_comb = {{4{p1_add_79686_comb[19]}}, p1_add_79686_comb} + {{4{p1_bit_slice_79687_comb[19]}}, p1_bit_slice_79687_comb};
  assign p1_add_80424_comb = {{4{p1_bit_slice_79688_comb[19]}}, p1_bit_slice_79688_comb} + {{4{p1_add_79689_comb[19]}}, p1_add_79689_comb};
  assign p1_add_80426_comb = {{4{p1_add_79690_comb[19]}}, p1_add_79690_comb} + {{4{p1_bit_slice_79691_comb[19]}}, p1_bit_slice_79691_comb};
  assign p1_add_80428_comb = {{4{p1_bit_slice_79692_comb[19]}}, p1_bit_slice_79692_comb} + {{4{p1_add_79693_comb[19]}}, p1_add_79693_comb};
  assign p1_add_80430_comb = {{4{p1_add_79694_comb[19]}}, p1_add_79694_comb} + {{4{p1_bit_slice_79695_comb[19]}}, p1_bit_slice_79695_comb};
  assign p1_concat_80432_comb = {p1_add_80112_comb, p1_smul_79186_comb[0]};
  assign p1_concat_80433_comb = {p1_add_80114_comb, p1_smul_79187_comb[0]};
  assign p1_concat_80434_comb = {p1_add_80116_comb, p1_smul_79192_comb[0]};
  assign p1_concat_80435_comb = {p1_add_80118_comb, p1_smul_79193_comb[0]};
  assign p1_concat_80436_comb = {p1_add_80120_comb, p1_smul_79198_comb[0]};
  assign p1_concat_80437_comb = {p1_add_80122_comb, p1_smul_79199_comb[0]};
  assign p1_concat_80438_comb = {p1_add_80124_comb, p1_smul_79204_comb[0]};
  assign p1_concat_80439_comb = {p1_add_80126_comb, p1_smul_79205_comb[0]};
  assign p1_concat_80440_comb = {p1_add_80128_comb, p1_smul_79210_comb[0]};
  assign p1_concat_80441_comb = {p1_add_80130_comb, p1_smul_79211_comb[0]};
  assign p1_concat_80442_comb = {p1_add_80132_comb, p1_smul_79216_comb[0]};
  assign p1_concat_80443_comb = {p1_add_80134_comb, p1_smul_79217_comb[0]};
  assign p1_concat_80444_comb = {p1_add_80136_comb, p1_smul_79222_comb[0]};
  assign p1_concat_80445_comb = {p1_add_80138_comb, p1_smul_79223_comb[0]};
  assign p1_concat_80446_comb = {p1_add_80140_comb, p1_smul_79228_comb[0]};
  assign p1_concat_80447_comb = {p1_add_80142_comb, p1_smul_79229_comb[0]};
  assign p1_concat_80448_comb = {p1_add_80144_comb, p1_smul_79234_comb[0]};
  assign p1_concat_80449_comb = {p1_add_80146_comb, p1_smul_79235_comb[0]};
  assign p1_concat_80450_comb = {p1_add_80148_comb, p1_smul_79240_comb[0]};
  assign p1_concat_80451_comb = {p1_add_80150_comb, p1_smul_79241_comb[0]};
  assign p1_concat_80452_comb = {p1_add_80152_comb, p1_smul_79246_comb[0]};
  assign p1_concat_80453_comb = {p1_add_80154_comb, p1_smul_79247_comb[0]};
  assign p1_concat_80454_comb = {p1_add_80156_comb, p1_smul_79252_comb[0]};
  assign p1_concat_80455_comb = {p1_add_80158_comb, p1_smul_79253_comb[0]};
  assign p1_concat_80456_comb = {p1_add_80160_comb, p1_smul_79258_comb[0]};
  assign p1_concat_80457_comb = {p1_add_80162_comb, p1_smul_79259_comb[0]};
  assign p1_concat_80458_comb = {p1_add_80164_comb, p1_smul_79264_comb[0]};
  assign p1_concat_80459_comb = {p1_add_80166_comb, p1_smul_79265_comb[0]};
  assign p1_concat_80460_comb = {p1_add_80168_comb, p1_smul_79270_comb[0]};
  assign p1_concat_80461_comb = {p1_add_80170_comb, p1_smul_79271_comb[0]};
  assign p1_concat_80462_comb = {p1_add_80172_comb, p1_smul_79276_comb[0]};
  assign p1_concat_80463_comb = {p1_add_80174_comb, p1_smul_79277_comb[0]};
  assign p1_sum__1572_comb = {{4{p1_concat_80176_comb[20]}}, p1_concat_80176_comb};
  assign p1_sum__1573_comb = {{4{p1_concat_80177_comb[20]}}, p1_concat_80177_comb};
  assign p1_sum__1574_comb = {{4{p1_concat_80178_comb[20]}}, p1_concat_80178_comb};
  assign p1_sum__1575_comb = {{4{p1_concat_80179_comb[20]}}, p1_concat_80179_comb};
  assign p1_sum__1544_comb = {{4{p1_concat_80180_comb[20]}}, p1_concat_80180_comb};
  assign p1_sum__1545_comb = {{4{p1_concat_80181_comb[20]}}, p1_concat_80181_comb};
  assign p1_sum__1546_comb = {{4{p1_concat_80182_comb[20]}}, p1_concat_80182_comb};
  assign p1_sum__1547_comb = {{4{p1_concat_80183_comb[20]}}, p1_concat_80183_comb};
  assign p1_sum__1516_comb = {{4{p1_concat_80184_comb[20]}}, p1_concat_80184_comb};
  assign p1_sum__1517_comb = {{4{p1_concat_80185_comb[20]}}, p1_concat_80185_comb};
  assign p1_sum__1518_comb = {{4{p1_concat_80186_comb[20]}}, p1_concat_80186_comb};
  assign p1_sum__1519_comb = {{4{p1_concat_80187_comb[20]}}, p1_concat_80187_comb};
  assign p1_sum__1488_comb = {{4{p1_concat_80188_comb[20]}}, p1_concat_80188_comb};
  assign p1_sum__1489_comb = {{4{p1_concat_80189_comb[20]}}, p1_concat_80189_comb};
  assign p1_sum__1490_comb = {{4{p1_concat_80190_comb[20]}}, p1_concat_80190_comb};
  assign p1_sum__1491_comb = {{4{p1_concat_80191_comb[20]}}, p1_concat_80191_comb};
  assign p1_sum__1460_comb = {{4{p1_concat_80192_comb[20]}}, p1_concat_80192_comb};
  assign p1_sum__1461_comb = {{4{p1_concat_80193_comb[20]}}, p1_concat_80193_comb};
  assign p1_sum__1462_comb = {{4{p1_concat_80194_comb[20]}}, p1_concat_80194_comb};
  assign p1_sum__1463_comb = {{4{p1_concat_80195_comb[20]}}, p1_concat_80195_comb};
  assign p1_sum__1432_comb = {{4{p1_concat_80196_comb[20]}}, p1_concat_80196_comb};
  assign p1_sum__1433_comb = {{4{p1_concat_80197_comb[20]}}, p1_concat_80197_comb};
  assign p1_sum__1434_comb = {{4{p1_concat_80198_comb[20]}}, p1_concat_80198_comb};
  assign p1_sum__1435_comb = {{4{p1_concat_80199_comb[20]}}, p1_concat_80199_comb};
  assign p1_sum__1404_comb = {{4{p1_concat_80200_comb[20]}}, p1_concat_80200_comb};
  assign p1_sum__1405_comb = {{4{p1_concat_80201_comb[20]}}, p1_concat_80201_comb};
  assign p1_sum__1406_comb = {{4{p1_concat_80202_comb[20]}}, p1_concat_80202_comb};
  assign p1_sum__1407_comb = {{4{p1_concat_80203_comb[20]}}, p1_concat_80203_comb};
  assign p1_sum__1376_comb = {{4{p1_concat_80204_comb[20]}}, p1_concat_80204_comb};
  assign p1_sum__1377_comb = {{4{p1_concat_80205_comb[20]}}, p1_concat_80205_comb};
  assign p1_sum__1378_comb = {{4{p1_concat_80206_comb[20]}}, p1_concat_80206_comb};
  assign p1_sum__1379_comb = {{4{p1_concat_80207_comb[20]}}, p1_concat_80207_comb};
  assign p1_sum__1568_comb = {{4{p1_add_80208_comb[20]}}, p1_add_80208_comb};
  assign p1_sum__1569_comb = {{4{p1_add_80209_comb[20]}}, p1_add_80209_comb};
  assign p1_sum__1570_comb = {{4{p1_add_80210_comb[20]}}, p1_add_80210_comb};
  assign p1_sum__1571_comb = {{4{p1_add_80211_comb[20]}}, p1_add_80211_comb};
  assign p1_sum__1540_comb = {{4{p1_add_80212_comb[20]}}, p1_add_80212_comb};
  assign p1_sum__1541_comb = {{4{p1_add_80213_comb[20]}}, p1_add_80213_comb};
  assign p1_sum__1542_comb = {{4{p1_add_80214_comb[20]}}, p1_add_80214_comb};
  assign p1_sum__1543_comb = {{4{p1_add_80215_comb[20]}}, p1_add_80215_comb};
  assign p1_sum__1512_comb = {{4{p1_add_80216_comb[20]}}, p1_add_80216_comb};
  assign p1_sum__1513_comb = {{4{p1_add_80217_comb[20]}}, p1_add_80217_comb};
  assign p1_sum__1514_comb = {{4{p1_add_80218_comb[20]}}, p1_add_80218_comb};
  assign p1_sum__1515_comb = {{4{p1_add_80219_comb[20]}}, p1_add_80219_comb};
  assign p1_sum__1484_comb = {{4{p1_add_80220_comb[20]}}, p1_add_80220_comb};
  assign p1_sum__1485_comb = {{4{p1_add_80221_comb[20]}}, p1_add_80221_comb};
  assign p1_sum__1486_comb = {{4{p1_add_80222_comb[20]}}, p1_add_80222_comb};
  assign p1_sum__1487_comb = {{4{p1_add_80223_comb[20]}}, p1_add_80223_comb};
  assign p1_sum__1456_comb = {{4{p1_add_80224_comb[20]}}, p1_add_80224_comb};
  assign p1_sum__1457_comb = {{4{p1_add_80225_comb[20]}}, p1_add_80225_comb};
  assign p1_sum__1458_comb = {{4{p1_add_80226_comb[20]}}, p1_add_80226_comb};
  assign p1_sum__1459_comb = {{4{p1_add_80227_comb[20]}}, p1_add_80227_comb};
  assign p1_sum__1428_comb = {{4{p1_add_80228_comb[20]}}, p1_add_80228_comb};
  assign p1_sum__1429_comb = {{4{p1_add_80229_comb[20]}}, p1_add_80229_comb};
  assign p1_sum__1430_comb = {{4{p1_add_80230_comb[20]}}, p1_add_80230_comb};
  assign p1_sum__1431_comb = {{4{p1_add_80231_comb[20]}}, p1_add_80231_comb};
  assign p1_sum__1400_comb = {{4{p1_add_80232_comb[20]}}, p1_add_80232_comb};
  assign p1_sum__1401_comb = {{4{p1_add_80233_comb[20]}}, p1_add_80233_comb};
  assign p1_sum__1402_comb = {{4{p1_add_80234_comb[20]}}, p1_add_80234_comb};
  assign p1_sum__1403_comb = {{4{p1_add_80235_comb[20]}}, p1_add_80235_comb};
  assign p1_sum__1372_comb = {{4{p1_add_80236_comb[20]}}, p1_add_80236_comb};
  assign p1_sum__1373_comb = {{4{p1_add_80237_comb[20]}}, p1_add_80237_comb};
  assign p1_sum__1374_comb = {{4{p1_add_80238_comb[20]}}, p1_add_80238_comb};
  assign p1_sum__1375_comb = {{4{p1_add_80239_comb[20]}}, p1_add_80239_comb};
  assign p1_sum__1564_comb = {{4{p1_concat_80240_comb[20]}}, p1_concat_80240_comb};
  assign p1_sum__1565_comb = {{4{p1_concat_80241_comb[20]}}, p1_concat_80241_comb};
  assign p1_sum__1566_comb = {{4{p1_concat_80242_comb[20]}}, p1_concat_80242_comb};
  assign p1_sum__1567_comb = {{4{p1_concat_80243_comb[20]}}, p1_concat_80243_comb};
  assign p1_sum__1536_comb = {{4{p1_concat_80244_comb[20]}}, p1_concat_80244_comb};
  assign p1_sum__1537_comb = {{4{p1_concat_80245_comb[20]}}, p1_concat_80245_comb};
  assign p1_sum__1538_comb = {{4{p1_concat_80246_comb[20]}}, p1_concat_80246_comb};
  assign p1_sum__1539_comb = {{4{p1_concat_80247_comb[20]}}, p1_concat_80247_comb};
  assign p1_sum__1508_comb = {{4{p1_concat_80248_comb[20]}}, p1_concat_80248_comb};
  assign p1_sum__1509_comb = {{4{p1_concat_80249_comb[20]}}, p1_concat_80249_comb};
  assign p1_sum__1510_comb = {{4{p1_concat_80250_comb[20]}}, p1_concat_80250_comb};
  assign p1_sum__1511_comb = {{4{p1_concat_80251_comb[20]}}, p1_concat_80251_comb};
  assign p1_sum__1480_comb = {{4{p1_concat_80252_comb[20]}}, p1_concat_80252_comb};
  assign p1_sum__1481_comb = {{4{p1_concat_80253_comb[20]}}, p1_concat_80253_comb};
  assign p1_sum__1482_comb = {{4{p1_concat_80254_comb[20]}}, p1_concat_80254_comb};
  assign p1_sum__1483_comb = {{4{p1_concat_80255_comb[20]}}, p1_concat_80255_comb};
  assign p1_sum__1452_comb = {{4{p1_concat_80256_comb[20]}}, p1_concat_80256_comb};
  assign p1_sum__1453_comb = {{4{p1_concat_80257_comb[20]}}, p1_concat_80257_comb};
  assign p1_sum__1454_comb = {{4{p1_concat_80258_comb[20]}}, p1_concat_80258_comb};
  assign p1_sum__1455_comb = {{4{p1_concat_80259_comb[20]}}, p1_concat_80259_comb};
  assign p1_sum__1424_comb = {{4{p1_concat_80260_comb[20]}}, p1_concat_80260_comb};
  assign p1_sum__1425_comb = {{4{p1_concat_80261_comb[20]}}, p1_concat_80261_comb};
  assign p1_sum__1426_comb = {{4{p1_concat_80262_comb[20]}}, p1_concat_80262_comb};
  assign p1_sum__1427_comb = {{4{p1_concat_80263_comb[20]}}, p1_concat_80263_comb};
  assign p1_sum__1396_comb = {{4{p1_concat_80264_comb[20]}}, p1_concat_80264_comb};
  assign p1_sum__1397_comb = {{4{p1_concat_80265_comb[20]}}, p1_concat_80265_comb};
  assign p1_sum__1398_comb = {{4{p1_concat_80266_comb[20]}}, p1_concat_80266_comb};
  assign p1_sum__1399_comb = {{4{p1_concat_80267_comb[20]}}, p1_concat_80267_comb};
  assign p1_sum__1368_comb = {{4{p1_concat_80268_comb[20]}}, p1_concat_80268_comb};
  assign p1_sum__1369_comb = {{4{p1_concat_80269_comb[20]}}, p1_concat_80269_comb};
  assign p1_sum__1370_comb = {{4{p1_concat_80270_comb[20]}}, p1_concat_80270_comb};
  assign p1_sum__1371_comb = {{4{p1_concat_80271_comb[20]}}, p1_concat_80271_comb};
  assign p1_concat_80560_comb = {p1_add_80272_comb, p1_smul_79472_comb[0]};
  assign p1_concat_80561_comb = {p1_add_80274_comb, p1_smul_79475_comb[0]};
  assign p1_concat_80562_comb = {p1_add_80276_comb, p1_smul_79478_comb[0]};
  assign p1_concat_80563_comb = {p1_add_80278_comb, p1_smul_79481_comb[0]};
  assign p1_concat_80564_comb = {p1_add_80280_comb, p1_smul_79482_comb[0]};
  assign p1_concat_80565_comb = {p1_add_80282_comb, p1_smul_79485_comb[0]};
  assign p1_concat_80566_comb = {p1_add_80284_comb, p1_smul_79488_comb[0]};
  assign p1_concat_80567_comb = {p1_add_80286_comb, p1_smul_79491_comb[0]};
  assign p1_concat_80568_comb = {p1_add_80288_comb, p1_smul_79492_comb[0]};
  assign p1_concat_80569_comb = {p1_add_80290_comb, p1_smul_79495_comb[0]};
  assign p1_concat_80570_comb = {p1_add_80292_comb, p1_smul_79498_comb[0]};
  assign p1_concat_80571_comb = {p1_add_80294_comb, p1_smul_79501_comb[0]};
  assign p1_concat_80572_comb = {p1_add_80296_comb, p1_smul_79502_comb[0]};
  assign p1_concat_80573_comb = {p1_add_80298_comb, p1_smul_79505_comb[0]};
  assign p1_concat_80574_comb = {p1_add_80300_comb, p1_smul_79508_comb[0]};
  assign p1_concat_80575_comb = {p1_add_80302_comb, p1_smul_79511_comb[0]};
  assign p1_concat_80576_comb = {p1_add_80304_comb, p1_smul_79512_comb[0]};
  assign p1_concat_80577_comb = {p1_add_80306_comb, p1_smul_79515_comb[0]};
  assign p1_concat_80578_comb = {p1_add_80308_comb, p1_smul_79518_comb[0]};
  assign p1_concat_80579_comb = {p1_add_80310_comb, p1_smul_79521_comb[0]};
  assign p1_concat_80580_comb = {p1_add_80312_comb, p1_smul_79522_comb[0]};
  assign p1_concat_80581_comb = {p1_add_80314_comb, p1_smul_79525_comb[0]};
  assign p1_concat_80582_comb = {p1_add_80316_comb, p1_smul_79528_comb[0]};
  assign p1_concat_80583_comb = {p1_add_80318_comb, p1_smul_79531_comb[0]};
  assign p1_concat_80584_comb = {p1_add_80320_comb, p1_smul_79532_comb[0]};
  assign p1_concat_80585_comb = {p1_add_80322_comb, p1_smul_79535_comb[0]};
  assign p1_concat_80586_comb = {p1_add_80324_comb, p1_smul_79538_comb[0]};
  assign p1_concat_80587_comb = {p1_add_80326_comb, p1_smul_79541_comb[0]};
  assign p1_concat_80588_comb = {p1_add_80328_comb, p1_smul_79542_comb[0]};
  assign p1_concat_80589_comb = {p1_add_80330_comb, p1_smul_79545_comb[0]};
  assign p1_concat_80590_comb = {p1_add_80332_comb, p1_smul_79548_comb[0]};
  assign p1_concat_80591_comb = {p1_add_80334_comb, p1_smul_79551_comb[0]};
  assign p1_add_80592_comb = {{4{p1_add_80016_comb[19]}}, p1_add_80016_comb} + {{4{p1_bit_slice_80017_comb[19]}}, p1_bit_slice_80017_comb};
  assign p1_add_80594_comb = {{4{p1_bit_slice_80018_comb[19]}}, p1_bit_slice_80018_comb} + {{4{p1_add_80019_comb[19]}}, p1_add_80019_comb};
  assign p1_add_80596_comb = {{4{p1_add_80020_comb[19]}}, p1_add_80020_comb} + {{4{p1_bit_slice_80021_comb[19]}}, p1_bit_slice_80021_comb};
  assign p1_add_80598_comb = {{4{p1_bit_slice_80022_comb[19]}}, p1_bit_slice_80022_comb} + {{4{p1_add_80023_comb[19]}}, p1_add_80023_comb};
  assign p1_add_80600_comb = {{4{p1_add_80024_comb[19]}}, p1_add_80024_comb} + {{4{p1_bit_slice_80025_comb[19]}}, p1_bit_slice_80025_comb};
  assign p1_add_80602_comb = {{4{p1_bit_slice_80026_comb[19]}}, p1_bit_slice_80026_comb} + {{4{p1_add_80027_comb[19]}}, p1_add_80027_comb};
  assign p1_add_80604_comb = {{4{p1_add_80028_comb[19]}}, p1_add_80028_comb} + {{4{p1_bit_slice_80029_comb[19]}}, p1_bit_slice_80029_comb};
  assign p1_add_80606_comb = {{4{p1_bit_slice_80030_comb[19]}}, p1_bit_slice_80030_comb} + {{4{p1_add_80031_comb[19]}}, p1_add_80031_comb};
  assign p1_add_80608_comb = {{4{p1_add_80032_comb[19]}}, p1_add_80032_comb} + {{4{p1_bit_slice_80033_comb[19]}}, p1_bit_slice_80033_comb};
  assign p1_add_80610_comb = {{4{p1_bit_slice_80034_comb[19]}}, p1_bit_slice_80034_comb} + {{4{p1_add_80035_comb[19]}}, p1_add_80035_comb};
  assign p1_add_80612_comb = {{4{p1_add_80036_comb[19]}}, p1_add_80036_comb} + {{4{p1_bit_slice_80037_comb[19]}}, p1_bit_slice_80037_comb};
  assign p1_add_80614_comb = {{4{p1_bit_slice_80038_comb[19]}}, p1_bit_slice_80038_comb} + {{4{p1_add_80039_comb[19]}}, p1_add_80039_comb};
  assign p1_add_80616_comb = {{4{p1_add_80040_comb[19]}}, p1_add_80040_comb} + {{4{p1_bit_slice_80041_comb[19]}}, p1_bit_slice_80041_comb};
  assign p1_add_80618_comb = {{4{p1_bit_slice_80042_comb[19]}}, p1_bit_slice_80042_comb} + {{4{p1_add_80043_comb[19]}}, p1_add_80043_comb};
  assign p1_add_80620_comb = {{4{p1_add_80044_comb[19]}}, p1_add_80044_comb} + {{4{p1_bit_slice_80045_comb[19]}}, p1_bit_slice_80045_comb};
  assign p1_add_80622_comb = {{4{p1_bit_slice_80046_comb[19]}}, p1_bit_slice_80046_comb} + {{4{p1_add_80047_comb[19]}}, p1_add_80047_comb};
  assign p1_add_80624_comb = {{11{p1_add_80048_comb[12]}}, p1_add_80048_comb} + {{11{p1_add_80049_comb[12]}}, p1_add_80049_comb};
  assign p1_add_80625_comb = {{11{p1_add_80050_comb[12]}}, p1_add_80050_comb} + {{11{p1_add_80051_comb[12]}}, p1_add_80051_comb};
  assign p1_add_80626_comb = {{11{p1_add_80052_comb[12]}}, p1_add_80052_comb} + {{11{p1_add_80053_comb[12]}}, p1_add_80053_comb};
  assign p1_add_80627_comb = {{11{p1_add_80054_comb[12]}}, p1_add_80054_comb} + {{11{p1_add_80055_comb[12]}}, p1_add_80055_comb};
  assign p1_add_80628_comb = {{11{p1_add_80056_comb[12]}}, p1_add_80056_comb} + {{11{p1_add_80057_comb[12]}}, p1_add_80057_comb};
  assign p1_add_80629_comb = {{11{p1_add_80058_comb[12]}}, p1_add_80058_comb} + {{11{p1_add_80059_comb[12]}}, p1_add_80059_comb};
  assign p1_add_80630_comb = {{11{p1_add_80060_comb[12]}}, p1_add_80060_comb} + {{11{p1_add_80061_comb[12]}}, p1_add_80061_comb};
  assign p1_add_80631_comb = {{11{p1_add_80062_comb[12]}}, p1_add_80062_comb} + {{11{p1_add_80063_comb[12]}}, p1_add_80063_comb};
  assign p1_add_80632_comb = {{11{p1_add_80064_comb[12]}}, p1_add_80064_comb} + {{11{p1_add_80065_comb[12]}}, p1_add_80065_comb};
  assign p1_add_80633_comb = {{11{p1_add_80066_comb[12]}}, p1_add_80066_comb} + {{11{p1_add_80067_comb[12]}}, p1_add_80067_comb};
  assign p1_add_80634_comb = {{11{p1_add_80068_comb[12]}}, p1_add_80068_comb} + {{11{p1_add_80069_comb[12]}}, p1_add_80069_comb};
  assign p1_add_80635_comb = {{11{p1_add_80070_comb[12]}}, p1_add_80070_comb} + {{11{p1_add_80071_comb[12]}}, p1_add_80071_comb};
  assign p1_add_80636_comb = {{11{p1_add_80072_comb[12]}}, p1_add_80072_comb} + {{11{p1_add_80073_comb[12]}}, p1_add_80073_comb};
  assign p1_add_80637_comb = {{11{p1_add_80074_comb[12]}}, p1_add_80074_comb} + {{11{p1_add_80075_comb[12]}}, p1_add_80075_comb};
  assign p1_add_80638_comb = {{11{p1_add_80076_comb[12]}}, p1_add_80076_comb} + {{11{p1_add_80077_comb[12]}}, p1_add_80077_comb};
  assign p1_add_80639_comb = {{11{p1_add_80078_comb[12]}}, p1_add_80078_comb} + {{11{p1_add_80079_comb[12]}}, p1_add_80079_comb};
  assign p1_sum__1246_comb = {p1_add_80400_comb, p1_add_79136_comb[0]};
  assign p1_sum__1247_comb = {p1_add_80402_comb, p1_add_79141_comb[0]};
  assign p1_sum__1232_comb = {p1_add_80404_comb, p1_add_79142_comb[0]};
  assign p1_sum__1233_comb = {p1_add_80406_comb, p1_add_79147_comb[0]};
  assign p1_sum__1218_comb = {p1_add_80408_comb, p1_add_79148_comb[0]};
  assign p1_sum__1219_comb = {p1_add_80410_comb, p1_add_79153_comb[0]};
  assign p1_sum__1204_comb = {p1_add_80412_comb, p1_add_79154_comb[0]};
  assign p1_sum__1205_comb = {p1_add_80414_comb, p1_add_79159_comb[0]};
  assign p1_sum__1190_comb = {p1_add_80416_comb, p1_add_79160_comb[0]};
  assign p1_sum__1191_comb = {p1_add_80418_comb, p1_add_79165_comb[0]};
  assign p1_sum__1176_comb = {p1_add_80420_comb, p1_add_79166_comb[0]};
  assign p1_sum__1177_comb = {p1_add_80422_comb, p1_add_79171_comb[0]};
  assign p1_sum__1162_comb = {p1_add_80424_comb, p1_add_79172_comb[0]};
  assign p1_sum__1163_comb = {p1_add_80426_comb, p1_add_79177_comb[0]};
  assign p1_sum__1148_comb = {p1_add_80428_comb, p1_add_79178_comb[0]};
  assign p1_sum__1149_comb = {p1_add_80430_comb, p1_add_79183_comb[0]};
  assign p1_sum__1242_comb = p1_sum__1572_comb + p1_sum__1573_comb;
  assign p1_sum__1243_comb = p1_sum__1574_comb + p1_sum__1575_comb;
  assign p1_sum__1228_comb = p1_sum__1544_comb + p1_sum__1545_comb;
  assign p1_sum__1229_comb = p1_sum__1546_comb + p1_sum__1547_comb;
  assign p1_sum__1214_comb = p1_sum__1516_comb + p1_sum__1517_comb;
  assign p1_sum__1215_comb = p1_sum__1518_comb + p1_sum__1519_comb;
  assign p1_sum__1200_comb = p1_sum__1488_comb + p1_sum__1489_comb;
  assign p1_sum__1201_comb = p1_sum__1490_comb + p1_sum__1491_comb;
  assign p1_sum__1186_comb = p1_sum__1460_comb + p1_sum__1461_comb;
  assign p1_sum__1187_comb = p1_sum__1462_comb + p1_sum__1463_comb;
  assign p1_sum__1172_comb = p1_sum__1432_comb + p1_sum__1433_comb;
  assign p1_sum__1173_comb = p1_sum__1434_comb + p1_sum__1435_comb;
  assign p1_sum__1158_comb = p1_sum__1404_comb + p1_sum__1405_comb;
  assign p1_sum__1159_comb = p1_sum__1406_comb + p1_sum__1407_comb;
  assign p1_sum__1144_comb = p1_sum__1376_comb + p1_sum__1377_comb;
  assign p1_sum__1145_comb = p1_sum__1378_comb + p1_sum__1379_comb;
  assign p1_sum__1240_comb = p1_sum__1568_comb + p1_sum__1569_comb;
  assign p1_sum__1241_comb = p1_sum__1570_comb + p1_sum__1571_comb;
  assign p1_sum__1226_comb = p1_sum__1540_comb + p1_sum__1541_comb;
  assign p1_sum__1227_comb = p1_sum__1542_comb + p1_sum__1543_comb;
  assign p1_sum__1212_comb = p1_sum__1512_comb + p1_sum__1513_comb;
  assign p1_sum__1213_comb = p1_sum__1514_comb + p1_sum__1515_comb;
  assign p1_sum__1198_comb = p1_sum__1484_comb + p1_sum__1485_comb;
  assign p1_sum__1199_comb = p1_sum__1486_comb + p1_sum__1487_comb;
  assign p1_sum__1184_comb = p1_sum__1456_comb + p1_sum__1457_comb;
  assign p1_sum__1185_comb = p1_sum__1458_comb + p1_sum__1459_comb;
  assign p1_sum__1170_comb = p1_sum__1428_comb + p1_sum__1429_comb;
  assign p1_sum__1171_comb = p1_sum__1430_comb + p1_sum__1431_comb;
  assign p1_sum__1156_comb = p1_sum__1400_comb + p1_sum__1401_comb;
  assign p1_sum__1157_comb = p1_sum__1402_comb + p1_sum__1403_comb;
  assign p1_sum__1142_comb = p1_sum__1372_comb + p1_sum__1373_comb;
  assign p1_sum__1143_comb = p1_sum__1374_comb + p1_sum__1375_comb;
  assign p1_sum__1238_comb = p1_sum__1564_comb + p1_sum__1565_comb;
  assign p1_sum__1239_comb = p1_sum__1566_comb + p1_sum__1567_comb;
  assign p1_sum__1224_comb = p1_sum__1536_comb + p1_sum__1537_comb;
  assign p1_sum__1225_comb = p1_sum__1538_comb + p1_sum__1539_comb;
  assign p1_sum__1210_comb = p1_sum__1508_comb + p1_sum__1509_comb;
  assign p1_sum__1211_comb = p1_sum__1510_comb + p1_sum__1511_comb;
  assign p1_sum__1196_comb = p1_sum__1480_comb + p1_sum__1481_comb;
  assign p1_sum__1197_comb = p1_sum__1482_comb + p1_sum__1483_comb;
  assign p1_sum__1182_comb = p1_sum__1452_comb + p1_sum__1453_comb;
  assign p1_sum__1183_comb = p1_sum__1454_comb + p1_sum__1455_comb;
  assign p1_sum__1168_comb = p1_sum__1424_comb + p1_sum__1425_comb;
  assign p1_sum__1169_comb = p1_sum__1426_comb + p1_sum__1427_comb;
  assign p1_sum__1154_comb = p1_sum__1396_comb + p1_sum__1397_comb;
  assign p1_sum__1155_comb = p1_sum__1398_comb + p1_sum__1399_comb;
  assign p1_sum__1140_comb = p1_sum__1368_comb + p1_sum__1369_comb;
  assign p1_sum__1141_comb = p1_sum__1370_comb + p1_sum__1371_comb;
  assign p1_sum__1234_comb = {p1_add_80592_comb, p1_add_79554_comb[0]};
  assign p1_sum__1235_comb = {p1_add_80594_comb, p1_add_79555_comb[0]};
  assign p1_sum__1220_comb = {p1_add_80596_comb, p1_add_79560_comb[0]};
  assign p1_sum__1221_comb = {p1_add_80598_comb, p1_add_79561_comb[0]};
  assign p1_sum__1206_comb = {p1_add_80600_comb, p1_add_79566_comb[0]};
  assign p1_sum__1207_comb = {p1_add_80602_comb, p1_add_79567_comb[0]};
  assign p1_sum__1192_comb = {p1_add_80604_comb, p1_add_79572_comb[0]};
  assign p1_sum__1193_comb = {p1_add_80606_comb, p1_add_79573_comb[0]};
  assign p1_sum__1178_comb = {p1_add_80608_comb, p1_add_79578_comb[0]};
  assign p1_sum__1179_comb = {p1_add_80610_comb, p1_add_79579_comb[0]};
  assign p1_sum__1164_comb = {p1_add_80612_comb, p1_add_79584_comb[0]};
  assign p1_sum__1165_comb = {p1_add_80614_comb, p1_add_79585_comb[0]};
  assign p1_sum__1150_comb = {p1_add_80616_comb, p1_add_79590_comb[0]};
  assign p1_sum__1151_comb = {p1_add_80618_comb, p1_add_79591_comb[0]};
  assign p1_sum__1136_comb = {p1_add_80620_comb, p1_add_79596_comb[0]};
  assign p1_sum__1137_comb = {p1_add_80622_comb, p1_add_79597_comb[0]};
  assign p1_add_80784_comb = p1_add_80624_comb + p1_add_80625_comb;
  assign p1_add_80786_comb = p1_add_80626_comb + p1_add_80627_comb;
  assign p1_add_80788_comb = p1_add_80628_comb + p1_add_80629_comb;
  assign p1_add_80790_comb = p1_add_80630_comb + p1_add_80631_comb;
  assign p1_add_80792_comb = p1_add_80632_comb + p1_add_80633_comb;
  assign p1_add_80794_comb = p1_add_80634_comb + p1_add_80635_comb;
  assign p1_add_80796_comb = p1_add_80636_comb + p1_add_80637_comb;
  assign p1_add_80798_comb = p1_add_80638_comb + p1_add_80639_comb;
  assign p1_sum__1079_comb = p1_sum__1246_comb + p1_sum__1247_comb;
  assign p1_sum__1072_comb = p1_sum__1232_comb + p1_sum__1233_comb;
  assign p1_sum__1065_comb = p1_sum__1218_comb + p1_sum__1219_comb;
  assign p1_sum__1058_comb = p1_sum__1204_comb + p1_sum__1205_comb;
  assign p1_sum__1051_comb = p1_sum__1190_comb + p1_sum__1191_comb;
  assign p1_sum__1044_comb = p1_sum__1176_comb + p1_sum__1177_comb;
  assign p1_sum__1037_comb = p1_sum__1162_comb + p1_sum__1163_comb;
  assign p1_sum__1030_comb = p1_sum__1148_comb + p1_sum__1149_comb;
  assign p1_add_80816_comb = {{4{p1_concat_80432_comb[19]}}, p1_concat_80432_comb} + {{4{p1_concat_80433_comb[19]}}, p1_concat_80433_comb};
  assign p1_add_80817_comb = {{4{p1_concat_80434_comb[19]}}, p1_concat_80434_comb} + {{4{p1_concat_80435_comb[19]}}, p1_concat_80435_comb};
  assign p1_add_80818_comb = {{4{p1_concat_80436_comb[19]}}, p1_concat_80436_comb} + {{4{p1_concat_80437_comb[19]}}, p1_concat_80437_comb};
  assign p1_add_80819_comb = {{4{p1_concat_80438_comb[19]}}, p1_concat_80438_comb} + {{4{p1_concat_80439_comb[19]}}, p1_concat_80439_comb};
  assign p1_add_80820_comb = {{4{p1_concat_80440_comb[19]}}, p1_concat_80440_comb} + {{4{p1_concat_80441_comb[19]}}, p1_concat_80441_comb};
  assign p1_add_80821_comb = {{4{p1_concat_80442_comb[19]}}, p1_concat_80442_comb} + {{4{p1_concat_80443_comb[19]}}, p1_concat_80443_comb};
  assign p1_add_80822_comb = {{4{p1_concat_80444_comb[19]}}, p1_concat_80444_comb} + {{4{p1_concat_80445_comb[19]}}, p1_concat_80445_comb};
  assign p1_add_80823_comb = {{4{p1_concat_80446_comb[19]}}, p1_concat_80446_comb} + {{4{p1_concat_80447_comb[19]}}, p1_concat_80447_comb};
  assign p1_add_80824_comb = {{4{p1_concat_80448_comb[19]}}, p1_concat_80448_comb} + {{4{p1_concat_80449_comb[19]}}, p1_concat_80449_comb};
  assign p1_add_80825_comb = {{4{p1_concat_80450_comb[19]}}, p1_concat_80450_comb} + {{4{p1_concat_80451_comb[19]}}, p1_concat_80451_comb};
  assign p1_add_80826_comb = {{4{p1_concat_80452_comb[19]}}, p1_concat_80452_comb} + {{4{p1_concat_80453_comb[19]}}, p1_concat_80453_comb};
  assign p1_add_80827_comb = {{4{p1_concat_80454_comb[19]}}, p1_concat_80454_comb} + {{4{p1_concat_80455_comb[19]}}, p1_concat_80455_comb};
  assign p1_add_80828_comb = {{4{p1_concat_80456_comb[19]}}, p1_concat_80456_comb} + {{4{p1_concat_80457_comb[19]}}, p1_concat_80457_comb};
  assign p1_add_80829_comb = {{4{p1_concat_80458_comb[19]}}, p1_concat_80458_comb} + {{4{p1_concat_80459_comb[19]}}, p1_concat_80459_comb};
  assign p1_add_80830_comb = {{4{p1_concat_80460_comb[19]}}, p1_concat_80460_comb} + {{4{p1_concat_80461_comb[19]}}, p1_concat_80461_comb};
  assign p1_add_80831_comb = {{4{p1_concat_80462_comb[19]}}, p1_concat_80462_comb} + {{4{p1_concat_80463_comb[19]}}, p1_concat_80463_comb};
  assign p1_sum__1077_comb = p1_sum__1242_comb + p1_sum__1243_comb;
  assign p1_sum__1070_comb = p1_sum__1228_comb + p1_sum__1229_comb;
  assign p1_sum__1063_comb = p1_sum__1214_comb + p1_sum__1215_comb;
  assign p1_sum__1056_comb = p1_sum__1200_comb + p1_sum__1201_comb;
  assign p1_sum__1049_comb = p1_sum__1186_comb + p1_sum__1187_comb;
  assign p1_sum__1042_comb = p1_sum__1172_comb + p1_sum__1173_comb;
  assign p1_sum__1035_comb = p1_sum__1158_comb + p1_sum__1159_comb;
  assign p1_sum__1028_comb = p1_sum__1144_comb + p1_sum__1145_comb;
  assign p1_sum__1076_comb = p1_sum__1240_comb + p1_sum__1241_comb;
  assign p1_sum__1069_comb = p1_sum__1226_comb + p1_sum__1227_comb;
  assign p1_sum__1062_comb = p1_sum__1212_comb + p1_sum__1213_comb;
  assign p1_sum__1055_comb = p1_sum__1198_comb + p1_sum__1199_comb;
  assign p1_sum__1048_comb = p1_sum__1184_comb + p1_sum__1185_comb;
  assign p1_sum__1041_comb = p1_sum__1170_comb + p1_sum__1171_comb;
  assign p1_sum__1034_comb = p1_sum__1156_comb + p1_sum__1157_comb;
  assign p1_sum__1027_comb = p1_sum__1142_comb + p1_sum__1143_comb;
  assign p1_sum__1075_comb = p1_sum__1238_comb + p1_sum__1239_comb;
  assign p1_sum__1068_comb = p1_sum__1224_comb + p1_sum__1225_comb;
  assign p1_sum__1061_comb = p1_sum__1210_comb + p1_sum__1211_comb;
  assign p1_sum__1054_comb = p1_sum__1196_comb + p1_sum__1197_comb;
  assign p1_sum__1047_comb = p1_sum__1182_comb + p1_sum__1183_comb;
  assign p1_sum__1040_comb = p1_sum__1168_comb + p1_sum__1169_comb;
  assign p1_sum__1033_comb = p1_sum__1154_comb + p1_sum__1155_comb;
  assign p1_sum__1026_comb = p1_sum__1140_comb + p1_sum__1141_comb;
  assign p1_add_80880_comb = {{4{p1_concat_80560_comb[19]}}, p1_concat_80560_comb} + {{4{p1_concat_80561_comb[19]}}, p1_concat_80561_comb};
  assign p1_add_80881_comb = {{4{p1_concat_80562_comb[19]}}, p1_concat_80562_comb} + {{4{p1_concat_80563_comb[19]}}, p1_concat_80563_comb};
  assign p1_add_80882_comb = {{4{p1_concat_80564_comb[19]}}, p1_concat_80564_comb} + {{4{p1_concat_80565_comb[19]}}, p1_concat_80565_comb};
  assign p1_add_80883_comb = {{4{p1_concat_80566_comb[19]}}, p1_concat_80566_comb} + {{4{p1_concat_80567_comb[19]}}, p1_concat_80567_comb};
  assign p1_add_80884_comb = {{4{p1_concat_80568_comb[19]}}, p1_concat_80568_comb} + {{4{p1_concat_80569_comb[19]}}, p1_concat_80569_comb};
  assign p1_add_80885_comb = {{4{p1_concat_80570_comb[19]}}, p1_concat_80570_comb} + {{4{p1_concat_80571_comb[19]}}, p1_concat_80571_comb};
  assign p1_add_80886_comb = {{4{p1_concat_80572_comb[19]}}, p1_concat_80572_comb} + {{4{p1_concat_80573_comb[19]}}, p1_concat_80573_comb};
  assign p1_add_80887_comb = {{4{p1_concat_80574_comb[19]}}, p1_concat_80574_comb} + {{4{p1_concat_80575_comb[19]}}, p1_concat_80575_comb};
  assign p1_add_80888_comb = {{4{p1_concat_80576_comb[19]}}, p1_concat_80576_comb} + {{4{p1_concat_80577_comb[19]}}, p1_concat_80577_comb};
  assign p1_add_80889_comb = {{4{p1_concat_80578_comb[19]}}, p1_concat_80578_comb} + {{4{p1_concat_80579_comb[19]}}, p1_concat_80579_comb};
  assign p1_add_80890_comb = {{4{p1_concat_80580_comb[19]}}, p1_concat_80580_comb} + {{4{p1_concat_80581_comb[19]}}, p1_concat_80581_comb};
  assign p1_add_80891_comb = {{4{p1_concat_80582_comb[19]}}, p1_concat_80582_comb} + {{4{p1_concat_80583_comb[19]}}, p1_concat_80583_comb};
  assign p1_add_80892_comb = {{4{p1_concat_80584_comb[19]}}, p1_concat_80584_comb} + {{4{p1_concat_80585_comb[19]}}, p1_concat_80585_comb};
  assign p1_add_80893_comb = {{4{p1_concat_80586_comb[19]}}, p1_concat_80586_comb} + {{4{p1_concat_80587_comb[19]}}, p1_concat_80587_comb};
  assign p1_add_80894_comb = {{4{p1_concat_80588_comb[19]}}, p1_concat_80588_comb} + {{4{p1_concat_80589_comb[19]}}, p1_concat_80589_comb};
  assign p1_add_80895_comb = {{4{p1_concat_80590_comb[19]}}, p1_concat_80590_comb} + {{4{p1_concat_80591_comb[19]}}, p1_concat_80591_comb};
  assign p1_sum__1073_comb = p1_sum__1234_comb + p1_sum__1235_comb;
  assign p1_sum__1066_comb = p1_sum__1220_comb + p1_sum__1221_comb;
  assign p1_sum__1059_comb = p1_sum__1206_comb + p1_sum__1207_comb;
  assign p1_sum__1052_comb = p1_sum__1192_comb + p1_sum__1193_comb;
  assign p1_sum__1045_comb = p1_sum__1178_comb + p1_sum__1179_comb;
  assign p1_sum__1038_comb = p1_sum__1164_comb + p1_sum__1165_comb;
  assign p1_sum__1031_comb = p1_sum__1150_comb + p1_sum__1151_comb;
  assign p1_sum__1024_comb = p1_sum__1136_comb + p1_sum__1137_comb;
  assign p1_umul_28632_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_80784_comb, 7'h5b);
  assign p1_umul_28634_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_80786_comb, 7'h5b);
  assign p1_umul_28636_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_80788_comb, 7'h5b);
  assign p1_umul_28638_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_80790_comb, 7'h5b);
  assign p1_umul_28640_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_80792_comb, 7'h5b);
  assign p1_umul_28642_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_80794_comb, 7'h5b);
  assign p1_umul_28644_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_80796_comb, 7'h5b);
  assign p1_umul_28646_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_80798_comb, 7'h5b);
  assign p1_add_80920_comb = p1_sum__1079_comb + 25'h000_0001;
  assign p1_add_80921_comb = p1_sum__1072_comb + 25'h000_0001;
  assign p1_add_80922_comb = p1_sum__1065_comb + 25'h000_0001;
  assign p1_add_80923_comb = p1_sum__1058_comb + 25'h000_0001;
  assign p1_add_80924_comb = p1_sum__1051_comb + 25'h000_0001;
  assign p1_add_80925_comb = p1_sum__1044_comb + 25'h000_0001;
  assign p1_add_80926_comb = p1_sum__1037_comb + 25'h000_0001;
  assign p1_add_80927_comb = p1_sum__1030_comb + 25'h000_0001;
  assign p1_add_80928_comb = p1_add_80816_comb + p1_add_80817_comb;
  assign p1_add_80929_comb = p1_add_80818_comb + p1_add_80819_comb;
  assign p1_add_80930_comb = p1_add_80820_comb + p1_add_80821_comb;
  assign p1_add_80931_comb = p1_add_80822_comb + p1_add_80823_comb;
  assign p1_add_80932_comb = p1_add_80824_comb + p1_add_80825_comb;
  assign p1_add_80933_comb = p1_add_80826_comb + p1_add_80827_comb;
  assign p1_add_80934_comb = p1_add_80828_comb + p1_add_80829_comb;
  assign p1_add_80935_comb = p1_add_80830_comb + p1_add_80831_comb;
  assign p1_add_80936_comb = p1_sum__1077_comb + 25'h000_0001;
  assign p1_add_80937_comb = p1_sum__1070_comb + 25'h000_0001;
  assign p1_add_80938_comb = p1_sum__1063_comb + 25'h000_0001;
  assign p1_add_80939_comb = p1_sum__1056_comb + 25'h000_0001;
  assign p1_add_80940_comb = p1_sum__1049_comb + 25'h000_0001;
  assign p1_add_80941_comb = p1_sum__1042_comb + 25'h000_0001;
  assign p1_add_80942_comb = p1_sum__1035_comb + 25'h000_0001;
  assign p1_add_80943_comb = p1_sum__1028_comb + 25'h000_0001;
  assign p1_add_80944_comb = p1_sum__1076_comb + 25'h000_0001;
  assign p1_add_80945_comb = p1_sum__1069_comb + 25'h000_0001;
  assign p1_add_80946_comb = p1_sum__1062_comb + 25'h000_0001;
  assign p1_add_80947_comb = p1_sum__1055_comb + 25'h000_0001;
  assign p1_add_80948_comb = p1_sum__1048_comb + 25'h000_0001;
  assign p1_add_80949_comb = p1_sum__1041_comb + 25'h000_0001;
  assign p1_add_80950_comb = p1_sum__1034_comb + 25'h000_0001;
  assign p1_add_80951_comb = p1_sum__1027_comb + 25'h000_0001;
  assign p1_add_80952_comb = p1_sum__1075_comb + 25'h000_0001;
  assign p1_add_80953_comb = p1_sum__1068_comb + 25'h000_0001;
  assign p1_add_80954_comb = p1_sum__1061_comb + 25'h000_0001;
  assign p1_add_80955_comb = p1_sum__1054_comb + 25'h000_0001;
  assign p1_add_80956_comb = p1_sum__1047_comb + 25'h000_0001;
  assign p1_add_80957_comb = p1_sum__1040_comb + 25'h000_0001;
  assign p1_add_80958_comb = p1_sum__1033_comb + 25'h000_0001;
  assign p1_add_80959_comb = p1_sum__1026_comb + 25'h000_0001;
  assign p1_add_80960_comb = p1_add_80880_comb + p1_add_80881_comb;
  assign p1_add_80961_comb = p1_add_80882_comb + p1_add_80883_comb;
  assign p1_add_80962_comb = p1_add_80884_comb + p1_add_80885_comb;
  assign p1_add_80963_comb = p1_add_80886_comb + p1_add_80887_comb;
  assign p1_add_80964_comb = p1_add_80888_comb + p1_add_80889_comb;
  assign p1_add_80965_comb = p1_add_80890_comb + p1_add_80891_comb;
  assign p1_add_80966_comb = p1_add_80892_comb + p1_add_80893_comb;
  assign p1_add_80967_comb = p1_add_80894_comb + p1_add_80895_comb;
  assign p1_add_80968_comb = p1_sum__1073_comb + 25'h000_0001;
  assign p1_add_80969_comb = p1_sum__1066_comb + 25'h000_0001;
  assign p1_add_80970_comb = p1_sum__1059_comb + 25'h000_0001;
  assign p1_add_80971_comb = p1_sum__1052_comb + 25'h000_0001;
  assign p1_add_80972_comb = p1_sum__1045_comb + 25'h000_0001;
  assign p1_add_80973_comb = p1_sum__1038_comb + 25'h000_0001;
  assign p1_add_80974_comb = p1_sum__1031_comb + 25'h000_0001;
  assign p1_add_80975_comb = p1_sum__1024_comb + 25'h000_0001;
  assign p1_bit_slice_80976_comb = p1_umul_28632_NarrowedMult__comb[23:7];
  assign p1_bit_slice_80977_comb = p1_umul_28634_NarrowedMult__comb[23:7];
  assign p1_bit_slice_80978_comb = p1_umul_28636_NarrowedMult__comb[23:7];
  assign p1_bit_slice_80979_comb = p1_umul_28638_NarrowedMult__comb[23:7];
  assign p1_bit_slice_80980_comb = p1_umul_28640_NarrowedMult__comb[23:7];
  assign p1_bit_slice_80981_comb = p1_umul_28642_NarrowedMult__comb[23:7];
  assign p1_bit_slice_80982_comb = p1_umul_28644_NarrowedMult__comb[23:7];
  assign p1_bit_slice_80983_comb = p1_umul_28646_NarrowedMult__comb[23:7];
  assign p1_bit_slice_80984_comb = p1_add_80920_comb[24:8];
  assign p1_bit_slice_80985_comb = p1_add_80921_comb[24:8];
  assign p1_bit_slice_80986_comb = p1_add_80922_comb[24:8];
  assign p1_bit_slice_80987_comb = p1_add_80923_comb[24:8];
  assign p1_bit_slice_80988_comb = p1_add_80924_comb[24:8];
  assign p1_bit_slice_80989_comb = p1_add_80925_comb[24:8];
  assign p1_bit_slice_80990_comb = p1_add_80926_comb[24:8];
  assign p1_bit_slice_80991_comb = p1_add_80927_comb[24:8];
  assign p1_bit_slice_80992_comb = p1_add_80928_comb[23:7];
  assign p1_bit_slice_80993_comb = p1_add_80929_comb[23:7];
  assign p1_bit_slice_80994_comb = p1_add_80930_comb[23:7];
  assign p1_bit_slice_80995_comb = p1_add_80931_comb[23:7];
  assign p1_bit_slice_80996_comb = p1_add_80932_comb[23:7];
  assign p1_bit_slice_80997_comb = p1_add_80933_comb[23:7];
  assign p1_bit_slice_80998_comb = p1_add_80934_comb[23:7];
  assign p1_bit_slice_80999_comb = p1_add_80935_comb[23:7];
  assign p1_bit_slice_81000_comb = p1_add_80936_comb[24:8];
  assign p1_bit_slice_81001_comb = p1_add_80937_comb[24:8];
  assign p1_bit_slice_81002_comb = p1_add_80938_comb[24:8];
  assign p1_bit_slice_81003_comb = p1_add_80939_comb[24:8];
  assign p1_bit_slice_81004_comb = p1_add_80940_comb[24:8];
  assign p1_bit_slice_81005_comb = p1_add_80941_comb[24:8];
  assign p1_bit_slice_81006_comb = p1_add_80942_comb[24:8];
  assign p1_bit_slice_81007_comb = p1_add_80943_comb[24:8];
  assign p1_bit_slice_81008_comb = p1_add_80944_comb[24:8];
  assign p1_bit_slice_81009_comb = p1_add_80945_comb[24:8];
  assign p1_bit_slice_81010_comb = p1_add_80946_comb[24:8];
  assign p1_bit_slice_81011_comb = p1_add_80947_comb[24:8];
  assign p1_bit_slice_81012_comb = p1_add_80948_comb[24:8];
  assign p1_bit_slice_81013_comb = p1_add_80949_comb[24:8];
  assign p1_bit_slice_81014_comb = p1_add_80950_comb[24:8];
  assign p1_bit_slice_81015_comb = p1_add_80951_comb[24:8];
  assign p1_bit_slice_81016_comb = p1_add_80952_comb[24:8];
  assign p1_bit_slice_81017_comb = p1_add_80953_comb[24:8];
  assign p1_bit_slice_81018_comb = p1_add_80954_comb[24:8];
  assign p1_bit_slice_81019_comb = p1_add_80955_comb[24:8];
  assign p1_bit_slice_81020_comb = p1_add_80956_comb[24:8];
  assign p1_bit_slice_81021_comb = p1_add_80957_comb[24:8];
  assign p1_bit_slice_81022_comb = p1_add_80958_comb[24:8];
  assign p1_bit_slice_81023_comb = p1_add_80959_comb[24:8];
  assign p1_bit_slice_81024_comb = p1_add_80960_comb[23:7];
  assign p1_bit_slice_81025_comb = p1_add_80961_comb[23:7];
  assign p1_bit_slice_81026_comb = p1_add_80962_comb[23:7];
  assign p1_bit_slice_81027_comb = p1_add_80963_comb[23:7];
  assign p1_bit_slice_81028_comb = p1_add_80964_comb[23:7];
  assign p1_bit_slice_81029_comb = p1_add_80965_comb[23:7];
  assign p1_bit_slice_81030_comb = p1_add_80966_comb[23:7];
  assign p1_bit_slice_81031_comb = p1_add_80967_comb[23:7];
  assign p1_bit_slice_81032_comb = p1_add_80968_comb[24:8];
  assign p1_bit_slice_81033_comb = p1_add_80969_comb[24:8];
  assign p1_bit_slice_81034_comb = p1_add_80970_comb[24:8];
  assign p1_bit_slice_81035_comb = p1_add_80971_comb[24:8];
  assign p1_bit_slice_81036_comb = p1_add_80972_comb[24:8];
  assign p1_bit_slice_81037_comb = p1_add_80973_comb[24:8];
  assign p1_bit_slice_81038_comb = p1_add_80974_comb[24:8];
  assign p1_bit_slice_81039_comb = p1_add_80975_comb[24:8];
  assign p1_add_81168_comb = {{1{p1_bit_slice_80976_comb[16]}}, p1_bit_slice_80976_comb} + 18'h0_0001;
  assign p1_add_81169_comb = {{1{p1_bit_slice_80977_comb[16]}}, p1_bit_slice_80977_comb} + 18'h0_0001;
  assign p1_add_81170_comb = {{1{p1_bit_slice_80978_comb[16]}}, p1_bit_slice_80978_comb} + 18'h0_0001;
  assign p1_add_81171_comb = {{1{p1_bit_slice_80979_comb[16]}}, p1_bit_slice_80979_comb} + 18'h0_0001;
  assign p1_add_81172_comb = {{1{p1_bit_slice_80980_comb[16]}}, p1_bit_slice_80980_comb} + 18'h0_0001;
  assign p1_add_81173_comb = {{1{p1_bit_slice_80981_comb[16]}}, p1_bit_slice_80981_comb} + 18'h0_0001;
  assign p1_add_81174_comb = {{1{p1_bit_slice_80982_comb[16]}}, p1_bit_slice_80982_comb} + 18'h0_0001;
  assign p1_add_81175_comb = {{1{p1_bit_slice_80983_comb[16]}}, p1_bit_slice_80983_comb} + 18'h0_0001;
  assign p1_add_81176_comb = {{1{p1_bit_slice_80984_comb[16]}}, p1_bit_slice_80984_comb} + 18'h0_0001;
  assign p1_add_81177_comb = {{1{p1_bit_slice_80985_comb[16]}}, p1_bit_slice_80985_comb} + 18'h0_0001;
  assign p1_add_81178_comb = {{1{p1_bit_slice_80986_comb[16]}}, p1_bit_slice_80986_comb} + 18'h0_0001;
  assign p1_add_81179_comb = {{1{p1_bit_slice_80987_comb[16]}}, p1_bit_slice_80987_comb} + 18'h0_0001;
  assign p1_add_81180_comb = {{1{p1_bit_slice_80988_comb[16]}}, p1_bit_slice_80988_comb} + 18'h0_0001;
  assign p1_add_81181_comb = {{1{p1_bit_slice_80989_comb[16]}}, p1_bit_slice_80989_comb} + 18'h0_0001;
  assign p1_add_81182_comb = {{1{p1_bit_slice_80990_comb[16]}}, p1_bit_slice_80990_comb} + 18'h0_0001;
  assign p1_add_81183_comb = {{1{p1_bit_slice_80991_comb[16]}}, p1_bit_slice_80991_comb} + 18'h0_0001;
  assign p1_add_81184_comb = {{1{p1_bit_slice_80992_comb[16]}}, p1_bit_slice_80992_comb} + 18'h0_0001;
  assign p1_add_81185_comb = {{1{p1_bit_slice_80993_comb[16]}}, p1_bit_slice_80993_comb} + 18'h0_0001;
  assign p1_add_81186_comb = {{1{p1_bit_slice_80994_comb[16]}}, p1_bit_slice_80994_comb} + 18'h0_0001;
  assign p1_add_81187_comb = {{1{p1_bit_slice_80995_comb[16]}}, p1_bit_slice_80995_comb} + 18'h0_0001;
  assign p1_add_81188_comb = {{1{p1_bit_slice_80996_comb[16]}}, p1_bit_slice_80996_comb} + 18'h0_0001;
  assign p1_add_81189_comb = {{1{p1_bit_slice_80997_comb[16]}}, p1_bit_slice_80997_comb} + 18'h0_0001;
  assign p1_add_81190_comb = {{1{p1_bit_slice_80998_comb[16]}}, p1_bit_slice_80998_comb} + 18'h0_0001;
  assign p1_add_81191_comb = {{1{p1_bit_slice_80999_comb[16]}}, p1_bit_slice_80999_comb} + 18'h0_0001;
  assign p1_add_81192_comb = {{1{p1_bit_slice_81000_comb[16]}}, p1_bit_slice_81000_comb} + 18'h0_0001;
  assign p1_add_81193_comb = {{1{p1_bit_slice_81001_comb[16]}}, p1_bit_slice_81001_comb} + 18'h0_0001;
  assign p1_add_81194_comb = {{1{p1_bit_slice_81002_comb[16]}}, p1_bit_slice_81002_comb} + 18'h0_0001;
  assign p1_add_81195_comb = {{1{p1_bit_slice_81003_comb[16]}}, p1_bit_slice_81003_comb} + 18'h0_0001;
  assign p1_add_81196_comb = {{1{p1_bit_slice_81004_comb[16]}}, p1_bit_slice_81004_comb} + 18'h0_0001;
  assign p1_add_81197_comb = {{1{p1_bit_slice_81005_comb[16]}}, p1_bit_slice_81005_comb} + 18'h0_0001;
  assign p1_add_81198_comb = {{1{p1_bit_slice_81006_comb[16]}}, p1_bit_slice_81006_comb} + 18'h0_0001;
  assign p1_add_81199_comb = {{1{p1_bit_slice_81007_comb[16]}}, p1_bit_slice_81007_comb} + 18'h0_0001;
  assign p1_add_81200_comb = {{1{p1_bit_slice_81008_comb[16]}}, p1_bit_slice_81008_comb} + 18'h0_0001;
  assign p1_add_81201_comb = {{1{p1_bit_slice_81009_comb[16]}}, p1_bit_slice_81009_comb} + 18'h0_0001;
  assign p1_add_81202_comb = {{1{p1_bit_slice_81010_comb[16]}}, p1_bit_slice_81010_comb} + 18'h0_0001;
  assign p1_add_81203_comb = {{1{p1_bit_slice_81011_comb[16]}}, p1_bit_slice_81011_comb} + 18'h0_0001;
  assign p1_add_81204_comb = {{1{p1_bit_slice_81012_comb[16]}}, p1_bit_slice_81012_comb} + 18'h0_0001;
  assign p1_add_81205_comb = {{1{p1_bit_slice_81013_comb[16]}}, p1_bit_slice_81013_comb} + 18'h0_0001;
  assign p1_add_81206_comb = {{1{p1_bit_slice_81014_comb[16]}}, p1_bit_slice_81014_comb} + 18'h0_0001;
  assign p1_add_81207_comb = {{1{p1_bit_slice_81015_comb[16]}}, p1_bit_slice_81015_comb} + 18'h0_0001;
  assign p1_add_81208_comb = {{1{p1_bit_slice_81016_comb[16]}}, p1_bit_slice_81016_comb} + 18'h0_0001;
  assign p1_add_81209_comb = {{1{p1_bit_slice_81017_comb[16]}}, p1_bit_slice_81017_comb} + 18'h0_0001;
  assign p1_add_81210_comb = {{1{p1_bit_slice_81018_comb[16]}}, p1_bit_slice_81018_comb} + 18'h0_0001;
  assign p1_add_81211_comb = {{1{p1_bit_slice_81019_comb[16]}}, p1_bit_slice_81019_comb} + 18'h0_0001;
  assign p1_add_81212_comb = {{1{p1_bit_slice_81020_comb[16]}}, p1_bit_slice_81020_comb} + 18'h0_0001;
  assign p1_add_81213_comb = {{1{p1_bit_slice_81021_comb[16]}}, p1_bit_slice_81021_comb} + 18'h0_0001;
  assign p1_add_81214_comb = {{1{p1_bit_slice_81022_comb[16]}}, p1_bit_slice_81022_comb} + 18'h0_0001;
  assign p1_add_81215_comb = {{1{p1_bit_slice_81023_comb[16]}}, p1_bit_slice_81023_comb} + 18'h0_0001;
  assign p1_add_81216_comb = {{1{p1_bit_slice_81024_comb[16]}}, p1_bit_slice_81024_comb} + 18'h0_0001;
  assign p1_add_81217_comb = {{1{p1_bit_slice_81025_comb[16]}}, p1_bit_slice_81025_comb} + 18'h0_0001;
  assign p1_add_81218_comb = {{1{p1_bit_slice_81026_comb[16]}}, p1_bit_slice_81026_comb} + 18'h0_0001;
  assign p1_add_81219_comb = {{1{p1_bit_slice_81027_comb[16]}}, p1_bit_slice_81027_comb} + 18'h0_0001;
  assign p1_add_81220_comb = {{1{p1_bit_slice_81028_comb[16]}}, p1_bit_slice_81028_comb} + 18'h0_0001;
  assign p1_add_81221_comb = {{1{p1_bit_slice_81029_comb[16]}}, p1_bit_slice_81029_comb} + 18'h0_0001;
  assign p1_add_81222_comb = {{1{p1_bit_slice_81030_comb[16]}}, p1_bit_slice_81030_comb} + 18'h0_0001;
  assign p1_add_81223_comb = {{1{p1_bit_slice_81031_comb[16]}}, p1_bit_slice_81031_comb} + 18'h0_0001;
  assign p1_add_81224_comb = {{1{p1_bit_slice_81032_comb[16]}}, p1_bit_slice_81032_comb} + 18'h0_0001;
  assign p1_add_81225_comb = {{1{p1_bit_slice_81033_comb[16]}}, p1_bit_slice_81033_comb} + 18'h0_0001;
  assign p1_add_81226_comb = {{1{p1_bit_slice_81034_comb[16]}}, p1_bit_slice_81034_comb} + 18'h0_0001;
  assign p1_add_81227_comb = {{1{p1_bit_slice_81035_comb[16]}}, p1_bit_slice_81035_comb} + 18'h0_0001;
  assign p1_add_81228_comb = {{1{p1_bit_slice_81036_comb[16]}}, p1_bit_slice_81036_comb} + 18'h0_0001;
  assign p1_add_81229_comb = {{1{p1_bit_slice_81037_comb[16]}}, p1_bit_slice_81037_comb} + 18'h0_0001;
  assign p1_add_81230_comb = {{1{p1_bit_slice_81038_comb[16]}}, p1_bit_slice_81038_comb} + 18'h0_0001;
  assign p1_add_81231_comb = {{1{p1_bit_slice_81039_comb[16]}}, p1_bit_slice_81039_comb} + 18'h0_0001;
  assign p1_clipped__136_comb = $signed(p1_add_81168_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81168_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81168_comb[12:1]);
  assign p1_clipped__152_comb = $signed(p1_add_81169_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81169_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81169_comb[12:1]);
  assign p1_clipped__168_comb = $signed(p1_add_81170_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81170_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81170_comb[12:1]);
  assign p1_clipped__184_comb = $signed(p1_add_81171_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81171_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81171_comb[12:1]);
  assign p1_clipped__200_comb = $signed(p1_add_81172_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81172_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81172_comb[12:1]);
  assign p1_clipped__216_comb = $signed(p1_add_81173_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81173_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81173_comb[12:1]);
  assign p1_clipped__232_comb = $signed(p1_add_81174_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81174_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81174_comb[12:1]);
  assign p1_clipped__248_comb = $signed(p1_add_81175_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81175_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81175_comb[12:1]);
  assign p1_clipped__137_comb = $signed(p1_add_81176_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81176_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81176_comb[12:1]);
  assign p1_clipped__153_comb = $signed(p1_add_81177_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81177_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81177_comb[12:1]);
  assign p1_clipped__169_comb = $signed(p1_add_81178_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81178_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81178_comb[12:1]);
  assign p1_clipped__185_comb = $signed(p1_add_81179_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81179_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81179_comb[12:1]);
  assign p1_clipped__201_comb = $signed(p1_add_81180_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81180_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81180_comb[12:1]);
  assign p1_clipped__217_comb = $signed(p1_add_81181_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81181_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81181_comb[12:1]);
  assign p1_clipped__233_comb = $signed(p1_add_81182_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81182_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81182_comb[12:1]);
  assign p1_clipped__249_comb = $signed(p1_add_81183_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81183_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81183_comb[12:1]);
  assign p1_clipped__138_comb = $signed(p1_add_81184_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81184_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81184_comb[12:1]);
  assign p1_clipped__154_comb = $signed(p1_add_81185_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81185_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81185_comb[12:1]);
  assign p1_clipped__170_comb = $signed(p1_add_81186_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81186_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81186_comb[12:1]);
  assign p1_clipped__186_comb = $signed(p1_add_81187_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81187_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81187_comb[12:1]);
  assign p1_clipped__202_comb = $signed(p1_add_81188_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81188_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81188_comb[12:1]);
  assign p1_clipped__218_comb = $signed(p1_add_81189_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81189_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81189_comb[12:1]);
  assign p1_clipped__234_comb = $signed(p1_add_81190_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81190_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81190_comb[12:1]);
  assign p1_clipped__250_comb = $signed(p1_add_81191_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81191_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81191_comb[12:1]);
  assign p1_clipped__139_comb = $signed(p1_add_81192_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81192_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81192_comb[12:1]);
  assign p1_clipped__155_comb = $signed(p1_add_81193_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81193_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81193_comb[12:1]);
  assign p1_clipped__171_comb = $signed(p1_add_81194_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81194_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81194_comb[12:1]);
  assign p1_clipped__187_comb = $signed(p1_add_81195_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81195_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81195_comb[12:1]);
  assign p1_clipped__203_comb = $signed(p1_add_81196_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81196_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81196_comb[12:1]);
  assign p1_clipped__219_comb = $signed(p1_add_81197_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81197_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81197_comb[12:1]);
  assign p1_clipped__235_comb = $signed(p1_add_81198_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81198_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81198_comb[12:1]);
  assign p1_clipped__251_comb = $signed(p1_add_81199_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81199_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81199_comb[12:1]);
  assign p1_clipped__140_comb = $signed(p1_add_81200_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81200_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81200_comb[12:1]);
  assign p1_clipped__156_comb = $signed(p1_add_81201_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81201_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81201_comb[12:1]);
  assign p1_clipped__172_comb = $signed(p1_add_81202_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81202_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81202_comb[12:1]);
  assign p1_clipped__188_comb = $signed(p1_add_81203_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81203_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81203_comb[12:1]);
  assign p1_clipped__204_comb = $signed(p1_add_81204_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81204_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81204_comb[12:1]);
  assign p1_clipped__220_comb = $signed(p1_add_81205_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81205_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81205_comb[12:1]);
  assign p1_clipped__236_comb = $signed(p1_add_81206_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81206_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81206_comb[12:1]);
  assign p1_clipped__252_comb = $signed(p1_add_81207_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81207_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81207_comb[12:1]);
  assign p1_clipped__141_comb = $signed(p1_add_81208_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81208_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81208_comb[12:1]);
  assign p1_clipped__157_comb = $signed(p1_add_81209_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81209_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81209_comb[12:1]);
  assign p1_clipped__173_comb = $signed(p1_add_81210_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81210_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81210_comb[12:1]);
  assign p1_clipped__189_comb = $signed(p1_add_81211_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81211_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81211_comb[12:1]);
  assign p1_clipped__205_comb = $signed(p1_add_81212_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81212_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81212_comb[12:1]);
  assign p1_clipped__221_comb = $signed(p1_add_81213_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81213_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81213_comb[12:1]);
  assign p1_clipped__237_comb = $signed(p1_add_81214_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81214_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81214_comb[12:1]);
  assign p1_clipped__253_comb = $signed(p1_add_81215_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81215_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81215_comb[12:1]);
  assign p1_clipped__142_comb = $signed(p1_add_81216_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81216_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81216_comb[12:1]);
  assign p1_clipped__158_comb = $signed(p1_add_81217_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81217_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81217_comb[12:1]);
  assign p1_clipped__174_comb = $signed(p1_add_81218_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81218_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81218_comb[12:1]);
  assign p1_clipped__190_comb = $signed(p1_add_81219_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81219_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81219_comb[12:1]);
  assign p1_clipped__206_comb = $signed(p1_add_81220_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81220_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81220_comb[12:1]);
  assign p1_clipped__222_comb = $signed(p1_add_81221_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81221_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81221_comb[12:1]);
  assign p1_clipped__238_comb = $signed(p1_add_81222_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81222_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81222_comb[12:1]);
  assign p1_clipped__254_comb = $signed(p1_add_81223_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81223_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81223_comb[12:1]);
  assign p1_clipped__143_comb = $signed(p1_add_81224_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81224_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81224_comb[12:1]);
  assign p1_clipped__159_comb = $signed(p1_add_81225_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81225_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81225_comb[12:1]);
  assign p1_clipped__175_comb = $signed(p1_add_81226_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81226_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81226_comb[12:1]);
  assign p1_clipped__191_comb = $signed(p1_add_81227_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81227_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81227_comb[12:1]);
  assign p1_clipped__207_comb = $signed(p1_add_81228_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81228_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81228_comb[12:1]);
  assign p1_clipped__223_comb = $signed(p1_add_81229_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81229_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81229_comb[12:1]);
  assign p1_clipped__239_comb = $signed(p1_add_81230_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81230_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81230_comb[12:1]);
  assign p1_clipped__255_comb = $signed(p1_add_81231_comb[17:1]) < $signed(17'h1_f800) ? 12'h800 : ($signed(p1_add_81231_comb[17:1]) > $signed(17'h0_07ff) ? 12'h7ff : p1_add_81231_comb[12:1]);
  assign p1_array_81872_comb[0] = p1_clipped__136_comb;
  assign p1_array_81872_comb[1] = p1_clipped__152_comb;
  assign p1_array_81872_comb[2] = p1_clipped__168_comb;
  assign p1_array_81872_comb[3] = p1_clipped__184_comb;
  assign p1_array_81872_comb[4] = p1_clipped__200_comb;
  assign p1_array_81872_comb[5] = p1_clipped__216_comb;
  assign p1_array_81872_comb[6] = p1_clipped__232_comb;
  assign p1_array_81872_comb[7] = p1_clipped__248_comb;
  assign p1_array_81873_comb[0] = p1_clipped__137_comb;
  assign p1_array_81873_comb[1] = p1_clipped__153_comb;
  assign p1_array_81873_comb[2] = p1_clipped__169_comb;
  assign p1_array_81873_comb[3] = p1_clipped__185_comb;
  assign p1_array_81873_comb[4] = p1_clipped__201_comb;
  assign p1_array_81873_comb[5] = p1_clipped__217_comb;
  assign p1_array_81873_comb[6] = p1_clipped__233_comb;
  assign p1_array_81873_comb[7] = p1_clipped__249_comb;
  assign p1_array_81874_comb[0] = p1_clipped__138_comb;
  assign p1_array_81874_comb[1] = p1_clipped__154_comb;
  assign p1_array_81874_comb[2] = p1_clipped__170_comb;
  assign p1_array_81874_comb[3] = p1_clipped__186_comb;
  assign p1_array_81874_comb[4] = p1_clipped__202_comb;
  assign p1_array_81874_comb[5] = p1_clipped__218_comb;
  assign p1_array_81874_comb[6] = p1_clipped__234_comb;
  assign p1_array_81874_comb[7] = p1_clipped__250_comb;
  assign p1_array_81875_comb[0] = p1_clipped__139_comb;
  assign p1_array_81875_comb[1] = p1_clipped__155_comb;
  assign p1_array_81875_comb[2] = p1_clipped__171_comb;
  assign p1_array_81875_comb[3] = p1_clipped__187_comb;
  assign p1_array_81875_comb[4] = p1_clipped__203_comb;
  assign p1_array_81875_comb[5] = p1_clipped__219_comb;
  assign p1_array_81875_comb[6] = p1_clipped__235_comb;
  assign p1_array_81875_comb[7] = p1_clipped__251_comb;
  assign p1_array_81876_comb[0] = p1_clipped__140_comb;
  assign p1_array_81876_comb[1] = p1_clipped__156_comb;
  assign p1_array_81876_comb[2] = p1_clipped__172_comb;
  assign p1_array_81876_comb[3] = p1_clipped__188_comb;
  assign p1_array_81876_comb[4] = p1_clipped__204_comb;
  assign p1_array_81876_comb[5] = p1_clipped__220_comb;
  assign p1_array_81876_comb[6] = p1_clipped__236_comb;
  assign p1_array_81876_comb[7] = p1_clipped__252_comb;
  assign p1_array_81877_comb[0] = p1_clipped__141_comb;
  assign p1_array_81877_comb[1] = p1_clipped__157_comb;
  assign p1_array_81877_comb[2] = p1_clipped__173_comb;
  assign p1_array_81877_comb[3] = p1_clipped__189_comb;
  assign p1_array_81877_comb[4] = p1_clipped__205_comb;
  assign p1_array_81877_comb[5] = p1_clipped__221_comb;
  assign p1_array_81877_comb[6] = p1_clipped__237_comb;
  assign p1_array_81877_comb[7] = p1_clipped__253_comb;
  assign p1_array_81878_comb[0] = p1_clipped__142_comb;
  assign p1_array_81878_comb[1] = p1_clipped__158_comb;
  assign p1_array_81878_comb[2] = p1_clipped__174_comb;
  assign p1_array_81878_comb[3] = p1_clipped__190_comb;
  assign p1_array_81878_comb[4] = p1_clipped__206_comb;
  assign p1_array_81878_comb[5] = p1_clipped__222_comb;
  assign p1_array_81878_comb[6] = p1_clipped__238_comb;
  assign p1_array_81878_comb[7] = p1_clipped__254_comb;
  assign p1_array_81879_comb[0] = p1_clipped__143_comb;
  assign p1_array_81879_comb[1] = p1_clipped__159_comb;
  assign p1_array_81879_comb[2] = p1_clipped__175_comb;
  assign p1_array_81879_comb[3] = p1_clipped__191_comb;
  assign p1_array_81879_comb[4] = p1_clipped__207_comb;
  assign p1_array_81879_comb[5] = p1_clipped__223_comb;
  assign p1_array_81879_comb[6] = p1_clipped__239_comb;
  assign p1_array_81879_comb[7] = p1_clipped__255_comb;
  assign p1_col_transformed_comb[0][0] = p1_array_81872_comb[0];
  assign p1_col_transformed_comb[0][1] = p1_array_81872_comb[1];
  assign p1_col_transformed_comb[0][2] = p1_array_81872_comb[2];
  assign p1_col_transformed_comb[0][3] = p1_array_81872_comb[3];
  assign p1_col_transformed_comb[0][4] = p1_array_81872_comb[4];
  assign p1_col_transformed_comb[0][5] = p1_array_81872_comb[5];
  assign p1_col_transformed_comb[0][6] = p1_array_81872_comb[6];
  assign p1_col_transformed_comb[0][7] = p1_array_81872_comb[7];
  assign p1_col_transformed_comb[1][0] = p1_array_81873_comb[0];
  assign p1_col_transformed_comb[1][1] = p1_array_81873_comb[1];
  assign p1_col_transformed_comb[1][2] = p1_array_81873_comb[2];
  assign p1_col_transformed_comb[1][3] = p1_array_81873_comb[3];
  assign p1_col_transformed_comb[1][4] = p1_array_81873_comb[4];
  assign p1_col_transformed_comb[1][5] = p1_array_81873_comb[5];
  assign p1_col_transformed_comb[1][6] = p1_array_81873_comb[6];
  assign p1_col_transformed_comb[1][7] = p1_array_81873_comb[7];
  assign p1_col_transformed_comb[2][0] = p1_array_81874_comb[0];
  assign p1_col_transformed_comb[2][1] = p1_array_81874_comb[1];
  assign p1_col_transformed_comb[2][2] = p1_array_81874_comb[2];
  assign p1_col_transformed_comb[2][3] = p1_array_81874_comb[3];
  assign p1_col_transformed_comb[2][4] = p1_array_81874_comb[4];
  assign p1_col_transformed_comb[2][5] = p1_array_81874_comb[5];
  assign p1_col_transformed_comb[2][6] = p1_array_81874_comb[6];
  assign p1_col_transformed_comb[2][7] = p1_array_81874_comb[7];
  assign p1_col_transformed_comb[3][0] = p1_array_81875_comb[0];
  assign p1_col_transformed_comb[3][1] = p1_array_81875_comb[1];
  assign p1_col_transformed_comb[3][2] = p1_array_81875_comb[2];
  assign p1_col_transformed_comb[3][3] = p1_array_81875_comb[3];
  assign p1_col_transformed_comb[3][4] = p1_array_81875_comb[4];
  assign p1_col_transformed_comb[3][5] = p1_array_81875_comb[5];
  assign p1_col_transformed_comb[3][6] = p1_array_81875_comb[6];
  assign p1_col_transformed_comb[3][7] = p1_array_81875_comb[7];
  assign p1_col_transformed_comb[4][0] = p1_array_81876_comb[0];
  assign p1_col_transformed_comb[4][1] = p1_array_81876_comb[1];
  assign p1_col_transformed_comb[4][2] = p1_array_81876_comb[2];
  assign p1_col_transformed_comb[4][3] = p1_array_81876_comb[3];
  assign p1_col_transformed_comb[4][4] = p1_array_81876_comb[4];
  assign p1_col_transformed_comb[4][5] = p1_array_81876_comb[5];
  assign p1_col_transformed_comb[4][6] = p1_array_81876_comb[6];
  assign p1_col_transformed_comb[4][7] = p1_array_81876_comb[7];
  assign p1_col_transformed_comb[5][0] = p1_array_81877_comb[0];
  assign p1_col_transformed_comb[5][1] = p1_array_81877_comb[1];
  assign p1_col_transformed_comb[5][2] = p1_array_81877_comb[2];
  assign p1_col_transformed_comb[5][3] = p1_array_81877_comb[3];
  assign p1_col_transformed_comb[5][4] = p1_array_81877_comb[4];
  assign p1_col_transformed_comb[5][5] = p1_array_81877_comb[5];
  assign p1_col_transformed_comb[5][6] = p1_array_81877_comb[6];
  assign p1_col_transformed_comb[5][7] = p1_array_81877_comb[7];
  assign p1_col_transformed_comb[6][0] = p1_array_81878_comb[0];
  assign p1_col_transformed_comb[6][1] = p1_array_81878_comb[1];
  assign p1_col_transformed_comb[6][2] = p1_array_81878_comb[2];
  assign p1_col_transformed_comb[6][3] = p1_array_81878_comb[3];
  assign p1_col_transformed_comb[6][4] = p1_array_81878_comb[4];
  assign p1_col_transformed_comb[6][5] = p1_array_81878_comb[5];
  assign p1_col_transformed_comb[6][6] = p1_array_81878_comb[6];
  assign p1_col_transformed_comb[6][7] = p1_array_81878_comb[7];
  assign p1_col_transformed_comb[7][0] = p1_array_81879_comb[0];
  assign p1_col_transformed_comb[7][1] = p1_array_81879_comb[1];
  assign p1_col_transformed_comb[7][2] = p1_array_81879_comb[2];
  assign p1_col_transformed_comb[7][3] = p1_array_81879_comb[3];
  assign p1_col_transformed_comb[7][4] = p1_array_81879_comb[4];
  assign p1_col_transformed_comb[7][5] = p1_array_81879_comb[5];
  assign p1_col_transformed_comb[7][6] = p1_array_81879_comb[6];
  assign p1_col_transformed_comb[7][7] = p1_array_81879_comb[7];

  // Registers for pipe stage 1:
  reg [11:0] p1_col_transformed[0:7][0:7];
  always @ (posedge clk) begin
    p1_col_transformed[0][0] <= p1_col_transformed_comb[0][0];
    p1_col_transformed[0][1] <= p1_col_transformed_comb[0][1];
    p1_col_transformed[0][2] <= p1_col_transformed_comb[0][2];
    p1_col_transformed[0][3] <= p1_col_transformed_comb[0][3];
    p1_col_transformed[0][4] <= p1_col_transformed_comb[0][4];
    p1_col_transformed[0][5] <= p1_col_transformed_comb[0][5];
    p1_col_transformed[0][6] <= p1_col_transformed_comb[0][6];
    p1_col_transformed[0][7] <= p1_col_transformed_comb[0][7];
    p1_col_transformed[1][0] <= p1_col_transformed_comb[1][0];
    p1_col_transformed[1][1] <= p1_col_transformed_comb[1][1];
    p1_col_transformed[1][2] <= p1_col_transformed_comb[1][2];
    p1_col_transformed[1][3] <= p1_col_transformed_comb[1][3];
    p1_col_transformed[1][4] <= p1_col_transformed_comb[1][4];
    p1_col_transformed[1][5] <= p1_col_transformed_comb[1][5];
    p1_col_transformed[1][6] <= p1_col_transformed_comb[1][6];
    p1_col_transformed[1][7] <= p1_col_transformed_comb[1][7];
    p1_col_transformed[2][0] <= p1_col_transformed_comb[2][0];
    p1_col_transformed[2][1] <= p1_col_transformed_comb[2][1];
    p1_col_transformed[2][2] <= p1_col_transformed_comb[2][2];
    p1_col_transformed[2][3] <= p1_col_transformed_comb[2][3];
    p1_col_transformed[2][4] <= p1_col_transformed_comb[2][4];
    p1_col_transformed[2][5] <= p1_col_transformed_comb[2][5];
    p1_col_transformed[2][6] <= p1_col_transformed_comb[2][6];
    p1_col_transformed[2][7] <= p1_col_transformed_comb[2][7];
    p1_col_transformed[3][0] <= p1_col_transformed_comb[3][0];
    p1_col_transformed[3][1] <= p1_col_transformed_comb[3][1];
    p1_col_transformed[3][2] <= p1_col_transformed_comb[3][2];
    p1_col_transformed[3][3] <= p1_col_transformed_comb[3][3];
    p1_col_transformed[3][4] <= p1_col_transformed_comb[3][4];
    p1_col_transformed[3][5] <= p1_col_transformed_comb[3][5];
    p1_col_transformed[3][6] <= p1_col_transformed_comb[3][6];
    p1_col_transformed[3][7] <= p1_col_transformed_comb[3][7];
    p1_col_transformed[4][0] <= p1_col_transformed_comb[4][0];
    p1_col_transformed[4][1] <= p1_col_transformed_comb[4][1];
    p1_col_transformed[4][2] <= p1_col_transformed_comb[4][2];
    p1_col_transformed[4][3] <= p1_col_transformed_comb[4][3];
    p1_col_transformed[4][4] <= p1_col_transformed_comb[4][4];
    p1_col_transformed[4][5] <= p1_col_transformed_comb[4][5];
    p1_col_transformed[4][6] <= p1_col_transformed_comb[4][6];
    p1_col_transformed[4][7] <= p1_col_transformed_comb[4][7];
    p1_col_transformed[5][0] <= p1_col_transformed_comb[5][0];
    p1_col_transformed[5][1] <= p1_col_transformed_comb[5][1];
    p1_col_transformed[5][2] <= p1_col_transformed_comb[5][2];
    p1_col_transformed[5][3] <= p1_col_transformed_comb[5][3];
    p1_col_transformed[5][4] <= p1_col_transformed_comb[5][4];
    p1_col_transformed[5][5] <= p1_col_transformed_comb[5][5];
    p1_col_transformed[5][6] <= p1_col_transformed_comb[5][6];
    p1_col_transformed[5][7] <= p1_col_transformed_comb[5][7];
    p1_col_transformed[6][0] <= p1_col_transformed_comb[6][0];
    p1_col_transformed[6][1] <= p1_col_transformed_comb[6][1];
    p1_col_transformed[6][2] <= p1_col_transformed_comb[6][2];
    p1_col_transformed[6][3] <= p1_col_transformed_comb[6][3];
    p1_col_transformed[6][4] <= p1_col_transformed_comb[6][4];
    p1_col_transformed[6][5] <= p1_col_transformed_comb[6][5];
    p1_col_transformed[6][6] <= p1_col_transformed_comb[6][6];
    p1_col_transformed[6][7] <= p1_col_transformed_comb[6][7];
    p1_col_transformed[7][0] <= p1_col_transformed_comb[7][0];
    p1_col_transformed[7][1] <= p1_col_transformed_comb[7][1];
    p1_col_transformed[7][2] <= p1_col_transformed_comb[7][2];
    p1_col_transformed[7][3] <= p1_col_transformed_comb[7][3];
    p1_col_transformed[7][4] <= p1_col_transformed_comb[7][4];
    p1_col_transformed[7][5] <= p1_col_transformed_comb[7][5];
    p1_col_transformed[7][6] <= p1_col_transformed_comb[7][6];
    p1_col_transformed[7][7] <= p1_col_transformed_comb[7][7];
  end
  assign out = {{p1_col_transformed[7][7], p1_col_transformed[7][6], p1_col_transformed[7][5], p1_col_transformed[7][4], p1_col_transformed[7][3], p1_col_transformed[7][2], p1_col_transformed[7][1], p1_col_transformed[7][0]}, {p1_col_transformed[6][7], p1_col_transformed[6][6], p1_col_transformed[6][5], p1_col_transformed[6][4], p1_col_transformed[6][3], p1_col_transformed[6][2], p1_col_transformed[6][1], p1_col_transformed[6][0]}, {p1_col_transformed[5][7], p1_col_transformed[5][6], p1_col_transformed[5][5], p1_col_transformed[5][4], p1_col_transformed[5][3], p1_col_transformed[5][2], p1_col_transformed[5][1], p1_col_transformed[5][0]}, {p1_col_transformed[4][7], p1_col_transformed[4][6], p1_col_transformed[4][5], p1_col_transformed[4][4], p1_col_transformed[4][3], p1_col_transformed[4][2], p1_col_transformed[4][1], p1_col_transformed[4][0]}, {p1_col_transformed[3][7], p1_col_transformed[3][6], p1_col_transformed[3][5], p1_col_transformed[3][4], p1_col_transformed[3][3], p1_col_transformed[3][2], p1_col_transformed[3][1], p1_col_transformed[3][0]}, {p1_col_transformed[2][7], p1_col_transformed[2][6], p1_col_transformed[2][5], p1_col_transformed[2][4], p1_col_transformed[2][3], p1_col_transformed[2][2], p1_col_transformed[2][1], p1_col_transformed[2][0]}, {p1_col_transformed[1][7], p1_col_transformed[1][6], p1_col_transformed[1][5], p1_col_transformed[1][4], p1_col_transformed[1][3], p1_col_transformed[1][2], p1_col_transformed[1][1], p1_col_transformed[1][0]}, {p1_col_transformed[0][7], p1_col_transformed[0][6], p1_col_transformed[0][5], p1_col_transformed[0][4], p1_col_transformed[0][3], p1_col_transformed[0][2], p1_col_transformed[0][1], p1_col_transformed[0][0]}};
endmodule
