module dct_2d_s12(
  input wire clk,
  input wire [767:0] x,
  output wire [767:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [17:0] smul18b_12b_x_6b (input reg [11:0] lhs, input reg [5:0] rhs);
    reg signed [11:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [17:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul18b_12b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [18:0] smul19b_12b_x_7b (input reg [11:0] lhs, input reg [6:0] rhs);
    reg signed [11:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [18:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul19b_12b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [20:0] smul21b_12b_x_9b (input reg [11:0] lhs, input reg [8:0] rhs);
    reg signed [11:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [20:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul21b_12b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [19:0] smul20b_12b_x_8b (input reg [11:0] lhs, input reg [7:0] rhs);
    reg signed [11:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [19:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul20b_12b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_7b (input reg [31:0] lhs, input reg [6:0] rhs);
    begin
      umul32b_32b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [11:0] x_unflattened[0:7][0:7];
  assign x_unflattened[0][0] = x[11:0];
  assign x_unflattened[0][1] = x[23:12];
  assign x_unflattened[0][2] = x[35:24];
  assign x_unflattened[0][3] = x[47:36];
  assign x_unflattened[0][4] = x[59:48];
  assign x_unflattened[0][5] = x[71:60];
  assign x_unflattened[0][6] = x[83:72];
  assign x_unflattened[0][7] = x[95:84];
  assign x_unflattened[1][0] = x[107:96];
  assign x_unflattened[1][1] = x[119:108];
  assign x_unflattened[1][2] = x[131:120];
  assign x_unflattened[1][3] = x[143:132];
  assign x_unflattened[1][4] = x[155:144];
  assign x_unflattened[1][5] = x[167:156];
  assign x_unflattened[1][6] = x[179:168];
  assign x_unflattened[1][7] = x[191:180];
  assign x_unflattened[2][0] = x[203:192];
  assign x_unflattened[2][1] = x[215:204];
  assign x_unflattened[2][2] = x[227:216];
  assign x_unflattened[2][3] = x[239:228];
  assign x_unflattened[2][4] = x[251:240];
  assign x_unflattened[2][5] = x[263:252];
  assign x_unflattened[2][6] = x[275:264];
  assign x_unflattened[2][7] = x[287:276];
  assign x_unflattened[3][0] = x[299:288];
  assign x_unflattened[3][1] = x[311:300];
  assign x_unflattened[3][2] = x[323:312];
  assign x_unflattened[3][3] = x[335:324];
  assign x_unflattened[3][4] = x[347:336];
  assign x_unflattened[3][5] = x[359:348];
  assign x_unflattened[3][6] = x[371:360];
  assign x_unflattened[3][7] = x[383:372];
  assign x_unflattened[4][0] = x[395:384];
  assign x_unflattened[4][1] = x[407:396];
  assign x_unflattened[4][2] = x[419:408];
  assign x_unflattened[4][3] = x[431:420];
  assign x_unflattened[4][4] = x[443:432];
  assign x_unflattened[4][5] = x[455:444];
  assign x_unflattened[4][6] = x[467:456];
  assign x_unflattened[4][7] = x[479:468];
  assign x_unflattened[5][0] = x[491:480];
  assign x_unflattened[5][1] = x[503:492];
  assign x_unflattened[5][2] = x[515:504];
  assign x_unflattened[5][3] = x[527:516];
  assign x_unflattened[5][4] = x[539:528];
  assign x_unflattened[5][5] = x[551:540];
  assign x_unflattened[5][6] = x[563:552];
  assign x_unflattened[5][7] = x[575:564];
  assign x_unflattened[6][0] = x[587:576];
  assign x_unflattened[6][1] = x[599:588];
  assign x_unflattened[6][2] = x[611:600];
  assign x_unflattened[6][3] = x[623:612];
  assign x_unflattened[6][4] = x[635:624];
  assign x_unflattened[6][5] = x[647:636];
  assign x_unflattened[6][6] = x[659:648];
  assign x_unflattened[6][7] = x[671:660];
  assign x_unflattened[7][0] = x[683:672];
  assign x_unflattened[7][1] = x[695:684];
  assign x_unflattened[7][2] = x[707:696];
  assign x_unflattened[7][3] = x[719:708];
  assign x_unflattened[7][4] = x[731:720];
  assign x_unflattened[7][5] = x[743:732];
  assign x_unflattened[7][6] = x[755:744];
  assign x_unflattened[7][7] = x[767:756];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [11:0] p0_x[0:7][0:7];
  always @ (posedge clk) begin
    p0_x[0][0] <= x_unflattened[0][0];
    p0_x[0][1] <= x_unflattened[0][1];
    p0_x[0][2] <= x_unflattened[0][2];
    p0_x[0][3] <= x_unflattened[0][3];
    p0_x[0][4] <= x_unflattened[0][4];
    p0_x[0][5] <= x_unflattened[0][5];
    p0_x[0][6] <= x_unflattened[0][6];
    p0_x[0][7] <= x_unflattened[0][7];
    p0_x[1][0] <= x_unflattened[1][0];
    p0_x[1][1] <= x_unflattened[1][1];
    p0_x[1][2] <= x_unflattened[1][2];
    p0_x[1][3] <= x_unflattened[1][3];
    p0_x[1][4] <= x_unflattened[1][4];
    p0_x[1][5] <= x_unflattened[1][5];
    p0_x[1][6] <= x_unflattened[1][6];
    p0_x[1][7] <= x_unflattened[1][7];
    p0_x[2][0] <= x_unflattened[2][0];
    p0_x[2][1] <= x_unflattened[2][1];
    p0_x[2][2] <= x_unflattened[2][2];
    p0_x[2][3] <= x_unflattened[2][3];
    p0_x[2][4] <= x_unflattened[2][4];
    p0_x[2][5] <= x_unflattened[2][5];
    p0_x[2][6] <= x_unflattened[2][6];
    p0_x[2][7] <= x_unflattened[2][7];
    p0_x[3][0] <= x_unflattened[3][0];
    p0_x[3][1] <= x_unflattened[3][1];
    p0_x[3][2] <= x_unflattened[3][2];
    p0_x[3][3] <= x_unflattened[3][3];
    p0_x[3][4] <= x_unflattened[3][4];
    p0_x[3][5] <= x_unflattened[3][5];
    p0_x[3][6] <= x_unflattened[3][6];
    p0_x[3][7] <= x_unflattened[3][7];
    p0_x[4][0] <= x_unflattened[4][0];
    p0_x[4][1] <= x_unflattened[4][1];
    p0_x[4][2] <= x_unflattened[4][2];
    p0_x[4][3] <= x_unflattened[4][3];
    p0_x[4][4] <= x_unflattened[4][4];
    p0_x[4][5] <= x_unflattened[4][5];
    p0_x[4][6] <= x_unflattened[4][6];
    p0_x[4][7] <= x_unflattened[4][7];
    p0_x[5][0] <= x_unflattened[5][0];
    p0_x[5][1] <= x_unflattened[5][1];
    p0_x[5][2] <= x_unflattened[5][2];
    p0_x[5][3] <= x_unflattened[5][3];
    p0_x[5][4] <= x_unflattened[5][4];
    p0_x[5][5] <= x_unflattened[5][5];
    p0_x[5][6] <= x_unflattened[5][6];
    p0_x[5][7] <= x_unflattened[5][7];
    p0_x[6][0] <= x_unflattened[6][0];
    p0_x[6][1] <= x_unflattened[6][1];
    p0_x[6][2] <= x_unflattened[6][2];
    p0_x[6][3] <= x_unflattened[6][3];
    p0_x[6][4] <= x_unflattened[6][4];
    p0_x[6][5] <= x_unflattened[6][5];
    p0_x[6][6] <= x_unflattened[6][6];
    p0_x[6][7] <= x_unflattened[6][7];
    p0_x[7][0] <= x_unflattened[7][0];
    p0_x[7][1] <= x_unflattened[7][1];
    p0_x[7][2] <= x_unflattened[7][2];
    p0_x[7][3] <= x_unflattened[7][3];
    p0_x[7][4] <= x_unflattened[7][4];
    p0_x[7][5] <= x_unflattened[7][5];
    p0_x[7][6] <= x_unflattened[7][6];
    p0_x[7][7] <= x_unflattened[7][7];
  end

  // ===== Pipe stage 1:
  wire [11:0] p1_array_index_66799_comb;
  wire [11:0] p1_array_index_66801_comb;
  wire [11:0] p1_array_index_66803_comb;
  wire [11:0] p1_array_index_66805_comb;
  wire [11:0] p1_array_index_66807_comb;
  wire [11:0] p1_array_index_66809_comb;
  wire [11:0] p1_array_index_66811_comb;
  wire [11:0] p1_array_index_66813_comb;
  wire [11:0] p1_array_index_66815_comb;
  wire [11:0] p1_array_index_66817_comb;
  wire [11:0] p1_array_index_66819_comb;
  wire [11:0] p1_array_index_66821_comb;
  wire [11:0] p1_array_index_66831_comb;
  wire [11:0] p1_array_index_66835_comb;
  wire [11:0] p1_array_index_66837_comb;
  wire [11:0] p1_array_index_66841_comb;
  wire [11:0] p1_array_index_66847_comb;
  wire [11:0] p1_array_index_66849_comb;
  wire [11:0] p1_array_index_66851_comb;
  wire [11:0] p1_array_index_66853_comb;
  wire [11:0] p1_array_index_66855_comb;
  wire [11:0] p1_array_index_66857_comb;
  wire [11:0] p1_array_index_66859_comb;
  wire [11:0] p1_array_index_66861_comb;
  wire [11:0] p1_array_index_66863_comb;
  wire [11:0] p1_array_index_66865_comb;
  wire [11:0] p1_array_index_66867_comb;
  wire [11:0] p1_array_index_66869_comb;
  wire [11:0] p1_array_index_66871_comb;
  wire [11:0] p1_array_index_66873_comb;
  wire [11:0] p1_array_index_66875_comb;
  wire [11:0] p1_array_index_66877_comb;
  wire [11:0] p1_array_index_66879_comb;
  wire [11:0] p1_array_index_66881_comb;
  wire [11:0] p1_array_index_66883_comb;
  wire [11:0] p1_array_index_66885_comb;
  wire [11:0] p1_array_index_66887_comb;
  wire [11:0] p1_array_index_66889_comb;
  wire [11:0] p1_array_index_66891_comb;
  wire [11:0] p1_array_index_66893_comb;
  wire [11:0] p1_array_index_66911_comb;
  wire [11:0] p1_array_index_66915_comb;
  wire [11:0] p1_array_index_66917_comb;
  wire [11:0] p1_array_index_66921_comb;
  wire [11:0] p1_array_index_66923_comb;
  wire [11:0] p1_array_index_66927_comb;
  wire [11:0] p1_array_index_66929_comb;
  wire [11:0] p1_array_index_66933_comb;
  wire [11:0] p1_array_index_66943_comb;
  wire [11:0] p1_array_index_66945_comb;
  wire [11:0] p1_array_index_66947_comb;
  wire [11:0] p1_array_index_66949_comb;
  wire [11:0] p1_array_index_66951_comb;
  wire [11:0] p1_array_index_66953_comb;
  wire [11:0] p1_array_index_66955_comb;
  wire [11:0] p1_array_index_66957_comb;
  wire [11:0] p1_array_index_66959_comb;
  wire [11:0] p1_array_index_66961_comb;
  wire [11:0] p1_array_index_66963_comb;
  wire [11:0] p1_array_index_66965_comb;
  wire [11:0] p1_array_index_66975_comb;
  wire [11:0] p1_array_index_66979_comb;
  wire [11:0] p1_array_index_66981_comb;
  wire [11:0] p1_array_index_66985_comb;
  wire [17:0] p1_smul_27786_NarrowedMult__comb;
  wire [17:0] p1_smul_27788_NarrowedMult__comb;
  wire [17:0] p1_smul_27802_NarrowedMult__comb;
  wire [17:0] p1_smul_27804_NarrowedMult__comb;
  wire [18:0] p1_smul_27910_NarrowedMult__comb;
  wire [18:0] p1_smul_27912_NarrowedMult__comb;
  wire [18:0] p1_smul_27918_NarrowedMult__comb;
  wire [18:0] p1_smul_27920_NarrowedMult__comb;
  wire [18:0] p1_smul_27926_NarrowedMult__comb;
  wire [18:0] p1_smul_27928_NarrowedMult__comb;
  wire [18:0] p1_smul_27934_NarrowedMult__comb;
  wire [18:0] p1_smul_27936_NarrowedMult__comb;
  wire [17:0] p1_smul_28038_NarrowedMult__comb;
  wire [17:0] p1_smul_28048_NarrowedMult__comb;
  wire [17:0] p1_smul_28054_NarrowedMult__comb;
  wire [17:0] p1_smul_28064_NarrowedMult__comb;
  wire [17:0] p1_smul_28296_NarrowedMult__comb;
  wire [17:0] p1_smul_28302_NarrowedMult__comb;
  wire [17:0] p1_smul_28312_NarrowedMult__comb;
  wire [17:0] p1_smul_28318_NarrowedMult__comb;
  wire [18:0] p1_smul_28420_NarrowedMult__comb;
  wire [18:0] p1_smul_28424_NarrowedMult__comb;
  wire [18:0] p1_smul_28430_NarrowedMult__comb;
  wire [18:0] p1_smul_28434_NarrowedMult__comb;
  wire [18:0] p1_smul_28436_NarrowedMult__comb;
  wire [18:0] p1_smul_28440_NarrowedMult__comb;
  wire [18:0] p1_smul_28446_NarrowedMult__comb;
  wire [18:0] p1_smul_28450_NarrowedMult__comb;
  wire [17:0] p1_smul_28548_NarrowedMult__comb;
  wire [17:0] p1_smul_28562_NarrowedMult__comb;
  wire [17:0] p1_smul_28564_NarrowedMult__comb;
  wire [17:0] p1_smul_28578_NarrowedMult__comb;
  wire [17:0] p1_smul_27754_NarrowedMult__comb;
  wire [17:0] p1_smul_27756_NarrowedMult__comb;
  wire [17:0] p1_smul_27770_NarrowedMult__comb;
  wire [17:0] p1_smul_27772_NarrowedMult__comb;
  wire [17:0] p1_smul_27818_NarrowedMult__comb;
  wire [17:0] p1_smul_27820_NarrowedMult__comb;
  wire [17:0] p1_smul_27834_NarrowedMult__comb;
  wire [17:0] p1_smul_27836_NarrowedMult__comb;
  wire [18:0] p1_smul_27878_NarrowedMult__comb;
  wire [18:0] p1_smul_27880_NarrowedMult__comb;
  wire [18:0] p1_smul_27886_NarrowedMult__comb;
  wire [18:0] p1_smul_27888_NarrowedMult__comb;
  wire [18:0] p1_smul_27894_NarrowedMult__comb;
  wire [18:0] p1_smul_27896_NarrowedMult__comb;
  wire [18:0] p1_smul_27902_NarrowedMult__comb;
  wire [18:0] p1_smul_27904_NarrowedMult__comb;
  wire [18:0] p1_smul_27942_NarrowedMult__comb;
  wire [18:0] p1_smul_27944_NarrowedMult__comb;
  wire [18:0] p1_smul_27950_NarrowedMult__comb;
  wire [18:0] p1_smul_27952_NarrowedMult__comb;
  wire [18:0] p1_smul_27958_NarrowedMult__comb;
  wire [18:0] p1_smul_27960_NarrowedMult__comb;
  wire [18:0] p1_smul_27966_NarrowedMult__comb;
  wire [18:0] p1_smul_27968_NarrowedMult__comb;
  wire [17:0] p1_smul_28006_NarrowedMult__comb;
  wire [17:0] p1_smul_28016_NarrowedMult__comb;
  wire [17:0] p1_smul_28022_NarrowedMult__comb;
  wire [17:0] p1_smul_28032_NarrowedMult__comb;
  wire [17:0] p1_smul_28070_NarrowedMult__comb;
  wire [17:0] p1_smul_28080_NarrowedMult__comb;
  wire [17:0] p1_smul_28086_NarrowedMult__comb;
  wire [17:0] p1_smul_28096_NarrowedMult__comb;
  wire [17:0] p1_smul_28264_NarrowedMult__comb;
  wire [17:0] p1_smul_28270_NarrowedMult__comb;
  wire [17:0] p1_smul_28280_NarrowedMult__comb;
  wire [17:0] p1_smul_28286_NarrowedMult__comb;
  wire [17:0] p1_smul_28328_NarrowedMult__comb;
  wire [17:0] p1_smul_28334_NarrowedMult__comb;
  wire [17:0] p1_smul_28344_NarrowedMult__comb;
  wire [17:0] p1_smul_28350_NarrowedMult__comb;
  wire [18:0] p1_smul_28388_NarrowedMult__comb;
  wire [18:0] p1_smul_28392_NarrowedMult__comb;
  wire [18:0] p1_smul_28398_NarrowedMult__comb;
  wire [18:0] p1_smul_28402_NarrowedMult__comb;
  wire [18:0] p1_smul_28404_NarrowedMult__comb;
  wire [18:0] p1_smul_28408_NarrowedMult__comb;
  wire [18:0] p1_smul_28414_NarrowedMult__comb;
  wire [18:0] p1_smul_28418_NarrowedMult__comb;
  wire [18:0] p1_smul_28452_NarrowedMult__comb;
  wire [18:0] p1_smul_28456_NarrowedMult__comb;
  wire [18:0] p1_smul_28462_NarrowedMult__comb;
  wire [18:0] p1_smul_28466_NarrowedMult__comb;
  wire [18:0] p1_smul_28468_NarrowedMult__comb;
  wire [18:0] p1_smul_28472_NarrowedMult__comb;
  wire [18:0] p1_smul_28478_NarrowedMult__comb;
  wire [18:0] p1_smul_28482_NarrowedMult__comb;
  wire [17:0] p1_smul_28516_NarrowedMult__comb;
  wire [17:0] p1_smul_28530_NarrowedMult__comb;
  wire [17:0] p1_smul_28532_NarrowedMult__comb;
  wire [17:0] p1_smul_28546_NarrowedMult__comb;
  wire [17:0] p1_smul_28580_NarrowedMult__comb;
  wire [17:0] p1_smul_28594_NarrowedMult__comb;
  wire [17:0] p1_smul_28596_NarrowedMult__comb;
  wire [17:0] p1_smul_28610_NarrowedMult__comb;
  wire [17:0] p1_smul_27738_NarrowedMult__comb;
  wire [17:0] p1_smul_27740_NarrowedMult__comb;
  wire [17:0] p1_smul_27850_NarrowedMult__comb;
  wire [17:0] p1_smul_27852_NarrowedMult__comb;
  wire [18:0] p1_smul_27862_NarrowedMult__comb;
  wire [18:0] p1_smul_27864_NarrowedMult__comb;
  wire [18:0] p1_smul_27870_NarrowedMult__comb;
  wire [18:0] p1_smul_27872_NarrowedMult__comb;
  wire [18:0] p1_smul_27974_NarrowedMult__comb;
  wire [18:0] p1_smul_27976_NarrowedMult__comb;
  wire [18:0] p1_smul_27982_NarrowedMult__comb;
  wire [18:0] p1_smul_27984_NarrowedMult__comb;
  wire [17:0] p1_smul_27990_NarrowedMult__comb;
  wire [17:0] p1_smul_28000_NarrowedMult__comb;
  wire [17:0] p1_smul_28102_NarrowedMult__comb;
  wire [17:0] p1_smul_28112_NarrowedMult__comb;
  wire [17:0] p1_smul_28248_NarrowedMult__comb;
  wire [17:0] p1_smul_28254_NarrowedMult__comb;
  wire [17:0] p1_smul_28360_NarrowedMult__comb;
  wire [17:0] p1_smul_28366_NarrowedMult__comb;
  wire [18:0] p1_smul_28372_NarrowedMult__comb;
  wire [18:0] p1_smul_28376_NarrowedMult__comb;
  wire [18:0] p1_smul_28382_NarrowedMult__comb;
  wire [18:0] p1_smul_28386_NarrowedMult__comb;
  wire [18:0] p1_smul_28484_NarrowedMult__comb;
  wire [18:0] p1_smul_28488_NarrowedMult__comb;
  wire [18:0] p1_smul_28494_NarrowedMult__comb;
  wire [18:0] p1_smul_28498_NarrowedMult__comb;
  wire [17:0] p1_smul_28500_NarrowedMult__comb;
  wire [17:0] p1_smul_28514_NarrowedMult__comb;
  wire [17:0] p1_smul_28612_NarrowedMult__comb;
  wire [17:0] p1_smul_28626_NarrowedMult__comb;
  wire [20:0] p1_smul_67439_comb;
  wire [20:0] p1_smul_67440_comb;
  wire [19:0] p1_smul_27784_NarrowedMult__comb;
  wire [19:0] p1_smul_27790_NarrowedMult__comb;
  wire [20:0] p1_smul_67447_comb;
  wire [20:0] p1_smul_67448_comb;
  wire [20:0] p1_smul_67449_comb;
  wire [20:0] p1_smul_67450_comb;
  wire [19:0] p1_smul_27800_NarrowedMult__comb;
  wire [19:0] p1_smul_27806_NarrowedMult__comb;
  wire [20:0] p1_smul_67457_comb;
  wire [20:0] p1_smul_67458_comb;
  wire [18:0] p1_smul_27908_NarrowedMult__comb;
  wire [18:0] p1_smul_27914_NarrowedMult__comb;
  wire [18:0] p1_smul_27916_NarrowedMult__comb;
  wire [18:0] p1_smul_27922_NarrowedMult__comb;
  wire [18:0] p1_smul_27924_NarrowedMult__comb;
  wire [18:0] p1_smul_27930_NarrowedMult__comb;
  wire [18:0] p1_smul_27932_NarrowedMult__comb;
  wire [18:0] p1_smul_27938_NarrowedMult__comb;
  wire [20:0] p1_smul_67483_comb;
  wire [20:0] p1_smul_67486_comb;
  wire [19:0] p1_smul_28042_NarrowedMult__comb;
  wire [19:0] p1_smul_28044_NarrowedMult__comb;
  wire [20:0] p1_smul_67489_comb;
  wire [20:0] p1_smul_67492_comb;
  wire [20:0] p1_smul_67493_comb;
  wire [20:0] p1_smul_67496_comb;
  wire [19:0] p1_smul_28058_NarrowedMult__comb;
  wire [19:0] p1_smul_28060_NarrowedMult__comb;
  wire [20:0] p1_smul_67499_comb;
  wire [20:0] p1_smul_67502_comb;
  wire [20:0] p1_smul_67503_comb;
  wire [20:0] p1_smul_67504_comb;
  wire [20:0] p1_smul_67505_comb;
  wire [20:0] p1_smul_67506_comb;
  wire [20:0] p1_smul_67507_comb;
  wire [20:0] p1_smul_67508_comb;
  wire [20:0] p1_smul_67509_comb;
  wire [20:0] p1_smul_67510_comb;
  wire [20:0] p1_smul_67511_comb;
  wire [20:0] p1_smul_67512_comb;
  wire [20:0] p1_smul_67513_comb;
  wire [20:0] p1_smul_67514_comb;
  wire [20:0] p1_smul_67515_comb;
  wire [20:0] p1_smul_67516_comb;
  wire [20:0] p1_smul_67517_comb;
  wire [20:0] p1_smul_67518_comb;
  wire [19:0] p1_smul_28292_NarrowedMult__comb;
  wire [20:0] p1_smul_67520_comb;
  wire [20:0] p1_smul_67523_comb;
  wire [20:0] p1_smul_67524_comb;
  wire [20:0] p1_smul_67527_comb;
  wire [19:0] p1_smul_28306_NarrowedMult__comb;
  wire [19:0] p1_smul_28308_NarrowedMult__comb;
  wire [20:0] p1_smul_67530_comb;
  wire [20:0] p1_smul_67533_comb;
  wire [20:0] p1_smul_67534_comb;
  wire [20:0] p1_smul_67537_comb;
  wire [19:0] p1_smul_28322_NarrowedMult__comb;
  wire [18:0] p1_smul_28422_NarrowedMult__comb;
  wire [18:0] p1_smul_28426_NarrowedMult__comb;
  wire [18:0] p1_smul_28428_NarrowedMult__comb;
  wire [18:0] p1_smul_28432_NarrowedMult__comb;
  wire [18:0] p1_smul_28438_NarrowedMult__comb;
  wire [18:0] p1_smul_28442_NarrowedMult__comb;
  wire [18:0] p1_smul_28444_NarrowedMult__comb;
  wire [18:0] p1_smul_28448_NarrowedMult__comb;
  wire [19:0] p1_smul_28550_NarrowedMult__comb;
  wire [20:0] p1_smul_67566_comb;
  wire [20:0] p1_smul_67567_comb;
  wire [20:0] p1_smul_67568_comb;
  wire [20:0] p1_smul_67569_comb;
  wire [19:0] p1_smul_28560_NarrowedMult__comb;
  wire [19:0] p1_smul_28566_NarrowedMult__comb;
  wire [20:0] p1_smul_67576_comb;
  wire [20:0] p1_smul_67577_comb;
  wire [20:0] p1_smul_67578_comb;
  wire [20:0] p1_smul_67579_comb;
  wire [19:0] p1_smul_28576_NarrowedMult__comb;
  wire [20:0] p1_smul_67583_comb;
  wire [20:0] p1_smul_67584_comb;
  wire [19:0] p1_smul_27752_NarrowedMult__comb;
  wire [19:0] p1_smul_27758_NarrowedMult__comb;
  wire [20:0] p1_smul_67591_comb;
  wire [20:0] p1_smul_67592_comb;
  wire [20:0] p1_smul_67593_comb;
  wire [20:0] p1_smul_67594_comb;
  wire [19:0] p1_smul_27768_NarrowedMult__comb;
  wire [19:0] p1_smul_27774_NarrowedMult__comb;
  wire [20:0] p1_smul_67601_comb;
  wire [20:0] p1_smul_67602_comb;
  wire [20:0] p1_smul_67603_comb;
  wire [20:0] p1_smul_67604_comb;
  wire [19:0] p1_smul_27816_NarrowedMult__comb;
  wire [19:0] p1_smul_27822_NarrowedMult__comb;
  wire [20:0] p1_smul_67611_comb;
  wire [20:0] p1_smul_67612_comb;
  wire [20:0] p1_smul_67613_comb;
  wire [20:0] p1_smul_67614_comb;
  wire [19:0] p1_smul_27832_NarrowedMult__comb;
  wire [19:0] p1_smul_27838_NarrowedMult__comb;
  wire [20:0] p1_smul_67621_comb;
  wire [20:0] p1_smul_67622_comb;
  wire [18:0] p1_smul_27876_NarrowedMult__comb;
  wire [18:0] p1_smul_27882_NarrowedMult__comb;
  wire [18:0] p1_smul_27884_NarrowedMult__comb;
  wire [18:0] p1_smul_27890_NarrowedMult__comb;
  wire [18:0] p1_smul_27892_NarrowedMult__comb;
  wire [18:0] p1_smul_27898_NarrowedMult__comb;
  wire [18:0] p1_smul_27900_NarrowedMult__comb;
  wire [18:0] p1_smul_27906_NarrowedMult__comb;
  wire [18:0] p1_smul_27940_NarrowedMult__comb;
  wire [18:0] p1_smul_27946_NarrowedMult__comb;
  wire [18:0] p1_smul_27948_NarrowedMult__comb;
  wire [18:0] p1_smul_27954_NarrowedMult__comb;
  wire [18:0] p1_smul_27956_NarrowedMult__comb;
  wire [18:0] p1_smul_27962_NarrowedMult__comb;
  wire [18:0] p1_smul_27964_NarrowedMult__comb;
  wire [18:0] p1_smul_27970_NarrowedMult__comb;
  wire [20:0] p1_smul_67671_comb;
  wire [20:0] p1_smul_67674_comb;
  wire [19:0] p1_smul_28010_NarrowedMult__comb;
  wire [19:0] p1_smul_28012_NarrowedMult__comb;
  wire [20:0] p1_smul_67677_comb;
  wire [20:0] p1_smul_67680_comb;
  wire [20:0] p1_smul_67681_comb;
  wire [20:0] p1_smul_67684_comb;
  wire [19:0] p1_smul_28026_NarrowedMult__comb;
  wire [19:0] p1_smul_28028_NarrowedMult__comb;
  wire [20:0] p1_smul_67687_comb;
  wire [20:0] p1_smul_67690_comb;
  wire [20:0] p1_smul_67691_comb;
  wire [20:0] p1_smul_67694_comb;
  wire [19:0] p1_smul_28074_NarrowedMult__comb;
  wire [19:0] p1_smul_28076_NarrowedMult__comb;
  wire [20:0] p1_smul_67697_comb;
  wire [20:0] p1_smul_67700_comb;
  wire [20:0] p1_smul_67701_comb;
  wire [20:0] p1_smul_67704_comb;
  wire [19:0] p1_smul_28090_NarrowedMult__comb;
  wire [19:0] p1_smul_28092_NarrowedMult__comb;
  wire [20:0] p1_smul_67707_comb;
  wire [20:0] p1_smul_67710_comb;
  wire [20:0] p1_smul_67711_comb;
  wire [20:0] p1_smul_67712_comb;
  wire [20:0] p1_smul_67713_comb;
  wire [20:0] p1_smul_67714_comb;
  wire [20:0] p1_smul_67715_comb;
  wire [20:0] p1_smul_67716_comb;
  wire [20:0] p1_smul_67717_comb;
  wire [20:0] p1_smul_67718_comb;
  wire [20:0] p1_smul_67719_comb;
  wire [20:0] p1_smul_67720_comb;
  wire [20:0] p1_smul_67721_comb;
  wire [20:0] p1_smul_67722_comb;
  wire [20:0] p1_smul_67723_comb;
  wire [20:0] p1_smul_67724_comb;
  wire [20:0] p1_smul_67725_comb;
  wire [20:0] p1_smul_67726_comb;
  wire [20:0] p1_smul_67727_comb;
  wire [20:0] p1_smul_67728_comb;
  wire [20:0] p1_smul_67729_comb;
  wire [20:0] p1_smul_67730_comb;
  wire [20:0] p1_smul_67731_comb;
  wire [20:0] p1_smul_67732_comb;
  wire [20:0] p1_smul_67733_comb;
  wire [20:0] p1_smul_67734_comb;
  wire [20:0] p1_smul_67735_comb;
  wire [20:0] p1_smul_67736_comb;
  wire [20:0] p1_smul_67737_comb;
  wire [20:0] p1_smul_67738_comb;
  wire [20:0] p1_smul_67739_comb;
  wire [20:0] p1_smul_67740_comb;
  wire [20:0] p1_smul_67741_comb;
  wire [20:0] p1_smul_67742_comb;
  wire [19:0] p1_smul_28260_NarrowedMult__comb;
  wire [20:0] p1_smul_67744_comb;
  wire [20:0] p1_smul_67747_comb;
  wire [20:0] p1_smul_67748_comb;
  wire [20:0] p1_smul_67751_comb;
  wire [19:0] p1_smul_28274_NarrowedMult__comb;
  wire [19:0] p1_smul_28276_NarrowedMult__comb;
  wire [20:0] p1_smul_67754_comb;
  wire [20:0] p1_smul_67757_comb;
  wire [20:0] p1_smul_67758_comb;
  wire [20:0] p1_smul_67761_comb;
  wire [19:0] p1_smul_28290_NarrowedMult__comb;
  wire [19:0] p1_smul_28324_NarrowedMult__comb;
  wire [20:0] p1_smul_67764_comb;
  wire [20:0] p1_smul_67767_comb;
  wire [20:0] p1_smul_67768_comb;
  wire [20:0] p1_smul_67771_comb;
  wire [19:0] p1_smul_28338_NarrowedMult__comb;
  wire [19:0] p1_smul_28340_NarrowedMult__comb;
  wire [20:0] p1_smul_67774_comb;
  wire [20:0] p1_smul_67777_comb;
  wire [20:0] p1_smul_67778_comb;
  wire [20:0] p1_smul_67781_comb;
  wire [19:0] p1_smul_28354_NarrowedMult__comb;
  wire [18:0] p1_smul_28390_NarrowedMult__comb;
  wire [18:0] p1_smul_28394_NarrowedMult__comb;
  wire [18:0] p1_smul_28396_NarrowedMult__comb;
  wire [18:0] p1_smul_28400_NarrowedMult__comb;
  wire [18:0] p1_smul_28406_NarrowedMult__comb;
  wire [18:0] p1_smul_28410_NarrowedMult__comb;
  wire [18:0] p1_smul_28412_NarrowedMult__comb;
  wire [18:0] p1_smul_28416_NarrowedMult__comb;
  wire [18:0] p1_smul_28454_NarrowedMult__comb;
  wire [18:0] p1_smul_28458_NarrowedMult__comb;
  wire [18:0] p1_smul_28460_NarrowedMult__comb;
  wire [18:0] p1_smul_28464_NarrowedMult__comb;
  wire [18:0] p1_smul_28470_NarrowedMult__comb;
  wire [18:0] p1_smul_28474_NarrowedMult__comb;
  wire [18:0] p1_smul_28476_NarrowedMult__comb;
  wire [18:0] p1_smul_28480_NarrowedMult__comb;
  wire [19:0] p1_smul_28518_NarrowedMult__comb;
  wire [20:0] p1_smul_67834_comb;
  wire [20:0] p1_smul_67835_comb;
  wire [20:0] p1_smul_67836_comb;
  wire [20:0] p1_smul_67837_comb;
  wire [19:0] p1_smul_28528_NarrowedMult__comb;
  wire [19:0] p1_smul_28534_NarrowedMult__comb;
  wire [20:0] p1_smul_67844_comb;
  wire [20:0] p1_smul_67845_comb;
  wire [20:0] p1_smul_67846_comb;
  wire [20:0] p1_smul_67847_comb;
  wire [19:0] p1_smul_28544_NarrowedMult__comb;
  wire [19:0] p1_smul_28582_NarrowedMult__comb;
  wire [20:0] p1_smul_67854_comb;
  wire [20:0] p1_smul_67855_comb;
  wire [20:0] p1_smul_67856_comb;
  wire [20:0] p1_smul_67857_comb;
  wire [19:0] p1_smul_28592_NarrowedMult__comb;
  wire [19:0] p1_smul_28598_NarrowedMult__comb;
  wire [20:0] p1_smul_67864_comb;
  wire [20:0] p1_smul_67865_comb;
  wire [20:0] p1_smul_67866_comb;
  wire [20:0] p1_smul_67867_comb;
  wire [19:0] p1_smul_28608_NarrowedMult__comb;
  wire [20:0] p1_smul_67871_comb;
  wire [20:0] p1_smul_67872_comb;
  wire [19:0] p1_smul_27736_NarrowedMult__comb;
  wire [19:0] p1_smul_27742_NarrowedMult__comb;
  wire [20:0] p1_smul_67879_comb;
  wire [20:0] p1_smul_67880_comb;
  wire [20:0] p1_smul_67881_comb;
  wire [20:0] p1_smul_67882_comb;
  wire [19:0] p1_smul_27848_NarrowedMult__comb;
  wire [19:0] p1_smul_27854_NarrowedMult__comb;
  wire [20:0] p1_smul_67889_comb;
  wire [20:0] p1_smul_67890_comb;
  wire [18:0] p1_smul_27860_NarrowedMult__comb;
  wire [18:0] p1_smul_27866_NarrowedMult__comb;
  wire [18:0] p1_smul_27868_NarrowedMult__comb;
  wire [18:0] p1_smul_27874_NarrowedMult__comb;
  wire [18:0] p1_smul_27972_NarrowedMult__comb;
  wire [18:0] p1_smul_27978_NarrowedMult__comb;
  wire [18:0] p1_smul_27980_NarrowedMult__comb;
  wire [18:0] p1_smul_27986_NarrowedMult__comb;
  wire [20:0] p1_smul_67915_comb;
  wire [20:0] p1_smul_67918_comb;
  wire [19:0] p1_smul_27994_NarrowedMult__comb;
  wire [19:0] p1_smul_27996_NarrowedMult__comb;
  wire [20:0] p1_smul_67921_comb;
  wire [20:0] p1_smul_67924_comb;
  wire [20:0] p1_smul_67925_comb;
  wire [20:0] p1_smul_67928_comb;
  wire [19:0] p1_smul_28106_NarrowedMult__comb;
  wire [19:0] p1_smul_28108_NarrowedMult__comb;
  wire [20:0] p1_smul_67931_comb;
  wire [20:0] p1_smul_67934_comb;
  wire [20:0] p1_smul_67935_comb;
  wire [20:0] p1_smul_67936_comb;
  wire [20:0] p1_smul_67937_comb;
  wire [20:0] p1_smul_67938_comb;
  wire [20:0] p1_smul_67939_comb;
  wire [20:0] p1_smul_67940_comb;
  wire [20:0] p1_smul_67941_comb;
  wire [20:0] p1_smul_67942_comb;
  wire [20:0] p1_smul_67943_comb;
  wire [20:0] p1_smul_67944_comb;
  wire [20:0] p1_smul_67945_comb;
  wire [20:0] p1_smul_67946_comb;
  wire [20:0] p1_smul_67947_comb;
  wire [20:0] p1_smul_67948_comb;
  wire [20:0] p1_smul_67949_comb;
  wire [20:0] p1_smul_67950_comb;
  wire [19:0] p1_smul_28244_NarrowedMult__comb;
  wire [20:0] p1_smul_67952_comb;
  wire [20:0] p1_smul_67955_comb;
  wire [20:0] p1_smul_67956_comb;
  wire [20:0] p1_smul_67959_comb;
  wire [19:0] p1_smul_28258_NarrowedMult__comb;
  wire [19:0] p1_smul_28356_NarrowedMult__comb;
  wire [20:0] p1_smul_67962_comb;
  wire [20:0] p1_smul_67965_comb;
  wire [20:0] p1_smul_67966_comb;
  wire [20:0] p1_smul_67969_comb;
  wire [19:0] p1_smul_28370_NarrowedMult__comb;
  wire [18:0] p1_smul_28374_NarrowedMult__comb;
  wire [18:0] p1_smul_28378_NarrowedMult__comb;
  wire [18:0] p1_smul_28380_NarrowedMult__comb;
  wire [18:0] p1_smul_28384_NarrowedMult__comb;
  wire [18:0] p1_smul_28486_NarrowedMult__comb;
  wire [18:0] p1_smul_28490_NarrowedMult__comb;
  wire [18:0] p1_smul_28492_NarrowedMult__comb;
  wire [18:0] p1_smul_28496_NarrowedMult__comb;
  wire [19:0] p1_smul_28502_NarrowedMult__comb;
  wire [20:0] p1_smul_67998_comb;
  wire [20:0] p1_smul_67999_comb;
  wire [20:0] p1_smul_68000_comb;
  wire [20:0] p1_smul_68001_comb;
  wire [19:0] p1_smul_28512_NarrowedMult__comb;
  wire [19:0] p1_smul_28614_NarrowedMult__comb;
  wire [20:0] p1_smul_68008_comb;
  wire [20:0] p1_smul_68009_comb;
  wire [20:0] p1_smul_68010_comb;
  wire [20:0] p1_smul_68011_comb;
  wire [19:0] p1_smul_28624_NarrowedMult__comb;
  wire [12:0] p1_add_68847_comb;
  wire [12:0] p1_add_68848_comb;
  wire [12:0] p1_add_68849_comb;
  wire [12:0] p1_add_68850_comb;
  wire [12:0] p1_add_68851_comb;
  wire [12:0] p1_add_68852_comb;
  wire [12:0] p1_add_68853_comb;
  wire [12:0] p1_add_68854_comb;
  wire [12:0] p1_add_68967_comb;
  wire [12:0] p1_add_68968_comb;
  wire [12:0] p1_add_68969_comb;
  wire [12:0] p1_add_68970_comb;
  wire [12:0] p1_add_68971_comb;
  wire [12:0] p1_add_68972_comb;
  wire [12:0] p1_add_68973_comb;
  wire [12:0] p1_add_68974_comb;
  wire [12:0] p1_add_68975_comb;
  wire [12:0] p1_add_68976_comb;
  wire [12:0] p1_add_68977_comb;
  wire [12:0] p1_add_68978_comb;
  wire [12:0] p1_add_68979_comb;
  wire [12:0] p1_add_68980_comb;
  wire [12:0] p1_add_68981_comb;
  wire [12:0] p1_add_68982_comb;
  wire [12:0] p1_add_69207_comb;
  wire [12:0] p1_add_69208_comb;
  wire [12:0] p1_add_69209_comb;
  wire [12:0] p1_add_69210_comb;
  wire [12:0] p1_add_69211_comb;
  wire [12:0] p1_add_69212_comb;
  wire [12:0] p1_add_69213_comb;
  wire [12:0] p1_add_69214_comb;
  wire [11:0] p1_add_68037_comb;
  wire [11:0] p1_add_68038_comb;
  wire [11:0] p1_add_68051_comb;
  wire [11:0] p1_add_68052_comb;
  wire [12:0] p1_add_68061_comb;
  wire [12:0] p1_add_68062_comb;
  wire [12:0] p1_add_68067_comb;
  wire [12:0] p1_add_68068_comb;
  wire [12:0] p1_add_68073_comb;
  wire [12:0] p1_add_68074_comb;
  wire [12:0] p1_add_68079_comb;
  wire [12:0] p1_add_68080_comb;
  wire [11:0] p1_add_68085_comb;
  wire [11:0] p1_add_68094_comb;
  wire [11:0] p1_add_68099_comb;
  wire [11:0] p1_add_68108_comb;
  wire [11:0] p1_add_68147_comb;
  wire [11:0] p1_add_68152_comb;
  wire [11:0] p1_add_68161_comb;
  wire [11:0] p1_add_68166_comb;
  wire [12:0] p1_add_68171_comb;
  wire [12:0] p1_add_68174_comb;
  wire [12:0] p1_add_68179_comb;
  wire [12:0] p1_add_68182_comb;
  wire [12:0] p1_add_68183_comb;
  wire [12:0] p1_add_68186_comb;
  wire [12:0] p1_add_68191_comb;
  wire [12:0] p1_add_68194_comb;
  wire [11:0] p1_add_68195_comb;
  wire [11:0] p1_add_68208_comb;
  wire [11:0] p1_add_68209_comb;
  wire [11:0] p1_add_68222_comb;
  wire [11:0] p1_add_68261_comb;
  wire [11:0] p1_add_68262_comb;
  wire [11:0] p1_add_68275_comb;
  wire [11:0] p1_add_68276_comb;
  wire [11:0] p1_add_68289_comb;
  wire [11:0] p1_add_68290_comb;
  wire [11:0] p1_add_68303_comb;
  wire [11:0] p1_add_68304_comb;
  wire [12:0] p1_add_68313_comb;
  wire [12:0] p1_add_68314_comb;
  wire [12:0] p1_add_68319_comb;
  wire [12:0] p1_add_68320_comb;
  wire [12:0] p1_add_68325_comb;
  wire [12:0] p1_add_68326_comb;
  wire [12:0] p1_add_68331_comb;
  wire [12:0] p1_add_68332_comb;
  wire [12:0] p1_add_68337_comb;
  wire [12:0] p1_add_68338_comb;
  wire [12:0] p1_add_68343_comb;
  wire [12:0] p1_add_68344_comb;
  wire [12:0] p1_add_68349_comb;
  wire [12:0] p1_add_68350_comb;
  wire [12:0] p1_add_68355_comb;
  wire [12:0] p1_add_68356_comb;
  wire [11:0] p1_add_68361_comb;
  wire [11:0] p1_add_68370_comb;
  wire [11:0] p1_add_68375_comb;
  wire [11:0] p1_add_68384_comb;
  wire [11:0] p1_add_68389_comb;
  wire [11:0] p1_add_68398_comb;
  wire [11:0] p1_add_68403_comb;
  wire [11:0] p1_add_68412_comb;
  wire [11:0] p1_add_68483_comb;
  wire [11:0] p1_add_68488_comb;
  wire [11:0] p1_add_68497_comb;
  wire [11:0] p1_add_68502_comb;
  wire [11:0] p1_add_68511_comb;
  wire [11:0] p1_add_68516_comb;
  wire [11:0] p1_add_68525_comb;
  wire [11:0] p1_add_68530_comb;
  wire [12:0] p1_add_68535_comb;
  wire [12:0] p1_add_68538_comb;
  wire [12:0] p1_add_68543_comb;
  wire [12:0] p1_add_68546_comb;
  wire [12:0] p1_add_68547_comb;
  wire [12:0] p1_add_68550_comb;
  wire [12:0] p1_add_68555_comb;
  wire [12:0] p1_add_68558_comb;
  wire [12:0] p1_add_68559_comb;
  wire [12:0] p1_add_68562_comb;
  wire [12:0] p1_add_68567_comb;
  wire [12:0] p1_add_68570_comb;
  wire [12:0] p1_add_68571_comb;
  wire [12:0] p1_add_68574_comb;
  wire [12:0] p1_add_68579_comb;
  wire [12:0] p1_add_68582_comb;
  wire [11:0] p1_add_68583_comb;
  wire [11:0] p1_add_68596_comb;
  wire [11:0] p1_add_68597_comb;
  wire [11:0] p1_add_68610_comb;
  wire [11:0] p1_add_68611_comb;
  wire [11:0] p1_add_68624_comb;
  wire [11:0] p1_add_68625_comb;
  wire [11:0] p1_add_68638_comb;
  wire [11:0] p1_add_68661_comb;
  wire [11:0] p1_add_68662_comb;
  wire [11:0] p1_add_68675_comb;
  wire [11:0] p1_add_68676_comb;
  wire [12:0] p1_add_68685_comb;
  wire [12:0] p1_add_68686_comb;
  wire [12:0] p1_add_68691_comb;
  wire [12:0] p1_add_68692_comb;
  wire [12:0] p1_add_68697_comb;
  wire [12:0] p1_add_68698_comb;
  wire [12:0] p1_add_68703_comb;
  wire [12:0] p1_add_68704_comb;
  wire [11:0] p1_add_68709_comb;
  wire [11:0] p1_add_68718_comb;
  wire [11:0] p1_add_68723_comb;
  wire [11:0] p1_add_68732_comb;
  wire [11:0] p1_add_68771_comb;
  wire [11:0] p1_add_68776_comb;
  wire [11:0] p1_add_68785_comb;
  wire [11:0] p1_add_68790_comb;
  wire [12:0] p1_add_68795_comb;
  wire [12:0] p1_add_68798_comb;
  wire [12:0] p1_add_68803_comb;
  wire [12:0] p1_add_68806_comb;
  wire [12:0] p1_add_68807_comb;
  wire [12:0] p1_add_68810_comb;
  wire [12:0] p1_add_68815_comb;
  wire [12:0] p1_add_68818_comb;
  wire [11:0] p1_add_68819_comb;
  wire [11:0] p1_add_68832_comb;
  wire [11:0] p1_add_68833_comb;
  wire [11:0] p1_add_68846_comb;
  wire [31:0] p1_sum__961_comb;
  wire [31:0] p1_sum__962_comb;
  wire [31:0] p1_sum__963_comb;
  wire [31:0] p1_sum__964_comb;
  wire [31:0] p1_sum__926_comb;
  wire [31:0] p1_sum__927_comb;
  wire [31:0] p1_sum__928_comb;
  wire [31:0] p1_sum__929_comb;
  wire [31:0] p1_sum__1010_comb;
  wire [31:0] p1_sum__1011_comb;
  wire [31:0] p1_sum__1012_comb;
  wire [31:0] p1_sum__1013_comb;
  wire [31:0] p1_sum__989_comb;
  wire [31:0] p1_sum__990_comb;
  wire [31:0] p1_sum__991_comb;
  wire [31:0] p1_sum__992_comb;
  wire [31:0] p1_sum__884_comb;
  wire [31:0] p1_sum__885_comb;
  wire [31:0] p1_sum__886_comb;
  wire [31:0] p1_sum__887_comb;
  wire [31:0] p1_sum__835_comb;
  wire [31:0] p1_sum__836_comb;
  wire [31:0] p1_sum__837_comb;
  wire [31:0] p1_sum__838_comb;
  wire [31:0] p1_sum__1017_comb;
  wire [31:0] p1_sum__1018_comb;
  wire [31:0] p1_sum__1019_comb;
  wire [31:0] p1_sum__1020_comb;
  wire [31:0] p1_sum__779_comb;
  wire [31:0] p1_sum__780_comb;
  wire [31:0] p1_sum__781_comb;
  wire [31:0] p1_sum__782_comb;
  wire [13:0] p1_add_68855_comb;
  wire [13:0] p1_add_68856_comb;
  wire [13:0] p1_add_68857_comb;
  wire [10:0] p1_bit_slice_68858_comb;
  wire [10:0] p1_bit_slice_68859_comb;
  wire [13:0] p1_add_68860_comb;
  wire [13:0] p1_add_68861_comb;
  wire [13:0] p1_add_68862_comb;
  wire [13:0] p1_add_68863_comb;
  wire [13:0] p1_add_68864_comb;
  wire [13:0] p1_add_68865_comb;
  wire [10:0] p1_bit_slice_68866_comb;
  wire [10:0] p1_bit_slice_68867_comb;
  wire [13:0] p1_add_68868_comb;
  wire [13:0] p1_add_68869_comb;
  wire [13:0] p1_add_68870_comb;
  wire [13:0] p1_add_68871_comb;
  wire [11:0] p1_bit_slice_68872_comb;
  wire [11:0] p1_bit_slice_68873_comb;
  wire [13:0] p1_add_68874_comb;
  wire [13:0] p1_add_68875_comb;
  wire [11:0] p1_bit_slice_68876_comb;
  wire [11:0] p1_bit_slice_68877_comb;
  wire [13:0] p1_add_68878_comb;
  wire [13:0] p1_add_68879_comb;
  wire [11:0] p1_bit_slice_68880_comb;
  wire [11:0] p1_bit_slice_68881_comb;
  wire [13:0] p1_add_68882_comb;
  wire [13:0] p1_add_68883_comb;
  wire [11:0] p1_bit_slice_68884_comb;
  wire [11:0] p1_bit_slice_68885_comb;
  wire [13:0] p1_add_68886_comb;
  wire [13:0] p1_add_68887_comb;
  wire [10:0] p1_bit_slice_68888_comb;
  wire [13:0] p1_add_68889_comb;
  wire [13:0] p1_add_68890_comb;
  wire [13:0] p1_add_68891_comb;
  wire [13:0] p1_add_68892_comb;
  wire [10:0] p1_bit_slice_68893_comb;
  wire [13:0] p1_add_68894_comb;
  wire [13:0] p1_add_68895_comb;
  wire [10:0] p1_bit_slice_68896_comb;
  wire [13:0] p1_add_68897_comb;
  wire [13:0] p1_add_68898_comb;
  wire [13:0] p1_add_68899_comb;
  wire [13:0] p1_add_68900_comb;
  wire [10:0] p1_bit_slice_68901_comb;
  wire [13:0] p1_add_68902_comb;
  wire [13:0] p1_add_68903_comb;
  wire [13:0] p1_add_68904_comb;
  wire [13:0] p1_add_68905_comb;
  wire [13:0] p1_add_68906_comb;
  wire [13:0] p1_add_68907_comb;
  wire [13:0] p1_add_68908_comb;
  wire [13:0] p1_add_68909_comb;
  wire [13:0] p1_add_68910_comb;
  wire [13:0] p1_add_68911_comb;
  wire [13:0] p1_add_68912_comb;
  wire [13:0] p1_add_68913_comb;
  wire [13:0] p1_add_68914_comb;
  wire [13:0] p1_add_68915_comb;
  wire [13:0] p1_add_68916_comb;
  wire [13:0] p1_add_68917_comb;
  wire [13:0] p1_add_68918_comb;
  wire [13:0] p1_add_68919_comb;
  wire [13:0] p1_add_68920_comb;
  wire [10:0] p1_bit_slice_68921_comb;
  wire [13:0] p1_add_68922_comb;
  wire [13:0] p1_add_68923_comb;
  wire [10:0] p1_bit_slice_68924_comb;
  wire [13:0] p1_add_68925_comb;
  wire [13:0] p1_add_68926_comb;
  wire [13:0] p1_add_68927_comb;
  wire [13:0] p1_add_68928_comb;
  wire [10:0] p1_bit_slice_68929_comb;
  wire [13:0] p1_add_68930_comb;
  wire [13:0] p1_add_68931_comb;
  wire [10:0] p1_bit_slice_68932_comb;
  wire [13:0] p1_add_68933_comb;
  wire [13:0] p1_add_68934_comb;
  wire [11:0] p1_bit_slice_68935_comb;
  wire [13:0] p1_add_68936_comb;
  wire [11:0] p1_bit_slice_68937_comb;
  wire [13:0] p1_add_68938_comb;
  wire [13:0] p1_add_68939_comb;
  wire [11:0] p1_bit_slice_68940_comb;
  wire [13:0] p1_add_68941_comb;
  wire [11:0] p1_bit_slice_68942_comb;
  wire [11:0] p1_bit_slice_68943_comb;
  wire [13:0] p1_add_68944_comb;
  wire [11:0] p1_bit_slice_68945_comb;
  wire [13:0] p1_add_68946_comb;
  wire [13:0] p1_add_68947_comb;
  wire [11:0] p1_bit_slice_68948_comb;
  wire [13:0] p1_add_68949_comb;
  wire [11:0] p1_bit_slice_68950_comb;
  wire [10:0] p1_bit_slice_68951_comb;
  wire [13:0] p1_add_68952_comb;
  wire [13:0] p1_add_68953_comb;
  wire [13:0] p1_add_68954_comb;
  wire [13:0] p1_add_68955_comb;
  wire [13:0] p1_add_68956_comb;
  wire [13:0] p1_add_68957_comb;
  wire [10:0] p1_bit_slice_68958_comb;
  wire [10:0] p1_bit_slice_68959_comb;
  wire [13:0] p1_add_68960_comb;
  wire [13:0] p1_add_68961_comb;
  wire [13:0] p1_add_68962_comb;
  wire [13:0] p1_add_68963_comb;
  wire [13:0] p1_add_68964_comb;
  wire [13:0] p1_add_68965_comb;
  wire [10:0] p1_bit_slice_68966_comb;
  wire [13:0] p1_add_68983_comb;
  wire [13:0] p1_add_68984_comb;
  wire [13:0] p1_add_68985_comb;
  wire [10:0] p1_bit_slice_68986_comb;
  wire [10:0] p1_bit_slice_68987_comb;
  wire [13:0] p1_add_68988_comb;
  wire [13:0] p1_add_68989_comb;
  wire [13:0] p1_add_68990_comb;
  wire [13:0] p1_add_68991_comb;
  wire [13:0] p1_add_68992_comb;
  wire [13:0] p1_add_68993_comb;
  wire [10:0] p1_bit_slice_68994_comb;
  wire [10:0] p1_bit_slice_68995_comb;
  wire [13:0] p1_add_68996_comb;
  wire [13:0] p1_add_68997_comb;
  wire [13:0] p1_add_68998_comb;
  wire [13:0] p1_add_68999_comb;
  wire [13:0] p1_add_69000_comb;
  wire [13:0] p1_add_69001_comb;
  wire [10:0] p1_bit_slice_69002_comb;
  wire [10:0] p1_bit_slice_69003_comb;
  wire [13:0] p1_add_69004_comb;
  wire [13:0] p1_add_69005_comb;
  wire [13:0] p1_add_69006_comb;
  wire [13:0] p1_add_69007_comb;
  wire [13:0] p1_add_69008_comb;
  wire [13:0] p1_add_69009_comb;
  wire [10:0] p1_bit_slice_69010_comb;
  wire [10:0] p1_bit_slice_69011_comb;
  wire [13:0] p1_add_69012_comb;
  wire [13:0] p1_add_69013_comb;
  wire [13:0] p1_add_69014_comb;
  wire [13:0] p1_add_69015_comb;
  wire [11:0] p1_bit_slice_69016_comb;
  wire [11:0] p1_bit_slice_69017_comb;
  wire [13:0] p1_add_69018_comb;
  wire [13:0] p1_add_69019_comb;
  wire [11:0] p1_bit_slice_69020_comb;
  wire [11:0] p1_bit_slice_69021_comb;
  wire [13:0] p1_add_69022_comb;
  wire [13:0] p1_add_69023_comb;
  wire [11:0] p1_bit_slice_69024_comb;
  wire [11:0] p1_bit_slice_69025_comb;
  wire [13:0] p1_add_69026_comb;
  wire [13:0] p1_add_69027_comb;
  wire [11:0] p1_bit_slice_69028_comb;
  wire [11:0] p1_bit_slice_69029_comb;
  wire [13:0] p1_add_69030_comb;
  wire [13:0] p1_add_69031_comb;
  wire [11:0] p1_bit_slice_69032_comb;
  wire [11:0] p1_bit_slice_69033_comb;
  wire [13:0] p1_add_69034_comb;
  wire [13:0] p1_add_69035_comb;
  wire [11:0] p1_bit_slice_69036_comb;
  wire [11:0] p1_bit_slice_69037_comb;
  wire [13:0] p1_add_69038_comb;
  wire [13:0] p1_add_69039_comb;
  wire [11:0] p1_bit_slice_69040_comb;
  wire [11:0] p1_bit_slice_69041_comb;
  wire [13:0] p1_add_69042_comb;
  wire [13:0] p1_add_69043_comb;
  wire [11:0] p1_bit_slice_69044_comb;
  wire [11:0] p1_bit_slice_69045_comb;
  wire [13:0] p1_add_69046_comb;
  wire [13:0] p1_add_69047_comb;
  wire [10:0] p1_bit_slice_69048_comb;
  wire [13:0] p1_add_69049_comb;
  wire [13:0] p1_add_69050_comb;
  wire [13:0] p1_add_69051_comb;
  wire [13:0] p1_add_69052_comb;
  wire [10:0] p1_bit_slice_69053_comb;
  wire [13:0] p1_add_69054_comb;
  wire [13:0] p1_add_69055_comb;
  wire [10:0] p1_bit_slice_69056_comb;
  wire [13:0] p1_add_69057_comb;
  wire [13:0] p1_add_69058_comb;
  wire [13:0] p1_add_69059_comb;
  wire [13:0] p1_add_69060_comb;
  wire [10:0] p1_bit_slice_69061_comb;
  wire [13:0] p1_add_69062_comb;
  wire [13:0] p1_add_69063_comb;
  wire [10:0] p1_bit_slice_69064_comb;
  wire [13:0] p1_add_69065_comb;
  wire [13:0] p1_add_69066_comb;
  wire [13:0] p1_add_69067_comb;
  wire [13:0] p1_add_69068_comb;
  wire [10:0] p1_bit_slice_69069_comb;
  wire [13:0] p1_add_69070_comb;
  wire [13:0] p1_add_69071_comb;
  wire [10:0] p1_bit_slice_69072_comb;
  wire [13:0] p1_add_69073_comb;
  wire [13:0] p1_add_69074_comb;
  wire [13:0] p1_add_69075_comb;
  wire [13:0] p1_add_69076_comb;
  wire [10:0] p1_bit_slice_69077_comb;
  wire [13:0] p1_add_69078_comb;
  wire [13:0] p1_add_69079_comb;
  wire [13:0] p1_add_69080_comb;
  wire [13:0] p1_add_69081_comb;
  wire [13:0] p1_add_69082_comb;
  wire [13:0] p1_add_69083_comb;
  wire [13:0] p1_add_69084_comb;
  wire [13:0] p1_add_69085_comb;
  wire [13:0] p1_add_69086_comb;
  wire [13:0] p1_add_69087_comb;
  wire [13:0] p1_add_69088_comb;
  wire [13:0] p1_add_69089_comb;
  wire [13:0] p1_add_69090_comb;
  wire [13:0] p1_add_69091_comb;
  wire [13:0] p1_add_69092_comb;
  wire [13:0] p1_add_69093_comb;
  wire [13:0] p1_add_69094_comb;
  wire [13:0] p1_add_69095_comb;
  wire [13:0] p1_add_69096_comb;
  wire [13:0] p1_add_69097_comb;
  wire [13:0] p1_add_69098_comb;
  wire [13:0] p1_add_69099_comb;
  wire [13:0] p1_add_69100_comb;
  wire [13:0] p1_add_69101_comb;
  wire [13:0] p1_add_69102_comb;
  wire [13:0] p1_add_69103_comb;
  wire [13:0] p1_add_69104_comb;
  wire [13:0] p1_add_69105_comb;
  wire [13:0] p1_add_69106_comb;
  wire [13:0] p1_add_69107_comb;
  wire [13:0] p1_add_69108_comb;
  wire [13:0] p1_add_69109_comb;
  wire [13:0] p1_add_69110_comb;
  wire [13:0] p1_add_69111_comb;
  wire [13:0] p1_add_69112_comb;
  wire [10:0] p1_bit_slice_69113_comb;
  wire [13:0] p1_add_69114_comb;
  wire [13:0] p1_add_69115_comb;
  wire [10:0] p1_bit_slice_69116_comb;
  wire [13:0] p1_add_69117_comb;
  wire [13:0] p1_add_69118_comb;
  wire [13:0] p1_add_69119_comb;
  wire [13:0] p1_add_69120_comb;
  wire [10:0] p1_bit_slice_69121_comb;
  wire [13:0] p1_add_69122_comb;
  wire [13:0] p1_add_69123_comb;
  wire [10:0] p1_bit_slice_69124_comb;
  wire [13:0] p1_add_69125_comb;
  wire [13:0] p1_add_69126_comb;
  wire [13:0] p1_add_69127_comb;
  wire [13:0] p1_add_69128_comb;
  wire [10:0] p1_bit_slice_69129_comb;
  wire [13:0] p1_add_69130_comb;
  wire [13:0] p1_add_69131_comb;
  wire [10:0] p1_bit_slice_69132_comb;
  wire [13:0] p1_add_69133_comb;
  wire [13:0] p1_add_69134_comb;
  wire [13:0] p1_add_69135_comb;
  wire [13:0] p1_add_69136_comb;
  wire [10:0] p1_bit_slice_69137_comb;
  wire [13:0] p1_add_69138_comb;
  wire [13:0] p1_add_69139_comb;
  wire [10:0] p1_bit_slice_69140_comb;
  wire [13:0] p1_add_69141_comb;
  wire [13:0] p1_add_69142_comb;
  wire [11:0] p1_bit_slice_69143_comb;
  wire [13:0] p1_add_69144_comb;
  wire [11:0] p1_bit_slice_69145_comb;
  wire [13:0] p1_add_69146_comb;
  wire [13:0] p1_add_69147_comb;
  wire [11:0] p1_bit_slice_69148_comb;
  wire [13:0] p1_add_69149_comb;
  wire [11:0] p1_bit_slice_69150_comb;
  wire [11:0] p1_bit_slice_69151_comb;
  wire [13:0] p1_add_69152_comb;
  wire [11:0] p1_bit_slice_69153_comb;
  wire [13:0] p1_add_69154_comb;
  wire [13:0] p1_add_69155_comb;
  wire [11:0] p1_bit_slice_69156_comb;
  wire [13:0] p1_add_69157_comb;
  wire [11:0] p1_bit_slice_69158_comb;
  wire [11:0] p1_bit_slice_69159_comb;
  wire [13:0] p1_add_69160_comb;
  wire [11:0] p1_bit_slice_69161_comb;
  wire [13:0] p1_add_69162_comb;
  wire [13:0] p1_add_69163_comb;
  wire [11:0] p1_bit_slice_69164_comb;
  wire [13:0] p1_add_69165_comb;
  wire [11:0] p1_bit_slice_69166_comb;
  wire [11:0] p1_bit_slice_69167_comb;
  wire [13:0] p1_add_69168_comb;
  wire [11:0] p1_bit_slice_69169_comb;
  wire [13:0] p1_add_69170_comb;
  wire [13:0] p1_add_69171_comb;
  wire [11:0] p1_bit_slice_69172_comb;
  wire [13:0] p1_add_69173_comb;
  wire [11:0] p1_bit_slice_69174_comb;
  wire [10:0] p1_bit_slice_69175_comb;
  wire [13:0] p1_add_69176_comb;
  wire [13:0] p1_add_69177_comb;
  wire [13:0] p1_add_69178_comb;
  wire [13:0] p1_add_69179_comb;
  wire [13:0] p1_add_69180_comb;
  wire [13:0] p1_add_69181_comb;
  wire [10:0] p1_bit_slice_69182_comb;
  wire [10:0] p1_bit_slice_69183_comb;
  wire [13:0] p1_add_69184_comb;
  wire [13:0] p1_add_69185_comb;
  wire [13:0] p1_add_69186_comb;
  wire [13:0] p1_add_69187_comb;
  wire [13:0] p1_add_69188_comb;
  wire [13:0] p1_add_69189_comb;
  wire [10:0] p1_bit_slice_69190_comb;
  wire [10:0] p1_bit_slice_69191_comb;
  wire [13:0] p1_add_69192_comb;
  wire [13:0] p1_add_69193_comb;
  wire [13:0] p1_add_69194_comb;
  wire [13:0] p1_add_69195_comb;
  wire [13:0] p1_add_69196_comb;
  wire [13:0] p1_add_69197_comb;
  wire [10:0] p1_bit_slice_69198_comb;
  wire [10:0] p1_bit_slice_69199_comb;
  wire [13:0] p1_add_69200_comb;
  wire [13:0] p1_add_69201_comb;
  wire [13:0] p1_add_69202_comb;
  wire [13:0] p1_add_69203_comb;
  wire [13:0] p1_add_69204_comb;
  wire [13:0] p1_add_69205_comb;
  wire [10:0] p1_bit_slice_69206_comb;
  wire [13:0] p1_add_69215_comb;
  wire [13:0] p1_add_69216_comb;
  wire [13:0] p1_add_69217_comb;
  wire [10:0] p1_bit_slice_69218_comb;
  wire [10:0] p1_bit_slice_69219_comb;
  wire [13:0] p1_add_69220_comb;
  wire [13:0] p1_add_69221_comb;
  wire [13:0] p1_add_69222_comb;
  wire [13:0] p1_add_69223_comb;
  wire [13:0] p1_add_69224_comb;
  wire [13:0] p1_add_69225_comb;
  wire [10:0] p1_bit_slice_69226_comb;
  wire [10:0] p1_bit_slice_69227_comb;
  wire [13:0] p1_add_69228_comb;
  wire [13:0] p1_add_69229_comb;
  wire [13:0] p1_add_69230_comb;
  wire [13:0] p1_add_69231_comb;
  wire [11:0] p1_bit_slice_69232_comb;
  wire [11:0] p1_bit_slice_69233_comb;
  wire [13:0] p1_add_69234_comb;
  wire [13:0] p1_add_69235_comb;
  wire [11:0] p1_bit_slice_69236_comb;
  wire [11:0] p1_bit_slice_69237_comb;
  wire [13:0] p1_add_69238_comb;
  wire [13:0] p1_add_69239_comb;
  wire [11:0] p1_bit_slice_69240_comb;
  wire [11:0] p1_bit_slice_69241_comb;
  wire [13:0] p1_add_69242_comb;
  wire [13:0] p1_add_69243_comb;
  wire [11:0] p1_bit_slice_69244_comb;
  wire [11:0] p1_bit_slice_69245_comb;
  wire [13:0] p1_add_69246_comb;
  wire [13:0] p1_add_69247_comb;
  wire [10:0] p1_bit_slice_69248_comb;
  wire [13:0] p1_add_69249_comb;
  wire [13:0] p1_add_69250_comb;
  wire [13:0] p1_add_69251_comb;
  wire [13:0] p1_add_69252_comb;
  wire [10:0] p1_bit_slice_69253_comb;
  wire [13:0] p1_add_69254_comb;
  wire [13:0] p1_add_69255_comb;
  wire [10:0] p1_bit_slice_69256_comb;
  wire [13:0] p1_add_69257_comb;
  wire [13:0] p1_add_69258_comb;
  wire [13:0] p1_add_69259_comb;
  wire [13:0] p1_add_69260_comb;
  wire [10:0] p1_bit_slice_69261_comb;
  wire [13:0] p1_add_69262_comb;
  wire [13:0] p1_add_69263_comb;
  wire [13:0] p1_add_69264_comb;
  wire [13:0] p1_add_69265_comb;
  wire [13:0] p1_add_69266_comb;
  wire [13:0] p1_add_69267_comb;
  wire [13:0] p1_add_69268_comb;
  wire [13:0] p1_add_69269_comb;
  wire [13:0] p1_add_69270_comb;
  wire [13:0] p1_add_69271_comb;
  wire [13:0] p1_add_69272_comb;
  wire [13:0] p1_add_69273_comb;
  wire [13:0] p1_add_69274_comb;
  wire [13:0] p1_add_69275_comb;
  wire [13:0] p1_add_69276_comb;
  wire [13:0] p1_add_69277_comb;
  wire [13:0] p1_add_69278_comb;
  wire [13:0] p1_add_69279_comb;
  wire [13:0] p1_add_69280_comb;
  wire [10:0] p1_bit_slice_69281_comb;
  wire [13:0] p1_add_69282_comb;
  wire [13:0] p1_add_69283_comb;
  wire [10:0] p1_bit_slice_69284_comb;
  wire [13:0] p1_add_69285_comb;
  wire [13:0] p1_add_69286_comb;
  wire [13:0] p1_add_69287_comb;
  wire [13:0] p1_add_69288_comb;
  wire [10:0] p1_bit_slice_69289_comb;
  wire [13:0] p1_add_69290_comb;
  wire [13:0] p1_add_69291_comb;
  wire [10:0] p1_bit_slice_69292_comb;
  wire [13:0] p1_add_69293_comb;
  wire [13:0] p1_add_69294_comb;
  wire [11:0] p1_bit_slice_69295_comb;
  wire [13:0] p1_add_69296_comb;
  wire [11:0] p1_bit_slice_69297_comb;
  wire [13:0] p1_add_69298_comb;
  wire [13:0] p1_add_69299_comb;
  wire [11:0] p1_bit_slice_69300_comb;
  wire [13:0] p1_add_69301_comb;
  wire [11:0] p1_bit_slice_69302_comb;
  wire [11:0] p1_bit_slice_69303_comb;
  wire [13:0] p1_add_69304_comb;
  wire [11:0] p1_bit_slice_69305_comb;
  wire [13:0] p1_add_69306_comb;
  wire [13:0] p1_add_69307_comb;
  wire [11:0] p1_bit_slice_69308_comb;
  wire [13:0] p1_add_69309_comb;
  wire [11:0] p1_bit_slice_69310_comb;
  wire [10:0] p1_bit_slice_69311_comb;
  wire [13:0] p1_add_69312_comb;
  wire [13:0] p1_add_69313_comb;
  wire [13:0] p1_add_69314_comb;
  wire [13:0] p1_add_69315_comb;
  wire [13:0] p1_add_69316_comb;
  wire [13:0] p1_add_69317_comb;
  wire [10:0] p1_bit_slice_69318_comb;
  wire [10:0] p1_bit_slice_69319_comb;
  wire [13:0] p1_add_69320_comb;
  wire [13:0] p1_add_69321_comb;
  wire [13:0] p1_add_69322_comb;
  wire [13:0] p1_add_69323_comb;
  wire [13:0] p1_add_69324_comb;
  wire [13:0] p1_add_69325_comb;
  wire [10:0] p1_bit_slice_69326_comb;
  wire [31:0] p1_sum__965_comb;
  wire [31:0] p1_sum__966_comb;
  wire [31:0] p1_sum__930_comb;
  wire [31:0] p1_sum__931_comb;
  wire [31:0] p1_sum__1014_comb;
  wire [31:0] p1_sum__1015_comb;
  wire [31:0] p1_sum__993_comb;
  wire [31:0] p1_sum__994_comb;
  wire [31:0] p1_sum__888_comb;
  wire [31:0] p1_sum__889_comb;
  wire [31:0] p1_sum__839_comb;
  wire [31:0] p1_sum__840_comb;
  wire [31:0] p1_sum__1021_comb;
  wire [31:0] p1_sum__1022_comb;
  wire [31:0] p1_sum__783_comb;
  wire [31:0] p1_sum__784_comb;
  wire [31:0] p1_sum__967_comb;
  wire [31:0] p1_sum__932_comb;
  wire [31:0] p1_sum__1016_comb;
  wire [31:0] p1_sum__995_comb;
  wire [31:0] p1_sum__890_comb;
  wire [31:0] p1_sum__841_comb;
  wire [31:0] p1_sum__1023_comb;
  wire [31:0] p1_sum__785_comb;
  wire [12:0] p1_add_69811_comb;
  wire [12:0] p1_add_69812_comb;
  wire [12:0] p1_add_69813_comb;
  wire [12:0] p1_add_69814_comb;
  wire [12:0] p1_add_69815_comb;
  wire [12:0] p1_add_69816_comb;
  wire [12:0] p1_add_69817_comb;
  wire [12:0] p1_add_69818_comb;
  wire [12:0] p1_add_69819_comb;
  wire [12:0] p1_add_69820_comb;
  wire [12:0] p1_add_69821_comb;
  wire [12:0] p1_add_69822_comb;
  wire [12:0] p1_add_69823_comb;
  wire [12:0] p1_add_69824_comb;
  wire [12:0] p1_add_69825_comb;
  wire [12:0] p1_add_69826_comb;
  wire [12:0] p1_add_69827_comb;
  wire [12:0] p1_add_69828_comb;
  wire [12:0] p1_add_69829_comb;
  wire [12:0] p1_add_69830_comb;
  wire [12:0] p1_add_69831_comb;
  wire [12:0] p1_add_69832_comb;
  wire [12:0] p1_add_69833_comb;
  wire [12:0] p1_add_69834_comb;
  wire [12:0] p1_add_69835_comb;
  wire [12:0] p1_add_69836_comb;
  wire [12:0] p1_add_69837_comb;
  wire [12:0] p1_add_69838_comb;
  wire [12:0] p1_add_69839_comb;
  wire [12:0] p1_add_69840_comb;
  wire [12:0] p1_add_69841_comb;
  wire [12:0] p1_add_69842_comb;
  wire [12:0] p1_add_69843_comb;
  wire [12:0] p1_add_69844_comb;
  wire [12:0] p1_add_69845_comb;
  wire [12:0] p1_add_69846_comb;
  wire [12:0] p1_add_69847_comb;
  wire [12:0] p1_add_69848_comb;
  wire [12:0] p1_add_69849_comb;
  wire [12:0] p1_add_69850_comb;
  wire [12:0] p1_add_69851_comb;
  wire [12:0] p1_add_69852_comb;
  wire [12:0] p1_add_69853_comb;
  wire [12:0] p1_add_69854_comb;
  wire [12:0] p1_add_69855_comb;
  wire [12:0] p1_add_69856_comb;
  wire [12:0] p1_add_69857_comb;
  wire [12:0] p1_add_69858_comb;
  wire [12:0] p1_add_69859_comb;
  wire [12:0] p1_add_69860_comb;
  wire [12:0] p1_add_69861_comb;
  wire [12:0] p1_add_69862_comb;
  wire [12:0] p1_add_69863_comb;
  wire [12:0] p1_add_69864_comb;
  wire [12:0] p1_add_69865_comb;
  wire [12:0] p1_add_69866_comb;
  wire [12:0] p1_add_69875_comb;
  wire [12:0] p1_add_69876_comb;
  wire [12:0] p1_add_69877_comb;
  wire [12:0] p1_add_69878_comb;
  wire [12:0] p1_add_69879_comb;
  wire [12:0] p1_add_69880_comb;
  wire [12:0] p1_add_69881_comb;
  wire [12:0] p1_add_69882_comb;
  wire [12:0] p1_add_69883_comb;
  wire [12:0] p1_add_69884_comb;
  wire [12:0] p1_add_69885_comb;
  wire [12:0] p1_add_69886_comb;
  wire [12:0] p1_add_69887_comb;
  wire [12:0] p1_add_69888_comb;
  wire [12:0] p1_add_69889_comb;
  wire [12:0] p1_add_69890_comb;
  wire [12:0] p1_add_69891_comb;
  wire [12:0] p1_add_69892_comb;
  wire [12:0] p1_add_69893_comb;
  wire [12:0] p1_add_69894_comb;
  wire [12:0] p1_add_69895_comb;
  wire [12:0] p1_add_69896_comb;
  wire [12:0] p1_add_69897_comb;
  wire [12:0] p1_add_69898_comb;
  wire [12:0] p1_add_69899_comb;
  wire [12:0] p1_add_69900_comb;
  wire [12:0] p1_add_69901_comb;
  wire [12:0] p1_add_69902_comb;
  wire [12:0] p1_add_69903_comb;
  wire [12:0] p1_add_69904_comb;
  wire [12:0] p1_add_69905_comb;
  wire [12:0] p1_add_69906_comb;
  wire [12:0] p1_add_69907_comb;
  wire [12:0] p1_add_69908_comb;
  wire [12:0] p1_add_69909_comb;
  wire [12:0] p1_add_69910_comb;
  wire [12:0] p1_add_69911_comb;
  wire [12:0] p1_add_69912_comb;
  wire [12:0] p1_add_69913_comb;
  wire [12:0] p1_add_69914_comb;
  wire [12:0] p1_add_69915_comb;
  wire [12:0] p1_add_69916_comb;
  wire [12:0] p1_add_69917_comb;
  wire [12:0] p1_add_69918_comb;
  wire [12:0] p1_add_69919_comb;
  wire [12:0] p1_add_69920_comb;
  wire [12:0] p1_add_69921_comb;
  wire [12:0] p1_add_69922_comb;
  wire [12:0] p1_add_69923_comb;
  wire [12:0] p1_add_69924_comb;
  wire [12:0] p1_add_69925_comb;
  wire [12:0] p1_add_69926_comb;
  wire [12:0] p1_add_69927_comb;
  wire [12:0] p1_add_69928_comb;
  wire [12:0] p1_add_69929_comb;
  wire [12:0] p1_add_69930_comb;
  wire [12:0] p1_add_69931_comb;
  wire [12:0] p1_add_69932_comb;
  wire [12:0] p1_add_69933_comb;
  wire [12:0] p1_add_69934_comb;
  wire [12:0] p1_add_69935_comb;
  wire [12:0] p1_add_69936_comb;
  wire [12:0] p1_add_69937_comb;
  wire [12:0] p1_add_69938_comb;
  wire [12:0] p1_add_69939_comb;
  wire [12:0] p1_add_69940_comb;
  wire [12:0] p1_add_69941_comb;
  wire [12:0] p1_add_69942_comb;
  wire [12:0] p1_add_69943_comb;
  wire [12:0] p1_add_69944_comb;
  wire [12:0] p1_add_69945_comb;
  wire [12:0] p1_add_69946_comb;
  wire [12:0] p1_add_69947_comb;
  wire [12:0] p1_add_69948_comb;
  wire [12:0] p1_add_69949_comb;
  wire [12:0] p1_add_69950_comb;
  wire [12:0] p1_add_69951_comb;
  wire [12:0] p1_add_69952_comb;
  wire [12:0] p1_add_69953_comb;
  wire [12:0] p1_add_69954_comb;
  wire [12:0] p1_add_69955_comb;
  wire [12:0] p1_add_69956_comb;
  wire [12:0] p1_add_69957_comb;
  wire [12:0] p1_add_69958_comb;
  wire [12:0] p1_add_69959_comb;
  wire [12:0] p1_add_69960_comb;
  wire [12:0] p1_add_69961_comb;
  wire [12:0] p1_add_69962_comb;
  wire [12:0] p1_add_69963_comb;
  wire [12:0] p1_add_69964_comb;
  wire [12:0] p1_add_69965_comb;
  wire [12:0] p1_add_69966_comb;
  wire [12:0] p1_add_69967_comb;
  wire [12:0] p1_add_69968_comb;
  wire [12:0] p1_add_69969_comb;
  wire [12:0] p1_add_69970_comb;
  wire [12:0] p1_add_69971_comb;
  wire [12:0] p1_add_69972_comb;
  wire [12:0] p1_add_69973_comb;
  wire [12:0] p1_add_69974_comb;
  wire [12:0] p1_add_69975_comb;
  wire [12:0] p1_add_69976_comb;
  wire [12:0] p1_add_69977_comb;
  wire [12:0] p1_add_69978_comb;
  wire [12:0] p1_add_69979_comb;
  wire [12:0] p1_add_69980_comb;
  wire [12:0] p1_add_69981_comb;
  wire [12:0] p1_add_69982_comb;
  wire [12:0] p1_add_69983_comb;
  wire [12:0] p1_add_69984_comb;
  wire [12:0] p1_add_69985_comb;
  wire [12:0] p1_add_69986_comb;
  wire [12:0] p1_add_69991_comb;
  wire [12:0] p1_add_69992_comb;
  wire [12:0] p1_add_69993_comb;
  wire [12:0] p1_add_69994_comb;
  wire [12:0] p1_add_69995_comb;
  wire [12:0] p1_add_69996_comb;
  wire [12:0] p1_add_69997_comb;
  wire [12:0] p1_add_69998_comb;
  wire [12:0] p1_add_69999_comb;
  wire [12:0] p1_add_70000_comb;
  wire [12:0] p1_add_70001_comb;
  wire [12:0] p1_add_70002_comb;
  wire [12:0] p1_add_70003_comb;
  wire [12:0] p1_add_70004_comb;
  wire [12:0] p1_add_70005_comb;
  wire [12:0] p1_add_70006_comb;
  wire [12:0] p1_add_70007_comb;
  wire [12:0] p1_add_70008_comb;
  wire [12:0] p1_add_70009_comb;
  wire [12:0] p1_add_70010_comb;
  wire [12:0] p1_add_70011_comb;
  wire [12:0] p1_add_70012_comb;
  wire [12:0] p1_add_70013_comb;
  wire [12:0] p1_add_70014_comb;
  wire [12:0] p1_add_70015_comb;
  wire [12:0] p1_add_70016_comb;
  wire [12:0] p1_add_70017_comb;
  wire [12:0] p1_add_70018_comb;
  wire [12:0] p1_add_70019_comb;
  wire [12:0] p1_add_70020_comb;
  wire [12:0] p1_add_70021_comb;
  wire [12:0] p1_add_70022_comb;
  wire [12:0] p1_add_70023_comb;
  wire [12:0] p1_add_70024_comb;
  wire [12:0] p1_add_70025_comb;
  wire [12:0] p1_add_70026_comb;
  wire [12:0] p1_add_70027_comb;
  wire [12:0] p1_add_70028_comb;
  wire [12:0] p1_add_70029_comb;
  wire [12:0] p1_add_70030_comb;
  wire [12:0] p1_add_70031_comb;
  wire [12:0] p1_add_70032_comb;
  wire [12:0] p1_add_70033_comb;
  wire [12:0] p1_add_70034_comb;
  wire [12:0] p1_add_70035_comb;
  wire [12:0] p1_add_70036_comb;
  wire [12:0] p1_add_70037_comb;
  wire [12:0] p1_add_70038_comb;
  wire [12:0] p1_add_70039_comb;
  wire [12:0] p1_add_70040_comb;
  wire [12:0] p1_add_70041_comb;
  wire [12:0] p1_add_70042_comb;
  wire [12:0] p1_add_70043_comb;
  wire [12:0] p1_add_70044_comb;
  wire [12:0] p1_add_70045_comb;
  wire [12:0] p1_add_70046_comb;
  wire [31:0] p1_umul_70287_comb;
  wire [31:0] p1_umul_70288_comb;
  wire [31:0] p1_umul_70317_comb;
  wire [31:0] p1_umul_70318_comb;
  wire [31:0] p1_umul_70319_comb;
  wire [31:0] p1_umul_70320_comb;
  wire [31:0] p1_umul_70377_comb;
  wire [31:0] p1_umul_70378_comb;
  wire [24:0] p1_sum__1768_comb;
  wire [24:0] p1_sum__1769_comb;
  wire [24:0] p1_sum__1770_comb;
  wire [24:0] p1_sum__1771_comb;
  wire [24:0] p1_sum__1748_comb;
  wire [24:0] p1_sum__1749_comb;
  wire [24:0] p1_sum__1750_comb;
  wire [24:0] p1_sum__1751_comb;
  wire [24:0] p1_sum__1752_comb;
  wire [24:0] p1_sum__1753_comb;
  wire [24:0] p1_sum__1754_comb;
  wire [24:0] p1_sum__1755_comb;
  wire [24:0] p1_sum__1728_comb;
  wire [24:0] p1_sum__1729_comb;
  wire [24:0] p1_sum__1730_comb;
  wire [24:0] p1_sum__1731_comb;
  wire [24:0] p1_sum__1732_comb;
  wire [24:0] p1_sum__1733_comb;
  wire [24:0] p1_sum__1734_comb;
  wire [24:0] p1_sum__1735_comb;
  wire [24:0] p1_sum__1704_comb;
  wire [24:0] p1_sum__1705_comb;
  wire [24:0] p1_sum__1706_comb;
  wire [24:0] p1_sum__1707_comb;
  wire [24:0] p1_sum__1708_comb;
  wire [24:0] p1_sum__1709_comb;
  wire [24:0] p1_sum__1710_comb;
  wire [24:0] p1_sum__1711_comb;
  wire [24:0] p1_sum__1680_comb;
  wire [24:0] p1_sum__1681_comb;
  wire [24:0] p1_sum__1682_comb;
  wire [24:0] p1_sum__1683_comb;
  wire [24:0] p1_sum__1684_comb;
  wire [24:0] p1_sum__1685_comb;
  wire [24:0] p1_sum__1686_comb;
  wire [24:0] p1_sum__1687_comb;
  wire [24:0] p1_sum__1656_comb;
  wire [24:0] p1_sum__1657_comb;
  wire [24:0] p1_sum__1658_comb;
  wire [24:0] p1_sum__1659_comb;
  wire [24:0] p1_sum__1660_comb;
  wire [24:0] p1_sum__1661_comb;
  wire [24:0] p1_sum__1662_comb;
  wire [24:0] p1_sum__1663_comb;
  wire [24:0] p1_sum__1636_comb;
  wire [24:0] p1_sum__1637_comb;
  wire [24:0] p1_sum__1638_comb;
  wire [24:0] p1_sum__1639_comb;
  wire [24:0] p1_sum__1640_comb;
  wire [24:0] p1_sum__1641_comb;
  wire [24:0] p1_sum__1642_comb;
  wire [24:0] p1_sum__1643_comb;
  wire [24:0] p1_sum__1620_comb;
  wire [24:0] p1_sum__1621_comb;
  wire [24:0] p1_sum__1622_comb;
  wire [24:0] p1_sum__1623_comb;
  wire [24:0] p1_sum__1796_comb;
  wire [24:0] p1_sum__1797_comb;
  wire [24:0] p1_sum__1798_comb;
  wire [24:0] p1_sum__1799_comb;
  wire [24:0] p1_sum__1784_comb;
  wire [24:0] p1_sum__1785_comb;
  wire [24:0] p1_sum__1786_comb;
  wire [24:0] p1_sum__1787_comb;
  wire [24:0] p1_sum__1724_comb;
  wire [24:0] p1_sum__1725_comb;
  wire [24:0] p1_sum__1726_comb;
  wire [24:0] p1_sum__1727_comb;
  wire [24:0] p1_sum__1696_comb;
  wire [24:0] p1_sum__1697_comb;
  wire [24:0] p1_sum__1698_comb;
  wire [24:0] p1_sum__1699_comb;
  wire [24:0] p1_sum__1788_comb;
  wire [24:0] p1_sum__1789_comb;
  wire [24:0] p1_sum__1790_comb;
  wire [24:0] p1_sum__1791_comb;
  wire [24:0] p1_sum__1772_comb;
  wire [24:0] p1_sum__1773_comb;
  wire [24:0] p1_sum__1774_comb;
  wire [24:0] p1_sum__1775_comb;
  wire [24:0] p1_sum__1700_comb;
  wire [24:0] p1_sum__1701_comb;
  wire [24:0] p1_sum__1702_comb;
  wire [24:0] p1_sum__1703_comb;
  wire [24:0] p1_sum__1672_comb;
  wire [24:0] p1_sum__1673_comb;
  wire [24:0] p1_sum__1674_comb;
  wire [24:0] p1_sum__1675_comb;
  wire [24:0] p1_sum__1776_comb;
  wire [24:0] p1_sum__1777_comb;
  wire [24:0] p1_sum__1778_comb;
  wire [24:0] p1_sum__1779_comb;
  wire [24:0] p1_sum__1756_comb;
  wire [24:0] p1_sum__1757_comb;
  wire [24:0] p1_sum__1758_comb;
  wire [24:0] p1_sum__1759_comb;
  wire [24:0] p1_sum__1676_comb;
  wire [24:0] p1_sum__1677_comb;
  wire [24:0] p1_sum__1678_comb;
  wire [24:0] p1_sum__1679_comb;
  wire [24:0] p1_sum__1648_comb;
  wire [24:0] p1_sum__1649_comb;
  wire [24:0] p1_sum__1650_comb;
  wire [24:0] p1_sum__1651_comb;
  wire [24:0] p1_sum__1760_comb;
  wire [24:0] p1_sum__1761_comb;
  wire [24:0] p1_sum__1762_comb;
  wire [24:0] p1_sum__1763_comb;
  wire [24:0] p1_sum__1736_comb;
  wire [24:0] p1_sum__1737_comb;
  wire [24:0] p1_sum__1738_comb;
  wire [24:0] p1_sum__1739_comb;
  wire [24:0] p1_sum__1652_comb;
  wire [24:0] p1_sum__1653_comb;
  wire [24:0] p1_sum__1654_comb;
  wire [24:0] p1_sum__1655_comb;
  wire [24:0] p1_sum__1628_comb;
  wire [24:0] p1_sum__1629_comb;
  wire [24:0] p1_sum__1630_comb;
  wire [24:0] p1_sum__1631_comb;
  wire [24:0] p1_sum__1740_comb;
  wire [24:0] p1_sum__1741_comb;
  wire [24:0] p1_sum__1742_comb;
  wire [24:0] p1_sum__1743_comb;
  wire [24:0] p1_sum__1712_comb;
  wire [24:0] p1_sum__1713_comb;
  wire [24:0] p1_sum__1714_comb;
  wire [24:0] p1_sum__1715_comb;
  wire [24:0] p1_sum__1632_comb;
  wire [24:0] p1_sum__1633_comb;
  wire [24:0] p1_sum__1634_comb;
  wire [24:0] p1_sum__1635_comb;
  wire [24:0] p1_sum__1612_comb;
  wire [24:0] p1_sum__1613_comb;
  wire [24:0] p1_sum__1614_comb;
  wire [24:0] p1_sum__1615_comb;
  wire [24:0] p1_sum__1716_comb;
  wire [24:0] p1_sum__1717_comb;
  wire [24:0] p1_sum__1718_comb;
  wire [24:0] p1_sum__1719_comb;
  wire [24:0] p1_sum__1688_comb;
  wire [24:0] p1_sum__1689_comb;
  wire [24:0] p1_sum__1690_comb;
  wire [24:0] p1_sum__1691_comb;
  wire [24:0] p1_sum__1616_comb;
  wire [24:0] p1_sum__1617_comb;
  wire [24:0] p1_sum__1618_comb;
  wire [24:0] p1_sum__1619_comb;
  wire [24:0] p1_sum__1600_comb;
  wire [24:0] p1_sum__1601_comb;
  wire [24:0] p1_sum__1602_comb;
  wire [24:0] p1_sum__1603_comb;
  wire [24:0] p1_sum__1692_comb;
  wire [24:0] p1_sum__1693_comb;
  wire [24:0] p1_sum__1694_comb;
  wire [24:0] p1_sum__1695_comb;
  wire [24:0] p1_sum__1664_comb;
  wire [24:0] p1_sum__1665_comb;
  wire [24:0] p1_sum__1666_comb;
  wire [24:0] p1_sum__1667_comb;
  wire [24:0] p1_sum__1604_comb;
  wire [24:0] p1_sum__1605_comb;
  wire [24:0] p1_sum__1606_comb;
  wire [24:0] p1_sum__1607_comb;
  wire [24:0] p1_sum__1592_comb;
  wire [24:0] p1_sum__1593_comb;
  wire [24:0] p1_sum__1594_comb;
  wire [24:0] p1_sum__1595_comb;
  wire [24:0] p1_sum__1804_comb;
  wire [24:0] p1_sum__1805_comb;
  wire [24:0] p1_sum__1806_comb;
  wire [24:0] p1_sum__1807_comb;
  wire [24:0] p1_sum__1668_comb;
  wire [24:0] p1_sum__1669_comb;
  wire [24:0] p1_sum__1670_comb;
  wire [24:0] p1_sum__1671_comb;
  wire [24:0] p1_sum__1800_comb;
  wire [24:0] p1_sum__1801_comb;
  wire [24:0] p1_sum__1802_comb;
  wire [24:0] p1_sum__1803_comb;
  wire [24:0] p1_sum__1644_comb;
  wire [24:0] p1_sum__1645_comb;
  wire [24:0] p1_sum__1646_comb;
  wire [24:0] p1_sum__1647_comb;
  wire [24:0] p1_sum__1792_comb;
  wire [24:0] p1_sum__1793_comb;
  wire [24:0] p1_sum__1794_comb;
  wire [24:0] p1_sum__1795_comb;
  wire [24:0] p1_sum__1624_comb;
  wire [24:0] p1_sum__1625_comb;
  wire [24:0] p1_sum__1626_comb;
  wire [24:0] p1_sum__1627_comb;
  wire [24:0] p1_sum__1780_comb;
  wire [24:0] p1_sum__1781_comb;
  wire [24:0] p1_sum__1782_comb;
  wire [24:0] p1_sum__1783_comb;
  wire [24:0] p1_sum__1608_comb;
  wire [24:0] p1_sum__1609_comb;
  wire [24:0] p1_sum__1610_comb;
  wire [24:0] p1_sum__1611_comb;
  wire [24:0] p1_sum__1764_comb;
  wire [24:0] p1_sum__1765_comb;
  wire [24:0] p1_sum__1766_comb;
  wire [24:0] p1_sum__1767_comb;
  wire [24:0] p1_sum__1596_comb;
  wire [24:0] p1_sum__1597_comb;
  wire [24:0] p1_sum__1598_comb;
  wire [24:0] p1_sum__1599_comb;
  wire [24:0] p1_sum__1744_comb;
  wire [24:0] p1_sum__1745_comb;
  wire [24:0] p1_sum__1746_comb;
  wire [24:0] p1_sum__1747_comb;
  wire [24:0] p1_sum__1588_comb;
  wire [24:0] p1_sum__1589_comb;
  wire [24:0] p1_sum__1590_comb;
  wire [24:0] p1_sum__1591_comb;
  wire [24:0] p1_sum__1720_comb;
  wire [24:0] p1_sum__1721_comb;
  wire [24:0] p1_sum__1722_comb;
  wire [24:0] p1_sum__1723_comb;
  wire [24:0] p1_sum__1584_comb;
  wire [24:0] p1_sum__1585_comb;
  wire [24:0] p1_sum__1586_comb;
  wire [24:0] p1_sum__1587_comb;
  wire [24:0] p1_sum__1340_comb;
  wire [24:0] p1_sum__1341_comb;
  wire [24:0] p1_sum__1330_comb;
  wire [24:0] p1_sum__1331_comb;
  wire [24:0] p1_sum__1332_comb;
  wire [24:0] p1_sum__1333_comb;
  wire [24:0] p1_sum__1320_comb;
  wire [24:0] p1_sum__1321_comb;
  wire [24:0] p1_sum__1322_comb;
  wire [24:0] p1_sum__1323_comb;
  wire [24:0] p1_sum__1308_comb;
  wire [24:0] p1_sum__1309_comb;
  wire [24:0] p1_sum__1310_comb;
  wire [24:0] p1_sum__1311_comb;
  wire [24:0] p1_sum__1296_comb;
  wire [24:0] p1_sum__1297_comb;
  wire [24:0] p1_sum__1298_comb;
  wire [24:0] p1_sum__1299_comb;
  wire [24:0] p1_sum__1284_comb;
  wire [24:0] p1_sum__1285_comb;
  wire [24:0] p1_sum__1286_comb;
  wire [24:0] p1_sum__1287_comb;
  wire [24:0] p1_sum__1274_comb;
  wire [24:0] p1_sum__1275_comb;
  wire [24:0] p1_sum__1276_comb;
  wire [24:0] p1_sum__1277_comb;
  wire [24:0] p1_sum__1266_comb;
  wire [24:0] p1_sum__1267_comb;
  wire [24:0] p1_sum__1354_comb;
  wire [24:0] p1_sum__1355_comb;
  wire [24:0] p1_sum__1348_comb;
  wire [24:0] p1_sum__1349_comb;
  wire [24:0] p1_sum__1318_comb;
  wire [24:0] p1_sum__1319_comb;
  wire [24:0] p1_sum__1304_comb;
  wire [24:0] p1_sum__1305_comb;
  wire [24:0] p1_sum__1350_comb;
  wire [24:0] p1_sum__1351_comb;
  wire [24:0] p1_sum__1342_comb;
  wire [24:0] p1_sum__1343_comb;
  wire [24:0] p1_sum__1306_comb;
  wire [24:0] p1_sum__1307_comb;
  wire [24:0] p1_sum__1292_comb;
  wire [24:0] p1_sum__1293_comb;
  wire [24:0] p1_sum__1344_comb;
  wire [24:0] p1_sum__1345_comb;
  wire [24:0] p1_sum__1334_comb;
  wire [24:0] p1_sum__1335_comb;
  wire [24:0] p1_sum__1294_comb;
  wire [24:0] p1_sum__1295_comb;
  wire [24:0] p1_sum__1280_comb;
  wire [24:0] p1_sum__1281_comb;
  wire [24:0] p1_sum__1336_comb;
  wire [24:0] p1_sum__1337_comb;
  wire [24:0] p1_sum__1324_comb;
  wire [24:0] p1_sum__1325_comb;
  wire [24:0] p1_sum__1282_comb;
  wire [24:0] p1_sum__1283_comb;
  wire [24:0] p1_sum__1270_comb;
  wire [24:0] p1_sum__1271_comb;
  wire [24:0] p1_sum__1326_comb;
  wire [24:0] p1_sum__1327_comb;
  wire [24:0] p1_sum__1312_comb;
  wire [24:0] p1_sum__1313_comb;
  wire [24:0] p1_sum__1272_comb;
  wire [24:0] p1_sum__1273_comb;
  wire [24:0] p1_sum__1262_comb;
  wire [24:0] p1_sum__1263_comb;
  wire [24:0] p1_sum__1314_comb;
  wire [24:0] p1_sum__1315_comb;
  wire [24:0] p1_sum__1300_comb;
  wire [24:0] p1_sum__1301_comb;
  wire [24:0] p1_sum__1264_comb;
  wire [24:0] p1_sum__1265_comb;
  wire [24:0] p1_sum__1256_comb;
  wire [24:0] p1_sum__1257_comb;
  wire [24:0] p1_sum__1302_comb;
  wire [24:0] p1_sum__1303_comb;
  wire [24:0] p1_sum__1288_comb;
  wire [24:0] p1_sum__1289_comb;
  wire [24:0] p1_sum__1258_comb;
  wire [24:0] p1_sum__1259_comb;
  wire [24:0] p1_sum__1252_comb;
  wire [24:0] p1_sum__1253_comb;
  wire [24:0] p1_sum__1358_comb;
  wire [24:0] p1_sum__1359_comb;
  wire [24:0] p1_sum__1290_comb;
  wire [24:0] p1_sum__1291_comb;
  wire [24:0] p1_sum__1356_comb;
  wire [24:0] p1_sum__1357_comb;
  wire [24:0] p1_sum__1278_comb;
  wire [24:0] p1_sum__1279_comb;
  wire [24:0] p1_sum__1352_comb;
  wire [24:0] p1_sum__1353_comb;
  wire [24:0] p1_sum__1268_comb;
  wire [24:0] p1_sum__1269_comb;
  wire [24:0] p1_sum__1346_comb;
  wire [24:0] p1_sum__1347_comb;
  wire [24:0] p1_sum__1260_comb;
  wire [24:0] p1_sum__1261_comb;
  wire [24:0] p1_sum__1338_comb;
  wire [24:0] p1_sum__1339_comb;
  wire [24:0] p1_sum__1254_comb;
  wire [24:0] p1_sum__1255_comb;
  wire [24:0] p1_sum__1328_comb;
  wire [24:0] p1_sum__1329_comb;
  wire [24:0] p1_sum__1250_comb;
  wire [24:0] p1_sum__1251_comb;
  wire [24:0] p1_sum__1316_comb;
  wire [24:0] p1_sum__1317_comb;
  wire [24:0] p1_sum__1248_comb;
  wire [24:0] p1_sum__1249_comb;
  wire [24:0] p1_add_70535_comb;
  wire [24:0] p1_add_70536_comb;
  wire [24:0] p1_add_70551_comb;
  wire [24:0] p1_add_70552_comb;
  wire [24:0] p1_add_70553_comb;
  wire [24:0] p1_add_70554_comb;
  wire [24:0] p1_add_70583_comb;
  wire [24:0] p1_add_70584_comb;
  wire [24:0] p1_sum__1126_comb;
  wire [24:0] p1_sum__1121_comb;
  wire [24:0] p1_sum__1122_comb;
  wire [24:0] p1_sum__1116_comb;
  wire [24:0] p1_sum__1117_comb;
  wire [24:0] p1_sum__1110_comb;
  wire [24:0] p1_sum__1111_comb;
  wire [24:0] p1_sum__1104_comb;
  wire [24:0] p1_sum__1105_comb;
  wire [24:0] p1_sum__1098_comb;
  wire [24:0] p1_sum__1099_comb;
  wire [24:0] p1_sum__1093_comb;
  wire [24:0] p1_sum__1094_comb;
  wire [24:0] p1_sum__1089_comb;
  wire [24:0] p1_sum__1133_comb;
  wire [24:0] p1_sum__1130_comb;
  wire [24:0] p1_sum__1115_comb;
  wire [24:0] p1_sum__1108_comb;
  wire [24:0] p1_sum__1131_comb;
  wire [24:0] p1_sum__1127_comb;
  wire [24:0] p1_sum__1109_comb;
  wire [24:0] p1_sum__1102_comb;
  wire [24:0] p1_sum__1128_comb;
  wire [24:0] p1_sum__1123_comb;
  wire [24:0] p1_sum__1103_comb;
  wire [24:0] p1_sum__1096_comb;
  wire [24:0] p1_sum__1124_comb;
  wire [24:0] p1_sum__1118_comb;
  wire [24:0] p1_sum__1097_comb;
  wire [24:0] p1_sum__1091_comb;
  wire [24:0] p1_sum__1119_comb;
  wire [24:0] p1_sum__1112_comb;
  wire [24:0] p1_sum__1092_comb;
  wire [24:0] p1_sum__1087_comb;
  wire [24:0] p1_sum__1113_comb;
  wire [24:0] p1_sum__1106_comb;
  wire [24:0] p1_sum__1088_comb;
  wire [24:0] p1_sum__1084_comb;
  wire [24:0] p1_sum__1107_comb;
  wire [24:0] p1_sum__1100_comb;
  wire [24:0] p1_sum__1085_comb;
  wire [24:0] p1_sum__1082_comb;
  wire [24:0] p1_sum__1135_comb;
  wire [24:0] p1_sum__1101_comb;
  wire [24:0] p1_sum__1134_comb;
  wire [24:0] p1_sum__1095_comb;
  wire [24:0] p1_sum__1132_comb;
  wire [24:0] p1_sum__1090_comb;
  wire [24:0] p1_sum__1129_comb;
  wire [24:0] p1_sum__1086_comb;
  wire [24:0] p1_sum__1125_comb;
  wire [24:0] p1_sum__1083_comb;
  wire [24:0] p1_sum__1120_comb;
  wire [24:0] p1_sum__1081_comb;
  wire [24:0] p1_sum__1114_comb;
  wire [24:0] p1_sum__1080_comb;
  wire [24:0] p1_add_70537_comb;
  wire [24:0] p1_add_70538_comb;
  wire [24:0] p1_add_70539_comb;
  wire [24:0] p1_add_70540_comb;
  wire [24:0] p1_add_70541_comb;
  wire [24:0] p1_add_70542_comb;
  wire [24:0] p1_add_70543_comb;
  wire [24:0] p1_add_70544_comb;
  wire [24:0] p1_add_70545_comb;
  wire [24:0] p1_add_70546_comb;
  wire [24:0] p1_add_70547_comb;
  wire [24:0] p1_add_70548_comb;
  wire [24:0] p1_add_70549_comb;
  wire [24:0] p1_add_70550_comb;
  wire [24:0] p1_add_70555_comb;
  wire [24:0] p1_add_70556_comb;
  wire [24:0] p1_add_70557_comb;
  wire [24:0] p1_add_70558_comb;
  wire [24:0] p1_add_70559_comb;
  wire [24:0] p1_add_70560_comb;
  wire [24:0] p1_add_70561_comb;
  wire [24:0] p1_add_70562_comb;
  wire [24:0] p1_add_70563_comb;
  wire [24:0] p1_add_70564_comb;
  wire [24:0] p1_add_70565_comb;
  wire [24:0] p1_add_70566_comb;
  wire [24:0] p1_add_70567_comb;
  wire [24:0] p1_add_70568_comb;
  wire [24:0] p1_add_70569_comb;
  wire [24:0] p1_add_70570_comb;
  wire [24:0] p1_add_70571_comb;
  wire [24:0] p1_add_70572_comb;
  wire [24:0] p1_add_70573_comb;
  wire [24:0] p1_add_70574_comb;
  wire [24:0] p1_add_70575_comb;
  wire [24:0] p1_add_70576_comb;
  wire [24:0] p1_add_70577_comb;
  wire [24:0] p1_add_70578_comb;
  wire [24:0] p1_add_70579_comb;
  wire [24:0] p1_add_70580_comb;
  wire [24:0] p1_add_70581_comb;
  wire [24:0] p1_add_70582_comb;
  wire [24:0] p1_add_70585_comb;
  wire [24:0] p1_add_70586_comb;
  wire [24:0] p1_add_70587_comb;
  wire [24:0] p1_add_70588_comb;
  wire [24:0] p1_add_70589_comb;
  wire [24:0] p1_add_70590_comb;
  wire [24:0] p1_add_70591_comb;
  wire [24:0] p1_add_70592_comb;
  wire [24:0] p1_add_70593_comb;
  wire [24:0] p1_add_70594_comb;
  wire [24:0] p1_add_70595_comb;
  wire [24:0] p1_add_70596_comb;
  wire [24:0] p1_add_70597_comb;
  wire [24:0] p1_add_70598_comb;
  wire p1_sgt_70616_comb;
  wire [11:0] p1_bit_slice_70617_comb;
  wire p1_sgt_70619_comb;
  wire [11:0] p1_bit_slice_70620_comb;
  wire p1_sgt_70622_comb;
  wire [11:0] p1_bit_slice_70623_comb;
  wire p1_sgt_70625_comb;
  wire [11:0] p1_bit_slice_70626_comb;
  wire p1_sgt_70628_comb;
  wire [11:0] p1_bit_slice_70629_comb;
  wire p1_sgt_70631_comb;
  wire [11:0] p1_bit_slice_70632_comb;
  wire p1_sgt_70634_comb;
  wire [11:0] p1_bit_slice_70635_comb;
  wire p1_sgt_70637_comb;
  wire [11:0] p1_bit_slice_70638_comb;
  wire p1_slt_70639_comb;
  wire p1_slt_70640_comb;
  wire p1_slt_70641_comb;
  wire p1_slt_70642_comb;
  wire p1_slt_70643_comb;
  wire p1_slt_70644_comb;
  wire p1_slt_70645_comb;
  wire p1_slt_70646_comb;
  assign p1_array_index_66799_comb = p0_x[3'h3][3'h3];
  assign p1_array_index_66801_comb = p0_x[3'h3][3'h4];
  assign p1_array_index_66803_comb = p0_x[3'h4][3'h3];
  assign p1_array_index_66805_comb = p0_x[3'h4][3'h4];
  assign p1_array_index_66807_comb = p0_x[3'h3][3'h1];
  assign p1_array_index_66809_comb = p0_x[3'h3][3'h2];
  assign p1_array_index_66811_comb = p0_x[3'h3][3'h5];
  assign p1_array_index_66813_comb = p0_x[3'h3][3'h6];
  assign p1_array_index_66815_comb = p0_x[3'h4][3'h1];
  assign p1_array_index_66817_comb = p0_x[3'h4][3'h2];
  assign p1_array_index_66819_comb = p0_x[3'h4][3'h5];
  assign p1_array_index_66821_comb = p0_x[3'h4][3'h6];
  assign p1_array_index_66831_comb = p0_x[3'h3][3'h0];
  assign p1_array_index_66835_comb = p0_x[3'h3][3'h7];
  assign p1_array_index_66837_comb = p0_x[3'h4][3'h0];
  assign p1_array_index_66841_comb = p0_x[3'h4][3'h7];
  assign p1_array_index_66847_comb = p0_x[3'h1][3'h3];
  assign p1_array_index_66849_comb = p0_x[3'h1][3'h4];
  assign p1_array_index_66851_comb = p0_x[3'h2][3'h3];
  assign p1_array_index_66853_comb = p0_x[3'h2][3'h4];
  assign p1_array_index_66855_comb = p0_x[3'h5][3'h3];
  assign p1_array_index_66857_comb = p0_x[3'h5][3'h4];
  assign p1_array_index_66859_comb = p0_x[3'h6][3'h3];
  assign p1_array_index_66861_comb = p0_x[3'h6][3'h4];
  assign p1_array_index_66863_comb = p0_x[3'h1][3'h1];
  assign p1_array_index_66865_comb = p0_x[3'h1][3'h2];
  assign p1_array_index_66867_comb = p0_x[3'h1][3'h5];
  assign p1_array_index_66869_comb = p0_x[3'h1][3'h6];
  assign p1_array_index_66871_comb = p0_x[3'h2][3'h1];
  assign p1_array_index_66873_comb = p0_x[3'h2][3'h2];
  assign p1_array_index_66875_comb = p0_x[3'h2][3'h5];
  assign p1_array_index_66877_comb = p0_x[3'h2][3'h6];
  assign p1_array_index_66879_comb = p0_x[3'h5][3'h1];
  assign p1_array_index_66881_comb = p0_x[3'h5][3'h2];
  assign p1_array_index_66883_comb = p0_x[3'h5][3'h5];
  assign p1_array_index_66885_comb = p0_x[3'h5][3'h6];
  assign p1_array_index_66887_comb = p0_x[3'h6][3'h1];
  assign p1_array_index_66889_comb = p0_x[3'h6][3'h2];
  assign p1_array_index_66891_comb = p0_x[3'h6][3'h5];
  assign p1_array_index_66893_comb = p0_x[3'h6][3'h6];
  assign p1_array_index_66911_comb = p0_x[3'h1][3'h0];
  assign p1_array_index_66915_comb = p0_x[3'h1][3'h7];
  assign p1_array_index_66917_comb = p0_x[3'h2][3'h0];
  assign p1_array_index_66921_comb = p0_x[3'h2][3'h7];
  assign p1_array_index_66923_comb = p0_x[3'h5][3'h0];
  assign p1_array_index_66927_comb = p0_x[3'h5][3'h7];
  assign p1_array_index_66929_comb = p0_x[3'h6][3'h0];
  assign p1_array_index_66933_comb = p0_x[3'h6][3'h7];
  assign p1_array_index_66943_comb = p0_x[3'h0][3'h3];
  assign p1_array_index_66945_comb = p0_x[3'h0][3'h4];
  assign p1_array_index_66947_comb = p0_x[3'h7][3'h3];
  assign p1_array_index_66949_comb = p0_x[3'h7][3'h4];
  assign p1_array_index_66951_comb = p0_x[3'h0][3'h1];
  assign p1_array_index_66953_comb = p0_x[3'h0][3'h2];
  assign p1_array_index_66955_comb = p0_x[3'h0][3'h5];
  assign p1_array_index_66957_comb = p0_x[3'h0][3'h6];
  assign p1_array_index_66959_comb = p0_x[3'h7][3'h1];
  assign p1_array_index_66961_comb = p0_x[3'h7][3'h2];
  assign p1_array_index_66963_comb = p0_x[3'h7][3'h5];
  assign p1_array_index_66965_comb = p0_x[3'h7][3'h6];
  assign p1_array_index_66975_comb = p0_x[3'h0][3'h0];
  assign p1_array_index_66979_comb = p0_x[3'h0][3'h7];
  assign p1_array_index_66981_comb = p0_x[3'h7][3'h0];
  assign p1_array_index_66985_comb = p0_x[3'h7][3'h7];
  assign p1_smul_27786_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66799_comb, 6'h19);
  assign p1_smul_27788_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66801_comb, 6'h27);
  assign p1_smul_27802_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66803_comb, 6'h19);
  assign p1_smul_27804_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66805_comb, 6'h27);
  assign p1_smul_27910_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66807_comb, 7'h31);
  assign p1_smul_27912_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66809_comb, 7'h4f);
  assign p1_smul_27918_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66811_comb, 7'h4f);
  assign p1_smul_27920_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66813_comb, 7'h31);
  assign p1_smul_27926_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66815_comb, 7'h31);
  assign p1_smul_27928_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66817_comb, 7'h4f);
  assign p1_smul_27934_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66819_comb, 7'h4f);
  assign p1_smul_27936_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66821_comb, 7'h31);
  assign p1_smul_28038_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66807_comb, 6'h27);
  assign p1_smul_28048_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66813_comb, 6'h19);
  assign p1_smul_28054_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66815_comb, 6'h27);
  assign p1_smul_28064_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66821_comb, 6'h19);
  assign p1_smul_28296_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66809_comb, 6'h27);
  assign p1_smul_28302_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66811_comb, 6'h27);
  assign p1_smul_28312_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66817_comb, 6'h27);
  assign p1_smul_28318_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66819_comb, 6'h27);
  assign p1_smul_28420_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66831_comb, 7'h31);
  assign p1_smul_28424_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66809_comb, 7'h31);
  assign p1_smul_28430_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66811_comb, 7'h31);
  assign p1_smul_28434_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66835_comb, 7'h31);
  assign p1_smul_28436_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66837_comb, 7'h31);
  assign p1_smul_28440_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66817_comb, 7'h31);
  assign p1_smul_28446_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66819_comb, 7'h31);
  assign p1_smul_28450_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66841_comb, 7'h31);
  assign p1_smul_28548_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66831_comb, 6'h19);
  assign p1_smul_28562_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66835_comb, 6'h19);
  assign p1_smul_28564_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66837_comb, 6'h19);
  assign p1_smul_28578_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66841_comb, 6'h19);
  assign p1_smul_27754_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66847_comb, 6'h19);
  assign p1_smul_27756_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66849_comb, 6'h27);
  assign p1_smul_27770_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66851_comb, 6'h19);
  assign p1_smul_27772_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66853_comb, 6'h27);
  assign p1_smul_27818_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66855_comb, 6'h19);
  assign p1_smul_27820_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66857_comb, 6'h27);
  assign p1_smul_27834_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66859_comb, 6'h19);
  assign p1_smul_27836_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66861_comb, 6'h27);
  assign p1_smul_27878_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66863_comb, 7'h31);
  assign p1_smul_27880_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66865_comb, 7'h4f);
  assign p1_smul_27886_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66867_comb, 7'h4f);
  assign p1_smul_27888_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66869_comb, 7'h31);
  assign p1_smul_27894_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66871_comb, 7'h31);
  assign p1_smul_27896_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66873_comb, 7'h4f);
  assign p1_smul_27902_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66875_comb, 7'h4f);
  assign p1_smul_27904_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66877_comb, 7'h31);
  assign p1_smul_27942_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66879_comb, 7'h31);
  assign p1_smul_27944_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66881_comb, 7'h4f);
  assign p1_smul_27950_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66883_comb, 7'h4f);
  assign p1_smul_27952_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66885_comb, 7'h31);
  assign p1_smul_27958_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66887_comb, 7'h31);
  assign p1_smul_27960_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66889_comb, 7'h4f);
  assign p1_smul_27966_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66891_comb, 7'h4f);
  assign p1_smul_27968_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66893_comb, 7'h31);
  assign p1_smul_28006_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66863_comb, 6'h27);
  assign p1_smul_28016_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66869_comb, 6'h19);
  assign p1_smul_28022_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66871_comb, 6'h27);
  assign p1_smul_28032_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66877_comb, 6'h19);
  assign p1_smul_28070_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66879_comb, 6'h27);
  assign p1_smul_28080_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66885_comb, 6'h19);
  assign p1_smul_28086_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66887_comb, 6'h27);
  assign p1_smul_28096_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66893_comb, 6'h19);
  assign p1_smul_28264_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66865_comb, 6'h27);
  assign p1_smul_28270_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66867_comb, 6'h27);
  assign p1_smul_28280_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66873_comb, 6'h27);
  assign p1_smul_28286_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66875_comb, 6'h27);
  assign p1_smul_28328_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66881_comb, 6'h27);
  assign p1_smul_28334_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66883_comb, 6'h27);
  assign p1_smul_28344_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66889_comb, 6'h27);
  assign p1_smul_28350_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66891_comb, 6'h27);
  assign p1_smul_28388_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66911_comb, 7'h31);
  assign p1_smul_28392_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66865_comb, 7'h31);
  assign p1_smul_28398_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66867_comb, 7'h31);
  assign p1_smul_28402_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66915_comb, 7'h31);
  assign p1_smul_28404_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66917_comb, 7'h31);
  assign p1_smul_28408_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66873_comb, 7'h31);
  assign p1_smul_28414_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66875_comb, 7'h31);
  assign p1_smul_28418_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66921_comb, 7'h31);
  assign p1_smul_28452_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66923_comb, 7'h31);
  assign p1_smul_28456_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66881_comb, 7'h31);
  assign p1_smul_28462_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66883_comb, 7'h31);
  assign p1_smul_28466_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66927_comb, 7'h31);
  assign p1_smul_28468_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66929_comb, 7'h31);
  assign p1_smul_28472_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66889_comb, 7'h31);
  assign p1_smul_28478_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66891_comb, 7'h31);
  assign p1_smul_28482_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66933_comb, 7'h31);
  assign p1_smul_28516_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66911_comb, 6'h19);
  assign p1_smul_28530_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66915_comb, 6'h19);
  assign p1_smul_28532_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66917_comb, 6'h19);
  assign p1_smul_28546_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66921_comb, 6'h19);
  assign p1_smul_28580_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66923_comb, 6'h19);
  assign p1_smul_28594_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66927_comb, 6'h19);
  assign p1_smul_28596_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66929_comb, 6'h19);
  assign p1_smul_28610_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66933_comb, 6'h19);
  assign p1_smul_27738_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66943_comb, 6'h19);
  assign p1_smul_27740_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66945_comb, 6'h27);
  assign p1_smul_27850_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66947_comb, 6'h19);
  assign p1_smul_27852_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66949_comb, 6'h27);
  assign p1_smul_27862_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66951_comb, 7'h31);
  assign p1_smul_27864_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66953_comb, 7'h4f);
  assign p1_smul_27870_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66955_comb, 7'h4f);
  assign p1_smul_27872_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66957_comb, 7'h31);
  assign p1_smul_27974_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66959_comb, 7'h31);
  assign p1_smul_27976_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66961_comb, 7'h4f);
  assign p1_smul_27982_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66963_comb, 7'h4f);
  assign p1_smul_27984_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66965_comb, 7'h31);
  assign p1_smul_27990_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66951_comb, 6'h27);
  assign p1_smul_28000_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66957_comb, 6'h19);
  assign p1_smul_28102_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66959_comb, 6'h27);
  assign p1_smul_28112_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66965_comb, 6'h19);
  assign p1_smul_28248_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66953_comb, 6'h27);
  assign p1_smul_28254_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66955_comb, 6'h27);
  assign p1_smul_28360_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66961_comb, 6'h27);
  assign p1_smul_28366_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66963_comb, 6'h27);
  assign p1_smul_28372_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66975_comb, 7'h31);
  assign p1_smul_28376_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66953_comb, 7'h31);
  assign p1_smul_28382_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66955_comb, 7'h31);
  assign p1_smul_28386_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66979_comb, 7'h31);
  assign p1_smul_28484_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66981_comb, 7'h31);
  assign p1_smul_28488_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66961_comb, 7'h31);
  assign p1_smul_28494_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66963_comb, 7'h31);
  assign p1_smul_28498_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66985_comb, 7'h31);
  assign p1_smul_28500_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66975_comb, 6'h19);
  assign p1_smul_28514_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66979_comb, 6'h19);
  assign p1_smul_28612_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66981_comb, 6'h19);
  assign p1_smul_28626_NarrowedMult__comb = smul18b_12b_x_6b(p1_array_index_66985_comb, 6'h19);
  assign p1_smul_67439_comb = smul21b_12b_x_9b(p1_array_index_66831_comb, 9'h0fb);
  assign p1_smul_67440_comb = smul21b_12b_x_9b(p1_array_index_66807_comb, 9'h0d5);
  assign p1_smul_27784_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66809_comb, 8'h47);
  assign p1_smul_27790_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66811_comb, 8'hb9);
  assign p1_smul_67447_comb = smul21b_12b_x_9b(p1_array_index_66813_comb, 9'h12b);
  assign p1_smul_67448_comb = smul21b_12b_x_9b(p1_array_index_66835_comb, 9'h105);
  assign p1_smul_67449_comb = smul21b_12b_x_9b(p1_array_index_66837_comb, 9'h0fb);
  assign p1_smul_67450_comb = smul21b_12b_x_9b(p1_array_index_66815_comb, 9'h0d5);
  assign p1_smul_27800_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66817_comb, 8'h47);
  assign p1_smul_27806_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66819_comb, 8'hb9);
  assign p1_smul_67457_comb = smul21b_12b_x_9b(p1_array_index_66821_comb, 9'h12b);
  assign p1_smul_67458_comb = smul21b_12b_x_9b(p1_array_index_66841_comb, 9'h105);
  assign p1_smul_27908_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66831_comb, 7'h3b);
  assign p1_smul_27914_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66799_comb, 7'h45);
  assign p1_smul_27916_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66801_comb, 7'h45);
  assign p1_smul_27922_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66835_comb, 7'h3b);
  assign p1_smul_27924_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66837_comb, 7'h3b);
  assign p1_smul_27930_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66803_comb, 7'h45);
  assign p1_smul_27932_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66805_comb, 7'h45);
  assign p1_smul_27938_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66841_comb, 7'h3b);
  assign p1_smul_67483_comb = smul21b_12b_x_9b(p1_array_index_66831_comb, 9'h0d5);
  assign p1_smul_67486_comb = smul21b_12b_x_9b(p1_array_index_66809_comb, 9'h105);
  assign p1_smul_28042_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66799_comb, 8'hb9);
  assign p1_smul_28044_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66801_comb, 8'h47);
  assign p1_smul_67489_comb = smul21b_12b_x_9b(p1_array_index_66811_comb, 9'h0fb);
  assign p1_smul_67492_comb = smul21b_12b_x_9b(p1_array_index_66835_comb, 9'h12b);
  assign p1_smul_67493_comb = smul21b_12b_x_9b(p1_array_index_66837_comb, 9'h0d5);
  assign p1_smul_67496_comb = smul21b_12b_x_9b(p1_array_index_66817_comb, 9'h105);
  assign p1_smul_28058_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66803_comb, 8'hb9);
  assign p1_smul_28060_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66805_comb, 8'h47);
  assign p1_smul_67499_comb = smul21b_12b_x_9b(p1_array_index_66819_comb, 9'h0fb);
  assign p1_smul_67502_comb = smul21b_12b_x_9b(p1_array_index_66841_comb, 9'h12b);
  assign p1_smul_67503_comb = smul21b_12b_x_9b(p1_array_index_66831_comb, 9'h0b5);
  assign p1_smul_67504_comb = smul21b_12b_x_9b(p1_array_index_66807_comb, 9'h14b);
  assign p1_smul_67505_comb = smul21b_12b_x_9b(p1_array_index_66809_comb, 9'h14b);
  assign p1_smul_67506_comb = smul21b_12b_x_9b(p1_array_index_66799_comb, 9'h0b5);
  assign p1_smul_67507_comb = smul21b_12b_x_9b(p1_array_index_66801_comb, 9'h0b5);
  assign p1_smul_67508_comb = smul21b_12b_x_9b(p1_array_index_66811_comb, 9'h14b);
  assign p1_smul_67509_comb = smul21b_12b_x_9b(p1_array_index_66813_comb, 9'h14b);
  assign p1_smul_67510_comb = smul21b_12b_x_9b(p1_array_index_66835_comb, 9'h0b5);
  assign p1_smul_67511_comb = smul21b_12b_x_9b(p1_array_index_66837_comb, 9'h0b5);
  assign p1_smul_67512_comb = smul21b_12b_x_9b(p1_array_index_66815_comb, 9'h14b);
  assign p1_smul_67513_comb = smul21b_12b_x_9b(p1_array_index_66817_comb, 9'h14b);
  assign p1_smul_67514_comb = smul21b_12b_x_9b(p1_array_index_66803_comb, 9'h0b5);
  assign p1_smul_67515_comb = smul21b_12b_x_9b(p1_array_index_66805_comb, 9'h0b5);
  assign p1_smul_67516_comb = smul21b_12b_x_9b(p1_array_index_66819_comb, 9'h14b);
  assign p1_smul_67517_comb = smul21b_12b_x_9b(p1_array_index_66821_comb, 9'h14b);
  assign p1_smul_67518_comb = smul21b_12b_x_9b(p1_array_index_66841_comb, 9'h0b5);
  assign p1_smul_28292_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66831_comb, 8'h47);
  assign p1_smul_67520_comb = smul21b_12b_x_9b(p1_array_index_66807_comb, 9'h105);
  assign p1_smul_67523_comb = smul21b_12b_x_9b(p1_array_index_66799_comb, 9'h0d5);
  assign p1_smul_67524_comb = smul21b_12b_x_9b(p1_array_index_66801_comb, 9'h0d5);
  assign p1_smul_67527_comb = smul21b_12b_x_9b(p1_array_index_66813_comb, 9'h105);
  assign p1_smul_28306_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66835_comb, 8'h47);
  assign p1_smul_28308_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66837_comb, 8'h47);
  assign p1_smul_67530_comb = smul21b_12b_x_9b(p1_array_index_66815_comb, 9'h105);
  assign p1_smul_67533_comb = smul21b_12b_x_9b(p1_array_index_66803_comb, 9'h0d5);
  assign p1_smul_67534_comb = smul21b_12b_x_9b(p1_array_index_66805_comb, 9'h0d5);
  assign p1_smul_67537_comb = smul21b_12b_x_9b(p1_array_index_66821_comb, 9'h105);
  assign p1_smul_28322_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66841_comb, 8'h47);
  assign p1_smul_28422_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66807_comb, 7'h45);
  assign p1_smul_28426_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66799_comb, 7'h3b);
  assign p1_smul_28428_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66801_comb, 7'h3b);
  assign p1_smul_28432_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66813_comb, 7'h45);
  assign p1_smul_28438_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66815_comb, 7'h45);
  assign p1_smul_28442_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66803_comb, 7'h3b);
  assign p1_smul_28444_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66805_comb, 7'h3b);
  assign p1_smul_28448_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66821_comb, 7'h45);
  assign p1_smul_28550_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66807_comb, 8'hb9);
  assign p1_smul_67566_comb = smul21b_12b_x_9b(p1_array_index_66809_comb, 9'h0d5);
  assign p1_smul_67567_comb = smul21b_12b_x_9b(p1_array_index_66799_comb, 9'h105);
  assign p1_smul_67568_comb = smul21b_12b_x_9b(p1_array_index_66801_comb, 9'h105);
  assign p1_smul_67569_comb = smul21b_12b_x_9b(p1_array_index_66811_comb, 9'h0d5);
  assign p1_smul_28560_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66813_comb, 8'hb9);
  assign p1_smul_28566_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66815_comb, 8'hb9);
  assign p1_smul_67576_comb = smul21b_12b_x_9b(p1_array_index_66817_comb, 9'h0d5);
  assign p1_smul_67577_comb = smul21b_12b_x_9b(p1_array_index_66803_comb, 9'h105);
  assign p1_smul_67578_comb = smul21b_12b_x_9b(p1_array_index_66805_comb, 9'h105);
  assign p1_smul_67579_comb = smul21b_12b_x_9b(p1_array_index_66819_comb, 9'h0d5);
  assign p1_smul_28576_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66821_comb, 8'hb9);
  assign p1_smul_67583_comb = smul21b_12b_x_9b(p1_array_index_66911_comb, 9'h0fb);
  assign p1_smul_67584_comb = smul21b_12b_x_9b(p1_array_index_66863_comb, 9'h0d5);
  assign p1_smul_27752_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66865_comb, 8'h47);
  assign p1_smul_27758_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66867_comb, 8'hb9);
  assign p1_smul_67591_comb = smul21b_12b_x_9b(p1_array_index_66869_comb, 9'h12b);
  assign p1_smul_67592_comb = smul21b_12b_x_9b(p1_array_index_66915_comb, 9'h105);
  assign p1_smul_67593_comb = smul21b_12b_x_9b(p1_array_index_66917_comb, 9'h0fb);
  assign p1_smul_67594_comb = smul21b_12b_x_9b(p1_array_index_66871_comb, 9'h0d5);
  assign p1_smul_27768_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66873_comb, 8'h47);
  assign p1_smul_27774_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66875_comb, 8'hb9);
  assign p1_smul_67601_comb = smul21b_12b_x_9b(p1_array_index_66877_comb, 9'h12b);
  assign p1_smul_67602_comb = smul21b_12b_x_9b(p1_array_index_66921_comb, 9'h105);
  assign p1_smul_67603_comb = smul21b_12b_x_9b(p1_array_index_66923_comb, 9'h0fb);
  assign p1_smul_67604_comb = smul21b_12b_x_9b(p1_array_index_66879_comb, 9'h0d5);
  assign p1_smul_27816_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66881_comb, 8'h47);
  assign p1_smul_27822_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66883_comb, 8'hb9);
  assign p1_smul_67611_comb = smul21b_12b_x_9b(p1_array_index_66885_comb, 9'h12b);
  assign p1_smul_67612_comb = smul21b_12b_x_9b(p1_array_index_66927_comb, 9'h105);
  assign p1_smul_67613_comb = smul21b_12b_x_9b(p1_array_index_66929_comb, 9'h0fb);
  assign p1_smul_67614_comb = smul21b_12b_x_9b(p1_array_index_66887_comb, 9'h0d5);
  assign p1_smul_27832_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66889_comb, 8'h47);
  assign p1_smul_27838_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66891_comb, 8'hb9);
  assign p1_smul_67621_comb = smul21b_12b_x_9b(p1_array_index_66893_comb, 9'h12b);
  assign p1_smul_67622_comb = smul21b_12b_x_9b(p1_array_index_66933_comb, 9'h105);
  assign p1_smul_27876_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66911_comb, 7'h3b);
  assign p1_smul_27882_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66847_comb, 7'h45);
  assign p1_smul_27884_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66849_comb, 7'h45);
  assign p1_smul_27890_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66915_comb, 7'h3b);
  assign p1_smul_27892_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66917_comb, 7'h3b);
  assign p1_smul_27898_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66851_comb, 7'h45);
  assign p1_smul_27900_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66853_comb, 7'h45);
  assign p1_smul_27906_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66921_comb, 7'h3b);
  assign p1_smul_27940_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66923_comb, 7'h3b);
  assign p1_smul_27946_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66855_comb, 7'h45);
  assign p1_smul_27948_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66857_comb, 7'h45);
  assign p1_smul_27954_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66927_comb, 7'h3b);
  assign p1_smul_27956_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66929_comb, 7'h3b);
  assign p1_smul_27962_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66859_comb, 7'h45);
  assign p1_smul_27964_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66861_comb, 7'h45);
  assign p1_smul_27970_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66933_comb, 7'h3b);
  assign p1_smul_67671_comb = smul21b_12b_x_9b(p1_array_index_66911_comb, 9'h0d5);
  assign p1_smul_67674_comb = smul21b_12b_x_9b(p1_array_index_66865_comb, 9'h105);
  assign p1_smul_28010_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66847_comb, 8'hb9);
  assign p1_smul_28012_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66849_comb, 8'h47);
  assign p1_smul_67677_comb = smul21b_12b_x_9b(p1_array_index_66867_comb, 9'h0fb);
  assign p1_smul_67680_comb = smul21b_12b_x_9b(p1_array_index_66915_comb, 9'h12b);
  assign p1_smul_67681_comb = smul21b_12b_x_9b(p1_array_index_66917_comb, 9'h0d5);
  assign p1_smul_67684_comb = smul21b_12b_x_9b(p1_array_index_66873_comb, 9'h105);
  assign p1_smul_28026_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66851_comb, 8'hb9);
  assign p1_smul_28028_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66853_comb, 8'h47);
  assign p1_smul_67687_comb = smul21b_12b_x_9b(p1_array_index_66875_comb, 9'h0fb);
  assign p1_smul_67690_comb = smul21b_12b_x_9b(p1_array_index_66921_comb, 9'h12b);
  assign p1_smul_67691_comb = smul21b_12b_x_9b(p1_array_index_66923_comb, 9'h0d5);
  assign p1_smul_67694_comb = smul21b_12b_x_9b(p1_array_index_66881_comb, 9'h105);
  assign p1_smul_28074_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66855_comb, 8'hb9);
  assign p1_smul_28076_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66857_comb, 8'h47);
  assign p1_smul_67697_comb = smul21b_12b_x_9b(p1_array_index_66883_comb, 9'h0fb);
  assign p1_smul_67700_comb = smul21b_12b_x_9b(p1_array_index_66927_comb, 9'h12b);
  assign p1_smul_67701_comb = smul21b_12b_x_9b(p1_array_index_66929_comb, 9'h0d5);
  assign p1_smul_67704_comb = smul21b_12b_x_9b(p1_array_index_66889_comb, 9'h105);
  assign p1_smul_28090_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66859_comb, 8'hb9);
  assign p1_smul_28092_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66861_comb, 8'h47);
  assign p1_smul_67707_comb = smul21b_12b_x_9b(p1_array_index_66891_comb, 9'h0fb);
  assign p1_smul_67710_comb = smul21b_12b_x_9b(p1_array_index_66933_comb, 9'h12b);
  assign p1_smul_67711_comb = smul21b_12b_x_9b(p1_array_index_66911_comb, 9'h0b5);
  assign p1_smul_67712_comb = smul21b_12b_x_9b(p1_array_index_66863_comb, 9'h14b);
  assign p1_smul_67713_comb = smul21b_12b_x_9b(p1_array_index_66865_comb, 9'h14b);
  assign p1_smul_67714_comb = smul21b_12b_x_9b(p1_array_index_66847_comb, 9'h0b5);
  assign p1_smul_67715_comb = smul21b_12b_x_9b(p1_array_index_66849_comb, 9'h0b5);
  assign p1_smul_67716_comb = smul21b_12b_x_9b(p1_array_index_66867_comb, 9'h14b);
  assign p1_smul_67717_comb = smul21b_12b_x_9b(p1_array_index_66869_comb, 9'h14b);
  assign p1_smul_67718_comb = smul21b_12b_x_9b(p1_array_index_66915_comb, 9'h0b5);
  assign p1_smul_67719_comb = smul21b_12b_x_9b(p1_array_index_66917_comb, 9'h0b5);
  assign p1_smul_67720_comb = smul21b_12b_x_9b(p1_array_index_66871_comb, 9'h14b);
  assign p1_smul_67721_comb = smul21b_12b_x_9b(p1_array_index_66873_comb, 9'h14b);
  assign p1_smul_67722_comb = smul21b_12b_x_9b(p1_array_index_66851_comb, 9'h0b5);
  assign p1_smul_67723_comb = smul21b_12b_x_9b(p1_array_index_66853_comb, 9'h0b5);
  assign p1_smul_67724_comb = smul21b_12b_x_9b(p1_array_index_66875_comb, 9'h14b);
  assign p1_smul_67725_comb = smul21b_12b_x_9b(p1_array_index_66877_comb, 9'h14b);
  assign p1_smul_67726_comb = smul21b_12b_x_9b(p1_array_index_66921_comb, 9'h0b5);
  assign p1_smul_67727_comb = smul21b_12b_x_9b(p1_array_index_66923_comb, 9'h0b5);
  assign p1_smul_67728_comb = smul21b_12b_x_9b(p1_array_index_66879_comb, 9'h14b);
  assign p1_smul_67729_comb = smul21b_12b_x_9b(p1_array_index_66881_comb, 9'h14b);
  assign p1_smul_67730_comb = smul21b_12b_x_9b(p1_array_index_66855_comb, 9'h0b5);
  assign p1_smul_67731_comb = smul21b_12b_x_9b(p1_array_index_66857_comb, 9'h0b5);
  assign p1_smul_67732_comb = smul21b_12b_x_9b(p1_array_index_66883_comb, 9'h14b);
  assign p1_smul_67733_comb = smul21b_12b_x_9b(p1_array_index_66885_comb, 9'h14b);
  assign p1_smul_67734_comb = smul21b_12b_x_9b(p1_array_index_66927_comb, 9'h0b5);
  assign p1_smul_67735_comb = smul21b_12b_x_9b(p1_array_index_66929_comb, 9'h0b5);
  assign p1_smul_67736_comb = smul21b_12b_x_9b(p1_array_index_66887_comb, 9'h14b);
  assign p1_smul_67737_comb = smul21b_12b_x_9b(p1_array_index_66889_comb, 9'h14b);
  assign p1_smul_67738_comb = smul21b_12b_x_9b(p1_array_index_66859_comb, 9'h0b5);
  assign p1_smul_67739_comb = smul21b_12b_x_9b(p1_array_index_66861_comb, 9'h0b5);
  assign p1_smul_67740_comb = smul21b_12b_x_9b(p1_array_index_66891_comb, 9'h14b);
  assign p1_smul_67741_comb = smul21b_12b_x_9b(p1_array_index_66893_comb, 9'h14b);
  assign p1_smul_67742_comb = smul21b_12b_x_9b(p1_array_index_66933_comb, 9'h0b5);
  assign p1_smul_28260_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66911_comb, 8'h47);
  assign p1_smul_67744_comb = smul21b_12b_x_9b(p1_array_index_66863_comb, 9'h105);
  assign p1_smul_67747_comb = smul21b_12b_x_9b(p1_array_index_66847_comb, 9'h0d5);
  assign p1_smul_67748_comb = smul21b_12b_x_9b(p1_array_index_66849_comb, 9'h0d5);
  assign p1_smul_67751_comb = smul21b_12b_x_9b(p1_array_index_66869_comb, 9'h105);
  assign p1_smul_28274_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66915_comb, 8'h47);
  assign p1_smul_28276_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66917_comb, 8'h47);
  assign p1_smul_67754_comb = smul21b_12b_x_9b(p1_array_index_66871_comb, 9'h105);
  assign p1_smul_67757_comb = smul21b_12b_x_9b(p1_array_index_66851_comb, 9'h0d5);
  assign p1_smul_67758_comb = smul21b_12b_x_9b(p1_array_index_66853_comb, 9'h0d5);
  assign p1_smul_67761_comb = smul21b_12b_x_9b(p1_array_index_66877_comb, 9'h105);
  assign p1_smul_28290_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66921_comb, 8'h47);
  assign p1_smul_28324_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66923_comb, 8'h47);
  assign p1_smul_67764_comb = smul21b_12b_x_9b(p1_array_index_66879_comb, 9'h105);
  assign p1_smul_67767_comb = smul21b_12b_x_9b(p1_array_index_66855_comb, 9'h0d5);
  assign p1_smul_67768_comb = smul21b_12b_x_9b(p1_array_index_66857_comb, 9'h0d5);
  assign p1_smul_67771_comb = smul21b_12b_x_9b(p1_array_index_66885_comb, 9'h105);
  assign p1_smul_28338_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66927_comb, 8'h47);
  assign p1_smul_28340_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66929_comb, 8'h47);
  assign p1_smul_67774_comb = smul21b_12b_x_9b(p1_array_index_66887_comb, 9'h105);
  assign p1_smul_67777_comb = smul21b_12b_x_9b(p1_array_index_66859_comb, 9'h0d5);
  assign p1_smul_67778_comb = smul21b_12b_x_9b(p1_array_index_66861_comb, 9'h0d5);
  assign p1_smul_67781_comb = smul21b_12b_x_9b(p1_array_index_66893_comb, 9'h105);
  assign p1_smul_28354_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66933_comb, 8'h47);
  assign p1_smul_28390_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66863_comb, 7'h45);
  assign p1_smul_28394_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66847_comb, 7'h3b);
  assign p1_smul_28396_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66849_comb, 7'h3b);
  assign p1_smul_28400_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66869_comb, 7'h45);
  assign p1_smul_28406_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66871_comb, 7'h45);
  assign p1_smul_28410_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66851_comb, 7'h3b);
  assign p1_smul_28412_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66853_comb, 7'h3b);
  assign p1_smul_28416_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66877_comb, 7'h45);
  assign p1_smul_28454_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66879_comb, 7'h45);
  assign p1_smul_28458_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66855_comb, 7'h3b);
  assign p1_smul_28460_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66857_comb, 7'h3b);
  assign p1_smul_28464_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66885_comb, 7'h45);
  assign p1_smul_28470_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66887_comb, 7'h45);
  assign p1_smul_28474_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66859_comb, 7'h3b);
  assign p1_smul_28476_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66861_comb, 7'h3b);
  assign p1_smul_28480_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66893_comb, 7'h45);
  assign p1_smul_28518_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66863_comb, 8'hb9);
  assign p1_smul_67834_comb = smul21b_12b_x_9b(p1_array_index_66865_comb, 9'h0d5);
  assign p1_smul_67835_comb = smul21b_12b_x_9b(p1_array_index_66847_comb, 9'h105);
  assign p1_smul_67836_comb = smul21b_12b_x_9b(p1_array_index_66849_comb, 9'h105);
  assign p1_smul_67837_comb = smul21b_12b_x_9b(p1_array_index_66867_comb, 9'h0d5);
  assign p1_smul_28528_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66869_comb, 8'hb9);
  assign p1_smul_28534_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66871_comb, 8'hb9);
  assign p1_smul_67844_comb = smul21b_12b_x_9b(p1_array_index_66873_comb, 9'h0d5);
  assign p1_smul_67845_comb = smul21b_12b_x_9b(p1_array_index_66851_comb, 9'h105);
  assign p1_smul_67846_comb = smul21b_12b_x_9b(p1_array_index_66853_comb, 9'h105);
  assign p1_smul_67847_comb = smul21b_12b_x_9b(p1_array_index_66875_comb, 9'h0d5);
  assign p1_smul_28544_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66877_comb, 8'hb9);
  assign p1_smul_28582_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66879_comb, 8'hb9);
  assign p1_smul_67854_comb = smul21b_12b_x_9b(p1_array_index_66881_comb, 9'h0d5);
  assign p1_smul_67855_comb = smul21b_12b_x_9b(p1_array_index_66855_comb, 9'h105);
  assign p1_smul_67856_comb = smul21b_12b_x_9b(p1_array_index_66857_comb, 9'h105);
  assign p1_smul_67857_comb = smul21b_12b_x_9b(p1_array_index_66883_comb, 9'h0d5);
  assign p1_smul_28592_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66885_comb, 8'hb9);
  assign p1_smul_28598_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66887_comb, 8'hb9);
  assign p1_smul_67864_comb = smul21b_12b_x_9b(p1_array_index_66889_comb, 9'h0d5);
  assign p1_smul_67865_comb = smul21b_12b_x_9b(p1_array_index_66859_comb, 9'h105);
  assign p1_smul_67866_comb = smul21b_12b_x_9b(p1_array_index_66861_comb, 9'h105);
  assign p1_smul_67867_comb = smul21b_12b_x_9b(p1_array_index_66891_comb, 9'h0d5);
  assign p1_smul_28608_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66893_comb, 8'hb9);
  assign p1_smul_67871_comb = smul21b_12b_x_9b(p1_array_index_66975_comb, 9'h0fb);
  assign p1_smul_67872_comb = smul21b_12b_x_9b(p1_array_index_66951_comb, 9'h0d5);
  assign p1_smul_27736_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66953_comb, 8'h47);
  assign p1_smul_27742_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66955_comb, 8'hb9);
  assign p1_smul_67879_comb = smul21b_12b_x_9b(p1_array_index_66957_comb, 9'h12b);
  assign p1_smul_67880_comb = smul21b_12b_x_9b(p1_array_index_66979_comb, 9'h105);
  assign p1_smul_67881_comb = smul21b_12b_x_9b(p1_array_index_66981_comb, 9'h0fb);
  assign p1_smul_67882_comb = smul21b_12b_x_9b(p1_array_index_66959_comb, 9'h0d5);
  assign p1_smul_27848_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66961_comb, 8'h47);
  assign p1_smul_27854_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66963_comb, 8'hb9);
  assign p1_smul_67889_comb = smul21b_12b_x_9b(p1_array_index_66965_comb, 9'h12b);
  assign p1_smul_67890_comb = smul21b_12b_x_9b(p1_array_index_66985_comb, 9'h105);
  assign p1_smul_27860_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66975_comb, 7'h3b);
  assign p1_smul_27866_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66943_comb, 7'h45);
  assign p1_smul_27868_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66945_comb, 7'h45);
  assign p1_smul_27874_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66979_comb, 7'h3b);
  assign p1_smul_27972_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66981_comb, 7'h3b);
  assign p1_smul_27978_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66947_comb, 7'h45);
  assign p1_smul_27980_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66949_comb, 7'h45);
  assign p1_smul_27986_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66985_comb, 7'h3b);
  assign p1_smul_67915_comb = smul21b_12b_x_9b(p1_array_index_66975_comb, 9'h0d5);
  assign p1_smul_67918_comb = smul21b_12b_x_9b(p1_array_index_66953_comb, 9'h105);
  assign p1_smul_27994_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66943_comb, 8'hb9);
  assign p1_smul_27996_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66945_comb, 8'h47);
  assign p1_smul_67921_comb = smul21b_12b_x_9b(p1_array_index_66955_comb, 9'h0fb);
  assign p1_smul_67924_comb = smul21b_12b_x_9b(p1_array_index_66979_comb, 9'h12b);
  assign p1_smul_67925_comb = smul21b_12b_x_9b(p1_array_index_66981_comb, 9'h0d5);
  assign p1_smul_67928_comb = smul21b_12b_x_9b(p1_array_index_66961_comb, 9'h105);
  assign p1_smul_28106_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66947_comb, 8'hb9);
  assign p1_smul_28108_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66949_comb, 8'h47);
  assign p1_smul_67931_comb = smul21b_12b_x_9b(p1_array_index_66963_comb, 9'h0fb);
  assign p1_smul_67934_comb = smul21b_12b_x_9b(p1_array_index_66985_comb, 9'h12b);
  assign p1_smul_67935_comb = smul21b_12b_x_9b(p1_array_index_66975_comb, 9'h0b5);
  assign p1_smul_67936_comb = smul21b_12b_x_9b(p1_array_index_66951_comb, 9'h14b);
  assign p1_smul_67937_comb = smul21b_12b_x_9b(p1_array_index_66953_comb, 9'h14b);
  assign p1_smul_67938_comb = smul21b_12b_x_9b(p1_array_index_66943_comb, 9'h0b5);
  assign p1_smul_67939_comb = smul21b_12b_x_9b(p1_array_index_66945_comb, 9'h0b5);
  assign p1_smul_67940_comb = smul21b_12b_x_9b(p1_array_index_66955_comb, 9'h14b);
  assign p1_smul_67941_comb = smul21b_12b_x_9b(p1_array_index_66957_comb, 9'h14b);
  assign p1_smul_67942_comb = smul21b_12b_x_9b(p1_array_index_66979_comb, 9'h0b5);
  assign p1_smul_67943_comb = smul21b_12b_x_9b(p1_array_index_66981_comb, 9'h0b5);
  assign p1_smul_67944_comb = smul21b_12b_x_9b(p1_array_index_66959_comb, 9'h14b);
  assign p1_smul_67945_comb = smul21b_12b_x_9b(p1_array_index_66961_comb, 9'h14b);
  assign p1_smul_67946_comb = smul21b_12b_x_9b(p1_array_index_66947_comb, 9'h0b5);
  assign p1_smul_67947_comb = smul21b_12b_x_9b(p1_array_index_66949_comb, 9'h0b5);
  assign p1_smul_67948_comb = smul21b_12b_x_9b(p1_array_index_66963_comb, 9'h14b);
  assign p1_smul_67949_comb = smul21b_12b_x_9b(p1_array_index_66965_comb, 9'h14b);
  assign p1_smul_67950_comb = smul21b_12b_x_9b(p1_array_index_66985_comb, 9'h0b5);
  assign p1_smul_28244_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66975_comb, 8'h47);
  assign p1_smul_67952_comb = smul21b_12b_x_9b(p1_array_index_66951_comb, 9'h105);
  assign p1_smul_67955_comb = smul21b_12b_x_9b(p1_array_index_66943_comb, 9'h0d5);
  assign p1_smul_67956_comb = smul21b_12b_x_9b(p1_array_index_66945_comb, 9'h0d5);
  assign p1_smul_67959_comb = smul21b_12b_x_9b(p1_array_index_66957_comb, 9'h105);
  assign p1_smul_28258_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66979_comb, 8'h47);
  assign p1_smul_28356_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66981_comb, 8'h47);
  assign p1_smul_67962_comb = smul21b_12b_x_9b(p1_array_index_66959_comb, 9'h105);
  assign p1_smul_67965_comb = smul21b_12b_x_9b(p1_array_index_66947_comb, 9'h0d5);
  assign p1_smul_67966_comb = smul21b_12b_x_9b(p1_array_index_66949_comb, 9'h0d5);
  assign p1_smul_67969_comb = smul21b_12b_x_9b(p1_array_index_66965_comb, 9'h105);
  assign p1_smul_28370_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66985_comb, 8'h47);
  assign p1_smul_28374_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66951_comb, 7'h45);
  assign p1_smul_28378_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66943_comb, 7'h3b);
  assign p1_smul_28380_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66945_comb, 7'h3b);
  assign p1_smul_28384_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66957_comb, 7'h45);
  assign p1_smul_28486_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66959_comb, 7'h45);
  assign p1_smul_28490_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66947_comb, 7'h3b);
  assign p1_smul_28492_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66949_comb, 7'h3b);
  assign p1_smul_28496_NarrowedMult__comb = smul19b_12b_x_7b(p1_array_index_66965_comb, 7'h45);
  assign p1_smul_28502_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66951_comb, 8'hb9);
  assign p1_smul_67998_comb = smul21b_12b_x_9b(p1_array_index_66953_comb, 9'h0d5);
  assign p1_smul_67999_comb = smul21b_12b_x_9b(p1_array_index_66943_comb, 9'h105);
  assign p1_smul_68000_comb = smul21b_12b_x_9b(p1_array_index_66945_comb, 9'h105);
  assign p1_smul_68001_comb = smul21b_12b_x_9b(p1_array_index_66955_comb, 9'h0d5);
  assign p1_smul_28512_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66957_comb, 8'hb9);
  assign p1_smul_28614_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66959_comb, 8'hb9);
  assign p1_smul_68008_comb = smul21b_12b_x_9b(p1_array_index_66961_comb, 9'h0d5);
  assign p1_smul_68009_comb = smul21b_12b_x_9b(p1_array_index_66947_comb, 9'h105);
  assign p1_smul_68010_comb = smul21b_12b_x_9b(p1_array_index_66949_comb, 9'h105);
  assign p1_smul_68011_comb = smul21b_12b_x_9b(p1_array_index_66963_comb, 9'h0d5);
  assign p1_smul_28624_NarrowedMult__comb = smul20b_12b_x_8b(p1_array_index_66965_comb, 8'hb9);
  assign p1_add_68847_comb = {{1{p1_array_index_66831_comb[11]}}, p1_array_index_66831_comb} + {{1{p1_array_index_66807_comb[11]}}, p1_array_index_66807_comb};
  assign p1_add_68848_comb = {{1{p1_array_index_66809_comb[11]}}, p1_array_index_66809_comb} + {{1{p1_array_index_66799_comb[11]}}, p1_array_index_66799_comb};
  assign p1_add_68849_comb = {{1{p1_array_index_66801_comb[11]}}, p1_array_index_66801_comb} + {{1{p1_array_index_66811_comb[11]}}, p1_array_index_66811_comb};
  assign p1_add_68850_comb = {{1{p1_array_index_66813_comb[11]}}, p1_array_index_66813_comb} + {{1{p1_array_index_66835_comb[11]}}, p1_array_index_66835_comb};
  assign p1_add_68851_comb = {{1{p1_array_index_66837_comb[11]}}, p1_array_index_66837_comb} + {{1{p1_array_index_66815_comb[11]}}, p1_array_index_66815_comb};
  assign p1_add_68852_comb = {{1{p1_array_index_66817_comb[11]}}, p1_array_index_66817_comb} + {{1{p1_array_index_66803_comb[11]}}, p1_array_index_66803_comb};
  assign p1_add_68853_comb = {{1{p1_array_index_66805_comb[11]}}, p1_array_index_66805_comb} + {{1{p1_array_index_66819_comb[11]}}, p1_array_index_66819_comb};
  assign p1_add_68854_comb = {{1{p1_array_index_66821_comb[11]}}, p1_array_index_66821_comb} + {{1{p1_array_index_66841_comb[11]}}, p1_array_index_66841_comb};
  assign p1_add_68967_comb = {{1{p1_array_index_66911_comb[11]}}, p1_array_index_66911_comb} + {{1{p1_array_index_66863_comb[11]}}, p1_array_index_66863_comb};
  assign p1_add_68968_comb = {{1{p1_array_index_66865_comb[11]}}, p1_array_index_66865_comb} + {{1{p1_array_index_66847_comb[11]}}, p1_array_index_66847_comb};
  assign p1_add_68969_comb = {{1{p1_array_index_66849_comb[11]}}, p1_array_index_66849_comb} + {{1{p1_array_index_66867_comb[11]}}, p1_array_index_66867_comb};
  assign p1_add_68970_comb = {{1{p1_array_index_66869_comb[11]}}, p1_array_index_66869_comb} + {{1{p1_array_index_66915_comb[11]}}, p1_array_index_66915_comb};
  assign p1_add_68971_comb = {{1{p1_array_index_66917_comb[11]}}, p1_array_index_66917_comb} + {{1{p1_array_index_66871_comb[11]}}, p1_array_index_66871_comb};
  assign p1_add_68972_comb = {{1{p1_array_index_66873_comb[11]}}, p1_array_index_66873_comb} + {{1{p1_array_index_66851_comb[11]}}, p1_array_index_66851_comb};
  assign p1_add_68973_comb = {{1{p1_array_index_66853_comb[11]}}, p1_array_index_66853_comb} + {{1{p1_array_index_66875_comb[11]}}, p1_array_index_66875_comb};
  assign p1_add_68974_comb = {{1{p1_array_index_66877_comb[11]}}, p1_array_index_66877_comb} + {{1{p1_array_index_66921_comb[11]}}, p1_array_index_66921_comb};
  assign p1_add_68975_comb = {{1{p1_array_index_66923_comb[11]}}, p1_array_index_66923_comb} + {{1{p1_array_index_66879_comb[11]}}, p1_array_index_66879_comb};
  assign p1_add_68976_comb = {{1{p1_array_index_66881_comb[11]}}, p1_array_index_66881_comb} + {{1{p1_array_index_66855_comb[11]}}, p1_array_index_66855_comb};
  assign p1_add_68977_comb = {{1{p1_array_index_66857_comb[11]}}, p1_array_index_66857_comb} + {{1{p1_array_index_66883_comb[11]}}, p1_array_index_66883_comb};
  assign p1_add_68978_comb = {{1{p1_array_index_66885_comb[11]}}, p1_array_index_66885_comb} + {{1{p1_array_index_66927_comb[11]}}, p1_array_index_66927_comb};
  assign p1_add_68979_comb = {{1{p1_array_index_66929_comb[11]}}, p1_array_index_66929_comb} + {{1{p1_array_index_66887_comb[11]}}, p1_array_index_66887_comb};
  assign p1_add_68980_comb = {{1{p1_array_index_66889_comb[11]}}, p1_array_index_66889_comb} + {{1{p1_array_index_66859_comb[11]}}, p1_array_index_66859_comb};
  assign p1_add_68981_comb = {{1{p1_array_index_66861_comb[11]}}, p1_array_index_66861_comb} + {{1{p1_array_index_66891_comb[11]}}, p1_array_index_66891_comb};
  assign p1_add_68982_comb = {{1{p1_array_index_66893_comb[11]}}, p1_array_index_66893_comb} + {{1{p1_array_index_66933_comb[11]}}, p1_array_index_66933_comb};
  assign p1_add_69207_comb = {{1{p1_array_index_66975_comb[11]}}, p1_array_index_66975_comb} + {{1{p1_array_index_66951_comb[11]}}, p1_array_index_66951_comb};
  assign p1_add_69208_comb = {{1{p1_array_index_66953_comb[11]}}, p1_array_index_66953_comb} + {{1{p1_array_index_66943_comb[11]}}, p1_array_index_66943_comb};
  assign p1_add_69209_comb = {{1{p1_array_index_66945_comb[11]}}, p1_array_index_66945_comb} + {{1{p1_array_index_66955_comb[11]}}, p1_array_index_66955_comb};
  assign p1_add_69210_comb = {{1{p1_array_index_66957_comb[11]}}, p1_array_index_66957_comb} + {{1{p1_array_index_66979_comb[11]}}, p1_array_index_66979_comb};
  assign p1_add_69211_comb = {{1{p1_array_index_66981_comb[11]}}, p1_array_index_66981_comb} + {{1{p1_array_index_66959_comb[11]}}, p1_array_index_66959_comb};
  assign p1_add_69212_comb = {{1{p1_array_index_66961_comb[11]}}, p1_array_index_66961_comb} + {{1{p1_array_index_66947_comb[11]}}, p1_array_index_66947_comb};
  assign p1_add_69213_comb = {{1{p1_array_index_66949_comb[11]}}, p1_array_index_66949_comb} + {{1{p1_array_index_66963_comb[11]}}, p1_array_index_66963_comb};
  assign p1_add_69214_comb = {{1{p1_array_index_66965_comb[11]}}, p1_array_index_66965_comb} + {{1{p1_array_index_66985_comb[11]}}, p1_array_index_66985_comb};
  assign p1_add_68037_comb = p1_smul_27786_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68038_comb = p1_smul_27788_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68051_comb = p1_smul_27802_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68052_comb = p1_smul_27804_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68061_comb = p1_smul_27910_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68062_comb = p1_smul_27912_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68067_comb = p1_smul_27918_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68068_comb = p1_smul_27920_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68073_comb = p1_smul_27926_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68074_comb = p1_smul_27928_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68079_comb = p1_smul_27934_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68080_comb = p1_smul_27936_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68085_comb = p1_smul_28038_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68094_comb = p1_smul_28048_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68099_comb = p1_smul_28054_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68108_comb = p1_smul_28064_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68147_comb = p1_smul_28296_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68152_comb = p1_smul_28302_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68161_comb = p1_smul_28312_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68166_comb = p1_smul_28318_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68171_comb = p1_smul_28420_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68174_comb = p1_smul_28424_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68179_comb = p1_smul_28430_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68182_comb = p1_smul_28434_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68183_comb = p1_smul_28436_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68186_comb = p1_smul_28440_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68191_comb = p1_smul_28446_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68194_comb = p1_smul_28450_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68195_comb = p1_smul_28548_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68208_comb = p1_smul_28562_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68209_comb = p1_smul_28564_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68222_comb = p1_smul_28578_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68261_comb = p1_smul_27754_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68262_comb = p1_smul_27756_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68275_comb = p1_smul_27770_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68276_comb = p1_smul_27772_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68289_comb = p1_smul_27818_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68290_comb = p1_smul_27820_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68303_comb = p1_smul_27834_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68304_comb = p1_smul_27836_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68313_comb = p1_smul_27878_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68314_comb = p1_smul_27880_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68319_comb = p1_smul_27886_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68320_comb = p1_smul_27888_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68325_comb = p1_smul_27894_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68326_comb = p1_smul_27896_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68331_comb = p1_smul_27902_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68332_comb = p1_smul_27904_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68337_comb = p1_smul_27942_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68338_comb = p1_smul_27944_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68343_comb = p1_smul_27950_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68344_comb = p1_smul_27952_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68349_comb = p1_smul_27958_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68350_comb = p1_smul_27960_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68355_comb = p1_smul_27966_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68356_comb = p1_smul_27968_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68361_comb = p1_smul_28006_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68370_comb = p1_smul_28016_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68375_comb = p1_smul_28022_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68384_comb = p1_smul_28032_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68389_comb = p1_smul_28070_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68398_comb = p1_smul_28080_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68403_comb = p1_smul_28086_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68412_comb = p1_smul_28096_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68483_comb = p1_smul_28264_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68488_comb = p1_smul_28270_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68497_comb = p1_smul_28280_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68502_comb = p1_smul_28286_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68511_comb = p1_smul_28328_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68516_comb = p1_smul_28334_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68525_comb = p1_smul_28344_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68530_comb = p1_smul_28350_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68535_comb = p1_smul_28388_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68538_comb = p1_smul_28392_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68543_comb = p1_smul_28398_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68546_comb = p1_smul_28402_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68547_comb = p1_smul_28404_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68550_comb = p1_smul_28408_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68555_comb = p1_smul_28414_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68558_comb = p1_smul_28418_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68559_comb = p1_smul_28452_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68562_comb = p1_smul_28456_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68567_comb = p1_smul_28462_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68570_comb = p1_smul_28466_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68571_comb = p1_smul_28468_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68574_comb = p1_smul_28472_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68579_comb = p1_smul_28478_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68582_comb = p1_smul_28482_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68583_comb = p1_smul_28516_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68596_comb = p1_smul_28530_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68597_comb = p1_smul_28532_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68610_comb = p1_smul_28546_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68611_comb = p1_smul_28580_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68624_comb = p1_smul_28594_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68625_comb = p1_smul_28596_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68638_comb = p1_smul_28610_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68661_comb = p1_smul_27738_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68662_comb = p1_smul_27740_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68675_comb = p1_smul_27850_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68676_comb = p1_smul_27852_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68685_comb = p1_smul_27862_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68686_comb = p1_smul_27864_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68691_comb = p1_smul_27870_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68692_comb = p1_smul_27872_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68697_comb = p1_smul_27974_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68698_comb = p1_smul_27976_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68703_comb = p1_smul_27982_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68704_comb = p1_smul_27984_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68709_comb = p1_smul_27990_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68718_comb = p1_smul_28000_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68723_comb = p1_smul_28102_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68732_comb = p1_smul_28112_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68771_comb = p1_smul_28248_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68776_comb = p1_smul_28254_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68785_comb = p1_smul_28360_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68790_comb = p1_smul_28366_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68795_comb = p1_smul_28372_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68798_comb = p1_smul_28376_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68803_comb = p1_smul_28382_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68806_comb = p1_smul_28386_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68807_comb = p1_smul_28484_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68810_comb = p1_smul_28488_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68815_comb = p1_smul_28494_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68818_comb = p1_smul_28498_NarrowedMult__comb[18:6] + 13'h0001;
  assign p1_add_68819_comb = p1_smul_28500_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68832_comb = p1_smul_28514_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68833_comb = p1_smul_28612_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_add_68846_comb = p1_smul_28626_NarrowedMult__comb[17:6] + 12'h001;
  assign p1_sum__961_comb = {{19{p1_add_68847_comb[12]}}, p1_add_68847_comb};
  assign p1_sum__962_comb = {{19{p1_add_68848_comb[12]}}, p1_add_68848_comb};
  assign p1_sum__963_comb = {{19{p1_add_68849_comb[12]}}, p1_add_68849_comb};
  assign p1_sum__964_comb = {{19{p1_add_68850_comb[12]}}, p1_add_68850_comb};
  assign p1_sum__926_comb = {{19{p1_add_68851_comb[12]}}, p1_add_68851_comb};
  assign p1_sum__927_comb = {{19{p1_add_68852_comb[12]}}, p1_add_68852_comb};
  assign p1_sum__928_comb = {{19{p1_add_68853_comb[12]}}, p1_add_68853_comb};
  assign p1_sum__929_comb = {{19{p1_add_68854_comb[12]}}, p1_add_68854_comb};
  assign p1_sum__1010_comb = {{19{p1_add_68967_comb[12]}}, p1_add_68967_comb};
  assign p1_sum__1011_comb = {{19{p1_add_68968_comb[12]}}, p1_add_68968_comb};
  assign p1_sum__1012_comb = {{19{p1_add_68969_comb[12]}}, p1_add_68969_comb};
  assign p1_sum__1013_comb = {{19{p1_add_68970_comb[12]}}, p1_add_68970_comb};
  assign p1_sum__989_comb = {{19{p1_add_68971_comb[12]}}, p1_add_68971_comb};
  assign p1_sum__990_comb = {{19{p1_add_68972_comb[12]}}, p1_add_68972_comb};
  assign p1_sum__991_comb = {{19{p1_add_68973_comb[12]}}, p1_add_68973_comb};
  assign p1_sum__992_comb = {{19{p1_add_68974_comb[12]}}, p1_add_68974_comb};
  assign p1_sum__884_comb = {{19{p1_add_68975_comb[12]}}, p1_add_68975_comb};
  assign p1_sum__885_comb = {{19{p1_add_68976_comb[12]}}, p1_add_68976_comb};
  assign p1_sum__886_comb = {{19{p1_add_68977_comb[12]}}, p1_add_68977_comb};
  assign p1_sum__887_comb = {{19{p1_add_68978_comb[12]}}, p1_add_68978_comb};
  assign p1_sum__835_comb = {{19{p1_add_68979_comb[12]}}, p1_add_68979_comb};
  assign p1_sum__836_comb = {{19{p1_add_68980_comb[12]}}, p1_add_68980_comb};
  assign p1_sum__837_comb = {{19{p1_add_68981_comb[12]}}, p1_add_68981_comb};
  assign p1_sum__838_comb = {{19{p1_add_68982_comb[12]}}, p1_add_68982_comb};
  assign p1_sum__1017_comb = {{19{p1_add_69207_comb[12]}}, p1_add_69207_comb};
  assign p1_sum__1018_comb = {{19{p1_add_69208_comb[12]}}, p1_add_69208_comb};
  assign p1_sum__1019_comb = {{19{p1_add_69209_comb[12]}}, p1_add_69209_comb};
  assign p1_sum__1020_comb = {{19{p1_add_69210_comb[12]}}, p1_add_69210_comb};
  assign p1_sum__779_comb = {{19{p1_add_69211_comb[12]}}, p1_add_69211_comb};
  assign p1_sum__780_comb = {{19{p1_add_69212_comb[12]}}, p1_add_69212_comb};
  assign p1_sum__781_comb = {{19{p1_add_69213_comb[12]}}, p1_add_69213_comb};
  assign p1_sum__782_comb = {{19{p1_add_69214_comb[12]}}, p1_add_69214_comb};
  assign p1_add_68855_comb = p1_smul_67439_comb[20:7] + 14'h0001;
  assign p1_add_68856_comb = p1_smul_67440_comb[20:7] + 14'h0001;
  assign p1_add_68857_comb = p1_smul_27784_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_68858_comb = p1_add_68037_comb[11:1];
  assign p1_bit_slice_68859_comb = p1_add_68038_comb[11:1];
  assign p1_add_68860_comb = p1_smul_27790_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68861_comb = p1_smul_67447_comb[20:7] + 14'h0001;
  assign p1_add_68862_comb = p1_smul_67448_comb[20:7] + 14'h0001;
  assign p1_add_68863_comb = p1_smul_67449_comb[20:7] + 14'h0001;
  assign p1_add_68864_comb = p1_smul_67450_comb[20:7] + 14'h0001;
  assign p1_add_68865_comb = p1_smul_27800_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_68866_comb = p1_add_68051_comb[11:1];
  assign p1_bit_slice_68867_comb = p1_add_68052_comb[11:1];
  assign p1_add_68868_comb = p1_smul_27806_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68869_comb = p1_smul_67457_comb[20:7] + 14'h0001;
  assign p1_add_68870_comb = p1_smul_67458_comb[20:7] + 14'h0001;
  assign p1_add_68871_comb = p1_smul_27908_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68872_comb = p1_add_68061_comb[12:1];
  assign p1_bit_slice_68873_comb = p1_add_68062_comb[12:1];
  assign p1_add_68874_comb = p1_smul_27914_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_68875_comb = p1_smul_27916_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68876_comb = p1_add_68067_comb[12:1];
  assign p1_bit_slice_68877_comb = p1_add_68068_comb[12:1];
  assign p1_add_68878_comb = p1_smul_27922_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_68879_comb = p1_smul_27924_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68880_comb = p1_add_68073_comb[12:1];
  assign p1_bit_slice_68881_comb = p1_add_68074_comb[12:1];
  assign p1_add_68882_comb = p1_smul_27930_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_68883_comb = p1_smul_27932_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68884_comb = p1_add_68079_comb[12:1];
  assign p1_bit_slice_68885_comb = p1_add_68080_comb[12:1];
  assign p1_add_68886_comb = p1_smul_27938_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_68887_comb = p1_smul_67483_comb[20:7] + 14'h0001;
  assign p1_bit_slice_68888_comb = p1_add_68085_comb[11:1];
  assign p1_add_68889_comb = p1_smul_67486_comb[20:7] + 14'h0001;
  assign p1_add_68890_comb = p1_smul_28042_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68891_comb = p1_smul_28044_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68892_comb = p1_smul_67489_comb[20:7] + 14'h0001;
  assign p1_bit_slice_68893_comb = p1_add_68094_comb[11:1];
  assign p1_add_68894_comb = p1_smul_67492_comb[20:7] + 14'h0001;
  assign p1_add_68895_comb = p1_smul_67493_comb[20:7] + 14'h0001;
  assign p1_bit_slice_68896_comb = p1_add_68099_comb[11:1];
  assign p1_add_68897_comb = p1_smul_67496_comb[20:7] + 14'h0001;
  assign p1_add_68898_comb = p1_smul_28058_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68899_comb = p1_smul_28060_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68900_comb = p1_smul_67499_comb[20:7] + 14'h0001;
  assign p1_bit_slice_68901_comb = p1_add_68108_comb[11:1];
  assign p1_add_68902_comb = p1_smul_67502_comb[20:7] + 14'h0001;
  assign p1_add_68903_comb = p1_smul_67503_comb[20:7] + 14'h0001;
  assign p1_add_68904_comb = p1_smul_67504_comb[20:7] + 14'h0001;
  assign p1_add_68905_comb = p1_smul_67505_comb[20:7] + 14'h0001;
  assign p1_add_68906_comb = p1_smul_67506_comb[20:7] + 14'h0001;
  assign p1_add_68907_comb = p1_smul_67507_comb[20:7] + 14'h0001;
  assign p1_add_68908_comb = p1_smul_67508_comb[20:7] + 14'h0001;
  assign p1_add_68909_comb = p1_smul_67509_comb[20:7] + 14'h0001;
  assign p1_add_68910_comb = p1_smul_67510_comb[20:7] + 14'h0001;
  assign p1_add_68911_comb = p1_smul_67511_comb[20:7] + 14'h0001;
  assign p1_add_68912_comb = p1_smul_67512_comb[20:7] + 14'h0001;
  assign p1_add_68913_comb = p1_smul_67513_comb[20:7] + 14'h0001;
  assign p1_add_68914_comb = p1_smul_67514_comb[20:7] + 14'h0001;
  assign p1_add_68915_comb = p1_smul_67515_comb[20:7] + 14'h0001;
  assign p1_add_68916_comb = p1_smul_67516_comb[20:7] + 14'h0001;
  assign p1_add_68917_comb = p1_smul_67517_comb[20:7] + 14'h0001;
  assign p1_add_68918_comb = p1_smul_67518_comb[20:7] + 14'h0001;
  assign p1_add_68919_comb = p1_smul_28292_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68920_comb = p1_smul_67520_comb[20:7] + 14'h0001;
  assign p1_bit_slice_68921_comb = p1_add_68147_comb[11:1];
  assign p1_add_68922_comb = p1_smul_67523_comb[20:7] + 14'h0001;
  assign p1_add_68923_comb = p1_smul_67524_comb[20:7] + 14'h0001;
  assign p1_bit_slice_68924_comb = p1_add_68152_comb[11:1];
  assign p1_add_68925_comb = p1_smul_67527_comb[20:7] + 14'h0001;
  assign p1_add_68926_comb = p1_smul_28306_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68927_comb = p1_smul_28308_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68928_comb = p1_smul_67530_comb[20:7] + 14'h0001;
  assign p1_bit_slice_68929_comb = p1_add_68161_comb[11:1];
  assign p1_add_68930_comb = p1_smul_67533_comb[20:7] + 14'h0001;
  assign p1_add_68931_comb = p1_smul_67534_comb[20:7] + 14'h0001;
  assign p1_bit_slice_68932_comb = p1_add_68166_comb[11:1];
  assign p1_add_68933_comb = p1_smul_67537_comb[20:7] + 14'h0001;
  assign p1_add_68934_comb = p1_smul_28322_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_68935_comb = p1_add_68171_comb[12:1];
  assign p1_add_68936_comb = p1_smul_28422_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68937_comb = p1_add_68174_comb[12:1];
  assign p1_add_68938_comb = p1_smul_28426_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_68939_comb = p1_smul_28428_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68940_comb = p1_add_68179_comb[12:1];
  assign p1_add_68941_comb = p1_smul_28432_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68942_comb = p1_add_68182_comb[12:1];
  assign p1_bit_slice_68943_comb = p1_add_68183_comb[12:1];
  assign p1_add_68944_comb = p1_smul_28438_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68945_comb = p1_add_68186_comb[12:1];
  assign p1_add_68946_comb = p1_smul_28442_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_68947_comb = p1_smul_28444_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68948_comb = p1_add_68191_comb[12:1];
  assign p1_add_68949_comb = p1_smul_28448_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_68950_comb = p1_add_68194_comb[12:1];
  assign p1_bit_slice_68951_comb = p1_add_68195_comb[11:1];
  assign p1_add_68952_comb = p1_smul_28550_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68953_comb = p1_smul_67566_comb[20:7] + 14'h0001;
  assign p1_add_68954_comb = p1_smul_67567_comb[20:7] + 14'h0001;
  assign p1_add_68955_comb = p1_smul_67568_comb[20:7] + 14'h0001;
  assign p1_add_68956_comb = p1_smul_67569_comb[20:7] + 14'h0001;
  assign p1_add_68957_comb = p1_smul_28560_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_68958_comb = p1_add_68208_comb[11:1];
  assign p1_bit_slice_68959_comb = p1_add_68209_comb[11:1];
  assign p1_add_68960_comb = p1_smul_28566_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68961_comb = p1_smul_67576_comb[20:7] + 14'h0001;
  assign p1_add_68962_comb = p1_smul_67577_comb[20:7] + 14'h0001;
  assign p1_add_68963_comb = p1_smul_67578_comb[20:7] + 14'h0001;
  assign p1_add_68964_comb = p1_smul_67579_comb[20:7] + 14'h0001;
  assign p1_add_68965_comb = p1_smul_28576_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_68966_comb = p1_add_68222_comb[11:1];
  assign p1_add_68983_comb = p1_smul_67583_comb[20:7] + 14'h0001;
  assign p1_add_68984_comb = p1_smul_67584_comb[20:7] + 14'h0001;
  assign p1_add_68985_comb = p1_smul_27752_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_68986_comb = p1_add_68261_comb[11:1];
  assign p1_bit_slice_68987_comb = p1_add_68262_comb[11:1];
  assign p1_add_68988_comb = p1_smul_27758_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68989_comb = p1_smul_67591_comb[20:7] + 14'h0001;
  assign p1_add_68990_comb = p1_smul_67592_comb[20:7] + 14'h0001;
  assign p1_add_68991_comb = p1_smul_67593_comb[20:7] + 14'h0001;
  assign p1_add_68992_comb = p1_smul_67594_comb[20:7] + 14'h0001;
  assign p1_add_68993_comb = p1_smul_27768_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_68994_comb = p1_add_68275_comb[11:1];
  assign p1_bit_slice_68995_comb = p1_add_68276_comb[11:1];
  assign p1_add_68996_comb = p1_smul_27774_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_68997_comb = p1_smul_67601_comb[20:7] + 14'h0001;
  assign p1_add_68998_comb = p1_smul_67602_comb[20:7] + 14'h0001;
  assign p1_add_68999_comb = p1_smul_67603_comb[20:7] + 14'h0001;
  assign p1_add_69000_comb = p1_smul_67604_comb[20:7] + 14'h0001;
  assign p1_add_69001_comb = p1_smul_27816_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69002_comb = p1_add_68289_comb[11:1];
  assign p1_bit_slice_69003_comb = p1_add_68290_comb[11:1];
  assign p1_add_69004_comb = p1_smul_27822_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69005_comb = p1_smul_67611_comb[20:7] + 14'h0001;
  assign p1_add_69006_comb = p1_smul_67612_comb[20:7] + 14'h0001;
  assign p1_add_69007_comb = p1_smul_67613_comb[20:7] + 14'h0001;
  assign p1_add_69008_comb = p1_smul_67614_comb[20:7] + 14'h0001;
  assign p1_add_69009_comb = p1_smul_27832_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69010_comb = p1_add_68303_comb[11:1];
  assign p1_bit_slice_69011_comb = p1_add_68304_comb[11:1];
  assign p1_add_69012_comb = p1_smul_27838_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69013_comb = p1_smul_67621_comb[20:7] + 14'h0001;
  assign p1_add_69014_comb = p1_smul_67622_comb[20:7] + 14'h0001;
  assign p1_add_69015_comb = p1_smul_27876_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69016_comb = p1_add_68313_comb[12:1];
  assign p1_bit_slice_69017_comb = p1_add_68314_comb[12:1];
  assign p1_add_69018_comb = p1_smul_27882_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69019_comb = p1_smul_27884_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69020_comb = p1_add_68319_comb[12:1];
  assign p1_bit_slice_69021_comb = p1_add_68320_comb[12:1];
  assign p1_add_69022_comb = p1_smul_27890_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69023_comb = p1_smul_27892_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69024_comb = p1_add_68325_comb[12:1];
  assign p1_bit_slice_69025_comb = p1_add_68326_comb[12:1];
  assign p1_add_69026_comb = p1_smul_27898_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69027_comb = p1_smul_27900_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69028_comb = p1_add_68331_comb[12:1];
  assign p1_bit_slice_69029_comb = p1_add_68332_comb[12:1];
  assign p1_add_69030_comb = p1_smul_27906_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69031_comb = p1_smul_27940_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69032_comb = p1_add_68337_comb[12:1];
  assign p1_bit_slice_69033_comb = p1_add_68338_comb[12:1];
  assign p1_add_69034_comb = p1_smul_27946_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69035_comb = p1_smul_27948_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69036_comb = p1_add_68343_comb[12:1];
  assign p1_bit_slice_69037_comb = p1_add_68344_comb[12:1];
  assign p1_add_69038_comb = p1_smul_27954_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69039_comb = p1_smul_27956_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69040_comb = p1_add_68349_comb[12:1];
  assign p1_bit_slice_69041_comb = p1_add_68350_comb[12:1];
  assign p1_add_69042_comb = p1_smul_27962_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69043_comb = p1_smul_27964_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69044_comb = p1_add_68355_comb[12:1];
  assign p1_bit_slice_69045_comb = p1_add_68356_comb[12:1];
  assign p1_add_69046_comb = p1_smul_27970_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69047_comb = p1_smul_67671_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69048_comb = p1_add_68361_comb[11:1];
  assign p1_add_69049_comb = p1_smul_67674_comb[20:7] + 14'h0001;
  assign p1_add_69050_comb = p1_smul_28010_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69051_comb = p1_smul_28012_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69052_comb = p1_smul_67677_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69053_comb = p1_add_68370_comb[11:1];
  assign p1_add_69054_comb = p1_smul_67680_comb[20:7] + 14'h0001;
  assign p1_add_69055_comb = p1_smul_67681_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69056_comb = p1_add_68375_comb[11:1];
  assign p1_add_69057_comb = p1_smul_67684_comb[20:7] + 14'h0001;
  assign p1_add_69058_comb = p1_smul_28026_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69059_comb = p1_smul_28028_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69060_comb = p1_smul_67687_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69061_comb = p1_add_68384_comb[11:1];
  assign p1_add_69062_comb = p1_smul_67690_comb[20:7] + 14'h0001;
  assign p1_add_69063_comb = p1_smul_67691_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69064_comb = p1_add_68389_comb[11:1];
  assign p1_add_69065_comb = p1_smul_67694_comb[20:7] + 14'h0001;
  assign p1_add_69066_comb = p1_smul_28074_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69067_comb = p1_smul_28076_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69068_comb = p1_smul_67697_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69069_comb = p1_add_68398_comb[11:1];
  assign p1_add_69070_comb = p1_smul_67700_comb[20:7] + 14'h0001;
  assign p1_add_69071_comb = p1_smul_67701_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69072_comb = p1_add_68403_comb[11:1];
  assign p1_add_69073_comb = p1_smul_67704_comb[20:7] + 14'h0001;
  assign p1_add_69074_comb = p1_smul_28090_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69075_comb = p1_smul_28092_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69076_comb = p1_smul_67707_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69077_comb = p1_add_68412_comb[11:1];
  assign p1_add_69078_comb = p1_smul_67710_comb[20:7] + 14'h0001;
  assign p1_add_69079_comb = p1_smul_67711_comb[20:7] + 14'h0001;
  assign p1_add_69080_comb = p1_smul_67712_comb[20:7] + 14'h0001;
  assign p1_add_69081_comb = p1_smul_67713_comb[20:7] + 14'h0001;
  assign p1_add_69082_comb = p1_smul_67714_comb[20:7] + 14'h0001;
  assign p1_add_69083_comb = p1_smul_67715_comb[20:7] + 14'h0001;
  assign p1_add_69084_comb = p1_smul_67716_comb[20:7] + 14'h0001;
  assign p1_add_69085_comb = p1_smul_67717_comb[20:7] + 14'h0001;
  assign p1_add_69086_comb = p1_smul_67718_comb[20:7] + 14'h0001;
  assign p1_add_69087_comb = p1_smul_67719_comb[20:7] + 14'h0001;
  assign p1_add_69088_comb = p1_smul_67720_comb[20:7] + 14'h0001;
  assign p1_add_69089_comb = p1_smul_67721_comb[20:7] + 14'h0001;
  assign p1_add_69090_comb = p1_smul_67722_comb[20:7] + 14'h0001;
  assign p1_add_69091_comb = p1_smul_67723_comb[20:7] + 14'h0001;
  assign p1_add_69092_comb = p1_smul_67724_comb[20:7] + 14'h0001;
  assign p1_add_69093_comb = p1_smul_67725_comb[20:7] + 14'h0001;
  assign p1_add_69094_comb = p1_smul_67726_comb[20:7] + 14'h0001;
  assign p1_add_69095_comb = p1_smul_67727_comb[20:7] + 14'h0001;
  assign p1_add_69096_comb = p1_smul_67728_comb[20:7] + 14'h0001;
  assign p1_add_69097_comb = p1_smul_67729_comb[20:7] + 14'h0001;
  assign p1_add_69098_comb = p1_smul_67730_comb[20:7] + 14'h0001;
  assign p1_add_69099_comb = p1_smul_67731_comb[20:7] + 14'h0001;
  assign p1_add_69100_comb = p1_smul_67732_comb[20:7] + 14'h0001;
  assign p1_add_69101_comb = p1_smul_67733_comb[20:7] + 14'h0001;
  assign p1_add_69102_comb = p1_smul_67734_comb[20:7] + 14'h0001;
  assign p1_add_69103_comb = p1_smul_67735_comb[20:7] + 14'h0001;
  assign p1_add_69104_comb = p1_smul_67736_comb[20:7] + 14'h0001;
  assign p1_add_69105_comb = p1_smul_67737_comb[20:7] + 14'h0001;
  assign p1_add_69106_comb = p1_smul_67738_comb[20:7] + 14'h0001;
  assign p1_add_69107_comb = p1_smul_67739_comb[20:7] + 14'h0001;
  assign p1_add_69108_comb = p1_smul_67740_comb[20:7] + 14'h0001;
  assign p1_add_69109_comb = p1_smul_67741_comb[20:7] + 14'h0001;
  assign p1_add_69110_comb = p1_smul_67742_comb[20:7] + 14'h0001;
  assign p1_add_69111_comb = p1_smul_28260_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69112_comb = p1_smul_67744_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69113_comb = p1_add_68483_comb[11:1];
  assign p1_add_69114_comb = p1_smul_67747_comb[20:7] + 14'h0001;
  assign p1_add_69115_comb = p1_smul_67748_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69116_comb = p1_add_68488_comb[11:1];
  assign p1_add_69117_comb = p1_smul_67751_comb[20:7] + 14'h0001;
  assign p1_add_69118_comb = p1_smul_28274_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69119_comb = p1_smul_28276_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69120_comb = p1_smul_67754_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69121_comb = p1_add_68497_comb[11:1];
  assign p1_add_69122_comb = p1_smul_67757_comb[20:7] + 14'h0001;
  assign p1_add_69123_comb = p1_smul_67758_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69124_comb = p1_add_68502_comb[11:1];
  assign p1_add_69125_comb = p1_smul_67761_comb[20:7] + 14'h0001;
  assign p1_add_69126_comb = p1_smul_28290_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69127_comb = p1_smul_28324_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69128_comb = p1_smul_67764_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69129_comb = p1_add_68511_comb[11:1];
  assign p1_add_69130_comb = p1_smul_67767_comb[20:7] + 14'h0001;
  assign p1_add_69131_comb = p1_smul_67768_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69132_comb = p1_add_68516_comb[11:1];
  assign p1_add_69133_comb = p1_smul_67771_comb[20:7] + 14'h0001;
  assign p1_add_69134_comb = p1_smul_28338_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69135_comb = p1_smul_28340_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69136_comb = p1_smul_67774_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69137_comb = p1_add_68525_comb[11:1];
  assign p1_add_69138_comb = p1_smul_67777_comb[20:7] + 14'h0001;
  assign p1_add_69139_comb = p1_smul_67778_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69140_comb = p1_add_68530_comb[11:1];
  assign p1_add_69141_comb = p1_smul_67781_comb[20:7] + 14'h0001;
  assign p1_add_69142_comb = p1_smul_28354_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69143_comb = p1_add_68535_comb[12:1];
  assign p1_add_69144_comb = p1_smul_28390_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69145_comb = p1_add_68538_comb[12:1];
  assign p1_add_69146_comb = p1_smul_28394_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69147_comb = p1_smul_28396_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69148_comb = p1_add_68543_comb[12:1];
  assign p1_add_69149_comb = p1_smul_28400_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69150_comb = p1_add_68546_comb[12:1];
  assign p1_bit_slice_69151_comb = p1_add_68547_comb[12:1];
  assign p1_add_69152_comb = p1_smul_28406_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69153_comb = p1_add_68550_comb[12:1];
  assign p1_add_69154_comb = p1_smul_28410_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69155_comb = p1_smul_28412_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69156_comb = p1_add_68555_comb[12:1];
  assign p1_add_69157_comb = p1_smul_28416_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69158_comb = p1_add_68558_comb[12:1];
  assign p1_bit_slice_69159_comb = p1_add_68559_comb[12:1];
  assign p1_add_69160_comb = p1_smul_28454_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69161_comb = p1_add_68562_comb[12:1];
  assign p1_add_69162_comb = p1_smul_28458_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69163_comb = p1_smul_28460_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69164_comb = p1_add_68567_comb[12:1];
  assign p1_add_69165_comb = p1_smul_28464_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69166_comb = p1_add_68570_comb[12:1];
  assign p1_bit_slice_69167_comb = p1_add_68571_comb[12:1];
  assign p1_add_69168_comb = p1_smul_28470_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69169_comb = p1_add_68574_comb[12:1];
  assign p1_add_69170_comb = p1_smul_28474_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69171_comb = p1_smul_28476_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69172_comb = p1_add_68579_comb[12:1];
  assign p1_add_69173_comb = p1_smul_28480_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69174_comb = p1_add_68582_comb[12:1];
  assign p1_bit_slice_69175_comb = p1_add_68583_comb[11:1];
  assign p1_add_69176_comb = p1_smul_28518_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69177_comb = p1_smul_67834_comb[20:7] + 14'h0001;
  assign p1_add_69178_comb = p1_smul_67835_comb[20:7] + 14'h0001;
  assign p1_add_69179_comb = p1_smul_67836_comb[20:7] + 14'h0001;
  assign p1_add_69180_comb = p1_smul_67837_comb[20:7] + 14'h0001;
  assign p1_add_69181_comb = p1_smul_28528_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69182_comb = p1_add_68596_comb[11:1];
  assign p1_bit_slice_69183_comb = p1_add_68597_comb[11:1];
  assign p1_add_69184_comb = p1_smul_28534_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69185_comb = p1_smul_67844_comb[20:7] + 14'h0001;
  assign p1_add_69186_comb = p1_smul_67845_comb[20:7] + 14'h0001;
  assign p1_add_69187_comb = p1_smul_67846_comb[20:7] + 14'h0001;
  assign p1_add_69188_comb = p1_smul_67847_comb[20:7] + 14'h0001;
  assign p1_add_69189_comb = p1_smul_28544_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69190_comb = p1_add_68610_comb[11:1];
  assign p1_bit_slice_69191_comb = p1_add_68611_comb[11:1];
  assign p1_add_69192_comb = p1_smul_28582_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69193_comb = p1_smul_67854_comb[20:7] + 14'h0001;
  assign p1_add_69194_comb = p1_smul_67855_comb[20:7] + 14'h0001;
  assign p1_add_69195_comb = p1_smul_67856_comb[20:7] + 14'h0001;
  assign p1_add_69196_comb = p1_smul_67857_comb[20:7] + 14'h0001;
  assign p1_add_69197_comb = p1_smul_28592_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69198_comb = p1_add_68624_comb[11:1];
  assign p1_bit_slice_69199_comb = p1_add_68625_comb[11:1];
  assign p1_add_69200_comb = p1_smul_28598_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69201_comb = p1_smul_67864_comb[20:7] + 14'h0001;
  assign p1_add_69202_comb = p1_smul_67865_comb[20:7] + 14'h0001;
  assign p1_add_69203_comb = p1_smul_67866_comb[20:7] + 14'h0001;
  assign p1_add_69204_comb = p1_smul_67867_comb[20:7] + 14'h0001;
  assign p1_add_69205_comb = p1_smul_28608_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69206_comb = p1_add_68638_comb[11:1];
  assign p1_add_69215_comb = p1_smul_67871_comb[20:7] + 14'h0001;
  assign p1_add_69216_comb = p1_smul_67872_comb[20:7] + 14'h0001;
  assign p1_add_69217_comb = p1_smul_27736_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69218_comb = p1_add_68661_comb[11:1];
  assign p1_bit_slice_69219_comb = p1_add_68662_comb[11:1];
  assign p1_add_69220_comb = p1_smul_27742_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69221_comb = p1_smul_67879_comb[20:7] + 14'h0001;
  assign p1_add_69222_comb = p1_smul_67880_comb[20:7] + 14'h0001;
  assign p1_add_69223_comb = p1_smul_67881_comb[20:7] + 14'h0001;
  assign p1_add_69224_comb = p1_smul_67882_comb[20:7] + 14'h0001;
  assign p1_add_69225_comb = p1_smul_27848_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69226_comb = p1_add_68675_comb[11:1];
  assign p1_bit_slice_69227_comb = p1_add_68676_comb[11:1];
  assign p1_add_69228_comb = p1_smul_27854_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69229_comb = p1_smul_67889_comb[20:7] + 14'h0001;
  assign p1_add_69230_comb = p1_smul_67890_comb[20:7] + 14'h0001;
  assign p1_add_69231_comb = p1_smul_27860_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69232_comb = p1_add_68685_comb[12:1];
  assign p1_bit_slice_69233_comb = p1_add_68686_comb[12:1];
  assign p1_add_69234_comb = p1_smul_27866_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69235_comb = p1_smul_27868_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69236_comb = p1_add_68691_comb[12:1];
  assign p1_bit_slice_69237_comb = p1_add_68692_comb[12:1];
  assign p1_add_69238_comb = p1_smul_27874_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69239_comb = p1_smul_27972_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69240_comb = p1_add_68697_comb[12:1];
  assign p1_bit_slice_69241_comb = p1_add_68698_comb[12:1];
  assign p1_add_69242_comb = p1_smul_27978_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69243_comb = p1_smul_27980_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69244_comb = p1_add_68703_comb[12:1];
  assign p1_bit_slice_69245_comb = p1_add_68704_comb[12:1];
  assign p1_add_69246_comb = p1_smul_27986_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69247_comb = p1_smul_67915_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69248_comb = p1_add_68709_comb[11:1];
  assign p1_add_69249_comb = p1_smul_67918_comb[20:7] + 14'h0001;
  assign p1_add_69250_comb = p1_smul_27994_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69251_comb = p1_smul_27996_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69252_comb = p1_smul_67921_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69253_comb = p1_add_68718_comb[11:1];
  assign p1_add_69254_comb = p1_smul_67924_comb[20:7] + 14'h0001;
  assign p1_add_69255_comb = p1_smul_67925_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69256_comb = p1_add_68723_comb[11:1];
  assign p1_add_69257_comb = p1_smul_67928_comb[20:7] + 14'h0001;
  assign p1_add_69258_comb = p1_smul_28106_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69259_comb = p1_smul_28108_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69260_comb = p1_smul_67931_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69261_comb = p1_add_68732_comb[11:1];
  assign p1_add_69262_comb = p1_smul_67934_comb[20:7] + 14'h0001;
  assign p1_add_69263_comb = p1_smul_67935_comb[20:7] + 14'h0001;
  assign p1_add_69264_comb = p1_smul_67936_comb[20:7] + 14'h0001;
  assign p1_add_69265_comb = p1_smul_67937_comb[20:7] + 14'h0001;
  assign p1_add_69266_comb = p1_smul_67938_comb[20:7] + 14'h0001;
  assign p1_add_69267_comb = p1_smul_67939_comb[20:7] + 14'h0001;
  assign p1_add_69268_comb = p1_smul_67940_comb[20:7] + 14'h0001;
  assign p1_add_69269_comb = p1_smul_67941_comb[20:7] + 14'h0001;
  assign p1_add_69270_comb = p1_smul_67942_comb[20:7] + 14'h0001;
  assign p1_add_69271_comb = p1_smul_67943_comb[20:7] + 14'h0001;
  assign p1_add_69272_comb = p1_smul_67944_comb[20:7] + 14'h0001;
  assign p1_add_69273_comb = p1_smul_67945_comb[20:7] + 14'h0001;
  assign p1_add_69274_comb = p1_smul_67946_comb[20:7] + 14'h0001;
  assign p1_add_69275_comb = p1_smul_67947_comb[20:7] + 14'h0001;
  assign p1_add_69276_comb = p1_smul_67948_comb[20:7] + 14'h0001;
  assign p1_add_69277_comb = p1_smul_67949_comb[20:7] + 14'h0001;
  assign p1_add_69278_comb = p1_smul_67950_comb[20:7] + 14'h0001;
  assign p1_add_69279_comb = p1_smul_28244_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69280_comb = p1_smul_67952_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69281_comb = p1_add_68771_comb[11:1];
  assign p1_add_69282_comb = p1_smul_67955_comb[20:7] + 14'h0001;
  assign p1_add_69283_comb = p1_smul_67956_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69284_comb = p1_add_68776_comb[11:1];
  assign p1_add_69285_comb = p1_smul_67959_comb[20:7] + 14'h0001;
  assign p1_add_69286_comb = p1_smul_28258_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69287_comb = p1_smul_28356_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69288_comb = p1_smul_67962_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69289_comb = p1_add_68785_comb[11:1];
  assign p1_add_69290_comb = p1_smul_67965_comb[20:7] + 14'h0001;
  assign p1_add_69291_comb = p1_smul_67966_comb[20:7] + 14'h0001;
  assign p1_bit_slice_69292_comb = p1_add_68790_comb[11:1];
  assign p1_add_69293_comb = p1_smul_67969_comb[20:7] + 14'h0001;
  assign p1_add_69294_comb = p1_smul_28370_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69295_comb = p1_add_68795_comb[12:1];
  assign p1_add_69296_comb = p1_smul_28374_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69297_comb = p1_add_68798_comb[12:1];
  assign p1_add_69298_comb = p1_smul_28378_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69299_comb = p1_smul_28380_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69300_comb = p1_add_68803_comb[12:1];
  assign p1_add_69301_comb = p1_smul_28384_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69302_comb = p1_add_68806_comb[12:1];
  assign p1_bit_slice_69303_comb = p1_add_68807_comb[12:1];
  assign p1_add_69304_comb = p1_smul_28486_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69305_comb = p1_add_68810_comb[12:1];
  assign p1_add_69306_comb = p1_smul_28490_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_add_69307_comb = p1_smul_28492_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69308_comb = p1_add_68815_comb[12:1];
  assign p1_add_69309_comb = p1_smul_28496_NarrowedMult__comb[18:5] + 14'h0001;
  assign p1_bit_slice_69310_comb = p1_add_68818_comb[12:1];
  assign p1_bit_slice_69311_comb = p1_add_68819_comb[11:1];
  assign p1_add_69312_comb = p1_smul_28502_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69313_comb = p1_smul_67998_comb[20:7] + 14'h0001;
  assign p1_add_69314_comb = p1_smul_67999_comb[20:7] + 14'h0001;
  assign p1_add_69315_comb = p1_smul_68000_comb[20:7] + 14'h0001;
  assign p1_add_69316_comb = p1_smul_68001_comb[20:7] + 14'h0001;
  assign p1_add_69317_comb = p1_smul_28512_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69318_comb = p1_add_68832_comb[11:1];
  assign p1_bit_slice_69319_comb = p1_add_68833_comb[11:1];
  assign p1_add_69320_comb = p1_smul_28614_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_add_69321_comb = p1_smul_68008_comb[20:7] + 14'h0001;
  assign p1_add_69322_comb = p1_smul_68009_comb[20:7] + 14'h0001;
  assign p1_add_69323_comb = p1_smul_68010_comb[20:7] + 14'h0001;
  assign p1_add_69324_comb = p1_smul_68011_comb[20:7] + 14'h0001;
  assign p1_add_69325_comb = p1_smul_28624_NarrowedMult__comb[19:6] + 14'h0001;
  assign p1_bit_slice_69326_comb = p1_add_68846_comb[11:1];
  assign p1_sum__965_comb = p1_sum__961_comb + p1_sum__962_comb;
  assign p1_sum__966_comb = p1_sum__963_comb + p1_sum__964_comb;
  assign p1_sum__930_comb = p1_sum__926_comb + p1_sum__927_comb;
  assign p1_sum__931_comb = p1_sum__928_comb + p1_sum__929_comb;
  assign p1_sum__1014_comb = p1_sum__1010_comb + p1_sum__1011_comb;
  assign p1_sum__1015_comb = p1_sum__1012_comb + p1_sum__1013_comb;
  assign p1_sum__993_comb = p1_sum__989_comb + p1_sum__990_comb;
  assign p1_sum__994_comb = p1_sum__991_comb + p1_sum__992_comb;
  assign p1_sum__888_comb = p1_sum__884_comb + p1_sum__885_comb;
  assign p1_sum__889_comb = p1_sum__886_comb + p1_sum__887_comb;
  assign p1_sum__839_comb = p1_sum__835_comb + p1_sum__836_comb;
  assign p1_sum__840_comb = p1_sum__837_comb + p1_sum__838_comb;
  assign p1_sum__1021_comb = p1_sum__1017_comb + p1_sum__1018_comb;
  assign p1_sum__1022_comb = p1_sum__1019_comb + p1_sum__1020_comb;
  assign p1_sum__783_comb = p1_sum__779_comb + p1_sum__780_comb;
  assign p1_sum__784_comb = p1_sum__781_comb + p1_sum__782_comb;
  assign p1_sum__967_comb = p1_sum__965_comb + p1_sum__966_comb;
  assign p1_sum__932_comb = p1_sum__930_comb + p1_sum__931_comb;
  assign p1_sum__1016_comb = p1_sum__1014_comb + p1_sum__1015_comb;
  assign p1_sum__995_comb = p1_sum__993_comb + p1_sum__994_comb;
  assign p1_sum__890_comb = p1_sum__888_comb + p1_sum__889_comb;
  assign p1_sum__841_comb = p1_sum__839_comb + p1_sum__840_comb;
  assign p1_sum__1023_comb = p1_sum__1021_comb + p1_sum__1022_comb;
  assign p1_sum__785_comb = p1_sum__783_comb + p1_sum__784_comb;
  assign p1_add_69811_comb = p1_add_68855_comb[13:1] + p1_add_68856_comb[13:1];
  assign p1_add_69812_comb = p1_add_68857_comb[13:1] + {{2{p1_bit_slice_68858_comb[10]}}, p1_bit_slice_68858_comb};
  assign p1_add_69813_comb = {{2{p1_bit_slice_68859_comb[10]}}, p1_bit_slice_68859_comb} + p1_add_68860_comb[13:1];
  assign p1_add_69814_comb = p1_add_68861_comb[13:1] + p1_add_68862_comb[13:1];
  assign p1_add_69815_comb = p1_add_68863_comb[13:1] + p1_add_68864_comb[13:1];
  assign p1_add_69816_comb = p1_add_68865_comb[13:1] + {{2{p1_bit_slice_68866_comb[10]}}, p1_bit_slice_68866_comb};
  assign p1_add_69817_comb = {{2{p1_bit_slice_68867_comb[10]}}, p1_bit_slice_68867_comb} + p1_add_68868_comb[13:1];
  assign p1_add_69818_comb = p1_add_68869_comb[13:1] + p1_add_68870_comb[13:1];
  assign p1_add_69819_comb = p1_add_68871_comb[13:1] + {{1{p1_bit_slice_68872_comb[11]}}, p1_bit_slice_68872_comb};
  assign p1_add_69820_comb = {{1{p1_bit_slice_68873_comb[11]}}, p1_bit_slice_68873_comb} + p1_add_68874_comb[13:1];
  assign p1_add_69821_comb = p1_add_68875_comb[13:1] + {{1{p1_bit_slice_68876_comb[11]}}, p1_bit_slice_68876_comb};
  assign p1_add_69822_comb = {{1{p1_bit_slice_68877_comb[11]}}, p1_bit_slice_68877_comb} + p1_add_68878_comb[13:1];
  assign p1_add_69823_comb = p1_add_68879_comb[13:1] + {{1{p1_bit_slice_68880_comb[11]}}, p1_bit_slice_68880_comb};
  assign p1_add_69824_comb = {{1{p1_bit_slice_68881_comb[11]}}, p1_bit_slice_68881_comb} + p1_add_68882_comb[13:1];
  assign p1_add_69825_comb = p1_add_68883_comb[13:1] + {{1{p1_bit_slice_68884_comb[11]}}, p1_bit_slice_68884_comb};
  assign p1_add_69826_comb = {{1{p1_bit_slice_68885_comb[11]}}, p1_bit_slice_68885_comb} + p1_add_68886_comb[13:1];
  assign p1_add_69827_comb = p1_add_68887_comb[13:1] + {{2{p1_bit_slice_68888_comb[10]}}, p1_bit_slice_68888_comb};
  assign p1_add_69828_comb = p1_add_68889_comb[13:1] + p1_add_68890_comb[13:1];
  assign p1_add_69829_comb = p1_add_68891_comb[13:1] + p1_add_68892_comb[13:1];
  assign p1_add_69830_comb = {{2{p1_bit_slice_68893_comb[10]}}, p1_bit_slice_68893_comb} + p1_add_68894_comb[13:1];
  assign p1_add_69831_comb = p1_add_68895_comb[13:1] + {{2{p1_bit_slice_68896_comb[10]}}, p1_bit_slice_68896_comb};
  assign p1_add_69832_comb = p1_add_68897_comb[13:1] + p1_add_68898_comb[13:1];
  assign p1_add_69833_comb = p1_add_68899_comb[13:1] + p1_add_68900_comb[13:1];
  assign p1_add_69834_comb = {{2{p1_bit_slice_68901_comb[10]}}, p1_bit_slice_68901_comb} + p1_add_68902_comb[13:1];
  assign p1_add_69835_comb = p1_add_68903_comb[13:1] + p1_add_68904_comb[13:1];
  assign p1_add_69836_comb = p1_add_68905_comb[13:1] + p1_add_68906_comb[13:1];
  assign p1_add_69837_comb = p1_add_68907_comb[13:1] + p1_add_68908_comb[13:1];
  assign p1_add_69838_comb = p1_add_68909_comb[13:1] + p1_add_68910_comb[13:1];
  assign p1_add_69839_comb = p1_add_68911_comb[13:1] + p1_add_68912_comb[13:1];
  assign p1_add_69840_comb = p1_add_68913_comb[13:1] + p1_add_68914_comb[13:1];
  assign p1_add_69841_comb = p1_add_68915_comb[13:1] + p1_add_68916_comb[13:1];
  assign p1_add_69842_comb = p1_add_68917_comb[13:1] + p1_add_68918_comb[13:1];
  assign p1_add_69843_comb = p1_add_68919_comb[13:1] + p1_add_68920_comb[13:1];
  assign p1_add_69844_comb = {{2{p1_bit_slice_68921_comb[10]}}, p1_bit_slice_68921_comb} + p1_add_68922_comb[13:1];
  assign p1_add_69845_comb = p1_add_68923_comb[13:1] + {{2{p1_bit_slice_68924_comb[10]}}, p1_bit_slice_68924_comb};
  assign p1_add_69846_comb = p1_add_68925_comb[13:1] + p1_add_68926_comb[13:1];
  assign p1_add_69847_comb = p1_add_68927_comb[13:1] + p1_add_68928_comb[13:1];
  assign p1_add_69848_comb = {{2{p1_bit_slice_68929_comb[10]}}, p1_bit_slice_68929_comb} + p1_add_68930_comb[13:1];
  assign p1_add_69849_comb = p1_add_68931_comb[13:1] + {{2{p1_bit_slice_68932_comb[10]}}, p1_bit_slice_68932_comb};
  assign p1_add_69850_comb = p1_add_68933_comb[13:1] + p1_add_68934_comb[13:1];
  assign p1_add_69851_comb = {{1{p1_bit_slice_68935_comb[11]}}, p1_bit_slice_68935_comb} + p1_add_68936_comb[13:1];
  assign p1_add_69852_comb = {{1{p1_bit_slice_68937_comb[11]}}, p1_bit_slice_68937_comb} + p1_add_68938_comb[13:1];
  assign p1_add_69853_comb = p1_add_68939_comb[13:1] + {{1{p1_bit_slice_68940_comb[11]}}, p1_bit_slice_68940_comb};
  assign p1_add_69854_comb = p1_add_68941_comb[13:1] + {{1{p1_bit_slice_68942_comb[11]}}, p1_bit_slice_68942_comb};
  assign p1_add_69855_comb = {{1{p1_bit_slice_68943_comb[11]}}, p1_bit_slice_68943_comb} + p1_add_68944_comb[13:1];
  assign p1_add_69856_comb = {{1{p1_bit_slice_68945_comb[11]}}, p1_bit_slice_68945_comb} + p1_add_68946_comb[13:1];
  assign p1_add_69857_comb = p1_add_68947_comb[13:1] + {{1{p1_bit_slice_68948_comb[11]}}, p1_bit_slice_68948_comb};
  assign p1_add_69858_comb = p1_add_68949_comb[13:1] + {{1{p1_bit_slice_68950_comb[11]}}, p1_bit_slice_68950_comb};
  assign p1_add_69859_comb = {{2{p1_bit_slice_68951_comb[10]}}, p1_bit_slice_68951_comb} + p1_add_68952_comb[13:1];
  assign p1_add_69860_comb = p1_add_68953_comb[13:1] + p1_add_68954_comb[13:1];
  assign p1_add_69861_comb = p1_add_68955_comb[13:1] + p1_add_68956_comb[13:1];
  assign p1_add_69862_comb = p1_add_68957_comb[13:1] + {{2{p1_bit_slice_68958_comb[10]}}, p1_bit_slice_68958_comb};
  assign p1_add_69863_comb = {{2{p1_bit_slice_68959_comb[10]}}, p1_bit_slice_68959_comb} + p1_add_68960_comb[13:1];
  assign p1_add_69864_comb = p1_add_68961_comb[13:1] + p1_add_68962_comb[13:1];
  assign p1_add_69865_comb = p1_add_68963_comb[13:1] + p1_add_68964_comb[13:1];
  assign p1_add_69866_comb = p1_add_68965_comb[13:1] + {{2{p1_bit_slice_68966_comb[10]}}, p1_bit_slice_68966_comb};
  assign p1_add_69875_comb = p1_add_68983_comb[13:1] + p1_add_68984_comb[13:1];
  assign p1_add_69876_comb = p1_add_68985_comb[13:1] + {{2{p1_bit_slice_68986_comb[10]}}, p1_bit_slice_68986_comb};
  assign p1_add_69877_comb = {{2{p1_bit_slice_68987_comb[10]}}, p1_bit_slice_68987_comb} + p1_add_68988_comb[13:1];
  assign p1_add_69878_comb = p1_add_68989_comb[13:1] + p1_add_68990_comb[13:1];
  assign p1_add_69879_comb = p1_add_68991_comb[13:1] + p1_add_68992_comb[13:1];
  assign p1_add_69880_comb = p1_add_68993_comb[13:1] + {{2{p1_bit_slice_68994_comb[10]}}, p1_bit_slice_68994_comb};
  assign p1_add_69881_comb = {{2{p1_bit_slice_68995_comb[10]}}, p1_bit_slice_68995_comb} + p1_add_68996_comb[13:1];
  assign p1_add_69882_comb = p1_add_68997_comb[13:1] + p1_add_68998_comb[13:1];
  assign p1_add_69883_comb = p1_add_68999_comb[13:1] + p1_add_69000_comb[13:1];
  assign p1_add_69884_comb = p1_add_69001_comb[13:1] + {{2{p1_bit_slice_69002_comb[10]}}, p1_bit_slice_69002_comb};
  assign p1_add_69885_comb = {{2{p1_bit_slice_69003_comb[10]}}, p1_bit_slice_69003_comb} + p1_add_69004_comb[13:1];
  assign p1_add_69886_comb = p1_add_69005_comb[13:1] + p1_add_69006_comb[13:1];
  assign p1_add_69887_comb = p1_add_69007_comb[13:1] + p1_add_69008_comb[13:1];
  assign p1_add_69888_comb = p1_add_69009_comb[13:1] + {{2{p1_bit_slice_69010_comb[10]}}, p1_bit_slice_69010_comb};
  assign p1_add_69889_comb = {{2{p1_bit_slice_69011_comb[10]}}, p1_bit_slice_69011_comb} + p1_add_69012_comb[13:1];
  assign p1_add_69890_comb = p1_add_69013_comb[13:1] + p1_add_69014_comb[13:1];
  assign p1_add_69891_comb = p1_add_69015_comb[13:1] + {{1{p1_bit_slice_69016_comb[11]}}, p1_bit_slice_69016_comb};
  assign p1_add_69892_comb = {{1{p1_bit_slice_69017_comb[11]}}, p1_bit_slice_69017_comb} + p1_add_69018_comb[13:1];
  assign p1_add_69893_comb = p1_add_69019_comb[13:1] + {{1{p1_bit_slice_69020_comb[11]}}, p1_bit_slice_69020_comb};
  assign p1_add_69894_comb = {{1{p1_bit_slice_69021_comb[11]}}, p1_bit_slice_69021_comb} + p1_add_69022_comb[13:1];
  assign p1_add_69895_comb = p1_add_69023_comb[13:1] + {{1{p1_bit_slice_69024_comb[11]}}, p1_bit_slice_69024_comb};
  assign p1_add_69896_comb = {{1{p1_bit_slice_69025_comb[11]}}, p1_bit_slice_69025_comb} + p1_add_69026_comb[13:1];
  assign p1_add_69897_comb = p1_add_69027_comb[13:1] + {{1{p1_bit_slice_69028_comb[11]}}, p1_bit_slice_69028_comb};
  assign p1_add_69898_comb = {{1{p1_bit_slice_69029_comb[11]}}, p1_bit_slice_69029_comb} + p1_add_69030_comb[13:1];
  assign p1_add_69899_comb = p1_add_69031_comb[13:1] + {{1{p1_bit_slice_69032_comb[11]}}, p1_bit_slice_69032_comb};
  assign p1_add_69900_comb = {{1{p1_bit_slice_69033_comb[11]}}, p1_bit_slice_69033_comb} + p1_add_69034_comb[13:1];
  assign p1_add_69901_comb = p1_add_69035_comb[13:1] + {{1{p1_bit_slice_69036_comb[11]}}, p1_bit_slice_69036_comb};
  assign p1_add_69902_comb = {{1{p1_bit_slice_69037_comb[11]}}, p1_bit_slice_69037_comb} + p1_add_69038_comb[13:1];
  assign p1_add_69903_comb = p1_add_69039_comb[13:1] + {{1{p1_bit_slice_69040_comb[11]}}, p1_bit_slice_69040_comb};
  assign p1_add_69904_comb = {{1{p1_bit_slice_69041_comb[11]}}, p1_bit_slice_69041_comb} + p1_add_69042_comb[13:1];
  assign p1_add_69905_comb = p1_add_69043_comb[13:1] + {{1{p1_bit_slice_69044_comb[11]}}, p1_bit_slice_69044_comb};
  assign p1_add_69906_comb = {{1{p1_bit_slice_69045_comb[11]}}, p1_bit_slice_69045_comb} + p1_add_69046_comb[13:1];
  assign p1_add_69907_comb = p1_add_69047_comb[13:1] + {{2{p1_bit_slice_69048_comb[10]}}, p1_bit_slice_69048_comb};
  assign p1_add_69908_comb = p1_add_69049_comb[13:1] + p1_add_69050_comb[13:1];
  assign p1_add_69909_comb = p1_add_69051_comb[13:1] + p1_add_69052_comb[13:1];
  assign p1_add_69910_comb = {{2{p1_bit_slice_69053_comb[10]}}, p1_bit_slice_69053_comb} + p1_add_69054_comb[13:1];
  assign p1_add_69911_comb = p1_add_69055_comb[13:1] + {{2{p1_bit_slice_69056_comb[10]}}, p1_bit_slice_69056_comb};
  assign p1_add_69912_comb = p1_add_69057_comb[13:1] + p1_add_69058_comb[13:1];
  assign p1_add_69913_comb = p1_add_69059_comb[13:1] + p1_add_69060_comb[13:1];
  assign p1_add_69914_comb = {{2{p1_bit_slice_69061_comb[10]}}, p1_bit_slice_69061_comb} + p1_add_69062_comb[13:1];
  assign p1_add_69915_comb = p1_add_69063_comb[13:1] + {{2{p1_bit_slice_69064_comb[10]}}, p1_bit_slice_69064_comb};
  assign p1_add_69916_comb = p1_add_69065_comb[13:1] + p1_add_69066_comb[13:1];
  assign p1_add_69917_comb = p1_add_69067_comb[13:1] + p1_add_69068_comb[13:1];
  assign p1_add_69918_comb = {{2{p1_bit_slice_69069_comb[10]}}, p1_bit_slice_69069_comb} + p1_add_69070_comb[13:1];
  assign p1_add_69919_comb = p1_add_69071_comb[13:1] + {{2{p1_bit_slice_69072_comb[10]}}, p1_bit_slice_69072_comb};
  assign p1_add_69920_comb = p1_add_69073_comb[13:1] + p1_add_69074_comb[13:1];
  assign p1_add_69921_comb = p1_add_69075_comb[13:1] + p1_add_69076_comb[13:1];
  assign p1_add_69922_comb = {{2{p1_bit_slice_69077_comb[10]}}, p1_bit_slice_69077_comb} + p1_add_69078_comb[13:1];
  assign p1_add_69923_comb = p1_add_69079_comb[13:1] + p1_add_69080_comb[13:1];
  assign p1_add_69924_comb = p1_add_69081_comb[13:1] + p1_add_69082_comb[13:1];
  assign p1_add_69925_comb = p1_add_69083_comb[13:1] + p1_add_69084_comb[13:1];
  assign p1_add_69926_comb = p1_add_69085_comb[13:1] + p1_add_69086_comb[13:1];
  assign p1_add_69927_comb = p1_add_69087_comb[13:1] + p1_add_69088_comb[13:1];
  assign p1_add_69928_comb = p1_add_69089_comb[13:1] + p1_add_69090_comb[13:1];
  assign p1_add_69929_comb = p1_add_69091_comb[13:1] + p1_add_69092_comb[13:1];
  assign p1_add_69930_comb = p1_add_69093_comb[13:1] + p1_add_69094_comb[13:1];
  assign p1_add_69931_comb = p1_add_69095_comb[13:1] + p1_add_69096_comb[13:1];
  assign p1_add_69932_comb = p1_add_69097_comb[13:1] + p1_add_69098_comb[13:1];
  assign p1_add_69933_comb = p1_add_69099_comb[13:1] + p1_add_69100_comb[13:1];
  assign p1_add_69934_comb = p1_add_69101_comb[13:1] + p1_add_69102_comb[13:1];
  assign p1_add_69935_comb = p1_add_69103_comb[13:1] + p1_add_69104_comb[13:1];
  assign p1_add_69936_comb = p1_add_69105_comb[13:1] + p1_add_69106_comb[13:1];
  assign p1_add_69937_comb = p1_add_69107_comb[13:1] + p1_add_69108_comb[13:1];
  assign p1_add_69938_comb = p1_add_69109_comb[13:1] + p1_add_69110_comb[13:1];
  assign p1_add_69939_comb = p1_add_69111_comb[13:1] + p1_add_69112_comb[13:1];
  assign p1_add_69940_comb = {{2{p1_bit_slice_69113_comb[10]}}, p1_bit_slice_69113_comb} + p1_add_69114_comb[13:1];
  assign p1_add_69941_comb = p1_add_69115_comb[13:1] + {{2{p1_bit_slice_69116_comb[10]}}, p1_bit_slice_69116_comb};
  assign p1_add_69942_comb = p1_add_69117_comb[13:1] + p1_add_69118_comb[13:1];
  assign p1_add_69943_comb = p1_add_69119_comb[13:1] + p1_add_69120_comb[13:1];
  assign p1_add_69944_comb = {{2{p1_bit_slice_69121_comb[10]}}, p1_bit_slice_69121_comb} + p1_add_69122_comb[13:1];
  assign p1_add_69945_comb = p1_add_69123_comb[13:1] + {{2{p1_bit_slice_69124_comb[10]}}, p1_bit_slice_69124_comb};
  assign p1_add_69946_comb = p1_add_69125_comb[13:1] + p1_add_69126_comb[13:1];
  assign p1_add_69947_comb = p1_add_69127_comb[13:1] + p1_add_69128_comb[13:1];
  assign p1_add_69948_comb = {{2{p1_bit_slice_69129_comb[10]}}, p1_bit_slice_69129_comb} + p1_add_69130_comb[13:1];
  assign p1_add_69949_comb = p1_add_69131_comb[13:1] + {{2{p1_bit_slice_69132_comb[10]}}, p1_bit_slice_69132_comb};
  assign p1_add_69950_comb = p1_add_69133_comb[13:1] + p1_add_69134_comb[13:1];
  assign p1_add_69951_comb = p1_add_69135_comb[13:1] + p1_add_69136_comb[13:1];
  assign p1_add_69952_comb = {{2{p1_bit_slice_69137_comb[10]}}, p1_bit_slice_69137_comb} + p1_add_69138_comb[13:1];
  assign p1_add_69953_comb = p1_add_69139_comb[13:1] + {{2{p1_bit_slice_69140_comb[10]}}, p1_bit_slice_69140_comb};
  assign p1_add_69954_comb = p1_add_69141_comb[13:1] + p1_add_69142_comb[13:1];
  assign p1_add_69955_comb = {{1{p1_bit_slice_69143_comb[11]}}, p1_bit_slice_69143_comb} + p1_add_69144_comb[13:1];
  assign p1_add_69956_comb = {{1{p1_bit_slice_69145_comb[11]}}, p1_bit_slice_69145_comb} + p1_add_69146_comb[13:1];
  assign p1_add_69957_comb = p1_add_69147_comb[13:1] + {{1{p1_bit_slice_69148_comb[11]}}, p1_bit_slice_69148_comb};
  assign p1_add_69958_comb = p1_add_69149_comb[13:1] + {{1{p1_bit_slice_69150_comb[11]}}, p1_bit_slice_69150_comb};
  assign p1_add_69959_comb = {{1{p1_bit_slice_69151_comb[11]}}, p1_bit_slice_69151_comb} + p1_add_69152_comb[13:1];
  assign p1_add_69960_comb = {{1{p1_bit_slice_69153_comb[11]}}, p1_bit_slice_69153_comb} + p1_add_69154_comb[13:1];
  assign p1_add_69961_comb = p1_add_69155_comb[13:1] + {{1{p1_bit_slice_69156_comb[11]}}, p1_bit_slice_69156_comb};
  assign p1_add_69962_comb = p1_add_69157_comb[13:1] + {{1{p1_bit_slice_69158_comb[11]}}, p1_bit_slice_69158_comb};
  assign p1_add_69963_comb = {{1{p1_bit_slice_69159_comb[11]}}, p1_bit_slice_69159_comb} + p1_add_69160_comb[13:1];
  assign p1_add_69964_comb = {{1{p1_bit_slice_69161_comb[11]}}, p1_bit_slice_69161_comb} + p1_add_69162_comb[13:1];
  assign p1_add_69965_comb = p1_add_69163_comb[13:1] + {{1{p1_bit_slice_69164_comb[11]}}, p1_bit_slice_69164_comb};
  assign p1_add_69966_comb = p1_add_69165_comb[13:1] + {{1{p1_bit_slice_69166_comb[11]}}, p1_bit_slice_69166_comb};
  assign p1_add_69967_comb = {{1{p1_bit_slice_69167_comb[11]}}, p1_bit_slice_69167_comb} + p1_add_69168_comb[13:1];
  assign p1_add_69968_comb = {{1{p1_bit_slice_69169_comb[11]}}, p1_bit_slice_69169_comb} + p1_add_69170_comb[13:1];
  assign p1_add_69969_comb = p1_add_69171_comb[13:1] + {{1{p1_bit_slice_69172_comb[11]}}, p1_bit_slice_69172_comb};
  assign p1_add_69970_comb = p1_add_69173_comb[13:1] + {{1{p1_bit_slice_69174_comb[11]}}, p1_bit_slice_69174_comb};
  assign p1_add_69971_comb = {{2{p1_bit_slice_69175_comb[10]}}, p1_bit_slice_69175_comb} + p1_add_69176_comb[13:1];
  assign p1_add_69972_comb = p1_add_69177_comb[13:1] + p1_add_69178_comb[13:1];
  assign p1_add_69973_comb = p1_add_69179_comb[13:1] + p1_add_69180_comb[13:1];
  assign p1_add_69974_comb = p1_add_69181_comb[13:1] + {{2{p1_bit_slice_69182_comb[10]}}, p1_bit_slice_69182_comb};
  assign p1_add_69975_comb = {{2{p1_bit_slice_69183_comb[10]}}, p1_bit_slice_69183_comb} + p1_add_69184_comb[13:1];
  assign p1_add_69976_comb = p1_add_69185_comb[13:1] + p1_add_69186_comb[13:1];
  assign p1_add_69977_comb = p1_add_69187_comb[13:1] + p1_add_69188_comb[13:1];
  assign p1_add_69978_comb = p1_add_69189_comb[13:1] + {{2{p1_bit_slice_69190_comb[10]}}, p1_bit_slice_69190_comb};
  assign p1_add_69979_comb = {{2{p1_bit_slice_69191_comb[10]}}, p1_bit_slice_69191_comb} + p1_add_69192_comb[13:1];
  assign p1_add_69980_comb = p1_add_69193_comb[13:1] + p1_add_69194_comb[13:1];
  assign p1_add_69981_comb = p1_add_69195_comb[13:1] + p1_add_69196_comb[13:1];
  assign p1_add_69982_comb = p1_add_69197_comb[13:1] + {{2{p1_bit_slice_69198_comb[10]}}, p1_bit_slice_69198_comb};
  assign p1_add_69983_comb = {{2{p1_bit_slice_69199_comb[10]}}, p1_bit_slice_69199_comb} + p1_add_69200_comb[13:1];
  assign p1_add_69984_comb = p1_add_69201_comb[13:1] + p1_add_69202_comb[13:1];
  assign p1_add_69985_comb = p1_add_69203_comb[13:1] + p1_add_69204_comb[13:1];
  assign p1_add_69986_comb = p1_add_69205_comb[13:1] + {{2{p1_bit_slice_69206_comb[10]}}, p1_bit_slice_69206_comb};
  assign p1_add_69991_comb = p1_add_69215_comb[13:1] + p1_add_69216_comb[13:1];
  assign p1_add_69992_comb = p1_add_69217_comb[13:1] + {{2{p1_bit_slice_69218_comb[10]}}, p1_bit_slice_69218_comb};
  assign p1_add_69993_comb = {{2{p1_bit_slice_69219_comb[10]}}, p1_bit_slice_69219_comb} + p1_add_69220_comb[13:1];
  assign p1_add_69994_comb = p1_add_69221_comb[13:1] + p1_add_69222_comb[13:1];
  assign p1_add_69995_comb = p1_add_69223_comb[13:1] + p1_add_69224_comb[13:1];
  assign p1_add_69996_comb = p1_add_69225_comb[13:1] + {{2{p1_bit_slice_69226_comb[10]}}, p1_bit_slice_69226_comb};
  assign p1_add_69997_comb = {{2{p1_bit_slice_69227_comb[10]}}, p1_bit_slice_69227_comb} + p1_add_69228_comb[13:1];
  assign p1_add_69998_comb = p1_add_69229_comb[13:1] + p1_add_69230_comb[13:1];
  assign p1_add_69999_comb = p1_add_69231_comb[13:1] + {{1{p1_bit_slice_69232_comb[11]}}, p1_bit_slice_69232_comb};
  assign p1_add_70000_comb = {{1{p1_bit_slice_69233_comb[11]}}, p1_bit_slice_69233_comb} + p1_add_69234_comb[13:1];
  assign p1_add_70001_comb = p1_add_69235_comb[13:1] + {{1{p1_bit_slice_69236_comb[11]}}, p1_bit_slice_69236_comb};
  assign p1_add_70002_comb = {{1{p1_bit_slice_69237_comb[11]}}, p1_bit_slice_69237_comb} + p1_add_69238_comb[13:1];
  assign p1_add_70003_comb = p1_add_69239_comb[13:1] + {{1{p1_bit_slice_69240_comb[11]}}, p1_bit_slice_69240_comb};
  assign p1_add_70004_comb = {{1{p1_bit_slice_69241_comb[11]}}, p1_bit_slice_69241_comb} + p1_add_69242_comb[13:1];
  assign p1_add_70005_comb = p1_add_69243_comb[13:1] + {{1{p1_bit_slice_69244_comb[11]}}, p1_bit_slice_69244_comb};
  assign p1_add_70006_comb = {{1{p1_bit_slice_69245_comb[11]}}, p1_bit_slice_69245_comb} + p1_add_69246_comb[13:1];
  assign p1_add_70007_comb = p1_add_69247_comb[13:1] + {{2{p1_bit_slice_69248_comb[10]}}, p1_bit_slice_69248_comb};
  assign p1_add_70008_comb = p1_add_69249_comb[13:1] + p1_add_69250_comb[13:1];
  assign p1_add_70009_comb = p1_add_69251_comb[13:1] + p1_add_69252_comb[13:1];
  assign p1_add_70010_comb = {{2{p1_bit_slice_69253_comb[10]}}, p1_bit_slice_69253_comb} + p1_add_69254_comb[13:1];
  assign p1_add_70011_comb = p1_add_69255_comb[13:1] + {{2{p1_bit_slice_69256_comb[10]}}, p1_bit_slice_69256_comb};
  assign p1_add_70012_comb = p1_add_69257_comb[13:1] + p1_add_69258_comb[13:1];
  assign p1_add_70013_comb = p1_add_69259_comb[13:1] + p1_add_69260_comb[13:1];
  assign p1_add_70014_comb = {{2{p1_bit_slice_69261_comb[10]}}, p1_bit_slice_69261_comb} + p1_add_69262_comb[13:1];
  assign p1_add_70015_comb = p1_add_69263_comb[13:1] + p1_add_69264_comb[13:1];
  assign p1_add_70016_comb = p1_add_69265_comb[13:1] + p1_add_69266_comb[13:1];
  assign p1_add_70017_comb = p1_add_69267_comb[13:1] + p1_add_69268_comb[13:1];
  assign p1_add_70018_comb = p1_add_69269_comb[13:1] + p1_add_69270_comb[13:1];
  assign p1_add_70019_comb = p1_add_69271_comb[13:1] + p1_add_69272_comb[13:1];
  assign p1_add_70020_comb = p1_add_69273_comb[13:1] + p1_add_69274_comb[13:1];
  assign p1_add_70021_comb = p1_add_69275_comb[13:1] + p1_add_69276_comb[13:1];
  assign p1_add_70022_comb = p1_add_69277_comb[13:1] + p1_add_69278_comb[13:1];
  assign p1_add_70023_comb = p1_add_69279_comb[13:1] + p1_add_69280_comb[13:1];
  assign p1_add_70024_comb = {{2{p1_bit_slice_69281_comb[10]}}, p1_bit_slice_69281_comb} + p1_add_69282_comb[13:1];
  assign p1_add_70025_comb = p1_add_69283_comb[13:1] + {{2{p1_bit_slice_69284_comb[10]}}, p1_bit_slice_69284_comb};
  assign p1_add_70026_comb = p1_add_69285_comb[13:1] + p1_add_69286_comb[13:1];
  assign p1_add_70027_comb = p1_add_69287_comb[13:1] + p1_add_69288_comb[13:1];
  assign p1_add_70028_comb = {{2{p1_bit_slice_69289_comb[10]}}, p1_bit_slice_69289_comb} + p1_add_69290_comb[13:1];
  assign p1_add_70029_comb = p1_add_69291_comb[13:1] + {{2{p1_bit_slice_69292_comb[10]}}, p1_bit_slice_69292_comb};
  assign p1_add_70030_comb = p1_add_69293_comb[13:1] + p1_add_69294_comb[13:1];
  assign p1_add_70031_comb = {{1{p1_bit_slice_69295_comb[11]}}, p1_bit_slice_69295_comb} + p1_add_69296_comb[13:1];
  assign p1_add_70032_comb = {{1{p1_bit_slice_69297_comb[11]}}, p1_bit_slice_69297_comb} + p1_add_69298_comb[13:1];
  assign p1_add_70033_comb = p1_add_69299_comb[13:1] + {{1{p1_bit_slice_69300_comb[11]}}, p1_bit_slice_69300_comb};
  assign p1_add_70034_comb = p1_add_69301_comb[13:1] + {{1{p1_bit_slice_69302_comb[11]}}, p1_bit_slice_69302_comb};
  assign p1_add_70035_comb = {{1{p1_bit_slice_69303_comb[11]}}, p1_bit_slice_69303_comb} + p1_add_69304_comb[13:1];
  assign p1_add_70036_comb = {{1{p1_bit_slice_69305_comb[11]}}, p1_bit_slice_69305_comb} + p1_add_69306_comb[13:1];
  assign p1_add_70037_comb = p1_add_69307_comb[13:1] + {{1{p1_bit_slice_69308_comb[11]}}, p1_bit_slice_69308_comb};
  assign p1_add_70038_comb = p1_add_69309_comb[13:1] + {{1{p1_bit_slice_69310_comb[11]}}, p1_bit_slice_69310_comb};
  assign p1_add_70039_comb = {{2{p1_bit_slice_69311_comb[10]}}, p1_bit_slice_69311_comb} + p1_add_69312_comb[13:1];
  assign p1_add_70040_comb = p1_add_69313_comb[13:1] + p1_add_69314_comb[13:1];
  assign p1_add_70041_comb = p1_add_69315_comb[13:1] + p1_add_69316_comb[13:1];
  assign p1_add_70042_comb = p1_add_69317_comb[13:1] + {{2{p1_bit_slice_69318_comb[10]}}, p1_bit_slice_69318_comb};
  assign p1_add_70043_comb = {{2{p1_bit_slice_69319_comb[10]}}, p1_bit_slice_69319_comb} + p1_add_69320_comb[13:1];
  assign p1_add_70044_comb = p1_add_69321_comb[13:1] + p1_add_69322_comb[13:1];
  assign p1_add_70045_comb = p1_add_69323_comb[13:1] + p1_add_69324_comb[13:1];
  assign p1_add_70046_comb = p1_add_69325_comb[13:1] + {{2{p1_bit_slice_69326_comb[10]}}, p1_bit_slice_69326_comb};
  assign p1_umul_70287_comb = umul32b_32b_x_7b(p1_sum__967_comb, 7'h5b);
  assign p1_umul_70288_comb = umul32b_32b_x_7b(p1_sum__932_comb, 7'h5b);
  assign p1_umul_70317_comb = umul32b_32b_x_7b(p1_sum__1016_comb, 7'h5b);
  assign p1_umul_70318_comb = umul32b_32b_x_7b(p1_sum__995_comb, 7'h5b);
  assign p1_umul_70319_comb = umul32b_32b_x_7b(p1_sum__890_comb, 7'h5b);
  assign p1_umul_70320_comb = umul32b_32b_x_7b(p1_sum__841_comb, 7'h5b);
  assign p1_umul_70377_comb = umul32b_32b_x_7b(p1_sum__1023_comb, 7'h5b);
  assign p1_umul_70378_comb = umul32b_32b_x_7b(p1_sum__785_comb, 7'h5b);
  assign p1_sum__1768_comb = {{12{p1_add_69811_comb[12]}}, p1_add_69811_comb};
  assign p1_sum__1769_comb = {{12{p1_add_69812_comb[12]}}, p1_add_69812_comb};
  assign p1_sum__1770_comb = {{12{p1_add_69813_comb[12]}}, p1_add_69813_comb};
  assign p1_sum__1771_comb = {{12{p1_add_69814_comb[12]}}, p1_add_69814_comb};
  assign p1_sum__1748_comb = {{12{p1_add_69815_comb[12]}}, p1_add_69815_comb};
  assign p1_sum__1749_comb = {{12{p1_add_69816_comb[12]}}, p1_add_69816_comb};
  assign p1_sum__1750_comb = {{12{p1_add_69817_comb[12]}}, p1_add_69817_comb};
  assign p1_sum__1751_comb = {{12{p1_add_69818_comb[12]}}, p1_add_69818_comb};
  assign p1_sum__1752_comb = {{12{p1_add_69819_comb[12]}}, p1_add_69819_comb};
  assign p1_sum__1753_comb = {{12{p1_add_69820_comb[12]}}, p1_add_69820_comb};
  assign p1_sum__1754_comb = {{12{p1_add_69821_comb[12]}}, p1_add_69821_comb};
  assign p1_sum__1755_comb = {{12{p1_add_69822_comb[12]}}, p1_add_69822_comb};
  assign p1_sum__1728_comb = {{12{p1_add_69823_comb[12]}}, p1_add_69823_comb};
  assign p1_sum__1729_comb = {{12{p1_add_69824_comb[12]}}, p1_add_69824_comb};
  assign p1_sum__1730_comb = {{12{p1_add_69825_comb[12]}}, p1_add_69825_comb};
  assign p1_sum__1731_comb = {{12{p1_add_69826_comb[12]}}, p1_add_69826_comb};
  assign p1_sum__1732_comb = {{12{p1_add_69827_comb[12]}}, p1_add_69827_comb};
  assign p1_sum__1733_comb = {{12{p1_add_69828_comb[12]}}, p1_add_69828_comb};
  assign p1_sum__1734_comb = {{12{p1_add_69829_comb[12]}}, p1_add_69829_comb};
  assign p1_sum__1735_comb = {{12{p1_add_69830_comb[12]}}, p1_add_69830_comb};
  assign p1_sum__1704_comb = {{12{p1_add_69831_comb[12]}}, p1_add_69831_comb};
  assign p1_sum__1705_comb = {{12{p1_add_69832_comb[12]}}, p1_add_69832_comb};
  assign p1_sum__1706_comb = {{12{p1_add_69833_comb[12]}}, p1_add_69833_comb};
  assign p1_sum__1707_comb = {{12{p1_add_69834_comb[12]}}, p1_add_69834_comb};
  assign p1_sum__1708_comb = {{12{p1_add_69835_comb[12]}}, p1_add_69835_comb};
  assign p1_sum__1709_comb = {{12{p1_add_69836_comb[12]}}, p1_add_69836_comb};
  assign p1_sum__1710_comb = {{12{p1_add_69837_comb[12]}}, p1_add_69837_comb};
  assign p1_sum__1711_comb = {{12{p1_add_69838_comb[12]}}, p1_add_69838_comb};
  assign p1_sum__1680_comb = {{12{p1_add_69839_comb[12]}}, p1_add_69839_comb};
  assign p1_sum__1681_comb = {{12{p1_add_69840_comb[12]}}, p1_add_69840_comb};
  assign p1_sum__1682_comb = {{12{p1_add_69841_comb[12]}}, p1_add_69841_comb};
  assign p1_sum__1683_comb = {{12{p1_add_69842_comb[12]}}, p1_add_69842_comb};
  assign p1_sum__1684_comb = {{12{p1_add_69843_comb[12]}}, p1_add_69843_comb};
  assign p1_sum__1685_comb = {{12{p1_add_69844_comb[12]}}, p1_add_69844_comb};
  assign p1_sum__1686_comb = {{12{p1_add_69845_comb[12]}}, p1_add_69845_comb};
  assign p1_sum__1687_comb = {{12{p1_add_69846_comb[12]}}, p1_add_69846_comb};
  assign p1_sum__1656_comb = {{12{p1_add_69847_comb[12]}}, p1_add_69847_comb};
  assign p1_sum__1657_comb = {{12{p1_add_69848_comb[12]}}, p1_add_69848_comb};
  assign p1_sum__1658_comb = {{12{p1_add_69849_comb[12]}}, p1_add_69849_comb};
  assign p1_sum__1659_comb = {{12{p1_add_69850_comb[12]}}, p1_add_69850_comb};
  assign p1_sum__1660_comb = {{12{p1_add_69851_comb[12]}}, p1_add_69851_comb};
  assign p1_sum__1661_comb = {{12{p1_add_69852_comb[12]}}, p1_add_69852_comb};
  assign p1_sum__1662_comb = {{12{p1_add_69853_comb[12]}}, p1_add_69853_comb};
  assign p1_sum__1663_comb = {{12{p1_add_69854_comb[12]}}, p1_add_69854_comb};
  assign p1_sum__1636_comb = {{12{p1_add_69855_comb[12]}}, p1_add_69855_comb};
  assign p1_sum__1637_comb = {{12{p1_add_69856_comb[12]}}, p1_add_69856_comb};
  assign p1_sum__1638_comb = {{12{p1_add_69857_comb[12]}}, p1_add_69857_comb};
  assign p1_sum__1639_comb = {{12{p1_add_69858_comb[12]}}, p1_add_69858_comb};
  assign p1_sum__1640_comb = {{12{p1_add_69859_comb[12]}}, p1_add_69859_comb};
  assign p1_sum__1641_comb = {{12{p1_add_69860_comb[12]}}, p1_add_69860_comb};
  assign p1_sum__1642_comb = {{12{p1_add_69861_comb[12]}}, p1_add_69861_comb};
  assign p1_sum__1643_comb = {{12{p1_add_69862_comb[12]}}, p1_add_69862_comb};
  assign p1_sum__1620_comb = {{12{p1_add_69863_comb[12]}}, p1_add_69863_comb};
  assign p1_sum__1621_comb = {{12{p1_add_69864_comb[12]}}, p1_add_69864_comb};
  assign p1_sum__1622_comb = {{12{p1_add_69865_comb[12]}}, p1_add_69865_comb};
  assign p1_sum__1623_comb = {{12{p1_add_69866_comb[12]}}, p1_add_69866_comb};
  assign p1_sum__1796_comb = {{12{p1_add_69875_comb[12]}}, p1_add_69875_comb};
  assign p1_sum__1797_comb = {{12{p1_add_69876_comb[12]}}, p1_add_69876_comb};
  assign p1_sum__1798_comb = {{12{p1_add_69877_comb[12]}}, p1_add_69877_comb};
  assign p1_sum__1799_comb = {{12{p1_add_69878_comb[12]}}, p1_add_69878_comb};
  assign p1_sum__1784_comb = {{12{p1_add_69879_comb[12]}}, p1_add_69879_comb};
  assign p1_sum__1785_comb = {{12{p1_add_69880_comb[12]}}, p1_add_69880_comb};
  assign p1_sum__1786_comb = {{12{p1_add_69881_comb[12]}}, p1_add_69881_comb};
  assign p1_sum__1787_comb = {{12{p1_add_69882_comb[12]}}, p1_add_69882_comb};
  assign p1_sum__1724_comb = {{12{p1_add_69883_comb[12]}}, p1_add_69883_comb};
  assign p1_sum__1725_comb = {{12{p1_add_69884_comb[12]}}, p1_add_69884_comb};
  assign p1_sum__1726_comb = {{12{p1_add_69885_comb[12]}}, p1_add_69885_comb};
  assign p1_sum__1727_comb = {{12{p1_add_69886_comb[12]}}, p1_add_69886_comb};
  assign p1_sum__1696_comb = {{12{p1_add_69887_comb[12]}}, p1_add_69887_comb};
  assign p1_sum__1697_comb = {{12{p1_add_69888_comb[12]}}, p1_add_69888_comb};
  assign p1_sum__1698_comb = {{12{p1_add_69889_comb[12]}}, p1_add_69889_comb};
  assign p1_sum__1699_comb = {{12{p1_add_69890_comb[12]}}, p1_add_69890_comb};
  assign p1_sum__1788_comb = {{12{p1_add_69891_comb[12]}}, p1_add_69891_comb};
  assign p1_sum__1789_comb = {{12{p1_add_69892_comb[12]}}, p1_add_69892_comb};
  assign p1_sum__1790_comb = {{12{p1_add_69893_comb[12]}}, p1_add_69893_comb};
  assign p1_sum__1791_comb = {{12{p1_add_69894_comb[12]}}, p1_add_69894_comb};
  assign p1_sum__1772_comb = {{12{p1_add_69895_comb[12]}}, p1_add_69895_comb};
  assign p1_sum__1773_comb = {{12{p1_add_69896_comb[12]}}, p1_add_69896_comb};
  assign p1_sum__1774_comb = {{12{p1_add_69897_comb[12]}}, p1_add_69897_comb};
  assign p1_sum__1775_comb = {{12{p1_add_69898_comb[12]}}, p1_add_69898_comb};
  assign p1_sum__1700_comb = {{12{p1_add_69899_comb[12]}}, p1_add_69899_comb};
  assign p1_sum__1701_comb = {{12{p1_add_69900_comb[12]}}, p1_add_69900_comb};
  assign p1_sum__1702_comb = {{12{p1_add_69901_comb[12]}}, p1_add_69901_comb};
  assign p1_sum__1703_comb = {{12{p1_add_69902_comb[12]}}, p1_add_69902_comb};
  assign p1_sum__1672_comb = {{12{p1_add_69903_comb[12]}}, p1_add_69903_comb};
  assign p1_sum__1673_comb = {{12{p1_add_69904_comb[12]}}, p1_add_69904_comb};
  assign p1_sum__1674_comb = {{12{p1_add_69905_comb[12]}}, p1_add_69905_comb};
  assign p1_sum__1675_comb = {{12{p1_add_69906_comb[12]}}, p1_add_69906_comb};
  assign p1_sum__1776_comb = {{12{p1_add_69907_comb[12]}}, p1_add_69907_comb};
  assign p1_sum__1777_comb = {{12{p1_add_69908_comb[12]}}, p1_add_69908_comb};
  assign p1_sum__1778_comb = {{12{p1_add_69909_comb[12]}}, p1_add_69909_comb};
  assign p1_sum__1779_comb = {{12{p1_add_69910_comb[12]}}, p1_add_69910_comb};
  assign p1_sum__1756_comb = {{12{p1_add_69911_comb[12]}}, p1_add_69911_comb};
  assign p1_sum__1757_comb = {{12{p1_add_69912_comb[12]}}, p1_add_69912_comb};
  assign p1_sum__1758_comb = {{12{p1_add_69913_comb[12]}}, p1_add_69913_comb};
  assign p1_sum__1759_comb = {{12{p1_add_69914_comb[12]}}, p1_add_69914_comb};
  assign p1_sum__1676_comb = {{12{p1_add_69915_comb[12]}}, p1_add_69915_comb};
  assign p1_sum__1677_comb = {{12{p1_add_69916_comb[12]}}, p1_add_69916_comb};
  assign p1_sum__1678_comb = {{12{p1_add_69917_comb[12]}}, p1_add_69917_comb};
  assign p1_sum__1679_comb = {{12{p1_add_69918_comb[12]}}, p1_add_69918_comb};
  assign p1_sum__1648_comb = {{12{p1_add_69919_comb[12]}}, p1_add_69919_comb};
  assign p1_sum__1649_comb = {{12{p1_add_69920_comb[12]}}, p1_add_69920_comb};
  assign p1_sum__1650_comb = {{12{p1_add_69921_comb[12]}}, p1_add_69921_comb};
  assign p1_sum__1651_comb = {{12{p1_add_69922_comb[12]}}, p1_add_69922_comb};
  assign p1_sum__1760_comb = {{12{p1_add_69923_comb[12]}}, p1_add_69923_comb};
  assign p1_sum__1761_comb = {{12{p1_add_69924_comb[12]}}, p1_add_69924_comb};
  assign p1_sum__1762_comb = {{12{p1_add_69925_comb[12]}}, p1_add_69925_comb};
  assign p1_sum__1763_comb = {{12{p1_add_69926_comb[12]}}, p1_add_69926_comb};
  assign p1_sum__1736_comb = {{12{p1_add_69927_comb[12]}}, p1_add_69927_comb};
  assign p1_sum__1737_comb = {{12{p1_add_69928_comb[12]}}, p1_add_69928_comb};
  assign p1_sum__1738_comb = {{12{p1_add_69929_comb[12]}}, p1_add_69929_comb};
  assign p1_sum__1739_comb = {{12{p1_add_69930_comb[12]}}, p1_add_69930_comb};
  assign p1_sum__1652_comb = {{12{p1_add_69931_comb[12]}}, p1_add_69931_comb};
  assign p1_sum__1653_comb = {{12{p1_add_69932_comb[12]}}, p1_add_69932_comb};
  assign p1_sum__1654_comb = {{12{p1_add_69933_comb[12]}}, p1_add_69933_comb};
  assign p1_sum__1655_comb = {{12{p1_add_69934_comb[12]}}, p1_add_69934_comb};
  assign p1_sum__1628_comb = {{12{p1_add_69935_comb[12]}}, p1_add_69935_comb};
  assign p1_sum__1629_comb = {{12{p1_add_69936_comb[12]}}, p1_add_69936_comb};
  assign p1_sum__1630_comb = {{12{p1_add_69937_comb[12]}}, p1_add_69937_comb};
  assign p1_sum__1631_comb = {{12{p1_add_69938_comb[12]}}, p1_add_69938_comb};
  assign p1_sum__1740_comb = {{12{p1_add_69939_comb[12]}}, p1_add_69939_comb};
  assign p1_sum__1741_comb = {{12{p1_add_69940_comb[12]}}, p1_add_69940_comb};
  assign p1_sum__1742_comb = {{12{p1_add_69941_comb[12]}}, p1_add_69941_comb};
  assign p1_sum__1743_comb = {{12{p1_add_69942_comb[12]}}, p1_add_69942_comb};
  assign p1_sum__1712_comb = {{12{p1_add_69943_comb[12]}}, p1_add_69943_comb};
  assign p1_sum__1713_comb = {{12{p1_add_69944_comb[12]}}, p1_add_69944_comb};
  assign p1_sum__1714_comb = {{12{p1_add_69945_comb[12]}}, p1_add_69945_comb};
  assign p1_sum__1715_comb = {{12{p1_add_69946_comb[12]}}, p1_add_69946_comb};
  assign p1_sum__1632_comb = {{12{p1_add_69947_comb[12]}}, p1_add_69947_comb};
  assign p1_sum__1633_comb = {{12{p1_add_69948_comb[12]}}, p1_add_69948_comb};
  assign p1_sum__1634_comb = {{12{p1_add_69949_comb[12]}}, p1_add_69949_comb};
  assign p1_sum__1635_comb = {{12{p1_add_69950_comb[12]}}, p1_add_69950_comb};
  assign p1_sum__1612_comb = {{12{p1_add_69951_comb[12]}}, p1_add_69951_comb};
  assign p1_sum__1613_comb = {{12{p1_add_69952_comb[12]}}, p1_add_69952_comb};
  assign p1_sum__1614_comb = {{12{p1_add_69953_comb[12]}}, p1_add_69953_comb};
  assign p1_sum__1615_comb = {{12{p1_add_69954_comb[12]}}, p1_add_69954_comb};
  assign p1_sum__1716_comb = {{12{p1_add_69955_comb[12]}}, p1_add_69955_comb};
  assign p1_sum__1717_comb = {{12{p1_add_69956_comb[12]}}, p1_add_69956_comb};
  assign p1_sum__1718_comb = {{12{p1_add_69957_comb[12]}}, p1_add_69957_comb};
  assign p1_sum__1719_comb = {{12{p1_add_69958_comb[12]}}, p1_add_69958_comb};
  assign p1_sum__1688_comb = {{12{p1_add_69959_comb[12]}}, p1_add_69959_comb};
  assign p1_sum__1689_comb = {{12{p1_add_69960_comb[12]}}, p1_add_69960_comb};
  assign p1_sum__1690_comb = {{12{p1_add_69961_comb[12]}}, p1_add_69961_comb};
  assign p1_sum__1691_comb = {{12{p1_add_69962_comb[12]}}, p1_add_69962_comb};
  assign p1_sum__1616_comb = {{12{p1_add_69963_comb[12]}}, p1_add_69963_comb};
  assign p1_sum__1617_comb = {{12{p1_add_69964_comb[12]}}, p1_add_69964_comb};
  assign p1_sum__1618_comb = {{12{p1_add_69965_comb[12]}}, p1_add_69965_comb};
  assign p1_sum__1619_comb = {{12{p1_add_69966_comb[12]}}, p1_add_69966_comb};
  assign p1_sum__1600_comb = {{12{p1_add_69967_comb[12]}}, p1_add_69967_comb};
  assign p1_sum__1601_comb = {{12{p1_add_69968_comb[12]}}, p1_add_69968_comb};
  assign p1_sum__1602_comb = {{12{p1_add_69969_comb[12]}}, p1_add_69969_comb};
  assign p1_sum__1603_comb = {{12{p1_add_69970_comb[12]}}, p1_add_69970_comb};
  assign p1_sum__1692_comb = {{12{p1_add_69971_comb[12]}}, p1_add_69971_comb};
  assign p1_sum__1693_comb = {{12{p1_add_69972_comb[12]}}, p1_add_69972_comb};
  assign p1_sum__1694_comb = {{12{p1_add_69973_comb[12]}}, p1_add_69973_comb};
  assign p1_sum__1695_comb = {{12{p1_add_69974_comb[12]}}, p1_add_69974_comb};
  assign p1_sum__1664_comb = {{12{p1_add_69975_comb[12]}}, p1_add_69975_comb};
  assign p1_sum__1665_comb = {{12{p1_add_69976_comb[12]}}, p1_add_69976_comb};
  assign p1_sum__1666_comb = {{12{p1_add_69977_comb[12]}}, p1_add_69977_comb};
  assign p1_sum__1667_comb = {{12{p1_add_69978_comb[12]}}, p1_add_69978_comb};
  assign p1_sum__1604_comb = {{12{p1_add_69979_comb[12]}}, p1_add_69979_comb};
  assign p1_sum__1605_comb = {{12{p1_add_69980_comb[12]}}, p1_add_69980_comb};
  assign p1_sum__1606_comb = {{12{p1_add_69981_comb[12]}}, p1_add_69981_comb};
  assign p1_sum__1607_comb = {{12{p1_add_69982_comb[12]}}, p1_add_69982_comb};
  assign p1_sum__1592_comb = {{12{p1_add_69983_comb[12]}}, p1_add_69983_comb};
  assign p1_sum__1593_comb = {{12{p1_add_69984_comb[12]}}, p1_add_69984_comb};
  assign p1_sum__1594_comb = {{12{p1_add_69985_comb[12]}}, p1_add_69985_comb};
  assign p1_sum__1595_comb = {{12{p1_add_69986_comb[12]}}, p1_add_69986_comb};
  assign p1_sum__1804_comb = {{12{p1_add_69991_comb[12]}}, p1_add_69991_comb};
  assign p1_sum__1805_comb = {{12{p1_add_69992_comb[12]}}, p1_add_69992_comb};
  assign p1_sum__1806_comb = {{12{p1_add_69993_comb[12]}}, p1_add_69993_comb};
  assign p1_sum__1807_comb = {{12{p1_add_69994_comb[12]}}, p1_add_69994_comb};
  assign p1_sum__1668_comb = {{12{p1_add_69995_comb[12]}}, p1_add_69995_comb};
  assign p1_sum__1669_comb = {{12{p1_add_69996_comb[12]}}, p1_add_69996_comb};
  assign p1_sum__1670_comb = {{12{p1_add_69997_comb[12]}}, p1_add_69997_comb};
  assign p1_sum__1671_comb = {{12{p1_add_69998_comb[12]}}, p1_add_69998_comb};
  assign p1_sum__1800_comb = {{12{p1_add_69999_comb[12]}}, p1_add_69999_comb};
  assign p1_sum__1801_comb = {{12{p1_add_70000_comb[12]}}, p1_add_70000_comb};
  assign p1_sum__1802_comb = {{12{p1_add_70001_comb[12]}}, p1_add_70001_comb};
  assign p1_sum__1803_comb = {{12{p1_add_70002_comb[12]}}, p1_add_70002_comb};
  assign p1_sum__1644_comb = {{12{p1_add_70003_comb[12]}}, p1_add_70003_comb};
  assign p1_sum__1645_comb = {{12{p1_add_70004_comb[12]}}, p1_add_70004_comb};
  assign p1_sum__1646_comb = {{12{p1_add_70005_comb[12]}}, p1_add_70005_comb};
  assign p1_sum__1647_comb = {{12{p1_add_70006_comb[12]}}, p1_add_70006_comb};
  assign p1_sum__1792_comb = {{12{p1_add_70007_comb[12]}}, p1_add_70007_comb};
  assign p1_sum__1793_comb = {{12{p1_add_70008_comb[12]}}, p1_add_70008_comb};
  assign p1_sum__1794_comb = {{12{p1_add_70009_comb[12]}}, p1_add_70009_comb};
  assign p1_sum__1795_comb = {{12{p1_add_70010_comb[12]}}, p1_add_70010_comb};
  assign p1_sum__1624_comb = {{12{p1_add_70011_comb[12]}}, p1_add_70011_comb};
  assign p1_sum__1625_comb = {{12{p1_add_70012_comb[12]}}, p1_add_70012_comb};
  assign p1_sum__1626_comb = {{12{p1_add_70013_comb[12]}}, p1_add_70013_comb};
  assign p1_sum__1627_comb = {{12{p1_add_70014_comb[12]}}, p1_add_70014_comb};
  assign p1_sum__1780_comb = {{12{p1_add_70015_comb[12]}}, p1_add_70015_comb};
  assign p1_sum__1781_comb = {{12{p1_add_70016_comb[12]}}, p1_add_70016_comb};
  assign p1_sum__1782_comb = {{12{p1_add_70017_comb[12]}}, p1_add_70017_comb};
  assign p1_sum__1783_comb = {{12{p1_add_70018_comb[12]}}, p1_add_70018_comb};
  assign p1_sum__1608_comb = {{12{p1_add_70019_comb[12]}}, p1_add_70019_comb};
  assign p1_sum__1609_comb = {{12{p1_add_70020_comb[12]}}, p1_add_70020_comb};
  assign p1_sum__1610_comb = {{12{p1_add_70021_comb[12]}}, p1_add_70021_comb};
  assign p1_sum__1611_comb = {{12{p1_add_70022_comb[12]}}, p1_add_70022_comb};
  assign p1_sum__1764_comb = {{12{p1_add_70023_comb[12]}}, p1_add_70023_comb};
  assign p1_sum__1765_comb = {{12{p1_add_70024_comb[12]}}, p1_add_70024_comb};
  assign p1_sum__1766_comb = {{12{p1_add_70025_comb[12]}}, p1_add_70025_comb};
  assign p1_sum__1767_comb = {{12{p1_add_70026_comb[12]}}, p1_add_70026_comb};
  assign p1_sum__1596_comb = {{12{p1_add_70027_comb[12]}}, p1_add_70027_comb};
  assign p1_sum__1597_comb = {{12{p1_add_70028_comb[12]}}, p1_add_70028_comb};
  assign p1_sum__1598_comb = {{12{p1_add_70029_comb[12]}}, p1_add_70029_comb};
  assign p1_sum__1599_comb = {{12{p1_add_70030_comb[12]}}, p1_add_70030_comb};
  assign p1_sum__1744_comb = {{12{p1_add_70031_comb[12]}}, p1_add_70031_comb};
  assign p1_sum__1745_comb = {{12{p1_add_70032_comb[12]}}, p1_add_70032_comb};
  assign p1_sum__1746_comb = {{12{p1_add_70033_comb[12]}}, p1_add_70033_comb};
  assign p1_sum__1747_comb = {{12{p1_add_70034_comb[12]}}, p1_add_70034_comb};
  assign p1_sum__1588_comb = {{12{p1_add_70035_comb[12]}}, p1_add_70035_comb};
  assign p1_sum__1589_comb = {{12{p1_add_70036_comb[12]}}, p1_add_70036_comb};
  assign p1_sum__1590_comb = {{12{p1_add_70037_comb[12]}}, p1_add_70037_comb};
  assign p1_sum__1591_comb = {{12{p1_add_70038_comb[12]}}, p1_add_70038_comb};
  assign p1_sum__1720_comb = {{12{p1_add_70039_comb[12]}}, p1_add_70039_comb};
  assign p1_sum__1721_comb = {{12{p1_add_70040_comb[12]}}, p1_add_70040_comb};
  assign p1_sum__1722_comb = {{12{p1_add_70041_comb[12]}}, p1_add_70041_comb};
  assign p1_sum__1723_comb = {{12{p1_add_70042_comb[12]}}, p1_add_70042_comb};
  assign p1_sum__1584_comb = {{12{p1_add_70043_comb[12]}}, p1_add_70043_comb};
  assign p1_sum__1585_comb = {{12{p1_add_70044_comb[12]}}, p1_add_70044_comb};
  assign p1_sum__1586_comb = {{12{p1_add_70045_comb[12]}}, p1_add_70045_comb};
  assign p1_sum__1587_comb = {{12{p1_add_70046_comb[12]}}, p1_add_70046_comb};
  assign p1_sum__1340_comb = p1_sum__1768_comb + p1_sum__1769_comb;
  assign p1_sum__1341_comb = p1_sum__1770_comb + p1_sum__1771_comb;
  assign p1_sum__1330_comb = p1_sum__1748_comb + p1_sum__1749_comb;
  assign p1_sum__1331_comb = p1_sum__1750_comb + p1_sum__1751_comb;
  assign p1_sum__1332_comb = p1_sum__1752_comb + p1_sum__1753_comb;
  assign p1_sum__1333_comb = p1_sum__1754_comb + p1_sum__1755_comb;
  assign p1_sum__1320_comb = p1_sum__1728_comb + p1_sum__1729_comb;
  assign p1_sum__1321_comb = p1_sum__1730_comb + p1_sum__1731_comb;
  assign p1_sum__1322_comb = p1_sum__1732_comb + p1_sum__1733_comb;
  assign p1_sum__1323_comb = p1_sum__1734_comb + p1_sum__1735_comb;
  assign p1_sum__1308_comb = p1_sum__1704_comb + p1_sum__1705_comb;
  assign p1_sum__1309_comb = p1_sum__1706_comb + p1_sum__1707_comb;
  assign p1_sum__1310_comb = p1_sum__1708_comb + p1_sum__1709_comb;
  assign p1_sum__1311_comb = p1_sum__1710_comb + p1_sum__1711_comb;
  assign p1_sum__1296_comb = p1_sum__1680_comb + p1_sum__1681_comb;
  assign p1_sum__1297_comb = p1_sum__1682_comb + p1_sum__1683_comb;
  assign p1_sum__1298_comb = p1_sum__1684_comb + p1_sum__1685_comb;
  assign p1_sum__1299_comb = p1_sum__1686_comb + p1_sum__1687_comb;
  assign p1_sum__1284_comb = p1_sum__1656_comb + p1_sum__1657_comb;
  assign p1_sum__1285_comb = p1_sum__1658_comb + p1_sum__1659_comb;
  assign p1_sum__1286_comb = p1_sum__1660_comb + p1_sum__1661_comb;
  assign p1_sum__1287_comb = p1_sum__1662_comb + p1_sum__1663_comb;
  assign p1_sum__1274_comb = p1_sum__1636_comb + p1_sum__1637_comb;
  assign p1_sum__1275_comb = p1_sum__1638_comb + p1_sum__1639_comb;
  assign p1_sum__1276_comb = p1_sum__1640_comb + p1_sum__1641_comb;
  assign p1_sum__1277_comb = p1_sum__1642_comb + p1_sum__1643_comb;
  assign p1_sum__1266_comb = p1_sum__1620_comb + p1_sum__1621_comb;
  assign p1_sum__1267_comb = p1_sum__1622_comb + p1_sum__1623_comb;
  assign p1_sum__1354_comb = p1_sum__1796_comb + p1_sum__1797_comb;
  assign p1_sum__1355_comb = p1_sum__1798_comb + p1_sum__1799_comb;
  assign p1_sum__1348_comb = p1_sum__1784_comb + p1_sum__1785_comb;
  assign p1_sum__1349_comb = p1_sum__1786_comb + p1_sum__1787_comb;
  assign p1_sum__1318_comb = p1_sum__1724_comb + p1_sum__1725_comb;
  assign p1_sum__1319_comb = p1_sum__1726_comb + p1_sum__1727_comb;
  assign p1_sum__1304_comb = p1_sum__1696_comb + p1_sum__1697_comb;
  assign p1_sum__1305_comb = p1_sum__1698_comb + p1_sum__1699_comb;
  assign p1_sum__1350_comb = p1_sum__1788_comb + p1_sum__1789_comb;
  assign p1_sum__1351_comb = p1_sum__1790_comb + p1_sum__1791_comb;
  assign p1_sum__1342_comb = p1_sum__1772_comb + p1_sum__1773_comb;
  assign p1_sum__1343_comb = p1_sum__1774_comb + p1_sum__1775_comb;
  assign p1_sum__1306_comb = p1_sum__1700_comb + p1_sum__1701_comb;
  assign p1_sum__1307_comb = p1_sum__1702_comb + p1_sum__1703_comb;
  assign p1_sum__1292_comb = p1_sum__1672_comb + p1_sum__1673_comb;
  assign p1_sum__1293_comb = p1_sum__1674_comb + p1_sum__1675_comb;
  assign p1_sum__1344_comb = p1_sum__1776_comb + p1_sum__1777_comb;
  assign p1_sum__1345_comb = p1_sum__1778_comb + p1_sum__1779_comb;
  assign p1_sum__1334_comb = p1_sum__1756_comb + p1_sum__1757_comb;
  assign p1_sum__1335_comb = p1_sum__1758_comb + p1_sum__1759_comb;
  assign p1_sum__1294_comb = p1_sum__1676_comb + p1_sum__1677_comb;
  assign p1_sum__1295_comb = p1_sum__1678_comb + p1_sum__1679_comb;
  assign p1_sum__1280_comb = p1_sum__1648_comb + p1_sum__1649_comb;
  assign p1_sum__1281_comb = p1_sum__1650_comb + p1_sum__1651_comb;
  assign p1_sum__1336_comb = p1_sum__1760_comb + p1_sum__1761_comb;
  assign p1_sum__1337_comb = p1_sum__1762_comb + p1_sum__1763_comb;
  assign p1_sum__1324_comb = p1_sum__1736_comb + p1_sum__1737_comb;
  assign p1_sum__1325_comb = p1_sum__1738_comb + p1_sum__1739_comb;
  assign p1_sum__1282_comb = p1_sum__1652_comb + p1_sum__1653_comb;
  assign p1_sum__1283_comb = p1_sum__1654_comb + p1_sum__1655_comb;
  assign p1_sum__1270_comb = p1_sum__1628_comb + p1_sum__1629_comb;
  assign p1_sum__1271_comb = p1_sum__1630_comb + p1_sum__1631_comb;
  assign p1_sum__1326_comb = p1_sum__1740_comb + p1_sum__1741_comb;
  assign p1_sum__1327_comb = p1_sum__1742_comb + p1_sum__1743_comb;
  assign p1_sum__1312_comb = p1_sum__1712_comb + p1_sum__1713_comb;
  assign p1_sum__1313_comb = p1_sum__1714_comb + p1_sum__1715_comb;
  assign p1_sum__1272_comb = p1_sum__1632_comb + p1_sum__1633_comb;
  assign p1_sum__1273_comb = p1_sum__1634_comb + p1_sum__1635_comb;
  assign p1_sum__1262_comb = p1_sum__1612_comb + p1_sum__1613_comb;
  assign p1_sum__1263_comb = p1_sum__1614_comb + p1_sum__1615_comb;
  assign p1_sum__1314_comb = p1_sum__1716_comb + p1_sum__1717_comb;
  assign p1_sum__1315_comb = p1_sum__1718_comb + p1_sum__1719_comb;
  assign p1_sum__1300_comb = p1_sum__1688_comb + p1_sum__1689_comb;
  assign p1_sum__1301_comb = p1_sum__1690_comb + p1_sum__1691_comb;
  assign p1_sum__1264_comb = p1_sum__1616_comb + p1_sum__1617_comb;
  assign p1_sum__1265_comb = p1_sum__1618_comb + p1_sum__1619_comb;
  assign p1_sum__1256_comb = p1_sum__1600_comb + p1_sum__1601_comb;
  assign p1_sum__1257_comb = p1_sum__1602_comb + p1_sum__1603_comb;
  assign p1_sum__1302_comb = p1_sum__1692_comb + p1_sum__1693_comb;
  assign p1_sum__1303_comb = p1_sum__1694_comb + p1_sum__1695_comb;
  assign p1_sum__1288_comb = p1_sum__1664_comb + p1_sum__1665_comb;
  assign p1_sum__1289_comb = p1_sum__1666_comb + p1_sum__1667_comb;
  assign p1_sum__1258_comb = p1_sum__1604_comb + p1_sum__1605_comb;
  assign p1_sum__1259_comb = p1_sum__1606_comb + p1_sum__1607_comb;
  assign p1_sum__1252_comb = p1_sum__1592_comb + p1_sum__1593_comb;
  assign p1_sum__1253_comb = p1_sum__1594_comb + p1_sum__1595_comb;
  assign p1_sum__1358_comb = p1_sum__1804_comb + p1_sum__1805_comb;
  assign p1_sum__1359_comb = p1_sum__1806_comb + p1_sum__1807_comb;
  assign p1_sum__1290_comb = p1_sum__1668_comb + p1_sum__1669_comb;
  assign p1_sum__1291_comb = p1_sum__1670_comb + p1_sum__1671_comb;
  assign p1_sum__1356_comb = p1_sum__1800_comb + p1_sum__1801_comb;
  assign p1_sum__1357_comb = p1_sum__1802_comb + p1_sum__1803_comb;
  assign p1_sum__1278_comb = p1_sum__1644_comb + p1_sum__1645_comb;
  assign p1_sum__1279_comb = p1_sum__1646_comb + p1_sum__1647_comb;
  assign p1_sum__1352_comb = p1_sum__1792_comb + p1_sum__1793_comb;
  assign p1_sum__1353_comb = p1_sum__1794_comb + p1_sum__1795_comb;
  assign p1_sum__1268_comb = p1_sum__1624_comb + p1_sum__1625_comb;
  assign p1_sum__1269_comb = p1_sum__1626_comb + p1_sum__1627_comb;
  assign p1_sum__1346_comb = p1_sum__1780_comb + p1_sum__1781_comb;
  assign p1_sum__1347_comb = p1_sum__1782_comb + p1_sum__1783_comb;
  assign p1_sum__1260_comb = p1_sum__1608_comb + p1_sum__1609_comb;
  assign p1_sum__1261_comb = p1_sum__1610_comb + p1_sum__1611_comb;
  assign p1_sum__1338_comb = p1_sum__1764_comb + p1_sum__1765_comb;
  assign p1_sum__1339_comb = p1_sum__1766_comb + p1_sum__1767_comb;
  assign p1_sum__1254_comb = p1_sum__1596_comb + p1_sum__1597_comb;
  assign p1_sum__1255_comb = p1_sum__1598_comb + p1_sum__1599_comb;
  assign p1_sum__1328_comb = p1_sum__1744_comb + p1_sum__1745_comb;
  assign p1_sum__1329_comb = p1_sum__1746_comb + p1_sum__1747_comb;
  assign p1_sum__1250_comb = p1_sum__1588_comb + p1_sum__1589_comb;
  assign p1_sum__1251_comb = p1_sum__1590_comb + p1_sum__1591_comb;
  assign p1_sum__1316_comb = p1_sum__1720_comb + p1_sum__1721_comb;
  assign p1_sum__1317_comb = p1_sum__1722_comb + p1_sum__1723_comb;
  assign p1_sum__1248_comb = p1_sum__1584_comb + p1_sum__1585_comb;
  assign p1_sum__1249_comb = p1_sum__1586_comb + p1_sum__1587_comb;
  assign p1_add_70535_comb = p1_umul_70287_comb[31:7] + 25'h000_0001;
  assign p1_add_70536_comb = p1_umul_70288_comb[31:7] + 25'h000_0001;
  assign p1_add_70551_comb = p1_umul_70317_comb[31:7] + 25'h000_0001;
  assign p1_add_70552_comb = p1_umul_70318_comb[31:7] + 25'h000_0001;
  assign p1_add_70553_comb = p1_umul_70319_comb[31:7] + 25'h000_0001;
  assign p1_add_70554_comb = p1_umul_70320_comb[31:7] + 25'h000_0001;
  assign p1_add_70583_comb = p1_umul_70377_comb[31:7] + 25'h000_0001;
  assign p1_add_70584_comb = p1_umul_70378_comb[31:7] + 25'h000_0001;
  assign p1_sum__1126_comb = p1_sum__1340_comb + p1_sum__1341_comb;
  assign p1_sum__1121_comb = p1_sum__1330_comb + p1_sum__1331_comb;
  assign p1_sum__1122_comb = p1_sum__1332_comb + p1_sum__1333_comb;
  assign p1_sum__1116_comb = p1_sum__1320_comb + p1_sum__1321_comb;
  assign p1_sum__1117_comb = p1_sum__1322_comb + p1_sum__1323_comb;
  assign p1_sum__1110_comb = p1_sum__1308_comb + p1_sum__1309_comb;
  assign p1_sum__1111_comb = p1_sum__1310_comb + p1_sum__1311_comb;
  assign p1_sum__1104_comb = p1_sum__1296_comb + p1_sum__1297_comb;
  assign p1_sum__1105_comb = p1_sum__1298_comb + p1_sum__1299_comb;
  assign p1_sum__1098_comb = p1_sum__1284_comb + p1_sum__1285_comb;
  assign p1_sum__1099_comb = p1_sum__1286_comb + p1_sum__1287_comb;
  assign p1_sum__1093_comb = p1_sum__1274_comb + p1_sum__1275_comb;
  assign p1_sum__1094_comb = p1_sum__1276_comb + p1_sum__1277_comb;
  assign p1_sum__1089_comb = p1_sum__1266_comb + p1_sum__1267_comb;
  assign p1_sum__1133_comb = p1_sum__1354_comb + p1_sum__1355_comb;
  assign p1_sum__1130_comb = p1_sum__1348_comb + p1_sum__1349_comb;
  assign p1_sum__1115_comb = p1_sum__1318_comb + p1_sum__1319_comb;
  assign p1_sum__1108_comb = p1_sum__1304_comb + p1_sum__1305_comb;
  assign p1_sum__1131_comb = p1_sum__1350_comb + p1_sum__1351_comb;
  assign p1_sum__1127_comb = p1_sum__1342_comb + p1_sum__1343_comb;
  assign p1_sum__1109_comb = p1_sum__1306_comb + p1_sum__1307_comb;
  assign p1_sum__1102_comb = p1_sum__1292_comb + p1_sum__1293_comb;
  assign p1_sum__1128_comb = p1_sum__1344_comb + p1_sum__1345_comb;
  assign p1_sum__1123_comb = p1_sum__1334_comb + p1_sum__1335_comb;
  assign p1_sum__1103_comb = p1_sum__1294_comb + p1_sum__1295_comb;
  assign p1_sum__1096_comb = p1_sum__1280_comb + p1_sum__1281_comb;
  assign p1_sum__1124_comb = p1_sum__1336_comb + p1_sum__1337_comb;
  assign p1_sum__1118_comb = p1_sum__1324_comb + p1_sum__1325_comb;
  assign p1_sum__1097_comb = p1_sum__1282_comb + p1_sum__1283_comb;
  assign p1_sum__1091_comb = p1_sum__1270_comb + p1_sum__1271_comb;
  assign p1_sum__1119_comb = p1_sum__1326_comb + p1_sum__1327_comb;
  assign p1_sum__1112_comb = p1_sum__1312_comb + p1_sum__1313_comb;
  assign p1_sum__1092_comb = p1_sum__1272_comb + p1_sum__1273_comb;
  assign p1_sum__1087_comb = p1_sum__1262_comb + p1_sum__1263_comb;
  assign p1_sum__1113_comb = p1_sum__1314_comb + p1_sum__1315_comb;
  assign p1_sum__1106_comb = p1_sum__1300_comb + p1_sum__1301_comb;
  assign p1_sum__1088_comb = p1_sum__1264_comb + p1_sum__1265_comb;
  assign p1_sum__1084_comb = p1_sum__1256_comb + p1_sum__1257_comb;
  assign p1_sum__1107_comb = p1_sum__1302_comb + p1_sum__1303_comb;
  assign p1_sum__1100_comb = p1_sum__1288_comb + p1_sum__1289_comb;
  assign p1_sum__1085_comb = p1_sum__1258_comb + p1_sum__1259_comb;
  assign p1_sum__1082_comb = p1_sum__1252_comb + p1_sum__1253_comb;
  assign p1_sum__1135_comb = p1_sum__1358_comb + p1_sum__1359_comb;
  assign p1_sum__1101_comb = p1_sum__1290_comb + p1_sum__1291_comb;
  assign p1_sum__1134_comb = p1_sum__1356_comb + p1_sum__1357_comb;
  assign p1_sum__1095_comb = p1_sum__1278_comb + p1_sum__1279_comb;
  assign p1_sum__1132_comb = p1_sum__1352_comb + p1_sum__1353_comb;
  assign p1_sum__1090_comb = p1_sum__1268_comb + p1_sum__1269_comb;
  assign p1_sum__1129_comb = p1_sum__1346_comb + p1_sum__1347_comb;
  assign p1_sum__1086_comb = p1_sum__1260_comb + p1_sum__1261_comb;
  assign p1_sum__1125_comb = p1_sum__1338_comb + p1_sum__1339_comb;
  assign p1_sum__1083_comb = p1_sum__1254_comb + p1_sum__1255_comb;
  assign p1_sum__1120_comb = p1_sum__1328_comb + p1_sum__1329_comb;
  assign p1_sum__1081_comb = p1_sum__1250_comb + p1_sum__1251_comb;
  assign p1_sum__1114_comb = p1_sum__1316_comb + p1_sum__1317_comb;
  assign p1_sum__1080_comb = p1_sum__1248_comb + p1_sum__1249_comb;
  assign p1_add_70537_comb = p1_sum__1126_comb + 25'h000_0001;
  assign p1_add_70538_comb = p1_sum__1121_comb + 25'h000_0001;
  assign p1_add_70539_comb = p1_sum__1122_comb + 25'h000_0001;
  assign p1_add_70540_comb = p1_sum__1116_comb + 25'h000_0001;
  assign p1_add_70541_comb = p1_sum__1117_comb + 25'h000_0001;
  assign p1_add_70542_comb = p1_sum__1110_comb + 25'h000_0001;
  assign p1_add_70543_comb = p1_sum__1111_comb + 25'h000_0001;
  assign p1_add_70544_comb = p1_sum__1104_comb + 25'h000_0001;
  assign p1_add_70545_comb = p1_sum__1105_comb + 25'h000_0001;
  assign p1_add_70546_comb = p1_sum__1098_comb + 25'h000_0001;
  assign p1_add_70547_comb = p1_sum__1099_comb + 25'h000_0001;
  assign p1_add_70548_comb = p1_sum__1093_comb + 25'h000_0001;
  assign p1_add_70549_comb = p1_sum__1094_comb + 25'h000_0001;
  assign p1_add_70550_comb = p1_sum__1089_comb + 25'h000_0001;
  assign p1_add_70555_comb = p1_sum__1133_comb + 25'h000_0001;
  assign p1_add_70556_comb = p1_sum__1130_comb + 25'h000_0001;
  assign p1_add_70557_comb = p1_sum__1115_comb + 25'h000_0001;
  assign p1_add_70558_comb = p1_sum__1108_comb + 25'h000_0001;
  assign p1_add_70559_comb = p1_sum__1131_comb + 25'h000_0001;
  assign p1_add_70560_comb = p1_sum__1127_comb + 25'h000_0001;
  assign p1_add_70561_comb = p1_sum__1109_comb + 25'h000_0001;
  assign p1_add_70562_comb = p1_sum__1102_comb + 25'h000_0001;
  assign p1_add_70563_comb = p1_sum__1128_comb + 25'h000_0001;
  assign p1_add_70564_comb = p1_sum__1123_comb + 25'h000_0001;
  assign p1_add_70565_comb = p1_sum__1103_comb + 25'h000_0001;
  assign p1_add_70566_comb = p1_sum__1096_comb + 25'h000_0001;
  assign p1_add_70567_comb = p1_sum__1124_comb + 25'h000_0001;
  assign p1_add_70568_comb = p1_sum__1118_comb + 25'h000_0001;
  assign p1_add_70569_comb = p1_sum__1097_comb + 25'h000_0001;
  assign p1_add_70570_comb = p1_sum__1091_comb + 25'h000_0001;
  assign p1_add_70571_comb = p1_sum__1119_comb + 25'h000_0001;
  assign p1_add_70572_comb = p1_sum__1112_comb + 25'h000_0001;
  assign p1_add_70573_comb = p1_sum__1092_comb + 25'h000_0001;
  assign p1_add_70574_comb = p1_sum__1087_comb + 25'h000_0001;
  assign p1_add_70575_comb = p1_sum__1113_comb + 25'h000_0001;
  assign p1_add_70576_comb = p1_sum__1106_comb + 25'h000_0001;
  assign p1_add_70577_comb = p1_sum__1088_comb + 25'h000_0001;
  assign p1_add_70578_comb = p1_sum__1084_comb + 25'h000_0001;
  assign p1_add_70579_comb = p1_sum__1107_comb + 25'h000_0001;
  assign p1_add_70580_comb = p1_sum__1100_comb + 25'h000_0001;
  assign p1_add_70581_comb = p1_sum__1085_comb + 25'h000_0001;
  assign p1_add_70582_comb = p1_sum__1082_comb + 25'h000_0001;
  assign p1_add_70585_comb = p1_sum__1135_comb + 25'h000_0001;
  assign p1_add_70586_comb = p1_sum__1101_comb + 25'h000_0001;
  assign p1_add_70587_comb = p1_sum__1134_comb + 25'h000_0001;
  assign p1_add_70588_comb = p1_sum__1095_comb + 25'h000_0001;
  assign p1_add_70589_comb = p1_sum__1132_comb + 25'h000_0001;
  assign p1_add_70590_comb = p1_sum__1090_comb + 25'h000_0001;
  assign p1_add_70591_comb = p1_sum__1129_comb + 25'h000_0001;
  assign p1_add_70592_comb = p1_sum__1086_comb + 25'h000_0001;
  assign p1_add_70593_comb = p1_sum__1125_comb + 25'h000_0001;
  assign p1_add_70594_comb = p1_sum__1083_comb + 25'h000_0001;
  assign p1_add_70595_comb = p1_sum__1120_comb + 25'h000_0001;
  assign p1_add_70596_comb = p1_sum__1081_comb + 25'h000_0001;
  assign p1_add_70597_comb = p1_sum__1114_comb + 25'h000_0001;
  assign p1_add_70598_comb = p1_sum__1080_comb + 25'h000_0001;
  assign p1_sgt_70616_comb = $signed(p1_add_70535_comb[24:1]) > $signed(24'h00_07ff);
  assign p1_bit_slice_70617_comb = p1_add_70535_comb[12:1];
  assign p1_sgt_70619_comb = $signed(p1_add_70536_comb[24:1]) > $signed(24'h00_07ff);
  assign p1_bit_slice_70620_comb = p1_add_70536_comb[12:1];
  assign p1_sgt_70622_comb = $signed(p1_add_70551_comb[24:1]) > $signed(24'h00_07ff);
  assign p1_bit_slice_70623_comb = p1_add_70551_comb[12:1];
  assign p1_sgt_70625_comb = $signed(p1_add_70552_comb[24:1]) > $signed(24'h00_07ff);
  assign p1_bit_slice_70626_comb = p1_add_70552_comb[12:1];
  assign p1_sgt_70628_comb = $signed(p1_add_70553_comb[24:1]) > $signed(24'h00_07ff);
  assign p1_bit_slice_70629_comb = p1_add_70553_comb[12:1];
  assign p1_sgt_70631_comb = $signed(p1_add_70554_comb[24:1]) > $signed(24'h00_07ff);
  assign p1_bit_slice_70632_comb = p1_add_70554_comb[12:1];
  assign p1_sgt_70634_comb = $signed(p1_add_70583_comb[24:1]) > $signed(24'h00_07ff);
  assign p1_bit_slice_70635_comb = p1_add_70583_comb[12:1];
  assign p1_sgt_70637_comb = $signed(p1_add_70584_comb[24:1]) > $signed(24'h00_07ff);
  assign p1_bit_slice_70638_comb = p1_add_70584_comb[12:1];
  assign p1_slt_70639_comb = $signed(p1_add_70535_comb[24:1]) < $signed(24'hff_f800);
  assign p1_slt_70640_comb = $signed(p1_add_70536_comb[24:1]) < $signed(24'hff_f800);
  assign p1_slt_70641_comb = $signed(p1_add_70551_comb[24:1]) < $signed(24'hff_f800);
  assign p1_slt_70642_comb = $signed(p1_add_70552_comb[24:1]) < $signed(24'hff_f800);
  assign p1_slt_70643_comb = $signed(p1_add_70553_comb[24:1]) < $signed(24'hff_f800);
  assign p1_slt_70644_comb = $signed(p1_add_70554_comb[24:1]) < $signed(24'hff_f800);
  assign p1_slt_70645_comb = $signed(p1_add_70583_comb[24:1]) < $signed(24'hff_f800);
  assign p1_slt_70646_comb = $signed(p1_add_70584_comb[24:1]) < $signed(24'hff_f800);

  // Registers for pipe stage 1:
  reg [24:0] p1_add_70537;
  reg [24:0] p1_add_70538;
  reg [24:0] p1_add_70539;
  reg [24:0] p1_add_70540;
  reg [24:0] p1_add_70541;
  reg [24:0] p1_add_70542;
  reg [24:0] p1_add_70543;
  reg [24:0] p1_add_70544;
  reg [24:0] p1_add_70545;
  reg [24:0] p1_add_70546;
  reg [24:0] p1_add_70547;
  reg [24:0] p1_add_70548;
  reg [24:0] p1_add_70549;
  reg [24:0] p1_add_70550;
  reg [24:0] p1_add_70555;
  reg [24:0] p1_add_70556;
  reg [24:0] p1_add_70557;
  reg [24:0] p1_add_70558;
  reg [24:0] p1_add_70559;
  reg [24:0] p1_add_70560;
  reg [24:0] p1_add_70561;
  reg [24:0] p1_add_70562;
  reg [24:0] p1_add_70563;
  reg [24:0] p1_add_70564;
  reg [24:0] p1_add_70565;
  reg [24:0] p1_add_70566;
  reg [24:0] p1_add_70567;
  reg [24:0] p1_add_70568;
  reg [24:0] p1_add_70569;
  reg [24:0] p1_add_70570;
  reg [24:0] p1_add_70571;
  reg [24:0] p1_add_70572;
  reg [24:0] p1_add_70573;
  reg [24:0] p1_add_70574;
  reg [24:0] p1_add_70575;
  reg [24:0] p1_add_70576;
  reg [24:0] p1_add_70577;
  reg [24:0] p1_add_70578;
  reg [24:0] p1_add_70579;
  reg [24:0] p1_add_70580;
  reg [24:0] p1_add_70581;
  reg [24:0] p1_add_70582;
  reg [24:0] p1_add_70585;
  reg [24:0] p1_add_70586;
  reg [24:0] p1_add_70587;
  reg [24:0] p1_add_70588;
  reg [24:0] p1_add_70589;
  reg [24:0] p1_add_70590;
  reg [24:0] p1_add_70591;
  reg [24:0] p1_add_70592;
  reg [24:0] p1_add_70593;
  reg [24:0] p1_add_70594;
  reg [24:0] p1_add_70595;
  reg [24:0] p1_add_70596;
  reg [24:0] p1_add_70597;
  reg [24:0] p1_add_70598;
  reg p1_sgt_70616;
  reg [11:0] p1_bit_slice_70617;
  reg p1_sgt_70619;
  reg [11:0] p1_bit_slice_70620;
  reg p1_sgt_70622;
  reg [11:0] p1_bit_slice_70623;
  reg p1_sgt_70625;
  reg [11:0] p1_bit_slice_70626;
  reg p1_sgt_70628;
  reg [11:0] p1_bit_slice_70629;
  reg p1_sgt_70631;
  reg [11:0] p1_bit_slice_70632;
  reg p1_sgt_70634;
  reg [11:0] p1_bit_slice_70635;
  reg p1_sgt_70637;
  reg [11:0] p1_bit_slice_70638;
  reg p1_slt_70639;
  reg p1_slt_70640;
  reg p1_slt_70641;
  reg p1_slt_70642;
  reg p1_slt_70643;
  reg p1_slt_70644;
  reg p1_slt_70645;
  reg p1_slt_70646;
  always @ (posedge clk) begin
    p1_add_70537 <= p1_add_70537_comb;
    p1_add_70538 <= p1_add_70538_comb;
    p1_add_70539 <= p1_add_70539_comb;
    p1_add_70540 <= p1_add_70540_comb;
    p1_add_70541 <= p1_add_70541_comb;
    p1_add_70542 <= p1_add_70542_comb;
    p1_add_70543 <= p1_add_70543_comb;
    p1_add_70544 <= p1_add_70544_comb;
    p1_add_70545 <= p1_add_70545_comb;
    p1_add_70546 <= p1_add_70546_comb;
    p1_add_70547 <= p1_add_70547_comb;
    p1_add_70548 <= p1_add_70548_comb;
    p1_add_70549 <= p1_add_70549_comb;
    p1_add_70550 <= p1_add_70550_comb;
    p1_add_70555 <= p1_add_70555_comb;
    p1_add_70556 <= p1_add_70556_comb;
    p1_add_70557 <= p1_add_70557_comb;
    p1_add_70558 <= p1_add_70558_comb;
    p1_add_70559 <= p1_add_70559_comb;
    p1_add_70560 <= p1_add_70560_comb;
    p1_add_70561 <= p1_add_70561_comb;
    p1_add_70562 <= p1_add_70562_comb;
    p1_add_70563 <= p1_add_70563_comb;
    p1_add_70564 <= p1_add_70564_comb;
    p1_add_70565 <= p1_add_70565_comb;
    p1_add_70566 <= p1_add_70566_comb;
    p1_add_70567 <= p1_add_70567_comb;
    p1_add_70568 <= p1_add_70568_comb;
    p1_add_70569 <= p1_add_70569_comb;
    p1_add_70570 <= p1_add_70570_comb;
    p1_add_70571 <= p1_add_70571_comb;
    p1_add_70572 <= p1_add_70572_comb;
    p1_add_70573 <= p1_add_70573_comb;
    p1_add_70574 <= p1_add_70574_comb;
    p1_add_70575 <= p1_add_70575_comb;
    p1_add_70576 <= p1_add_70576_comb;
    p1_add_70577 <= p1_add_70577_comb;
    p1_add_70578 <= p1_add_70578_comb;
    p1_add_70579 <= p1_add_70579_comb;
    p1_add_70580 <= p1_add_70580_comb;
    p1_add_70581 <= p1_add_70581_comb;
    p1_add_70582 <= p1_add_70582_comb;
    p1_add_70585 <= p1_add_70585_comb;
    p1_add_70586 <= p1_add_70586_comb;
    p1_add_70587 <= p1_add_70587_comb;
    p1_add_70588 <= p1_add_70588_comb;
    p1_add_70589 <= p1_add_70589_comb;
    p1_add_70590 <= p1_add_70590_comb;
    p1_add_70591 <= p1_add_70591_comb;
    p1_add_70592 <= p1_add_70592_comb;
    p1_add_70593 <= p1_add_70593_comb;
    p1_add_70594 <= p1_add_70594_comb;
    p1_add_70595 <= p1_add_70595_comb;
    p1_add_70596 <= p1_add_70596_comb;
    p1_add_70597 <= p1_add_70597_comb;
    p1_add_70598 <= p1_add_70598_comb;
    p1_sgt_70616 <= p1_sgt_70616_comb;
    p1_bit_slice_70617 <= p1_bit_slice_70617_comb;
    p1_sgt_70619 <= p1_sgt_70619_comb;
    p1_bit_slice_70620 <= p1_bit_slice_70620_comb;
    p1_sgt_70622 <= p1_sgt_70622_comb;
    p1_bit_slice_70623 <= p1_bit_slice_70623_comb;
    p1_sgt_70625 <= p1_sgt_70625_comb;
    p1_bit_slice_70626 <= p1_bit_slice_70626_comb;
    p1_sgt_70628 <= p1_sgt_70628_comb;
    p1_bit_slice_70629 <= p1_bit_slice_70629_comb;
    p1_sgt_70631 <= p1_sgt_70631_comb;
    p1_bit_slice_70632 <= p1_bit_slice_70632_comb;
    p1_sgt_70634 <= p1_sgt_70634_comb;
    p1_bit_slice_70635 <= p1_bit_slice_70635_comb;
    p1_sgt_70637 <= p1_sgt_70637_comb;
    p1_bit_slice_70638 <= p1_bit_slice_70638_comb;
    p1_slt_70639 <= p1_slt_70639_comb;
    p1_slt_70640 <= p1_slt_70640_comb;
    p1_slt_70641 <= p1_slt_70641_comb;
    p1_slt_70642 <= p1_slt_70642_comb;
    p1_slt_70643 <= p1_slt_70643_comb;
    p1_slt_70644 <= p1_slt_70644_comb;
    p1_slt_70645 <= p1_slt_70645_comb;
    p1_slt_70646 <= p1_slt_70646_comb;
  end

  // ===== Pipe stage 2:
  wire [11:0] p2_clipped__56_comb;
  wire [11:0] p2_clipped__72_comb;
  wire [11:0] p2_clipped__24_comb;
  wire [11:0] p2_clipped__40_comb;
  wire [11:0] p2_clipped__88_comb;
  wire [11:0] p2_clipped__104_comb;
  wire [11:0] p2_clipped__8_comb;
  wire [11:0] p2_clipped__120_comb;
  wire [17:0] p2_smul_28634_NarrowedMult__comb;
  wire [17:0] p2_smul_28636_NarrowedMult__comb;
  wire [18:0] p2_smul_28758_NarrowedMult__comb;
  wire [18:0] p2_smul_28760_NarrowedMult__comb;
  wire [18:0] p2_smul_28766_NarrowedMult__comb;
  wire [18:0] p2_smul_28768_NarrowedMult__comb;
  wire [17:0] p2_smul_28886_NarrowedMult__comb;
  wire [17:0] p2_smul_28896_NarrowedMult__comb;
  wire [17:0] p2_smul_29144_NarrowedMult__comb;
  wire [17:0] p2_smul_29150_NarrowedMult__comb;
  wire [18:0] p2_smul_29268_NarrowedMult__comb;
  wire [18:0] p2_smul_29272_NarrowedMult__comb;
  wire [18:0] p2_smul_29278_NarrowedMult__comb;
  wire [18:0] p2_smul_29282_NarrowedMult__comb;
  wire [17:0] p2_smul_29396_NarrowedMult__comb;
  wire [17:0] p2_smul_29410_NarrowedMult__comb;
  wire [20:0] p2_smul_72231_comb;
  wire [20:0] p2_smul_72232_comb;
  wire [20:0] p2_smul_72233_comb;
  wire [20:0] p2_smul_72234_comb;
  wire [20:0] p2_smul_72235_comb;
  wire [20:0] p2_smul_72236_comb;
  wire [20:0] p2_smul_72237_comb;
  wire [20:0] p2_smul_72238_comb;
  wire [11:0] p2_clipped__9_comb;
  wire [11:0] p2_clipped__25_comb;
  wire [11:0] p2_clipped__41_comb;
  wire [11:0] p2_clipped__57_comb;
  wire [11:0] p2_clipped__73_comb;
  wire [11:0] p2_clipped__89_comb;
  wire [11:0] p2_clipped__105_comb;
  wire [11:0] p2_clipped__121_comb;
  wire [11:0] p2_clipped__10_comb;
  wire [11:0] p2_clipped__26_comb;
  wire [11:0] p2_clipped__42_comb;
  wire [11:0] p2_clipped__58_comb;
  wire [11:0] p2_clipped__74_comb;
  wire [11:0] p2_clipped__90_comb;
  wire [11:0] p2_clipped__106_comb;
  wire [11:0] p2_clipped__122_comb;
  wire [11:0] p2_clipped__11_comb;
  wire [11:0] p2_clipped__27_comb;
  wire [11:0] p2_clipped__43_comb;
  wire [11:0] p2_clipped__59_comb;
  wire [11:0] p2_clipped__75_comb;
  wire [11:0] p2_clipped__91_comb;
  wire [11:0] p2_clipped__107_comb;
  wire [11:0] p2_clipped__123_comb;
  wire [11:0] p2_clipped__12_comb;
  wire [11:0] p2_clipped__28_comb;
  wire [11:0] p2_clipped__44_comb;
  wire [11:0] p2_clipped__60_comb;
  wire [11:0] p2_clipped__76_comb;
  wire [11:0] p2_clipped__92_comb;
  wire [11:0] p2_clipped__108_comb;
  wire [11:0] p2_clipped__124_comb;
  wire [11:0] p2_clipped__13_comb;
  wire [11:0] p2_clipped__29_comb;
  wire [11:0] p2_clipped__45_comb;
  wire [11:0] p2_clipped__61_comb;
  wire [11:0] p2_clipped__77_comb;
  wire [11:0] p2_clipped__93_comb;
  wire [11:0] p2_clipped__109_comb;
  wire [11:0] p2_clipped__125_comb;
  wire [11:0] p2_clipped__14_comb;
  wire [11:0] p2_clipped__30_comb;
  wire [11:0] p2_clipped__46_comb;
  wire [11:0] p2_clipped__62_comb;
  wire [11:0] p2_clipped__78_comb;
  wire [11:0] p2_clipped__94_comb;
  wire [11:0] p2_clipped__110_comb;
  wire [11:0] p2_clipped__126_comb;
  wire [11:0] p2_clipped__15_comb;
  wire [11:0] p2_clipped__31_comb;
  wire [11:0] p2_clipped__47_comb;
  wire [11:0] p2_clipped__63_comb;
  wire [11:0] p2_clipped__79_comb;
  wire [11:0] p2_clipped__95_comb;
  wire [11:0] p2_clipped__111_comb;
  wire [11:0] p2_clipped__127_comb;
  wire [20:0] p2_smul_71975_comb;
  wire [20:0] p2_smul_71976_comb;
  wire [19:0] p2_smul_28632_NarrowedMult__comb;
  wire [19:0] p2_smul_28638_NarrowedMult__comb;
  wire [20:0] p2_smul_71983_comb;
  wire [20:0] p2_smul_71984_comb;
  wire [18:0] p2_smul_28756_NarrowedMult__comb;
  wire [18:0] p2_smul_28762_NarrowedMult__comb;
  wire [18:0] p2_smul_28764_NarrowedMult__comb;
  wire [18:0] p2_smul_28770_NarrowedMult__comb;
  wire [20:0] p2_smul_72151_comb;
  wire [20:0] p2_smul_72154_comb;
  wire [19:0] p2_smul_28890_NarrowedMult__comb;
  wire [19:0] p2_smul_28892_NarrowedMult__comb;
  wire [20:0] p2_smul_72157_comb;
  wire [20:0] p2_smul_72160_comb;
  wire [19:0] p2_smul_29140_NarrowedMult__comb;
  wire [20:0] p2_smul_72296_comb;
  wire [20:0] p2_smul_72299_comb;
  wire [20:0] p2_smul_72300_comb;
  wire [20:0] p2_smul_72303_comb;
  wire [19:0] p2_smul_29154_NarrowedMult__comb;
  wire [18:0] p2_smul_29270_NarrowedMult__comb;
  wire [18:0] p2_smul_29274_NarrowedMult__comb;
  wire [18:0] p2_smul_29276_NarrowedMult__comb;
  wire [18:0] p2_smul_29280_NarrowedMult__comb;
  wire [19:0] p2_smul_29398_NarrowedMult__comb;
  wire [20:0] p2_smul_72474_comb;
  wire [20:0] p2_smul_72475_comb;
  wire [20:0] p2_smul_72476_comb;
  wire [20:0] p2_smul_72477_comb;
  wire [19:0] p2_smul_29408_NarrowedMult__comb;
  wire [20:0] p2_smul_72239_comb;
  wire [20:0] p2_smul_72240_comb;
  wire [20:0] p2_smul_72241_comb;
  wire [20:0] p2_smul_72242_comb;
  wire [20:0] p2_smul_72243_comb;
  wire [20:0] p2_smul_72244_comb;
  wire [20:0] p2_smul_72245_comb;
  wire [20:0] p2_smul_72246_comb;
  wire [20:0] p2_smul_72247_comb;
  wire [20:0] p2_smul_72248_comb;
  wire [20:0] p2_smul_72249_comb;
  wire [20:0] p2_smul_72250_comb;
  wire [20:0] p2_smul_72251_comb;
  wire [20:0] p2_smul_72252_comb;
  wire [20:0] p2_smul_72253_comb;
  wire [20:0] p2_smul_72254_comb;
  wire [20:0] p2_smul_72255_comb;
  wire [20:0] p2_smul_72256_comb;
  wire [20:0] p2_smul_72257_comb;
  wire [20:0] p2_smul_72258_comb;
  wire [20:0] p2_smul_72259_comb;
  wire [20:0] p2_smul_72260_comb;
  wire [20:0] p2_smul_72261_comb;
  wire [20:0] p2_smul_72262_comb;
  wire [20:0] p2_smul_72263_comb;
  wire [20:0] p2_smul_72264_comb;
  wire [20:0] p2_smul_72265_comb;
  wire [20:0] p2_smul_72266_comb;
  wire [20:0] p2_smul_72267_comb;
  wire [20:0] p2_smul_72268_comb;
  wire [20:0] p2_smul_72269_comb;
  wire [20:0] p2_smul_72270_comb;
  wire [20:0] p2_smul_72271_comb;
  wire [20:0] p2_smul_72272_comb;
  wire [20:0] p2_smul_72273_comb;
  wire [20:0] p2_smul_72274_comb;
  wire [20:0] p2_smul_72275_comb;
  wire [20:0] p2_smul_72276_comb;
  wire [20:0] p2_smul_72277_comb;
  wire [20:0] p2_smul_72278_comb;
  wire [20:0] p2_smul_72279_comb;
  wire [20:0] p2_smul_72280_comb;
  wire [20:0] p2_smul_72281_comb;
  wire [20:0] p2_smul_72282_comb;
  wire [20:0] p2_smul_72283_comb;
  wire [20:0] p2_smul_72284_comb;
  wire [20:0] p2_smul_72285_comb;
  wire [20:0] p2_smul_72286_comb;
  wire [20:0] p2_smul_72287_comb;
  wire [20:0] p2_smul_72288_comb;
  wire [20:0] p2_smul_72289_comb;
  wire [20:0] p2_smul_72290_comb;
  wire [20:0] p2_smul_72291_comb;
  wire [20:0] p2_smul_72292_comb;
  wire [20:0] p2_smul_72293_comb;
  wire [20:0] p2_smul_72294_comb;
  wire [11:0] p2_add_72621_comb;
  wire [11:0] p2_add_72622_comb;
  wire [12:0] p2_add_72729_comb;
  wire [12:0] p2_add_72730_comb;
  wire [12:0] p2_add_72735_comb;
  wire [12:0] p2_add_72736_comb;
  wire [11:0] p2_add_72825_comb;
  wire [11:0] p2_add_72834_comb;
  wire [11:0] p2_add_73067_comb;
  wire [11:0] p2_add_73072_comb;
  wire [12:0] p2_add_73175_comb;
  wire [12:0] p2_add_73178_comb;
  wire [12:0] p2_add_73183_comb;
  wire [12:0] p2_add_73186_comb;
  wire [11:0] p2_add_73271_comb;
  wire [11:0] p2_add_73284_comb;
  wire [12:0] p2_add_73383_comb;
  wire [12:0] p2_add_73384_comb;
  wire [12:0] p2_add_73385_comb;
  wire [12:0] p2_add_73386_comb;
  wire [13:0] p2_add_73607_comb;
  wire [13:0] p2_add_73608_comb;
  wire [13:0] p2_add_73609_comb;
  wire [13:0] p2_add_73610_comb;
  wire [13:0] p2_add_73611_comb;
  wire [13:0] p2_add_73612_comb;
  wire [13:0] p2_add_73613_comb;
  wire [13:0] p2_add_73614_comb;
  wire [17:0] p2_smul_28650_NarrowedMult__comb;
  wire [17:0] p2_smul_28652_NarrowedMult__comb;
  wire [17:0] p2_smul_28666_NarrowedMult__comb;
  wire [17:0] p2_smul_28668_NarrowedMult__comb;
  wire [17:0] p2_smul_28682_NarrowedMult__comb;
  wire [17:0] p2_smul_28684_NarrowedMult__comb;
  wire [17:0] p2_smul_28698_NarrowedMult__comb;
  wire [17:0] p2_smul_28700_NarrowedMult__comb;
  wire [17:0] p2_smul_28714_NarrowedMult__comb;
  wire [17:0] p2_smul_28716_NarrowedMult__comb;
  wire [17:0] p2_smul_28730_NarrowedMult__comb;
  wire [17:0] p2_smul_28732_NarrowedMult__comb;
  wire [17:0] p2_smul_28746_NarrowedMult__comb;
  wire [17:0] p2_smul_28748_NarrowedMult__comb;
  wire [18:0] p2_smul_28774_NarrowedMult__comb;
  wire [18:0] p2_smul_28776_NarrowedMult__comb;
  wire [18:0] p2_smul_28782_NarrowedMult__comb;
  wire [18:0] p2_smul_28784_NarrowedMult__comb;
  wire [18:0] p2_smul_28790_NarrowedMult__comb;
  wire [18:0] p2_smul_28792_NarrowedMult__comb;
  wire [18:0] p2_smul_28798_NarrowedMult__comb;
  wire [18:0] p2_smul_28800_NarrowedMult__comb;
  wire [18:0] p2_smul_28806_NarrowedMult__comb;
  wire [18:0] p2_smul_28808_NarrowedMult__comb;
  wire [18:0] p2_smul_28814_NarrowedMult__comb;
  wire [18:0] p2_smul_28816_NarrowedMult__comb;
  wire [18:0] p2_smul_28822_NarrowedMult__comb;
  wire [18:0] p2_smul_28824_NarrowedMult__comb;
  wire [18:0] p2_smul_28830_NarrowedMult__comb;
  wire [18:0] p2_smul_28832_NarrowedMult__comb;
  wire [18:0] p2_smul_28838_NarrowedMult__comb;
  wire [18:0] p2_smul_28840_NarrowedMult__comb;
  wire [18:0] p2_smul_28846_NarrowedMult__comb;
  wire [18:0] p2_smul_28848_NarrowedMult__comb;
  wire [18:0] p2_smul_28854_NarrowedMult__comb;
  wire [18:0] p2_smul_28856_NarrowedMult__comb;
  wire [18:0] p2_smul_28862_NarrowedMult__comb;
  wire [18:0] p2_smul_28864_NarrowedMult__comb;
  wire [18:0] p2_smul_28870_NarrowedMult__comb;
  wire [18:0] p2_smul_28872_NarrowedMult__comb;
  wire [18:0] p2_smul_28878_NarrowedMult__comb;
  wire [18:0] p2_smul_28880_NarrowedMult__comb;
  wire [17:0] p2_smul_28902_NarrowedMult__comb;
  wire [17:0] p2_smul_28912_NarrowedMult__comb;
  wire [17:0] p2_smul_28918_NarrowedMult__comb;
  wire [17:0] p2_smul_28928_NarrowedMult__comb;
  wire [17:0] p2_smul_28934_NarrowedMult__comb;
  wire [17:0] p2_smul_28944_NarrowedMult__comb;
  wire [17:0] p2_smul_28950_NarrowedMult__comb;
  wire [17:0] p2_smul_28960_NarrowedMult__comb;
  wire [17:0] p2_smul_28966_NarrowedMult__comb;
  wire [17:0] p2_smul_28976_NarrowedMult__comb;
  wire [17:0] p2_smul_28982_NarrowedMult__comb;
  wire [17:0] p2_smul_28992_NarrowedMult__comb;
  wire [17:0] p2_smul_28998_NarrowedMult__comb;
  wire [17:0] p2_smul_29008_NarrowedMult__comb;
  wire [17:0] p2_smul_29160_NarrowedMult__comb;
  wire [17:0] p2_smul_29166_NarrowedMult__comb;
  wire [17:0] p2_smul_29176_NarrowedMult__comb;
  wire [17:0] p2_smul_29182_NarrowedMult__comb;
  wire [17:0] p2_smul_29192_NarrowedMult__comb;
  wire [17:0] p2_smul_29198_NarrowedMult__comb;
  wire [17:0] p2_smul_29208_NarrowedMult__comb;
  wire [17:0] p2_smul_29214_NarrowedMult__comb;
  wire [17:0] p2_smul_29224_NarrowedMult__comb;
  wire [17:0] p2_smul_29230_NarrowedMult__comb;
  wire [17:0] p2_smul_29240_NarrowedMult__comb;
  wire [17:0] p2_smul_29246_NarrowedMult__comb;
  wire [17:0] p2_smul_29256_NarrowedMult__comb;
  wire [17:0] p2_smul_29262_NarrowedMult__comb;
  wire [18:0] p2_smul_29284_NarrowedMult__comb;
  wire [18:0] p2_smul_29288_NarrowedMult__comb;
  wire [18:0] p2_smul_29294_NarrowedMult__comb;
  wire [18:0] p2_smul_29298_NarrowedMult__comb;
  wire [18:0] p2_smul_29300_NarrowedMult__comb;
  wire [18:0] p2_smul_29304_NarrowedMult__comb;
  wire [18:0] p2_smul_29310_NarrowedMult__comb;
  wire [18:0] p2_smul_29314_NarrowedMult__comb;
  wire [18:0] p2_smul_29316_NarrowedMult__comb;
  wire [18:0] p2_smul_29320_NarrowedMult__comb;
  wire [18:0] p2_smul_29326_NarrowedMult__comb;
  wire [18:0] p2_smul_29330_NarrowedMult__comb;
  wire [18:0] p2_smul_29332_NarrowedMult__comb;
  wire [18:0] p2_smul_29336_NarrowedMult__comb;
  wire [18:0] p2_smul_29342_NarrowedMult__comb;
  wire [18:0] p2_smul_29346_NarrowedMult__comb;
  wire [18:0] p2_smul_29348_NarrowedMult__comb;
  wire [18:0] p2_smul_29352_NarrowedMult__comb;
  wire [18:0] p2_smul_29358_NarrowedMult__comb;
  wire [18:0] p2_smul_29362_NarrowedMult__comb;
  wire [18:0] p2_smul_29364_NarrowedMult__comb;
  wire [18:0] p2_smul_29368_NarrowedMult__comb;
  wire [18:0] p2_smul_29374_NarrowedMult__comb;
  wire [18:0] p2_smul_29378_NarrowedMult__comb;
  wire [18:0] p2_smul_29380_NarrowedMult__comb;
  wire [18:0] p2_smul_29384_NarrowedMult__comb;
  wire [18:0] p2_smul_29390_NarrowedMult__comb;
  wire [18:0] p2_smul_29394_NarrowedMult__comb;
  wire [17:0] p2_smul_29412_NarrowedMult__comb;
  wire [17:0] p2_smul_29426_NarrowedMult__comb;
  wire [17:0] p2_smul_29428_NarrowedMult__comb;
  wire [17:0] p2_smul_29442_NarrowedMult__comb;
  wire [17:0] p2_smul_29444_NarrowedMult__comb;
  wire [17:0] p2_smul_29458_NarrowedMult__comb;
  wire [17:0] p2_smul_29460_NarrowedMult__comb;
  wire [17:0] p2_smul_29474_NarrowedMult__comb;
  wire [17:0] p2_smul_29476_NarrowedMult__comb;
  wire [17:0] p2_smul_29490_NarrowedMult__comb;
  wire [17:0] p2_smul_29492_NarrowedMult__comb;
  wire [17:0] p2_smul_29506_NarrowedMult__comb;
  wire [17:0] p2_smul_29508_NarrowedMult__comb;
  wire [17:0] p2_smul_29522_NarrowedMult__comb;
  wire [12:0] p2_add_73387_comb;
  wire [12:0] p2_add_73388_comb;
  wire [12:0] p2_add_73389_comb;
  wire [12:0] p2_add_73390_comb;
  wire [12:0] p2_add_73391_comb;
  wire [12:0] p2_add_73392_comb;
  wire [12:0] p2_add_73393_comb;
  wire [12:0] p2_add_73394_comb;
  wire [12:0] p2_add_73395_comb;
  wire [12:0] p2_add_73396_comb;
  wire [12:0] p2_add_73397_comb;
  wire [12:0] p2_add_73398_comb;
  wire [12:0] p2_add_73399_comb;
  wire [12:0] p2_add_73400_comb;
  wire [12:0] p2_add_73401_comb;
  wire [12:0] p2_add_73402_comb;
  wire [12:0] p2_add_73403_comb;
  wire [12:0] p2_add_73404_comb;
  wire [12:0] p2_add_73405_comb;
  wire [12:0] p2_add_73406_comb;
  wire [12:0] p2_add_73407_comb;
  wire [12:0] p2_add_73408_comb;
  wire [12:0] p2_add_73409_comb;
  wire [12:0] p2_add_73410_comb;
  wire [12:0] p2_add_73411_comb;
  wire [12:0] p2_add_73412_comb;
  wire [12:0] p2_add_73413_comb;
  wire [12:0] p2_add_73414_comb;
  wire [13:0] p2_add_73415_comb;
  wire [13:0] p2_add_73416_comb;
  wire [13:0] p2_add_73417_comb;
  wire [10:0] p2_bit_slice_73418_comb;
  wire [10:0] p2_bit_slice_73419_comb;
  wire [13:0] p2_add_73420_comb;
  wire [13:0] p2_add_73421_comb;
  wire [13:0] p2_add_73422_comb;
  wire [13:0] p2_add_73479_comb;
  wire [11:0] p2_bit_slice_73480_comb;
  wire [11:0] p2_bit_slice_73481_comb;
  wire [13:0] p2_add_73482_comb;
  wire [13:0] p2_add_73483_comb;
  wire [11:0] p2_bit_slice_73484_comb;
  wire [11:0] p2_bit_slice_73485_comb;
  wire [13:0] p2_add_73486_comb;
  wire [13:0] p2_add_73543_comb;
  wire [10:0] p2_bit_slice_73544_comb;
  wire [13:0] p2_add_73545_comb;
  wire [13:0] p2_add_73546_comb;
  wire [13:0] p2_add_73547_comb;
  wire [13:0] p2_add_73548_comb;
  wire [10:0] p2_bit_slice_73549_comb;
  wire [13:0] p2_add_73550_comb;
  wire [13:0] p2_add_73671_comb;
  wire [13:0] p2_add_73672_comb;
  wire [10:0] p2_bit_slice_73673_comb;
  wire [13:0] p2_add_73674_comb;
  wire [13:0] p2_add_73675_comb;
  wire [10:0] p2_bit_slice_73676_comb;
  wire [13:0] p2_add_73677_comb;
  wire [13:0] p2_add_73678_comb;
  wire [11:0] p2_bit_slice_73735_comb;
  wire [13:0] p2_add_73736_comb;
  wire [11:0] p2_bit_slice_73737_comb;
  wire [13:0] p2_add_73738_comb;
  wire [13:0] p2_add_73739_comb;
  wire [11:0] p2_bit_slice_73740_comb;
  wire [13:0] p2_add_73741_comb;
  wire [11:0] p2_bit_slice_73742_comb;
  wire [10:0] p2_bit_slice_73799_comb;
  wire [13:0] p2_add_73800_comb;
  wire [13:0] p2_add_73801_comb;
  wire [13:0] p2_add_73802_comb;
  wire [13:0] p2_add_73803_comb;
  wire [13:0] p2_add_73804_comb;
  wire [13:0] p2_add_73805_comb;
  wire [10:0] p2_bit_slice_73806_comb;
  wire [31:0] p2_sum__520_comb;
  wire [31:0] p2_sum__521_comb;
  wire [31:0] p2_sum__522_comb;
  wire [31:0] p2_sum__523_comb;
  wire [20:0] p2_smul_71985_comb;
  wire [20:0] p2_smul_71986_comb;
  wire [19:0] p2_smul_28648_NarrowedMult__comb;
  wire [19:0] p2_smul_28654_NarrowedMult__comb;
  wire [20:0] p2_smul_71993_comb;
  wire [20:0] p2_smul_71994_comb;
  wire [20:0] p2_smul_71995_comb;
  wire [20:0] p2_smul_71996_comb;
  wire [19:0] p2_smul_28664_NarrowedMult__comb;
  wire [19:0] p2_smul_28670_NarrowedMult__comb;
  wire [20:0] p2_smul_72003_comb;
  wire [20:0] p2_smul_72004_comb;
  wire [20:0] p2_smul_72005_comb;
  wire [20:0] p2_smul_72006_comb;
  wire [19:0] p2_smul_28680_NarrowedMult__comb;
  wire [19:0] p2_smul_28686_NarrowedMult__comb;
  wire [20:0] p2_smul_72013_comb;
  wire [20:0] p2_smul_72014_comb;
  wire [20:0] p2_smul_72015_comb;
  wire [20:0] p2_smul_72016_comb;
  wire [19:0] p2_smul_28696_NarrowedMult__comb;
  wire [19:0] p2_smul_28702_NarrowedMult__comb;
  wire [20:0] p2_smul_72023_comb;
  wire [20:0] p2_smul_72024_comb;
  wire [20:0] p2_smul_72025_comb;
  wire [20:0] p2_smul_72026_comb;
  wire [19:0] p2_smul_28712_NarrowedMult__comb;
  wire [19:0] p2_smul_28718_NarrowedMult__comb;
  wire [20:0] p2_smul_72033_comb;
  wire [20:0] p2_smul_72034_comb;
  wire [20:0] p2_smul_72035_comb;
  wire [20:0] p2_smul_72036_comb;
  wire [19:0] p2_smul_28728_NarrowedMult__comb;
  wire [19:0] p2_smul_28734_NarrowedMult__comb;
  wire [20:0] p2_smul_72043_comb;
  wire [20:0] p2_smul_72044_comb;
  wire [20:0] p2_smul_72045_comb;
  wire [20:0] p2_smul_72046_comb;
  wire [19:0] p2_smul_28744_NarrowedMult__comb;
  wire [19:0] p2_smul_28750_NarrowedMult__comb;
  wire [20:0] p2_smul_72053_comb;
  wire [20:0] p2_smul_72054_comb;
  wire [18:0] p2_smul_28772_NarrowedMult__comb;
  wire [18:0] p2_smul_28778_NarrowedMult__comb;
  wire [18:0] p2_smul_28780_NarrowedMult__comb;
  wire [18:0] p2_smul_28786_NarrowedMult__comb;
  wire [18:0] p2_smul_28788_NarrowedMult__comb;
  wire [18:0] p2_smul_28794_NarrowedMult__comb;
  wire [18:0] p2_smul_28796_NarrowedMult__comb;
  wire [18:0] p2_smul_28802_NarrowedMult__comb;
  wire [18:0] p2_smul_28804_NarrowedMult__comb;
  wire [18:0] p2_smul_28810_NarrowedMult__comb;
  wire [18:0] p2_smul_28812_NarrowedMult__comb;
  wire [18:0] p2_smul_28818_NarrowedMult__comb;
  wire [18:0] p2_smul_28820_NarrowedMult__comb;
  wire [18:0] p2_smul_28826_NarrowedMult__comb;
  wire [18:0] p2_smul_28828_NarrowedMult__comb;
  wire [18:0] p2_smul_28834_NarrowedMult__comb;
  wire [18:0] p2_smul_28836_NarrowedMult__comb;
  wire [18:0] p2_smul_28842_NarrowedMult__comb;
  wire [18:0] p2_smul_28844_NarrowedMult__comb;
  wire [18:0] p2_smul_28850_NarrowedMult__comb;
  wire [18:0] p2_smul_28852_NarrowedMult__comb;
  wire [18:0] p2_smul_28858_NarrowedMult__comb;
  wire [18:0] p2_smul_28860_NarrowedMult__comb;
  wire [18:0] p2_smul_28866_NarrowedMult__comb;
  wire [18:0] p2_smul_28868_NarrowedMult__comb;
  wire [18:0] p2_smul_28874_NarrowedMult__comb;
  wire [18:0] p2_smul_28876_NarrowedMult__comb;
  wire [18:0] p2_smul_28882_NarrowedMult__comb;
  wire [20:0] p2_smul_72161_comb;
  wire [20:0] p2_smul_72164_comb;
  wire [19:0] p2_smul_28906_NarrowedMult__comb;
  wire [19:0] p2_smul_28908_NarrowedMult__comb;
  wire [20:0] p2_smul_72167_comb;
  wire [20:0] p2_smul_72170_comb;
  wire [20:0] p2_smul_72171_comb;
  wire [20:0] p2_smul_72174_comb;
  wire [19:0] p2_smul_28922_NarrowedMult__comb;
  wire [19:0] p2_smul_28924_NarrowedMult__comb;
  wire [20:0] p2_smul_72177_comb;
  wire [20:0] p2_smul_72180_comb;
  wire [20:0] p2_smul_72181_comb;
  wire [20:0] p2_smul_72184_comb;
  wire [19:0] p2_smul_28938_NarrowedMult__comb;
  wire [19:0] p2_smul_28940_NarrowedMult__comb;
  wire [20:0] p2_smul_72187_comb;
  wire [20:0] p2_smul_72190_comb;
  wire [20:0] p2_smul_72191_comb;
  wire [20:0] p2_smul_72194_comb;
  wire [19:0] p2_smul_28954_NarrowedMult__comb;
  wire [19:0] p2_smul_28956_NarrowedMult__comb;
  wire [20:0] p2_smul_72197_comb;
  wire [20:0] p2_smul_72200_comb;
  wire [20:0] p2_smul_72201_comb;
  wire [20:0] p2_smul_72204_comb;
  wire [19:0] p2_smul_28970_NarrowedMult__comb;
  wire [19:0] p2_smul_28972_NarrowedMult__comb;
  wire [20:0] p2_smul_72207_comb;
  wire [20:0] p2_smul_72210_comb;
  wire [20:0] p2_smul_72211_comb;
  wire [20:0] p2_smul_72214_comb;
  wire [19:0] p2_smul_28986_NarrowedMult__comb;
  wire [19:0] p2_smul_28988_NarrowedMult__comb;
  wire [20:0] p2_smul_72217_comb;
  wire [20:0] p2_smul_72220_comb;
  wire [20:0] p2_smul_72221_comb;
  wire [20:0] p2_smul_72224_comb;
  wire [19:0] p2_smul_29002_NarrowedMult__comb;
  wire [19:0] p2_smul_29004_NarrowedMult__comb;
  wire [20:0] p2_smul_72227_comb;
  wire [20:0] p2_smul_72230_comb;
  wire [19:0] p2_smul_29156_NarrowedMult__comb;
  wire [20:0] p2_smul_72306_comb;
  wire [20:0] p2_smul_72309_comb;
  wire [20:0] p2_smul_72310_comb;
  wire [20:0] p2_smul_72313_comb;
  wire [19:0] p2_smul_29170_NarrowedMult__comb;
  wire [19:0] p2_smul_29172_NarrowedMult__comb;
  wire [20:0] p2_smul_72316_comb;
  wire [20:0] p2_smul_72319_comb;
  wire [20:0] p2_smul_72320_comb;
  wire [20:0] p2_smul_72323_comb;
  wire [19:0] p2_smul_29186_NarrowedMult__comb;
  wire [19:0] p2_smul_29188_NarrowedMult__comb;
  wire [20:0] p2_smul_72326_comb;
  wire [20:0] p2_smul_72329_comb;
  wire [20:0] p2_smul_72330_comb;
  wire [20:0] p2_smul_72333_comb;
  wire [19:0] p2_smul_29202_NarrowedMult__comb;
  wire [19:0] p2_smul_29204_NarrowedMult__comb;
  wire [20:0] p2_smul_72336_comb;
  wire [20:0] p2_smul_72339_comb;
  wire [20:0] p2_smul_72340_comb;
  wire [20:0] p2_smul_72343_comb;
  wire [19:0] p2_smul_29218_NarrowedMult__comb;
  wire [19:0] p2_smul_29220_NarrowedMult__comb;
  wire [20:0] p2_smul_72346_comb;
  wire [20:0] p2_smul_72349_comb;
  wire [20:0] p2_smul_72350_comb;
  wire [20:0] p2_smul_72353_comb;
  wire [19:0] p2_smul_29234_NarrowedMult__comb;
  wire [19:0] p2_smul_29236_NarrowedMult__comb;
  wire [20:0] p2_smul_72356_comb;
  wire [20:0] p2_smul_72359_comb;
  wire [20:0] p2_smul_72360_comb;
  wire [20:0] p2_smul_72363_comb;
  wire [19:0] p2_smul_29250_NarrowedMult__comb;
  wire [19:0] p2_smul_29252_NarrowedMult__comb;
  wire [20:0] p2_smul_72366_comb;
  wire [20:0] p2_smul_72369_comb;
  wire [20:0] p2_smul_72370_comb;
  wire [20:0] p2_smul_72373_comb;
  wire [19:0] p2_smul_29266_NarrowedMult__comb;
  wire [18:0] p2_smul_29286_NarrowedMult__comb;
  wire [18:0] p2_smul_29290_NarrowedMult__comb;
  wire [18:0] p2_smul_29292_NarrowedMult__comb;
  wire [18:0] p2_smul_29296_NarrowedMult__comb;
  wire [18:0] p2_smul_29302_NarrowedMult__comb;
  wire [18:0] p2_smul_29306_NarrowedMult__comb;
  wire [18:0] p2_smul_29308_NarrowedMult__comb;
  wire [18:0] p2_smul_29312_NarrowedMult__comb;
  wire [18:0] p2_smul_29318_NarrowedMult__comb;
  wire [18:0] p2_smul_29322_NarrowedMult__comb;
  wire [18:0] p2_smul_29324_NarrowedMult__comb;
  wire [18:0] p2_smul_29328_NarrowedMult__comb;
  wire [18:0] p2_smul_29334_NarrowedMult__comb;
  wire [18:0] p2_smul_29338_NarrowedMult__comb;
  wire [18:0] p2_smul_29340_NarrowedMult__comb;
  wire [18:0] p2_smul_29344_NarrowedMult__comb;
  wire [18:0] p2_smul_29350_NarrowedMult__comb;
  wire [18:0] p2_smul_29354_NarrowedMult__comb;
  wire [18:0] p2_smul_29356_NarrowedMult__comb;
  wire [18:0] p2_smul_29360_NarrowedMult__comb;
  wire [18:0] p2_smul_29366_NarrowedMult__comb;
  wire [18:0] p2_smul_29370_NarrowedMult__comb;
  wire [18:0] p2_smul_29372_NarrowedMult__comb;
  wire [18:0] p2_smul_29376_NarrowedMult__comb;
  wire [18:0] p2_smul_29382_NarrowedMult__comb;
  wire [18:0] p2_smul_29386_NarrowedMult__comb;
  wire [18:0] p2_smul_29388_NarrowedMult__comb;
  wire [18:0] p2_smul_29392_NarrowedMult__comb;
  wire [19:0] p2_smul_29414_NarrowedMult__comb;
  wire [20:0] p2_smul_72484_comb;
  wire [20:0] p2_smul_72485_comb;
  wire [20:0] p2_smul_72486_comb;
  wire [20:0] p2_smul_72487_comb;
  wire [19:0] p2_smul_29424_NarrowedMult__comb;
  wire [19:0] p2_smul_29430_NarrowedMult__comb;
  wire [20:0] p2_smul_72494_comb;
  wire [20:0] p2_smul_72495_comb;
  wire [20:0] p2_smul_72496_comb;
  wire [20:0] p2_smul_72497_comb;
  wire [19:0] p2_smul_29440_NarrowedMult__comb;
  wire [19:0] p2_smul_29446_NarrowedMult__comb;
  wire [20:0] p2_smul_72504_comb;
  wire [20:0] p2_smul_72505_comb;
  wire [20:0] p2_smul_72506_comb;
  wire [20:0] p2_smul_72507_comb;
  wire [19:0] p2_smul_29456_NarrowedMult__comb;
  wire [19:0] p2_smul_29462_NarrowedMult__comb;
  wire [20:0] p2_smul_72514_comb;
  wire [20:0] p2_smul_72515_comb;
  wire [20:0] p2_smul_72516_comb;
  wire [20:0] p2_smul_72517_comb;
  wire [19:0] p2_smul_29472_NarrowedMult__comb;
  wire [19:0] p2_smul_29478_NarrowedMult__comb;
  wire [20:0] p2_smul_72524_comb;
  wire [20:0] p2_smul_72525_comb;
  wire [20:0] p2_smul_72526_comb;
  wire [20:0] p2_smul_72527_comb;
  wire [19:0] p2_smul_29488_NarrowedMult__comb;
  wire [19:0] p2_smul_29494_NarrowedMult__comb;
  wire [20:0] p2_smul_72534_comb;
  wire [20:0] p2_smul_72535_comb;
  wire [20:0] p2_smul_72536_comb;
  wire [20:0] p2_smul_72537_comb;
  wire [19:0] p2_smul_29504_NarrowedMult__comb;
  wire [19:0] p2_smul_29510_NarrowedMult__comb;
  wire [20:0] p2_smul_72544_comb;
  wire [20:0] p2_smul_72545_comb;
  wire [20:0] p2_smul_72546_comb;
  wire [20:0] p2_smul_72547_comb;
  wire [19:0] p2_smul_29520_NarrowedMult__comb;
  wire [13:0] p2_add_73615_comb;
  wire [13:0] p2_add_73616_comb;
  wire [13:0] p2_add_73617_comb;
  wire [13:0] p2_add_73618_comb;
  wire [13:0] p2_add_73619_comb;
  wire [13:0] p2_add_73620_comb;
  wire [13:0] p2_add_73621_comb;
  wire [13:0] p2_add_73622_comb;
  wire [13:0] p2_add_73623_comb;
  wire [13:0] p2_add_73624_comb;
  wire [13:0] p2_add_73625_comb;
  wire [13:0] p2_add_73626_comb;
  wire [13:0] p2_add_73627_comb;
  wire [13:0] p2_add_73628_comb;
  wire [13:0] p2_add_73629_comb;
  wire [13:0] p2_add_73630_comb;
  wire [13:0] p2_add_73631_comb;
  wire [13:0] p2_add_73632_comb;
  wire [13:0] p2_add_73633_comb;
  wire [13:0] p2_add_73634_comb;
  wire [13:0] p2_add_73635_comb;
  wire [13:0] p2_add_73636_comb;
  wire [13:0] p2_add_73637_comb;
  wire [13:0] p2_add_73638_comb;
  wire [13:0] p2_add_73639_comb;
  wire [13:0] p2_add_73640_comb;
  wire [13:0] p2_add_73641_comb;
  wire [13:0] p2_add_73642_comb;
  wire [13:0] p2_add_73643_comb;
  wire [13:0] p2_add_73644_comb;
  wire [13:0] p2_add_73645_comb;
  wire [13:0] p2_add_73646_comb;
  wire [13:0] p2_add_73647_comb;
  wire [13:0] p2_add_73648_comb;
  wire [13:0] p2_add_73649_comb;
  wire [13:0] p2_add_73650_comb;
  wire [13:0] p2_add_73651_comb;
  wire [13:0] p2_add_73652_comb;
  wire [13:0] p2_add_73653_comb;
  wire [13:0] p2_add_73654_comb;
  wire [13:0] p2_add_73655_comb;
  wire [13:0] p2_add_73656_comb;
  wire [13:0] p2_add_73657_comb;
  wire [13:0] p2_add_73658_comb;
  wire [13:0] p2_add_73659_comb;
  wire [13:0] p2_add_73660_comb;
  wire [13:0] p2_add_73661_comb;
  wire [13:0] p2_add_73662_comb;
  wire [13:0] p2_add_73663_comb;
  wire [13:0] p2_add_73664_comb;
  wire [13:0] p2_add_73665_comb;
  wire [13:0] p2_add_73666_comb;
  wire [13:0] p2_add_73667_comb;
  wire [13:0] p2_add_73668_comb;
  wire [13:0] p2_add_73669_comb;
  wire [13:0] p2_add_73670_comb;
  wire [31:0] p2_sum__464_comb;
  wire [31:0] p2_sum__465_comb;
  wire [31:0] p2_sum__466_comb;
  wire [31:0] p2_sum__467_comb;
  wire [31:0] p2_sum__408_comb;
  wire [31:0] p2_sum__409_comb;
  wire [31:0] p2_sum__410_comb;
  wire [31:0] p2_sum__411_comb;
  wire [31:0] p2_sum__352_comb;
  wire [31:0] p2_sum__353_comb;
  wire [31:0] p2_sum__354_comb;
  wire [31:0] p2_sum__355_comb;
  wire [31:0] p2_sum__296_comb;
  wire [31:0] p2_sum__297_comb;
  wire [31:0] p2_sum__298_comb;
  wire [31:0] p2_sum__299_comb;
  wire [31:0] p2_sum__240_comb;
  wire [31:0] p2_sum__241_comb;
  wire [31:0] p2_sum__242_comb;
  wire [31:0] p2_sum__243_comb;
  wire [31:0] p2_sum__184_comb;
  wire [31:0] p2_sum__185_comb;
  wire [31:0] p2_sum__186_comb;
  wire [31:0] p2_sum__187_comb;
  wire [31:0] p2_sum__128_comb;
  wire [31:0] p2_sum__129_comb;
  wire [31:0] p2_sum__130_comb;
  wire [31:0] p2_sum__131_comb;
  wire [31:0] p2_sum__524_comb;
  wire [31:0] p2_sum__525_comb;
  wire [12:0] p2_add_74455_comb;
  wire [12:0] p2_add_74456_comb;
  wire [12:0] p2_add_74457_comb;
  wire [12:0] p2_add_74458_comb;
  wire [11:0] p2_add_72635_comb;
  wire [11:0] p2_add_72636_comb;
  wire [11:0] p2_add_72649_comb;
  wire [11:0] p2_add_72650_comb;
  wire [11:0] p2_add_72663_comb;
  wire [11:0] p2_add_72664_comb;
  wire [11:0] p2_add_72677_comb;
  wire [11:0] p2_add_72678_comb;
  wire [11:0] p2_add_72691_comb;
  wire [11:0] p2_add_72692_comb;
  wire [11:0] p2_add_72705_comb;
  wire [11:0] p2_add_72706_comb;
  wire [11:0] p2_add_72719_comb;
  wire [11:0] p2_add_72720_comb;
  wire [12:0] p2_add_72741_comb;
  wire [12:0] p2_add_72742_comb;
  wire [12:0] p2_add_72747_comb;
  wire [12:0] p2_add_72748_comb;
  wire [12:0] p2_add_72753_comb;
  wire [12:0] p2_add_72754_comb;
  wire [12:0] p2_add_72759_comb;
  wire [12:0] p2_add_72760_comb;
  wire [12:0] p2_add_72765_comb;
  wire [12:0] p2_add_72766_comb;
  wire [12:0] p2_add_72771_comb;
  wire [12:0] p2_add_72772_comb;
  wire [12:0] p2_add_72777_comb;
  wire [12:0] p2_add_72778_comb;
  wire [12:0] p2_add_72783_comb;
  wire [12:0] p2_add_72784_comb;
  wire [12:0] p2_add_72789_comb;
  wire [12:0] p2_add_72790_comb;
  wire [12:0] p2_add_72795_comb;
  wire [12:0] p2_add_72796_comb;
  wire [12:0] p2_add_72801_comb;
  wire [12:0] p2_add_72802_comb;
  wire [12:0] p2_add_72807_comb;
  wire [12:0] p2_add_72808_comb;
  wire [12:0] p2_add_72813_comb;
  wire [12:0] p2_add_72814_comb;
  wire [12:0] p2_add_72819_comb;
  wire [12:0] p2_add_72820_comb;
  wire [11:0] p2_add_72839_comb;
  wire [11:0] p2_add_72848_comb;
  wire [11:0] p2_add_72853_comb;
  wire [11:0] p2_add_72862_comb;
  wire [11:0] p2_add_72867_comb;
  wire [11:0] p2_add_72876_comb;
  wire [11:0] p2_add_72881_comb;
  wire [11:0] p2_add_72890_comb;
  wire [11:0] p2_add_72895_comb;
  wire [11:0] p2_add_72904_comb;
  wire [11:0] p2_add_72909_comb;
  wire [11:0] p2_add_72918_comb;
  wire [11:0] p2_add_72923_comb;
  wire [11:0] p2_add_72932_comb;
  wire [11:0] p2_add_73081_comb;
  wire [11:0] p2_add_73086_comb;
  wire [11:0] p2_add_73095_comb;
  wire [11:0] p2_add_73100_comb;
  wire [11:0] p2_add_73109_comb;
  wire [11:0] p2_add_73114_comb;
  wire [11:0] p2_add_73123_comb;
  wire [11:0] p2_add_73128_comb;
  wire [11:0] p2_add_73137_comb;
  wire [11:0] p2_add_73142_comb;
  wire [11:0] p2_add_73151_comb;
  wire [11:0] p2_add_73156_comb;
  wire [11:0] p2_add_73165_comb;
  wire [11:0] p2_add_73170_comb;
  wire [12:0] p2_add_73187_comb;
  wire [12:0] p2_add_73190_comb;
  wire [12:0] p2_add_73195_comb;
  wire [12:0] p2_add_73198_comb;
  wire [12:0] p2_add_73199_comb;
  wire [12:0] p2_add_73202_comb;
  wire [12:0] p2_add_73207_comb;
  wire [12:0] p2_add_73210_comb;
  wire [12:0] p2_add_73211_comb;
  wire [12:0] p2_add_73214_comb;
  wire [12:0] p2_add_73219_comb;
  wire [12:0] p2_add_73222_comb;
  wire [12:0] p2_add_73223_comb;
  wire [12:0] p2_add_73226_comb;
  wire [12:0] p2_add_73231_comb;
  wire [12:0] p2_add_73234_comb;
  wire [12:0] p2_add_73235_comb;
  wire [12:0] p2_add_73238_comb;
  wire [12:0] p2_add_73243_comb;
  wire [12:0] p2_add_73246_comb;
  wire [12:0] p2_add_73247_comb;
  wire [12:0] p2_add_73250_comb;
  wire [12:0] p2_add_73255_comb;
  wire [12:0] p2_add_73258_comb;
  wire [12:0] p2_add_73259_comb;
  wire [12:0] p2_add_73262_comb;
  wire [12:0] p2_add_73267_comb;
  wire [12:0] p2_add_73270_comb;
  wire [11:0] p2_add_73285_comb;
  wire [11:0] p2_add_73298_comb;
  wire [11:0] p2_add_73299_comb;
  wire [11:0] p2_add_73312_comb;
  wire [11:0] p2_add_73313_comb;
  wire [11:0] p2_add_73326_comb;
  wire [11:0] p2_add_73327_comb;
  wire [11:0] p2_add_73340_comb;
  wire [11:0] p2_add_73341_comb;
  wire [11:0] p2_add_73354_comb;
  wire [11:0] p2_add_73355_comb;
  wire [11:0] p2_add_73368_comb;
  wire [11:0] p2_add_73369_comb;
  wire [11:0] p2_add_73382_comb;
  wire [31:0] p2_sum__468_comb;
  wire [31:0] p2_sum__469_comb;
  wire [31:0] p2_sum__412_comb;
  wire [31:0] p2_sum__413_comb;
  wire [31:0] p2_sum__356_comb;
  wire [31:0] p2_sum__357_comb;
  wire [31:0] p2_sum__300_comb;
  wire [31:0] p2_sum__301_comb;
  wire [31:0] p2_sum__244_comb;
  wire [31:0] p2_sum__245_comb;
  wire [31:0] p2_sum__188_comb;
  wire [31:0] p2_sum__189_comb;
  wire [31:0] p2_sum__132_comb;
  wire [31:0] p2_sum__133_comb;
  wire [12:0] p2_add_74359_comb;
  wire [12:0] p2_add_74360_comb;
  wire [12:0] p2_add_74361_comb;
  wire [12:0] p2_add_74362_comb;
  wire [12:0] p2_add_74391_comb;
  wire [12:0] p2_add_74392_comb;
  wire [12:0] p2_add_74393_comb;
  wire [12:0] p2_add_74394_comb;
  wire [12:0] p2_add_74423_comb;
  wire [12:0] p2_add_74424_comb;
  wire [12:0] p2_add_74425_comb;
  wire [12:0] p2_add_74426_comb;
  wire [12:0] p2_add_74487_comb;
  wire [12:0] p2_add_74488_comb;
  wire [12:0] p2_add_74489_comb;
  wire [12:0] p2_add_74490_comb;
  wire [12:0] p2_add_74519_comb;
  wire [12:0] p2_add_74520_comb;
  wire [12:0] p2_add_74521_comb;
  wire [12:0] p2_add_74522_comb;
  wire [12:0] p2_add_74551_comb;
  wire [12:0] p2_add_74552_comb;
  wire [12:0] p2_add_74553_comb;
  wire [12:0] p2_add_74554_comb;
  wire [31:0] p2_sum__526_comb;
  wire [24:0] p2_sum__1568_comb;
  wire [24:0] p2_sum__1569_comb;
  wire [24:0] p2_sum__1570_comb;
  wire [24:0] p2_sum__1571_comb;
  wire [13:0] p2_add_73423_comb;
  wire [13:0] p2_add_73424_comb;
  wire [13:0] p2_add_73425_comb;
  wire [10:0] p2_bit_slice_73426_comb;
  wire [10:0] p2_bit_slice_73427_comb;
  wire [13:0] p2_add_73428_comb;
  wire [13:0] p2_add_73429_comb;
  wire [13:0] p2_add_73430_comb;
  wire [13:0] p2_add_73431_comb;
  wire [13:0] p2_add_73432_comb;
  wire [13:0] p2_add_73433_comb;
  wire [10:0] p2_bit_slice_73434_comb;
  wire [10:0] p2_bit_slice_73435_comb;
  wire [13:0] p2_add_73436_comb;
  wire [13:0] p2_add_73437_comb;
  wire [13:0] p2_add_73438_comb;
  wire [13:0] p2_add_73439_comb;
  wire [13:0] p2_add_73440_comb;
  wire [13:0] p2_add_73441_comb;
  wire [10:0] p2_bit_slice_73442_comb;
  wire [10:0] p2_bit_slice_73443_comb;
  wire [13:0] p2_add_73444_comb;
  wire [13:0] p2_add_73445_comb;
  wire [13:0] p2_add_73446_comb;
  wire [13:0] p2_add_73447_comb;
  wire [13:0] p2_add_73448_comb;
  wire [13:0] p2_add_73449_comb;
  wire [10:0] p2_bit_slice_73450_comb;
  wire [10:0] p2_bit_slice_73451_comb;
  wire [13:0] p2_add_73452_comb;
  wire [13:0] p2_add_73453_comb;
  wire [13:0] p2_add_73454_comb;
  wire [13:0] p2_add_73455_comb;
  wire [13:0] p2_add_73456_comb;
  wire [13:0] p2_add_73457_comb;
  wire [10:0] p2_bit_slice_73458_comb;
  wire [10:0] p2_bit_slice_73459_comb;
  wire [13:0] p2_add_73460_comb;
  wire [13:0] p2_add_73461_comb;
  wire [13:0] p2_add_73462_comb;
  wire [13:0] p2_add_73463_comb;
  wire [13:0] p2_add_73464_comb;
  wire [13:0] p2_add_73465_comb;
  wire [10:0] p2_bit_slice_73466_comb;
  wire [10:0] p2_bit_slice_73467_comb;
  wire [13:0] p2_add_73468_comb;
  wire [13:0] p2_add_73469_comb;
  wire [13:0] p2_add_73470_comb;
  wire [13:0] p2_add_73471_comb;
  wire [13:0] p2_add_73472_comb;
  wire [13:0] p2_add_73473_comb;
  wire [10:0] p2_bit_slice_73474_comb;
  wire [10:0] p2_bit_slice_73475_comb;
  wire [13:0] p2_add_73476_comb;
  wire [13:0] p2_add_73477_comb;
  wire [13:0] p2_add_73478_comb;
  wire [13:0] p2_add_73487_comb;
  wire [11:0] p2_bit_slice_73488_comb;
  wire [11:0] p2_bit_slice_73489_comb;
  wire [13:0] p2_add_73490_comb;
  wire [13:0] p2_add_73491_comb;
  wire [11:0] p2_bit_slice_73492_comb;
  wire [11:0] p2_bit_slice_73493_comb;
  wire [13:0] p2_add_73494_comb;
  wire [13:0] p2_add_73495_comb;
  wire [11:0] p2_bit_slice_73496_comb;
  wire [11:0] p2_bit_slice_73497_comb;
  wire [13:0] p2_add_73498_comb;
  wire [13:0] p2_add_73499_comb;
  wire [11:0] p2_bit_slice_73500_comb;
  wire [11:0] p2_bit_slice_73501_comb;
  wire [13:0] p2_add_73502_comb;
  wire [13:0] p2_add_73503_comb;
  wire [11:0] p2_bit_slice_73504_comb;
  wire [11:0] p2_bit_slice_73505_comb;
  wire [13:0] p2_add_73506_comb;
  wire [13:0] p2_add_73507_comb;
  wire [11:0] p2_bit_slice_73508_comb;
  wire [11:0] p2_bit_slice_73509_comb;
  wire [13:0] p2_add_73510_comb;
  wire [13:0] p2_add_73511_comb;
  wire [11:0] p2_bit_slice_73512_comb;
  wire [11:0] p2_bit_slice_73513_comb;
  wire [13:0] p2_add_73514_comb;
  wire [13:0] p2_add_73515_comb;
  wire [11:0] p2_bit_slice_73516_comb;
  wire [11:0] p2_bit_slice_73517_comb;
  wire [13:0] p2_add_73518_comb;
  wire [13:0] p2_add_73519_comb;
  wire [11:0] p2_bit_slice_73520_comb;
  wire [11:0] p2_bit_slice_73521_comb;
  wire [13:0] p2_add_73522_comb;
  wire [13:0] p2_add_73523_comb;
  wire [11:0] p2_bit_slice_73524_comb;
  wire [11:0] p2_bit_slice_73525_comb;
  wire [13:0] p2_add_73526_comb;
  wire [13:0] p2_add_73527_comb;
  wire [11:0] p2_bit_slice_73528_comb;
  wire [11:0] p2_bit_slice_73529_comb;
  wire [13:0] p2_add_73530_comb;
  wire [13:0] p2_add_73531_comb;
  wire [11:0] p2_bit_slice_73532_comb;
  wire [11:0] p2_bit_slice_73533_comb;
  wire [13:0] p2_add_73534_comb;
  wire [13:0] p2_add_73535_comb;
  wire [11:0] p2_bit_slice_73536_comb;
  wire [11:0] p2_bit_slice_73537_comb;
  wire [13:0] p2_add_73538_comb;
  wire [13:0] p2_add_73539_comb;
  wire [11:0] p2_bit_slice_73540_comb;
  wire [11:0] p2_bit_slice_73541_comb;
  wire [13:0] p2_add_73542_comb;
  wire [13:0] p2_add_73551_comb;
  wire [10:0] p2_bit_slice_73552_comb;
  wire [13:0] p2_add_73553_comb;
  wire [13:0] p2_add_73554_comb;
  wire [13:0] p2_add_73555_comb;
  wire [13:0] p2_add_73556_comb;
  wire [10:0] p2_bit_slice_73557_comb;
  wire [13:0] p2_add_73558_comb;
  wire [13:0] p2_add_73559_comb;
  wire [10:0] p2_bit_slice_73560_comb;
  wire [13:0] p2_add_73561_comb;
  wire [13:0] p2_add_73562_comb;
  wire [13:0] p2_add_73563_comb;
  wire [13:0] p2_add_73564_comb;
  wire [10:0] p2_bit_slice_73565_comb;
  wire [13:0] p2_add_73566_comb;
  wire [13:0] p2_add_73567_comb;
  wire [10:0] p2_bit_slice_73568_comb;
  wire [13:0] p2_add_73569_comb;
  wire [13:0] p2_add_73570_comb;
  wire [13:0] p2_add_73571_comb;
  wire [13:0] p2_add_73572_comb;
  wire [10:0] p2_bit_slice_73573_comb;
  wire [13:0] p2_add_73574_comb;
  wire [13:0] p2_add_73575_comb;
  wire [10:0] p2_bit_slice_73576_comb;
  wire [13:0] p2_add_73577_comb;
  wire [13:0] p2_add_73578_comb;
  wire [13:0] p2_add_73579_comb;
  wire [13:0] p2_add_73580_comb;
  wire [10:0] p2_bit_slice_73581_comb;
  wire [13:0] p2_add_73582_comb;
  wire [13:0] p2_add_73583_comb;
  wire [10:0] p2_bit_slice_73584_comb;
  wire [13:0] p2_add_73585_comb;
  wire [13:0] p2_add_73586_comb;
  wire [13:0] p2_add_73587_comb;
  wire [13:0] p2_add_73588_comb;
  wire [10:0] p2_bit_slice_73589_comb;
  wire [13:0] p2_add_73590_comb;
  wire [13:0] p2_add_73591_comb;
  wire [10:0] p2_bit_slice_73592_comb;
  wire [13:0] p2_add_73593_comb;
  wire [13:0] p2_add_73594_comb;
  wire [13:0] p2_add_73595_comb;
  wire [13:0] p2_add_73596_comb;
  wire [10:0] p2_bit_slice_73597_comb;
  wire [13:0] p2_add_73598_comb;
  wire [13:0] p2_add_73599_comb;
  wire [10:0] p2_bit_slice_73600_comb;
  wire [13:0] p2_add_73601_comb;
  wire [13:0] p2_add_73602_comb;
  wire [13:0] p2_add_73603_comb;
  wire [13:0] p2_add_73604_comb;
  wire [10:0] p2_bit_slice_73605_comb;
  wire [13:0] p2_add_73606_comb;
  wire [13:0] p2_add_73679_comb;
  wire [13:0] p2_add_73680_comb;
  wire [10:0] p2_bit_slice_73681_comb;
  wire [13:0] p2_add_73682_comb;
  wire [13:0] p2_add_73683_comb;
  wire [10:0] p2_bit_slice_73684_comb;
  wire [13:0] p2_add_73685_comb;
  wire [13:0] p2_add_73686_comb;
  wire [13:0] p2_add_73687_comb;
  wire [13:0] p2_add_73688_comb;
  wire [10:0] p2_bit_slice_73689_comb;
  wire [13:0] p2_add_73690_comb;
  wire [13:0] p2_add_73691_comb;
  wire [10:0] p2_bit_slice_73692_comb;
  wire [13:0] p2_add_73693_comb;
  wire [13:0] p2_add_73694_comb;
  wire [13:0] p2_add_73695_comb;
  wire [13:0] p2_add_73696_comb;
  wire [10:0] p2_bit_slice_73697_comb;
  wire [13:0] p2_add_73698_comb;
  wire [13:0] p2_add_73699_comb;
  wire [10:0] p2_bit_slice_73700_comb;
  wire [13:0] p2_add_73701_comb;
  wire [13:0] p2_add_73702_comb;
  wire [13:0] p2_add_73703_comb;
  wire [13:0] p2_add_73704_comb;
  wire [10:0] p2_bit_slice_73705_comb;
  wire [13:0] p2_add_73706_comb;
  wire [13:0] p2_add_73707_comb;
  wire [10:0] p2_bit_slice_73708_comb;
  wire [13:0] p2_add_73709_comb;
  wire [13:0] p2_add_73710_comb;
  wire [13:0] p2_add_73711_comb;
  wire [13:0] p2_add_73712_comb;
  wire [10:0] p2_bit_slice_73713_comb;
  wire [13:0] p2_add_73714_comb;
  wire [13:0] p2_add_73715_comb;
  wire [10:0] p2_bit_slice_73716_comb;
  wire [13:0] p2_add_73717_comb;
  wire [13:0] p2_add_73718_comb;
  wire [13:0] p2_add_73719_comb;
  wire [13:0] p2_add_73720_comb;
  wire [10:0] p2_bit_slice_73721_comb;
  wire [13:0] p2_add_73722_comb;
  wire [13:0] p2_add_73723_comb;
  wire [10:0] p2_bit_slice_73724_comb;
  wire [13:0] p2_add_73725_comb;
  wire [13:0] p2_add_73726_comb;
  wire [13:0] p2_add_73727_comb;
  wire [13:0] p2_add_73728_comb;
  wire [10:0] p2_bit_slice_73729_comb;
  wire [13:0] p2_add_73730_comb;
  wire [13:0] p2_add_73731_comb;
  wire [10:0] p2_bit_slice_73732_comb;
  wire [13:0] p2_add_73733_comb;
  wire [13:0] p2_add_73734_comb;
  wire [11:0] p2_bit_slice_73743_comb;
  wire [13:0] p2_add_73744_comb;
  wire [11:0] p2_bit_slice_73745_comb;
  wire [13:0] p2_add_73746_comb;
  wire [13:0] p2_add_73747_comb;
  wire [11:0] p2_bit_slice_73748_comb;
  wire [13:0] p2_add_73749_comb;
  wire [11:0] p2_bit_slice_73750_comb;
  wire [11:0] p2_bit_slice_73751_comb;
  wire [13:0] p2_add_73752_comb;
  wire [11:0] p2_bit_slice_73753_comb;
  wire [13:0] p2_add_73754_comb;
  wire [13:0] p2_add_73755_comb;
  wire [11:0] p2_bit_slice_73756_comb;
  wire [13:0] p2_add_73757_comb;
  wire [11:0] p2_bit_slice_73758_comb;
  wire [11:0] p2_bit_slice_73759_comb;
  wire [13:0] p2_add_73760_comb;
  wire [11:0] p2_bit_slice_73761_comb;
  wire [13:0] p2_add_73762_comb;
  wire [13:0] p2_add_73763_comb;
  wire [11:0] p2_bit_slice_73764_comb;
  wire [13:0] p2_add_73765_comb;
  wire [11:0] p2_bit_slice_73766_comb;
  wire [11:0] p2_bit_slice_73767_comb;
  wire [13:0] p2_add_73768_comb;
  wire [11:0] p2_bit_slice_73769_comb;
  wire [13:0] p2_add_73770_comb;
  wire [13:0] p2_add_73771_comb;
  wire [11:0] p2_bit_slice_73772_comb;
  wire [13:0] p2_add_73773_comb;
  wire [11:0] p2_bit_slice_73774_comb;
  wire [11:0] p2_bit_slice_73775_comb;
  wire [13:0] p2_add_73776_comb;
  wire [11:0] p2_bit_slice_73777_comb;
  wire [13:0] p2_add_73778_comb;
  wire [13:0] p2_add_73779_comb;
  wire [11:0] p2_bit_slice_73780_comb;
  wire [13:0] p2_add_73781_comb;
  wire [11:0] p2_bit_slice_73782_comb;
  wire [11:0] p2_bit_slice_73783_comb;
  wire [13:0] p2_add_73784_comb;
  wire [11:0] p2_bit_slice_73785_comb;
  wire [13:0] p2_add_73786_comb;
  wire [13:0] p2_add_73787_comb;
  wire [11:0] p2_bit_slice_73788_comb;
  wire [13:0] p2_add_73789_comb;
  wire [11:0] p2_bit_slice_73790_comb;
  wire [11:0] p2_bit_slice_73791_comb;
  wire [13:0] p2_add_73792_comb;
  wire [11:0] p2_bit_slice_73793_comb;
  wire [13:0] p2_add_73794_comb;
  wire [13:0] p2_add_73795_comb;
  wire [11:0] p2_bit_slice_73796_comb;
  wire [13:0] p2_add_73797_comb;
  wire [11:0] p2_bit_slice_73798_comb;
  wire [10:0] p2_bit_slice_73807_comb;
  wire [13:0] p2_add_73808_comb;
  wire [13:0] p2_add_73809_comb;
  wire [13:0] p2_add_73810_comb;
  wire [13:0] p2_add_73811_comb;
  wire [13:0] p2_add_73812_comb;
  wire [13:0] p2_add_73813_comb;
  wire [10:0] p2_bit_slice_73814_comb;
  wire [10:0] p2_bit_slice_73815_comb;
  wire [13:0] p2_add_73816_comb;
  wire [13:0] p2_add_73817_comb;
  wire [13:0] p2_add_73818_comb;
  wire [13:0] p2_add_73819_comb;
  wire [13:0] p2_add_73820_comb;
  wire [13:0] p2_add_73821_comb;
  wire [10:0] p2_bit_slice_73822_comb;
  wire [10:0] p2_bit_slice_73823_comb;
  wire [13:0] p2_add_73824_comb;
  wire [13:0] p2_add_73825_comb;
  wire [13:0] p2_add_73826_comb;
  wire [13:0] p2_add_73827_comb;
  wire [13:0] p2_add_73828_comb;
  wire [13:0] p2_add_73829_comb;
  wire [10:0] p2_bit_slice_73830_comb;
  wire [10:0] p2_bit_slice_73831_comb;
  wire [13:0] p2_add_73832_comb;
  wire [13:0] p2_add_73833_comb;
  wire [13:0] p2_add_73834_comb;
  wire [13:0] p2_add_73835_comb;
  wire [13:0] p2_add_73836_comb;
  wire [13:0] p2_add_73837_comb;
  wire [10:0] p2_bit_slice_73838_comb;
  wire [10:0] p2_bit_slice_73839_comb;
  wire [13:0] p2_add_73840_comb;
  wire [13:0] p2_add_73841_comb;
  wire [13:0] p2_add_73842_comb;
  wire [13:0] p2_add_73843_comb;
  wire [13:0] p2_add_73844_comb;
  wire [13:0] p2_add_73845_comb;
  wire [10:0] p2_bit_slice_73846_comb;
  wire [10:0] p2_bit_slice_73847_comb;
  wire [13:0] p2_add_73848_comb;
  wire [13:0] p2_add_73849_comb;
  wire [13:0] p2_add_73850_comb;
  wire [13:0] p2_add_73851_comb;
  wire [13:0] p2_add_73852_comb;
  wire [13:0] p2_add_73853_comb;
  wire [10:0] p2_bit_slice_73854_comb;
  wire [10:0] p2_bit_slice_73855_comb;
  wire [13:0] p2_add_73856_comb;
  wire [13:0] p2_add_73857_comb;
  wire [13:0] p2_add_73858_comb;
  wire [13:0] p2_add_73859_comb;
  wire [13:0] p2_add_73860_comb;
  wire [13:0] p2_add_73861_comb;
  wire [10:0] p2_bit_slice_73862_comb;
  wire [12:0] p2_add_74459_comb;
  wire [12:0] p2_add_74460_comb;
  wire [12:0] p2_add_74461_comb;
  wire [12:0] p2_add_74462_comb;
  wire [12:0] p2_add_74463_comb;
  wire [12:0] p2_add_74464_comb;
  wire [12:0] p2_add_74465_comb;
  wire [12:0] p2_add_74466_comb;
  wire [12:0] p2_add_74467_comb;
  wire [12:0] p2_add_74468_comb;
  wire [12:0] p2_add_74469_comb;
  wire [12:0] p2_add_74470_comb;
  wire [12:0] p2_add_74471_comb;
  wire [12:0] p2_add_74472_comb;
  wire [12:0] p2_add_74473_comb;
  wire [12:0] p2_add_74474_comb;
  wire [12:0] p2_add_74475_comb;
  wire [12:0] p2_add_74476_comb;
  wire [12:0] p2_add_74477_comb;
  wire [12:0] p2_add_74478_comb;
  wire [12:0] p2_add_74479_comb;
  wire [12:0] p2_add_74480_comb;
  wire [12:0] p2_add_74481_comb;
  wire [12:0] p2_add_74482_comb;
  wire [12:0] p2_add_74483_comb;
  wire [12:0] p2_add_74484_comb;
  wire [12:0] p2_add_74485_comb;
  wire [12:0] p2_add_74486_comb;
  wire [31:0] p2_sum__470_comb;
  wire [31:0] p2_sum__414_comb;
  wire [31:0] p2_sum__358_comb;
  wire [31:0] p2_sum__302_comb;
  wire [31:0] p2_sum__246_comb;
  wire [31:0] p2_sum__190_comb;
  wire [31:0] p2_sum__134_comb;
  wire [24:0] p2_sum__1580_comb;
  wire [24:0] p2_sum__1581_comb;
  wire [24:0] p2_sum__1582_comb;
  wire [24:0] p2_sum__1583_comb;
  wire [24:0] p2_sum__1576_comb;
  wire [24:0] p2_sum__1577_comb;
  wire [24:0] p2_sum__1578_comb;
  wire [24:0] p2_sum__1579_comb;
  wire [24:0] p2_sum__1572_comb;
  wire [24:0] p2_sum__1573_comb;
  wire [24:0] p2_sum__1574_comb;
  wire [24:0] p2_sum__1575_comb;
  wire [24:0] p2_sum__1564_comb;
  wire [24:0] p2_sum__1565_comb;
  wire [24:0] p2_sum__1566_comb;
  wire [24:0] p2_sum__1567_comb;
  wire [24:0] p2_sum__1560_comb;
  wire [24:0] p2_sum__1561_comb;
  wire [24:0] p2_sum__1562_comb;
  wire [24:0] p2_sum__1563_comb;
  wire [24:0] p2_sum__1556_comb;
  wire [24:0] p2_sum__1557_comb;
  wire [24:0] p2_sum__1558_comb;
  wire [24:0] p2_sum__1559_comb;
  wire [31:0] p2_umul_74655_comb;
  wire [24:0] p2_sum__1240_comb;
  wire [24:0] p2_sum__1241_comb;
  wire [24:0] p2_sum__1540_comb;
  wire [24:0] p2_sum__1541_comb;
  wire [24:0] p2_sum__1542_comb;
  wire [24:0] p2_sum__1543_comb;
  wire [24:0] p2_sum__1512_comb;
  wire [24:0] p2_sum__1513_comb;
  wire [24:0] p2_sum__1514_comb;
  wire [24:0] p2_sum__1515_comb;
  wire [24:0] p2_sum__1484_comb;
  wire [24:0] p2_sum__1485_comb;
  wire [24:0] p2_sum__1486_comb;
  wire [24:0] p2_sum__1487_comb;
  wire [24:0] p2_sum__1456_comb;
  wire [24:0] p2_sum__1457_comb;
  wire [24:0] p2_sum__1458_comb;
  wire [24:0] p2_sum__1459_comb;
  wire [24:0] p2_sum__1428_comb;
  wire [24:0] p2_sum__1429_comb;
  wire [24:0] p2_sum__1430_comb;
  wire [24:0] p2_sum__1431_comb;
  wire [24:0] p2_sum__1400_comb;
  wire [24:0] p2_sum__1401_comb;
  wire [24:0] p2_sum__1402_comb;
  wire [24:0] p2_sum__1403_comb;
  wire [24:0] p2_sum__1372_comb;
  wire [24:0] p2_sum__1373_comb;
  wire [24:0] p2_sum__1374_comb;
  wire [24:0] p2_sum__1375_comb;
  wire [31:0] p2_umul_74656_comb;
  wire [31:0] p2_umul_74657_comb;
  wire [31:0] p2_umul_74658_comb;
  wire [31:0] p2_umul_74659_comb;
  wire [31:0] p2_umul_74660_comb;
  wire [31:0] p2_umul_74661_comb;
  wire [31:0] p2_umul_74662_comb;
  wire [24:0] p2_sum__1246_comb;
  wire [24:0] p2_sum__1247_comb;
  wire [24:0] p2_sum__1244_comb;
  wire [24:0] p2_sum__1245_comb;
  wire [24:0] p2_sum__1242_comb;
  wire [24:0] p2_sum__1243_comb;
  wire [24:0] p2_sum__1238_comb;
  wire [24:0] p2_sum__1239_comb;
  wire [24:0] p2_sum__1236_comb;
  wire [24:0] p2_sum__1237_comb;
  wire [24:0] p2_sum__1234_comb;
  wire [24:0] p2_sum__1235_comb;
  wire [24:0] p2_sum__1076_comb;
  wire [12:0] p2_add_74363_comb;
  wire [12:0] p2_add_74364_comb;
  wire [12:0] p2_add_74365_comb;
  wire [12:0] p2_add_74366_comb;
  wire [12:0] p2_add_74367_comb;
  wire [12:0] p2_add_74368_comb;
  wire [12:0] p2_add_74369_comb;
  wire [12:0] p2_add_74370_comb;
  wire [12:0] p2_add_74371_comb;
  wire [12:0] p2_add_74372_comb;
  wire [12:0] p2_add_74373_comb;
  wire [12:0] p2_add_74374_comb;
  wire [12:0] p2_add_74375_comb;
  wire [12:0] p2_add_74376_comb;
  wire [12:0] p2_add_74377_comb;
  wire [12:0] p2_add_74378_comb;
  wire [12:0] p2_add_74379_comb;
  wire [12:0] p2_add_74380_comb;
  wire [12:0] p2_add_74381_comb;
  wire [12:0] p2_add_74382_comb;
  wire [12:0] p2_add_74383_comb;
  wire [12:0] p2_add_74384_comb;
  wire [12:0] p2_add_74385_comb;
  wire [12:0] p2_add_74386_comb;
  wire [12:0] p2_add_74387_comb;
  wire [12:0] p2_add_74388_comb;
  wire [12:0] p2_add_74389_comb;
  wire [12:0] p2_add_74390_comb;
  wire [12:0] p2_add_74395_comb;
  wire [12:0] p2_add_74396_comb;
  wire [12:0] p2_add_74397_comb;
  wire [12:0] p2_add_74398_comb;
  wire [12:0] p2_add_74399_comb;
  wire [12:0] p2_add_74400_comb;
  wire [12:0] p2_add_74401_comb;
  wire [12:0] p2_add_74402_comb;
  wire [12:0] p2_add_74403_comb;
  wire [12:0] p2_add_74404_comb;
  wire [12:0] p2_add_74405_comb;
  wire [12:0] p2_add_74406_comb;
  wire [12:0] p2_add_74407_comb;
  wire [12:0] p2_add_74408_comb;
  wire [12:0] p2_add_74409_comb;
  wire [12:0] p2_add_74410_comb;
  wire [12:0] p2_add_74411_comb;
  wire [12:0] p2_add_74412_comb;
  wire [12:0] p2_add_74413_comb;
  wire [12:0] p2_add_74414_comb;
  wire [12:0] p2_add_74415_comb;
  wire [12:0] p2_add_74416_comb;
  wire [12:0] p2_add_74417_comb;
  wire [12:0] p2_add_74418_comb;
  wire [12:0] p2_add_74419_comb;
  wire [12:0] p2_add_74420_comb;
  wire [12:0] p2_add_74421_comb;
  wire [12:0] p2_add_74422_comb;
  wire [12:0] p2_add_74427_comb;
  wire [12:0] p2_add_74428_comb;
  wire [12:0] p2_add_74429_comb;
  wire [12:0] p2_add_74430_comb;
  wire [12:0] p2_add_74431_comb;
  wire [12:0] p2_add_74432_comb;
  wire [12:0] p2_add_74433_comb;
  wire [12:0] p2_add_74434_comb;
  wire [12:0] p2_add_74435_comb;
  wire [12:0] p2_add_74436_comb;
  wire [12:0] p2_add_74437_comb;
  wire [12:0] p2_add_74438_comb;
  wire [12:0] p2_add_74439_comb;
  wire [12:0] p2_add_74440_comb;
  wire [12:0] p2_add_74441_comb;
  wire [12:0] p2_add_74442_comb;
  wire [12:0] p2_add_74443_comb;
  wire [12:0] p2_add_74444_comb;
  wire [12:0] p2_add_74445_comb;
  wire [12:0] p2_add_74446_comb;
  wire [12:0] p2_add_74447_comb;
  wire [12:0] p2_add_74448_comb;
  wire [12:0] p2_add_74449_comb;
  wire [12:0] p2_add_74450_comb;
  wire [12:0] p2_add_74451_comb;
  wire [12:0] p2_add_74452_comb;
  wire [12:0] p2_add_74453_comb;
  wire [12:0] p2_add_74454_comb;
  wire [12:0] p2_add_74491_comb;
  wire [12:0] p2_add_74492_comb;
  wire [12:0] p2_add_74493_comb;
  wire [12:0] p2_add_74494_comb;
  wire [12:0] p2_add_74495_comb;
  wire [12:0] p2_add_74496_comb;
  wire [12:0] p2_add_74497_comb;
  wire [12:0] p2_add_74498_comb;
  wire [12:0] p2_add_74499_comb;
  wire [12:0] p2_add_74500_comb;
  wire [12:0] p2_add_74501_comb;
  wire [12:0] p2_add_74502_comb;
  wire [12:0] p2_add_74503_comb;
  wire [12:0] p2_add_74504_comb;
  wire [12:0] p2_add_74505_comb;
  wire [12:0] p2_add_74506_comb;
  wire [12:0] p2_add_74507_comb;
  wire [12:0] p2_add_74508_comb;
  wire [12:0] p2_add_74509_comb;
  wire [12:0] p2_add_74510_comb;
  wire [12:0] p2_add_74511_comb;
  wire [12:0] p2_add_74512_comb;
  wire [12:0] p2_add_74513_comb;
  wire [12:0] p2_add_74514_comb;
  wire [12:0] p2_add_74515_comb;
  wire [12:0] p2_add_74516_comb;
  wire [12:0] p2_add_74517_comb;
  wire [12:0] p2_add_74518_comb;
  wire [12:0] p2_add_74523_comb;
  wire [12:0] p2_add_74524_comb;
  wire [12:0] p2_add_74525_comb;
  wire [12:0] p2_add_74526_comb;
  wire [12:0] p2_add_74527_comb;
  wire [12:0] p2_add_74528_comb;
  wire [12:0] p2_add_74529_comb;
  wire [12:0] p2_add_74530_comb;
  wire [12:0] p2_add_74531_comb;
  wire [12:0] p2_add_74532_comb;
  wire [12:0] p2_add_74533_comb;
  wire [12:0] p2_add_74534_comb;
  wire [12:0] p2_add_74535_comb;
  wire [12:0] p2_add_74536_comb;
  wire [12:0] p2_add_74537_comb;
  wire [12:0] p2_add_74538_comb;
  wire [12:0] p2_add_74539_comb;
  wire [12:0] p2_add_74540_comb;
  wire [12:0] p2_add_74541_comb;
  wire [12:0] p2_add_74542_comb;
  wire [12:0] p2_add_74543_comb;
  wire [12:0] p2_add_74544_comb;
  wire [12:0] p2_add_74545_comb;
  wire [12:0] p2_add_74546_comb;
  wire [12:0] p2_add_74547_comb;
  wire [12:0] p2_add_74548_comb;
  wire [12:0] p2_add_74549_comb;
  wire [12:0] p2_add_74550_comb;
  wire [12:0] p2_add_74555_comb;
  wire [12:0] p2_add_74556_comb;
  wire [12:0] p2_add_74557_comb;
  wire [12:0] p2_add_74558_comb;
  wire [12:0] p2_add_74559_comb;
  wire [12:0] p2_add_74560_comb;
  wire [12:0] p2_add_74561_comb;
  wire [12:0] p2_add_74562_comb;
  wire [12:0] p2_add_74563_comb;
  wire [12:0] p2_add_74564_comb;
  wire [12:0] p2_add_74565_comb;
  wire [12:0] p2_add_74566_comb;
  wire [12:0] p2_add_74567_comb;
  wire [12:0] p2_add_74568_comb;
  wire [12:0] p2_add_74569_comb;
  wire [12:0] p2_add_74570_comb;
  wire [12:0] p2_add_74571_comb;
  wire [12:0] p2_add_74572_comb;
  wire [12:0] p2_add_74573_comb;
  wire [12:0] p2_add_74574_comb;
  wire [12:0] p2_add_74575_comb;
  wire [12:0] p2_add_74576_comb;
  wire [12:0] p2_add_74577_comb;
  wire [12:0] p2_add_74578_comb;
  wire [12:0] p2_add_74579_comb;
  wire [12:0] p2_add_74580_comb;
  wire [12:0] p2_add_74581_comb;
  wire [12:0] p2_add_74582_comb;
  wire [24:0] p2_sum__1226_comb;
  wire [24:0] p2_sum__1227_comb;
  wire [24:0] p2_sum__1212_comb;
  wire [24:0] p2_sum__1213_comb;
  wire [24:0] p2_sum__1198_comb;
  wire [24:0] p2_sum__1199_comb;
  wire [24:0] p2_sum__1184_comb;
  wire [24:0] p2_sum__1185_comb;
  wire [24:0] p2_sum__1170_comb;
  wire [24:0] p2_sum__1171_comb;
  wire [24:0] p2_sum__1156_comb;
  wire [24:0] p2_sum__1157_comb;
  wire [24:0] p2_sum__1142_comb;
  wire [24:0] p2_sum__1143_comb;
  wire [24:0] p2_bit_slice_74693_comb;
  wire [24:0] p2_bit_slice_74694_comb;
  wire [24:0] p2_bit_slice_74695_comb;
  wire [24:0] p2_bit_slice_74696_comb;
  wire [24:0] p2_bit_slice_74697_comb;
  wire [24:0] p2_bit_slice_74698_comb;
  wire [24:0] p2_bit_slice_74699_comb;
  wire [24:0] p2_sum__1079_comb;
  wire [24:0] p2_sum__1078_comb;
  wire [24:0] p2_sum__1077_comb;
  wire [24:0] p2_sum__1075_comb;
  wire [24:0] p2_sum__1074_comb;
  wire [24:0] p2_sum__1073_comb;
  wire [24:0] p2_add_74708_comb;
  wire [24:0] p2_add_74709_comb;
  assign p2_clipped__56_comb = p1_slt_70639 ? 12'h800 : (p1_sgt_70616 ? 12'h7ff : p1_bit_slice_70617);
  assign p2_clipped__72_comb = p1_slt_70640 ? 12'h800 : (p1_sgt_70619 ? 12'h7ff : p1_bit_slice_70620);
  assign p2_clipped__24_comb = p1_slt_70641 ? 12'h800 : (p1_sgt_70622 ? 12'h7ff : p1_bit_slice_70623);
  assign p2_clipped__40_comb = p1_slt_70642 ? 12'h800 : (p1_sgt_70625 ? 12'h7ff : p1_bit_slice_70626);
  assign p2_clipped__88_comb = p1_slt_70643 ? 12'h800 : (p1_sgt_70628 ? 12'h7ff : p1_bit_slice_70629);
  assign p2_clipped__104_comb = p1_slt_70644 ? 12'h800 : (p1_sgt_70631 ? 12'h7ff : p1_bit_slice_70632);
  assign p2_clipped__8_comb = p1_slt_70645 ? 12'h800 : (p1_sgt_70634 ? 12'h7ff : p1_bit_slice_70635);
  assign p2_clipped__120_comb = p1_slt_70646 ? 12'h800 : (p1_sgt_70637 ? 12'h7ff : p1_bit_slice_70638);
  assign p2_smul_28634_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__56_comb, 6'h19);
  assign p2_smul_28636_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__72_comb, 6'h27);
  assign p2_smul_28758_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__24_comb, 7'h31);
  assign p2_smul_28760_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__40_comb, 7'h4f);
  assign p2_smul_28766_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__88_comb, 7'h4f);
  assign p2_smul_28768_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__104_comb, 7'h31);
  assign p2_smul_28886_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__24_comb, 6'h27);
  assign p2_smul_28896_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__104_comb, 6'h19);
  assign p2_smul_29144_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__40_comb, 6'h27);
  assign p2_smul_29150_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__88_comb, 6'h27);
  assign p2_smul_29268_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__8_comb, 7'h31);
  assign p2_smul_29272_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__40_comb, 7'h31);
  assign p2_smul_29278_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__88_comb, 7'h31);
  assign p2_smul_29282_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__120_comb, 7'h31);
  assign p2_smul_29396_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__8_comb, 6'h19);
  assign p2_smul_29410_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__120_comb, 6'h19);
  assign p2_smul_72231_comb = smul21b_12b_x_9b(p2_clipped__8_comb, 9'h0b5);
  assign p2_smul_72232_comb = smul21b_12b_x_9b(p2_clipped__24_comb, 9'h14b);
  assign p2_smul_72233_comb = smul21b_12b_x_9b(p2_clipped__40_comb, 9'h14b);
  assign p2_smul_72234_comb = smul21b_12b_x_9b(p2_clipped__56_comb, 9'h0b5);
  assign p2_smul_72235_comb = smul21b_12b_x_9b(p2_clipped__72_comb, 9'h0b5);
  assign p2_smul_72236_comb = smul21b_12b_x_9b(p2_clipped__88_comb, 9'h14b);
  assign p2_smul_72237_comb = smul21b_12b_x_9b(p2_clipped__104_comb, 9'h14b);
  assign p2_smul_72238_comb = smul21b_12b_x_9b(p2_clipped__120_comb, 9'h0b5);
  assign p2_clipped__9_comb = $signed(p1_add_70585[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70585[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70585[12:1]);
  assign p2_clipped__25_comb = $signed(p1_add_70555[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70555[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70555[12:1]);
  assign p2_clipped__41_comb = $signed(p1_add_70556[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70556[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70556[12:1]);
  assign p2_clipped__57_comb = $signed(p1_add_70537[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70537[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70537[12:1]);
  assign p2_clipped__73_comb = $signed(p1_add_70538[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70538[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70538[12:1]);
  assign p2_clipped__89_comb = $signed(p1_add_70557[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70557[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70557[12:1]);
  assign p2_clipped__105_comb = $signed(p1_add_70558[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70558[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70558[12:1]);
  assign p2_clipped__121_comb = $signed(p1_add_70586[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70586[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70586[12:1]);
  assign p2_clipped__10_comb = $signed(p1_add_70587[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70587[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70587[12:1]);
  assign p2_clipped__26_comb = $signed(p1_add_70559[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70559[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70559[12:1]);
  assign p2_clipped__42_comb = $signed(p1_add_70560[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70560[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70560[12:1]);
  assign p2_clipped__58_comb = $signed(p1_add_70539[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70539[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70539[12:1]);
  assign p2_clipped__74_comb = $signed(p1_add_70540[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70540[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70540[12:1]);
  assign p2_clipped__90_comb = $signed(p1_add_70561[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70561[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70561[12:1]);
  assign p2_clipped__106_comb = $signed(p1_add_70562[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70562[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70562[12:1]);
  assign p2_clipped__122_comb = $signed(p1_add_70588[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70588[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70588[12:1]);
  assign p2_clipped__11_comb = $signed(p1_add_70589[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70589[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70589[12:1]);
  assign p2_clipped__27_comb = $signed(p1_add_70563[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70563[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70563[12:1]);
  assign p2_clipped__43_comb = $signed(p1_add_70564[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70564[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70564[12:1]);
  assign p2_clipped__59_comb = $signed(p1_add_70541[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70541[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70541[12:1]);
  assign p2_clipped__75_comb = $signed(p1_add_70542[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70542[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70542[12:1]);
  assign p2_clipped__91_comb = $signed(p1_add_70565[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70565[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70565[12:1]);
  assign p2_clipped__107_comb = $signed(p1_add_70566[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70566[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70566[12:1]);
  assign p2_clipped__123_comb = $signed(p1_add_70590[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70590[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70590[12:1]);
  assign p2_clipped__12_comb = $signed(p1_add_70591[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70591[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70591[12:1]);
  assign p2_clipped__28_comb = $signed(p1_add_70567[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70567[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70567[12:1]);
  assign p2_clipped__44_comb = $signed(p1_add_70568[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70568[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70568[12:1]);
  assign p2_clipped__60_comb = $signed(p1_add_70543[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70543[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70543[12:1]);
  assign p2_clipped__76_comb = $signed(p1_add_70544[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70544[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70544[12:1]);
  assign p2_clipped__92_comb = $signed(p1_add_70569[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70569[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70569[12:1]);
  assign p2_clipped__108_comb = $signed(p1_add_70570[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70570[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70570[12:1]);
  assign p2_clipped__124_comb = $signed(p1_add_70592[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70592[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70592[12:1]);
  assign p2_clipped__13_comb = $signed(p1_add_70593[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70593[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70593[12:1]);
  assign p2_clipped__29_comb = $signed(p1_add_70571[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70571[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70571[12:1]);
  assign p2_clipped__45_comb = $signed(p1_add_70572[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70572[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70572[12:1]);
  assign p2_clipped__61_comb = $signed(p1_add_70545[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70545[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70545[12:1]);
  assign p2_clipped__77_comb = $signed(p1_add_70546[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70546[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70546[12:1]);
  assign p2_clipped__93_comb = $signed(p1_add_70573[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70573[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70573[12:1]);
  assign p2_clipped__109_comb = $signed(p1_add_70574[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70574[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70574[12:1]);
  assign p2_clipped__125_comb = $signed(p1_add_70594[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70594[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70594[12:1]);
  assign p2_clipped__14_comb = $signed(p1_add_70595[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70595[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70595[12:1]);
  assign p2_clipped__30_comb = $signed(p1_add_70575[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70575[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70575[12:1]);
  assign p2_clipped__46_comb = $signed(p1_add_70576[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70576[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70576[12:1]);
  assign p2_clipped__62_comb = $signed(p1_add_70547[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70547[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70547[12:1]);
  assign p2_clipped__78_comb = $signed(p1_add_70548[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70548[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70548[12:1]);
  assign p2_clipped__94_comb = $signed(p1_add_70577[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70577[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70577[12:1]);
  assign p2_clipped__110_comb = $signed(p1_add_70578[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70578[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70578[12:1]);
  assign p2_clipped__126_comb = $signed(p1_add_70596[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70596[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70596[12:1]);
  assign p2_clipped__15_comb = $signed(p1_add_70597[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70597[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70597[12:1]);
  assign p2_clipped__31_comb = $signed(p1_add_70579[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70579[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70579[12:1]);
  assign p2_clipped__47_comb = $signed(p1_add_70580[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70580[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70580[12:1]);
  assign p2_clipped__63_comb = $signed(p1_add_70549[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70549[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70549[12:1]);
  assign p2_clipped__79_comb = $signed(p1_add_70550[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70550[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70550[12:1]);
  assign p2_clipped__95_comb = $signed(p1_add_70581[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70581[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70581[12:1]);
  assign p2_clipped__111_comb = $signed(p1_add_70582[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70582[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70582[12:1]);
  assign p2_clipped__127_comb = $signed(p1_add_70598[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p1_add_70598[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p1_add_70598[12:1]);
  assign p2_smul_71975_comb = smul21b_12b_x_9b(p2_clipped__8_comb, 9'h0fb);
  assign p2_smul_71976_comb = smul21b_12b_x_9b(p2_clipped__24_comb, 9'h0d5);
  assign p2_smul_28632_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__40_comb, 8'h47);
  assign p2_smul_28638_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__88_comb, 8'hb9);
  assign p2_smul_71983_comb = smul21b_12b_x_9b(p2_clipped__104_comb, 9'h12b);
  assign p2_smul_71984_comb = smul21b_12b_x_9b(p2_clipped__120_comb, 9'h105);
  assign p2_smul_28756_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__8_comb, 7'h3b);
  assign p2_smul_28762_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__56_comb, 7'h45);
  assign p2_smul_28764_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__72_comb, 7'h45);
  assign p2_smul_28770_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__120_comb, 7'h3b);
  assign p2_smul_72151_comb = smul21b_12b_x_9b(p2_clipped__8_comb, 9'h0d5);
  assign p2_smul_72154_comb = smul21b_12b_x_9b(p2_clipped__40_comb, 9'h105);
  assign p2_smul_28890_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__56_comb, 8'hb9);
  assign p2_smul_28892_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__72_comb, 8'h47);
  assign p2_smul_72157_comb = smul21b_12b_x_9b(p2_clipped__88_comb, 9'h0fb);
  assign p2_smul_72160_comb = smul21b_12b_x_9b(p2_clipped__120_comb, 9'h12b);
  assign p2_smul_29140_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__8_comb, 8'h47);
  assign p2_smul_72296_comb = smul21b_12b_x_9b(p2_clipped__24_comb, 9'h105);
  assign p2_smul_72299_comb = smul21b_12b_x_9b(p2_clipped__56_comb, 9'h0d5);
  assign p2_smul_72300_comb = smul21b_12b_x_9b(p2_clipped__72_comb, 9'h0d5);
  assign p2_smul_72303_comb = smul21b_12b_x_9b(p2_clipped__104_comb, 9'h105);
  assign p2_smul_29154_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__120_comb, 8'h47);
  assign p2_smul_29270_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__24_comb, 7'h45);
  assign p2_smul_29274_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__56_comb, 7'h3b);
  assign p2_smul_29276_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__72_comb, 7'h3b);
  assign p2_smul_29280_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__104_comb, 7'h45);
  assign p2_smul_29398_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__24_comb, 8'hb9);
  assign p2_smul_72474_comb = smul21b_12b_x_9b(p2_clipped__40_comb, 9'h0d5);
  assign p2_smul_72475_comb = smul21b_12b_x_9b(p2_clipped__56_comb, 9'h105);
  assign p2_smul_72476_comb = smul21b_12b_x_9b(p2_clipped__72_comb, 9'h105);
  assign p2_smul_72477_comb = smul21b_12b_x_9b(p2_clipped__88_comb, 9'h0d5);
  assign p2_smul_29408_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__104_comb, 8'hb9);
  assign p2_smul_72239_comb = smul21b_12b_x_9b(p2_clipped__9_comb, 9'h0b5);
  assign p2_smul_72240_comb = smul21b_12b_x_9b(p2_clipped__25_comb, 9'h14b);
  assign p2_smul_72241_comb = smul21b_12b_x_9b(p2_clipped__41_comb, 9'h14b);
  assign p2_smul_72242_comb = smul21b_12b_x_9b(p2_clipped__57_comb, 9'h0b5);
  assign p2_smul_72243_comb = smul21b_12b_x_9b(p2_clipped__73_comb, 9'h0b5);
  assign p2_smul_72244_comb = smul21b_12b_x_9b(p2_clipped__89_comb, 9'h14b);
  assign p2_smul_72245_comb = smul21b_12b_x_9b(p2_clipped__105_comb, 9'h14b);
  assign p2_smul_72246_comb = smul21b_12b_x_9b(p2_clipped__121_comb, 9'h0b5);
  assign p2_smul_72247_comb = smul21b_12b_x_9b(p2_clipped__10_comb, 9'h0b5);
  assign p2_smul_72248_comb = smul21b_12b_x_9b(p2_clipped__26_comb, 9'h14b);
  assign p2_smul_72249_comb = smul21b_12b_x_9b(p2_clipped__42_comb, 9'h14b);
  assign p2_smul_72250_comb = smul21b_12b_x_9b(p2_clipped__58_comb, 9'h0b5);
  assign p2_smul_72251_comb = smul21b_12b_x_9b(p2_clipped__74_comb, 9'h0b5);
  assign p2_smul_72252_comb = smul21b_12b_x_9b(p2_clipped__90_comb, 9'h14b);
  assign p2_smul_72253_comb = smul21b_12b_x_9b(p2_clipped__106_comb, 9'h14b);
  assign p2_smul_72254_comb = smul21b_12b_x_9b(p2_clipped__122_comb, 9'h0b5);
  assign p2_smul_72255_comb = smul21b_12b_x_9b(p2_clipped__11_comb, 9'h0b5);
  assign p2_smul_72256_comb = smul21b_12b_x_9b(p2_clipped__27_comb, 9'h14b);
  assign p2_smul_72257_comb = smul21b_12b_x_9b(p2_clipped__43_comb, 9'h14b);
  assign p2_smul_72258_comb = smul21b_12b_x_9b(p2_clipped__59_comb, 9'h0b5);
  assign p2_smul_72259_comb = smul21b_12b_x_9b(p2_clipped__75_comb, 9'h0b5);
  assign p2_smul_72260_comb = smul21b_12b_x_9b(p2_clipped__91_comb, 9'h14b);
  assign p2_smul_72261_comb = smul21b_12b_x_9b(p2_clipped__107_comb, 9'h14b);
  assign p2_smul_72262_comb = smul21b_12b_x_9b(p2_clipped__123_comb, 9'h0b5);
  assign p2_smul_72263_comb = smul21b_12b_x_9b(p2_clipped__12_comb, 9'h0b5);
  assign p2_smul_72264_comb = smul21b_12b_x_9b(p2_clipped__28_comb, 9'h14b);
  assign p2_smul_72265_comb = smul21b_12b_x_9b(p2_clipped__44_comb, 9'h14b);
  assign p2_smul_72266_comb = smul21b_12b_x_9b(p2_clipped__60_comb, 9'h0b5);
  assign p2_smul_72267_comb = smul21b_12b_x_9b(p2_clipped__76_comb, 9'h0b5);
  assign p2_smul_72268_comb = smul21b_12b_x_9b(p2_clipped__92_comb, 9'h14b);
  assign p2_smul_72269_comb = smul21b_12b_x_9b(p2_clipped__108_comb, 9'h14b);
  assign p2_smul_72270_comb = smul21b_12b_x_9b(p2_clipped__124_comb, 9'h0b5);
  assign p2_smul_72271_comb = smul21b_12b_x_9b(p2_clipped__13_comb, 9'h0b5);
  assign p2_smul_72272_comb = smul21b_12b_x_9b(p2_clipped__29_comb, 9'h14b);
  assign p2_smul_72273_comb = smul21b_12b_x_9b(p2_clipped__45_comb, 9'h14b);
  assign p2_smul_72274_comb = smul21b_12b_x_9b(p2_clipped__61_comb, 9'h0b5);
  assign p2_smul_72275_comb = smul21b_12b_x_9b(p2_clipped__77_comb, 9'h0b5);
  assign p2_smul_72276_comb = smul21b_12b_x_9b(p2_clipped__93_comb, 9'h14b);
  assign p2_smul_72277_comb = smul21b_12b_x_9b(p2_clipped__109_comb, 9'h14b);
  assign p2_smul_72278_comb = smul21b_12b_x_9b(p2_clipped__125_comb, 9'h0b5);
  assign p2_smul_72279_comb = smul21b_12b_x_9b(p2_clipped__14_comb, 9'h0b5);
  assign p2_smul_72280_comb = smul21b_12b_x_9b(p2_clipped__30_comb, 9'h14b);
  assign p2_smul_72281_comb = smul21b_12b_x_9b(p2_clipped__46_comb, 9'h14b);
  assign p2_smul_72282_comb = smul21b_12b_x_9b(p2_clipped__62_comb, 9'h0b5);
  assign p2_smul_72283_comb = smul21b_12b_x_9b(p2_clipped__78_comb, 9'h0b5);
  assign p2_smul_72284_comb = smul21b_12b_x_9b(p2_clipped__94_comb, 9'h14b);
  assign p2_smul_72285_comb = smul21b_12b_x_9b(p2_clipped__110_comb, 9'h14b);
  assign p2_smul_72286_comb = smul21b_12b_x_9b(p2_clipped__126_comb, 9'h0b5);
  assign p2_smul_72287_comb = smul21b_12b_x_9b(p2_clipped__15_comb, 9'h0b5);
  assign p2_smul_72288_comb = smul21b_12b_x_9b(p2_clipped__31_comb, 9'h14b);
  assign p2_smul_72289_comb = smul21b_12b_x_9b(p2_clipped__47_comb, 9'h14b);
  assign p2_smul_72290_comb = smul21b_12b_x_9b(p2_clipped__63_comb, 9'h0b5);
  assign p2_smul_72291_comb = smul21b_12b_x_9b(p2_clipped__79_comb, 9'h0b5);
  assign p2_smul_72292_comb = smul21b_12b_x_9b(p2_clipped__95_comb, 9'h14b);
  assign p2_smul_72293_comb = smul21b_12b_x_9b(p2_clipped__111_comb, 9'h14b);
  assign p2_smul_72294_comb = smul21b_12b_x_9b(p2_clipped__127_comb, 9'h0b5);
  assign p2_add_72621_comb = p2_smul_28634_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72622_comb = p2_smul_28636_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72729_comb = p2_smul_28758_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72730_comb = p2_smul_28760_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72735_comb = p2_smul_28766_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72736_comb = p2_smul_28768_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72825_comb = p2_smul_28886_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72834_comb = p2_smul_28896_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73067_comb = p2_smul_29144_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73072_comb = p2_smul_29150_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73175_comb = p2_smul_29268_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73178_comb = p2_smul_29272_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73183_comb = p2_smul_29278_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73186_comb = p2_smul_29282_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73271_comb = p2_smul_29396_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73284_comb = p2_smul_29410_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73383_comb = {{1{p2_clipped__8_comb[11]}}, p2_clipped__8_comb} + {{1{p2_clipped__24_comb[11]}}, p2_clipped__24_comb};
  assign p2_add_73384_comb = {{1{p2_clipped__40_comb[11]}}, p2_clipped__40_comb} + {{1{p2_clipped__56_comb[11]}}, p2_clipped__56_comb};
  assign p2_add_73385_comb = {{1{p2_clipped__72_comb[11]}}, p2_clipped__72_comb} + {{1{p2_clipped__88_comb[11]}}, p2_clipped__88_comb};
  assign p2_add_73386_comb = {{1{p2_clipped__104_comb[11]}}, p2_clipped__104_comb} + {{1{p2_clipped__120_comb[11]}}, p2_clipped__120_comb};
  assign p2_add_73607_comb = p2_smul_72231_comb[20:7] + 14'h0001;
  assign p2_add_73608_comb = p2_smul_72232_comb[20:7] + 14'h0001;
  assign p2_add_73609_comb = p2_smul_72233_comb[20:7] + 14'h0001;
  assign p2_add_73610_comb = p2_smul_72234_comb[20:7] + 14'h0001;
  assign p2_add_73611_comb = p2_smul_72235_comb[20:7] + 14'h0001;
  assign p2_add_73612_comb = p2_smul_72236_comb[20:7] + 14'h0001;
  assign p2_add_73613_comb = p2_smul_72237_comb[20:7] + 14'h0001;
  assign p2_add_73614_comb = p2_smul_72238_comb[20:7] + 14'h0001;
  assign p2_smul_28650_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__57_comb, 6'h19);
  assign p2_smul_28652_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__73_comb, 6'h27);
  assign p2_smul_28666_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__58_comb, 6'h19);
  assign p2_smul_28668_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__74_comb, 6'h27);
  assign p2_smul_28682_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__59_comb, 6'h19);
  assign p2_smul_28684_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__75_comb, 6'h27);
  assign p2_smul_28698_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__60_comb, 6'h19);
  assign p2_smul_28700_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__76_comb, 6'h27);
  assign p2_smul_28714_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__61_comb, 6'h19);
  assign p2_smul_28716_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__77_comb, 6'h27);
  assign p2_smul_28730_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__62_comb, 6'h19);
  assign p2_smul_28732_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__78_comb, 6'h27);
  assign p2_smul_28746_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__63_comb, 6'h19);
  assign p2_smul_28748_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__79_comb, 6'h27);
  assign p2_smul_28774_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__25_comb, 7'h31);
  assign p2_smul_28776_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__41_comb, 7'h4f);
  assign p2_smul_28782_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__89_comb, 7'h4f);
  assign p2_smul_28784_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__105_comb, 7'h31);
  assign p2_smul_28790_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__26_comb, 7'h31);
  assign p2_smul_28792_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__42_comb, 7'h4f);
  assign p2_smul_28798_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__90_comb, 7'h4f);
  assign p2_smul_28800_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__106_comb, 7'h31);
  assign p2_smul_28806_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__27_comb, 7'h31);
  assign p2_smul_28808_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__43_comb, 7'h4f);
  assign p2_smul_28814_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__91_comb, 7'h4f);
  assign p2_smul_28816_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__107_comb, 7'h31);
  assign p2_smul_28822_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__28_comb, 7'h31);
  assign p2_smul_28824_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__44_comb, 7'h4f);
  assign p2_smul_28830_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__92_comb, 7'h4f);
  assign p2_smul_28832_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__108_comb, 7'h31);
  assign p2_smul_28838_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__29_comb, 7'h31);
  assign p2_smul_28840_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__45_comb, 7'h4f);
  assign p2_smul_28846_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__93_comb, 7'h4f);
  assign p2_smul_28848_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__109_comb, 7'h31);
  assign p2_smul_28854_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__30_comb, 7'h31);
  assign p2_smul_28856_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__46_comb, 7'h4f);
  assign p2_smul_28862_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__94_comb, 7'h4f);
  assign p2_smul_28864_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__110_comb, 7'h31);
  assign p2_smul_28870_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__31_comb, 7'h31);
  assign p2_smul_28872_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__47_comb, 7'h4f);
  assign p2_smul_28878_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__95_comb, 7'h4f);
  assign p2_smul_28880_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__111_comb, 7'h31);
  assign p2_smul_28902_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__25_comb, 6'h27);
  assign p2_smul_28912_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__105_comb, 6'h19);
  assign p2_smul_28918_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__26_comb, 6'h27);
  assign p2_smul_28928_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__106_comb, 6'h19);
  assign p2_smul_28934_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__27_comb, 6'h27);
  assign p2_smul_28944_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__107_comb, 6'h19);
  assign p2_smul_28950_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__28_comb, 6'h27);
  assign p2_smul_28960_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__108_comb, 6'h19);
  assign p2_smul_28966_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__29_comb, 6'h27);
  assign p2_smul_28976_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__109_comb, 6'h19);
  assign p2_smul_28982_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__30_comb, 6'h27);
  assign p2_smul_28992_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__110_comb, 6'h19);
  assign p2_smul_28998_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__31_comb, 6'h27);
  assign p2_smul_29008_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__111_comb, 6'h19);
  assign p2_smul_29160_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__41_comb, 6'h27);
  assign p2_smul_29166_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__89_comb, 6'h27);
  assign p2_smul_29176_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__42_comb, 6'h27);
  assign p2_smul_29182_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__90_comb, 6'h27);
  assign p2_smul_29192_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__43_comb, 6'h27);
  assign p2_smul_29198_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__91_comb, 6'h27);
  assign p2_smul_29208_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__44_comb, 6'h27);
  assign p2_smul_29214_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__92_comb, 6'h27);
  assign p2_smul_29224_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__45_comb, 6'h27);
  assign p2_smul_29230_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__93_comb, 6'h27);
  assign p2_smul_29240_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__46_comb, 6'h27);
  assign p2_smul_29246_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__94_comb, 6'h27);
  assign p2_smul_29256_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__47_comb, 6'h27);
  assign p2_smul_29262_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__95_comb, 6'h27);
  assign p2_smul_29284_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__9_comb, 7'h31);
  assign p2_smul_29288_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__41_comb, 7'h31);
  assign p2_smul_29294_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__89_comb, 7'h31);
  assign p2_smul_29298_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__121_comb, 7'h31);
  assign p2_smul_29300_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__10_comb, 7'h31);
  assign p2_smul_29304_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__42_comb, 7'h31);
  assign p2_smul_29310_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__90_comb, 7'h31);
  assign p2_smul_29314_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__122_comb, 7'h31);
  assign p2_smul_29316_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__11_comb, 7'h31);
  assign p2_smul_29320_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__43_comb, 7'h31);
  assign p2_smul_29326_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__91_comb, 7'h31);
  assign p2_smul_29330_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__123_comb, 7'h31);
  assign p2_smul_29332_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__12_comb, 7'h31);
  assign p2_smul_29336_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__44_comb, 7'h31);
  assign p2_smul_29342_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__92_comb, 7'h31);
  assign p2_smul_29346_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__124_comb, 7'h31);
  assign p2_smul_29348_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__13_comb, 7'h31);
  assign p2_smul_29352_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__45_comb, 7'h31);
  assign p2_smul_29358_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__93_comb, 7'h31);
  assign p2_smul_29362_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__125_comb, 7'h31);
  assign p2_smul_29364_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__14_comb, 7'h31);
  assign p2_smul_29368_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__46_comb, 7'h31);
  assign p2_smul_29374_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__94_comb, 7'h31);
  assign p2_smul_29378_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__126_comb, 7'h31);
  assign p2_smul_29380_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__15_comb, 7'h31);
  assign p2_smul_29384_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__47_comb, 7'h31);
  assign p2_smul_29390_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__95_comb, 7'h31);
  assign p2_smul_29394_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__127_comb, 7'h31);
  assign p2_smul_29412_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__9_comb, 6'h19);
  assign p2_smul_29426_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__121_comb, 6'h19);
  assign p2_smul_29428_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__10_comb, 6'h19);
  assign p2_smul_29442_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__122_comb, 6'h19);
  assign p2_smul_29444_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__11_comb, 6'h19);
  assign p2_smul_29458_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__123_comb, 6'h19);
  assign p2_smul_29460_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__12_comb, 6'h19);
  assign p2_smul_29474_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__124_comb, 6'h19);
  assign p2_smul_29476_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__13_comb, 6'h19);
  assign p2_smul_29490_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__125_comb, 6'h19);
  assign p2_smul_29492_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__14_comb, 6'h19);
  assign p2_smul_29506_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__126_comb, 6'h19);
  assign p2_smul_29508_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__15_comb, 6'h19);
  assign p2_smul_29522_NarrowedMult__comb = smul18b_12b_x_6b(p2_clipped__127_comb, 6'h19);
  assign p2_add_73387_comb = {{1{p2_clipped__9_comb[11]}}, p2_clipped__9_comb} + {{1{p2_clipped__25_comb[11]}}, p2_clipped__25_comb};
  assign p2_add_73388_comb = {{1{p2_clipped__41_comb[11]}}, p2_clipped__41_comb} + {{1{p2_clipped__57_comb[11]}}, p2_clipped__57_comb};
  assign p2_add_73389_comb = {{1{p2_clipped__73_comb[11]}}, p2_clipped__73_comb} + {{1{p2_clipped__89_comb[11]}}, p2_clipped__89_comb};
  assign p2_add_73390_comb = {{1{p2_clipped__105_comb[11]}}, p2_clipped__105_comb} + {{1{p2_clipped__121_comb[11]}}, p2_clipped__121_comb};
  assign p2_add_73391_comb = {{1{p2_clipped__10_comb[11]}}, p2_clipped__10_comb} + {{1{p2_clipped__26_comb[11]}}, p2_clipped__26_comb};
  assign p2_add_73392_comb = {{1{p2_clipped__42_comb[11]}}, p2_clipped__42_comb} + {{1{p2_clipped__58_comb[11]}}, p2_clipped__58_comb};
  assign p2_add_73393_comb = {{1{p2_clipped__74_comb[11]}}, p2_clipped__74_comb} + {{1{p2_clipped__90_comb[11]}}, p2_clipped__90_comb};
  assign p2_add_73394_comb = {{1{p2_clipped__106_comb[11]}}, p2_clipped__106_comb} + {{1{p2_clipped__122_comb[11]}}, p2_clipped__122_comb};
  assign p2_add_73395_comb = {{1{p2_clipped__11_comb[11]}}, p2_clipped__11_comb} + {{1{p2_clipped__27_comb[11]}}, p2_clipped__27_comb};
  assign p2_add_73396_comb = {{1{p2_clipped__43_comb[11]}}, p2_clipped__43_comb} + {{1{p2_clipped__59_comb[11]}}, p2_clipped__59_comb};
  assign p2_add_73397_comb = {{1{p2_clipped__75_comb[11]}}, p2_clipped__75_comb} + {{1{p2_clipped__91_comb[11]}}, p2_clipped__91_comb};
  assign p2_add_73398_comb = {{1{p2_clipped__107_comb[11]}}, p2_clipped__107_comb} + {{1{p2_clipped__123_comb[11]}}, p2_clipped__123_comb};
  assign p2_add_73399_comb = {{1{p2_clipped__12_comb[11]}}, p2_clipped__12_comb} + {{1{p2_clipped__28_comb[11]}}, p2_clipped__28_comb};
  assign p2_add_73400_comb = {{1{p2_clipped__44_comb[11]}}, p2_clipped__44_comb} + {{1{p2_clipped__60_comb[11]}}, p2_clipped__60_comb};
  assign p2_add_73401_comb = {{1{p2_clipped__76_comb[11]}}, p2_clipped__76_comb} + {{1{p2_clipped__92_comb[11]}}, p2_clipped__92_comb};
  assign p2_add_73402_comb = {{1{p2_clipped__108_comb[11]}}, p2_clipped__108_comb} + {{1{p2_clipped__124_comb[11]}}, p2_clipped__124_comb};
  assign p2_add_73403_comb = {{1{p2_clipped__13_comb[11]}}, p2_clipped__13_comb} + {{1{p2_clipped__29_comb[11]}}, p2_clipped__29_comb};
  assign p2_add_73404_comb = {{1{p2_clipped__45_comb[11]}}, p2_clipped__45_comb} + {{1{p2_clipped__61_comb[11]}}, p2_clipped__61_comb};
  assign p2_add_73405_comb = {{1{p2_clipped__77_comb[11]}}, p2_clipped__77_comb} + {{1{p2_clipped__93_comb[11]}}, p2_clipped__93_comb};
  assign p2_add_73406_comb = {{1{p2_clipped__109_comb[11]}}, p2_clipped__109_comb} + {{1{p2_clipped__125_comb[11]}}, p2_clipped__125_comb};
  assign p2_add_73407_comb = {{1{p2_clipped__14_comb[11]}}, p2_clipped__14_comb} + {{1{p2_clipped__30_comb[11]}}, p2_clipped__30_comb};
  assign p2_add_73408_comb = {{1{p2_clipped__46_comb[11]}}, p2_clipped__46_comb} + {{1{p2_clipped__62_comb[11]}}, p2_clipped__62_comb};
  assign p2_add_73409_comb = {{1{p2_clipped__78_comb[11]}}, p2_clipped__78_comb} + {{1{p2_clipped__94_comb[11]}}, p2_clipped__94_comb};
  assign p2_add_73410_comb = {{1{p2_clipped__110_comb[11]}}, p2_clipped__110_comb} + {{1{p2_clipped__126_comb[11]}}, p2_clipped__126_comb};
  assign p2_add_73411_comb = {{1{p2_clipped__15_comb[11]}}, p2_clipped__15_comb} + {{1{p2_clipped__31_comb[11]}}, p2_clipped__31_comb};
  assign p2_add_73412_comb = {{1{p2_clipped__47_comb[11]}}, p2_clipped__47_comb} + {{1{p2_clipped__63_comb[11]}}, p2_clipped__63_comb};
  assign p2_add_73413_comb = {{1{p2_clipped__79_comb[11]}}, p2_clipped__79_comb} + {{1{p2_clipped__95_comb[11]}}, p2_clipped__95_comb};
  assign p2_add_73414_comb = {{1{p2_clipped__111_comb[11]}}, p2_clipped__111_comb} + {{1{p2_clipped__127_comb[11]}}, p2_clipped__127_comb};
  assign p2_add_73415_comb = p2_smul_71975_comb[20:7] + 14'h0001;
  assign p2_add_73416_comb = p2_smul_71976_comb[20:7] + 14'h0001;
  assign p2_add_73417_comb = p2_smul_28632_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73418_comb = p2_add_72621_comb[11:1];
  assign p2_bit_slice_73419_comb = p2_add_72622_comb[11:1];
  assign p2_add_73420_comb = p2_smul_28638_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73421_comb = p2_smul_71983_comb[20:7] + 14'h0001;
  assign p2_add_73422_comb = p2_smul_71984_comb[20:7] + 14'h0001;
  assign p2_add_73479_comb = p2_smul_28756_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73480_comb = p2_add_72729_comb[12:1];
  assign p2_bit_slice_73481_comb = p2_add_72730_comb[12:1];
  assign p2_add_73482_comb = p2_smul_28762_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73483_comb = p2_smul_28764_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73484_comb = p2_add_72735_comb[12:1];
  assign p2_bit_slice_73485_comb = p2_add_72736_comb[12:1];
  assign p2_add_73486_comb = p2_smul_28770_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73543_comb = p2_smul_72151_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73544_comb = p2_add_72825_comb[11:1];
  assign p2_add_73545_comb = p2_smul_72154_comb[20:7] + 14'h0001;
  assign p2_add_73546_comb = p2_smul_28890_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73547_comb = p2_smul_28892_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73548_comb = p2_smul_72157_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73549_comb = p2_add_72834_comb[11:1];
  assign p2_add_73550_comb = p2_smul_72160_comb[20:7] + 14'h0001;
  assign p2_add_73671_comb = p2_smul_29140_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73672_comb = p2_smul_72296_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73673_comb = p2_add_73067_comb[11:1];
  assign p2_add_73674_comb = p2_smul_72299_comb[20:7] + 14'h0001;
  assign p2_add_73675_comb = p2_smul_72300_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73676_comb = p2_add_73072_comb[11:1];
  assign p2_add_73677_comb = p2_smul_72303_comb[20:7] + 14'h0001;
  assign p2_add_73678_comb = p2_smul_29154_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73735_comb = p2_add_73175_comb[12:1];
  assign p2_add_73736_comb = p2_smul_29270_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73737_comb = p2_add_73178_comb[12:1];
  assign p2_add_73738_comb = p2_smul_29274_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73739_comb = p2_smul_29276_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73740_comb = p2_add_73183_comb[12:1];
  assign p2_add_73741_comb = p2_smul_29280_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73742_comb = p2_add_73186_comb[12:1];
  assign p2_bit_slice_73799_comb = p2_add_73271_comb[11:1];
  assign p2_add_73800_comb = p2_smul_29398_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73801_comb = p2_smul_72474_comb[20:7] + 14'h0001;
  assign p2_add_73802_comb = p2_smul_72475_comb[20:7] + 14'h0001;
  assign p2_add_73803_comb = p2_smul_72476_comb[20:7] + 14'h0001;
  assign p2_add_73804_comb = p2_smul_72477_comb[20:7] + 14'h0001;
  assign p2_add_73805_comb = p2_smul_29408_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73806_comb = p2_add_73284_comb[11:1];
  assign p2_sum__520_comb = {{19{p2_add_73383_comb[12]}}, p2_add_73383_comb};
  assign p2_sum__521_comb = {{19{p2_add_73384_comb[12]}}, p2_add_73384_comb};
  assign p2_sum__522_comb = {{19{p2_add_73385_comb[12]}}, p2_add_73385_comb};
  assign p2_sum__523_comb = {{19{p2_add_73386_comb[12]}}, p2_add_73386_comb};
  assign p2_smul_71985_comb = smul21b_12b_x_9b(p2_clipped__9_comb, 9'h0fb);
  assign p2_smul_71986_comb = smul21b_12b_x_9b(p2_clipped__25_comb, 9'h0d5);
  assign p2_smul_28648_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__41_comb, 8'h47);
  assign p2_smul_28654_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__89_comb, 8'hb9);
  assign p2_smul_71993_comb = smul21b_12b_x_9b(p2_clipped__105_comb, 9'h12b);
  assign p2_smul_71994_comb = smul21b_12b_x_9b(p2_clipped__121_comb, 9'h105);
  assign p2_smul_71995_comb = smul21b_12b_x_9b(p2_clipped__10_comb, 9'h0fb);
  assign p2_smul_71996_comb = smul21b_12b_x_9b(p2_clipped__26_comb, 9'h0d5);
  assign p2_smul_28664_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__42_comb, 8'h47);
  assign p2_smul_28670_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__90_comb, 8'hb9);
  assign p2_smul_72003_comb = smul21b_12b_x_9b(p2_clipped__106_comb, 9'h12b);
  assign p2_smul_72004_comb = smul21b_12b_x_9b(p2_clipped__122_comb, 9'h105);
  assign p2_smul_72005_comb = smul21b_12b_x_9b(p2_clipped__11_comb, 9'h0fb);
  assign p2_smul_72006_comb = smul21b_12b_x_9b(p2_clipped__27_comb, 9'h0d5);
  assign p2_smul_28680_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__43_comb, 8'h47);
  assign p2_smul_28686_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__91_comb, 8'hb9);
  assign p2_smul_72013_comb = smul21b_12b_x_9b(p2_clipped__107_comb, 9'h12b);
  assign p2_smul_72014_comb = smul21b_12b_x_9b(p2_clipped__123_comb, 9'h105);
  assign p2_smul_72015_comb = smul21b_12b_x_9b(p2_clipped__12_comb, 9'h0fb);
  assign p2_smul_72016_comb = smul21b_12b_x_9b(p2_clipped__28_comb, 9'h0d5);
  assign p2_smul_28696_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__44_comb, 8'h47);
  assign p2_smul_28702_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__92_comb, 8'hb9);
  assign p2_smul_72023_comb = smul21b_12b_x_9b(p2_clipped__108_comb, 9'h12b);
  assign p2_smul_72024_comb = smul21b_12b_x_9b(p2_clipped__124_comb, 9'h105);
  assign p2_smul_72025_comb = smul21b_12b_x_9b(p2_clipped__13_comb, 9'h0fb);
  assign p2_smul_72026_comb = smul21b_12b_x_9b(p2_clipped__29_comb, 9'h0d5);
  assign p2_smul_28712_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__45_comb, 8'h47);
  assign p2_smul_28718_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__93_comb, 8'hb9);
  assign p2_smul_72033_comb = smul21b_12b_x_9b(p2_clipped__109_comb, 9'h12b);
  assign p2_smul_72034_comb = smul21b_12b_x_9b(p2_clipped__125_comb, 9'h105);
  assign p2_smul_72035_comb = smul21b_12b_x_9b(p2_clipped__14_comb, 9'h0fb);
  assign p2_smul_72036_comb = smul21b_12b_x_9b(p2_clipped__30_comb, 9'h0d5);
  assign p2_smul_28728_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__46_comb, 8'h47);
  assign p2_smul_28734_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__94_comb, 8'hb9);
  assign p2_smul_72043_comb = smul21b_12b_x_9b(p2_clipped__110_comb, 9'h12b);
  assign p2_smul_72044_comb = smul21b_12b_x_9b(p2_clipped__126_comb, 9'h105);
  assign p2_smul_72045_comb = smul21b_12b_x_9b(p2_clipped__15_comb, 9'h0fb);
  assign p2_smul_72046_comb = smul21b_12b_x_9b(p2_clipped__31_comb, 9'h0d5);
  assign p2_smul_28744_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__47_comb, 8'h47);
  assign p2_smul_28750_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__95_comb, 8'hb9);
  assign p2_smul_72053_comb = smul21b_12b_x_9b(p2_clipped__111_comb, 9'h12b);
  assign p2_smul_72054_comb = smul21b_12b_x_9b(p2_clipped__127_comb, 9'h105);
  assign p2_smul_28772_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__9_comb, 7'h3b);
  assign p2_smul_28778_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__57_comb, 7'h45);
  assign p2_smul_28780_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__73_comb, 7'h45);
  assign p2_smul_28786_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__121_comb, 7'h3b);
  assign p2_smul_28788_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__10_comb, 7'h3b);
  assign p2_smul_28794_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__58_comb, 7'h45);
  assign p2_smul_28796_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__74_comb, 7'h45);
  assign p2_smul_28802_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__122_comb, 7'h3b);
  assign p2_smul_28804_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__11_comb, 7'h3b);
  assign p2_smul_28810_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__59_comb, 7'h45);
  assign p2_smul_28812_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__75_comb, 7'h45);
  assign p2_smul_28818_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__123_comb, 7'h3b);
  assign p2_smul_28820_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__12_comb, 7'h3b);
  assign p2_smul_28826_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__60_comb, 7'h45);
  assign p2_smul_28828_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__76_comb, 7'h45);
  assign p2_smul_28834_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__124_comb, 7'h3b);
  assign p2_smul_28836_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__13_comb, 7'h3b);
  assign p2_smul_28842_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__61_comb, 7'h45);
  assign p2_smul_28844_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__77_comb, 7'h45);
  assign p2_smul_28850_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__125_comb, 7'h3b);
  assign p2_smul_28852_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__14_comb, 7'h3b);
  assign p2_smul_28858_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__62_comb, 7'h45);
  assign p2_smul_28860_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__78_comb, 7'h45);
  assign p2_smul_28866_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__126_comb, 7'h3b);
  assign p2_smul_28868_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__15_comb, 7'h3b);
  assign p2_smul_28874_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__63_comb, 7'h45);
  assign p2_smul_28876_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__79_comb, 7'h45);
  assign p2_smul_28882_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__127_comb, 7'h3b);
  assign p2_smul_72161_comb = smul21b_12b_x_9b(p2_clipped__9_comb, 9'h0d5);
  assign p2_smul_72164_comb = smul21b_12b_x_9b(p2_clipped__41_comb, 9'h105);
  assign p2_smul_28906_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__57_comb, 8'hb9);
  assign p2_smul_28908_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__73_comb, 8'h47);
  assign p2_smul_72167_comb = smul21b_12b_x_9b(p2_clipped__89_comb, 9'h0fb);
  assign p2_smul_72170_comb = smul21b_12b_x_9b(p2_clipped__121_comb, 9'h12b);
  assign p2_smul_72171_comb = smul21b_12b_x_9b(p2_clipped__10_comb, 9'h0d5);
  assign p2_smul_72174_comb = smul21b_12b_x_9b(p2_clipped__42_comb, 9'h105);
  assign p2_smul_28922_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__58_comb, 8'hb9);
  assign p2_smul_28924_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__74_comb, 8'h47);
  assign p2_smul_72177_comb = smul21b_12b_x_9b(p2_clipped__90_comb, 9'h0fb);
  assign p2_smul_72180_comb = smul21b_12b_x_9b(p2_clipped__122_comb, 9'h12b);
  assign p2_smul_72181_comb = smul21b_12b_x_9b(p2_clipped__11_comb, 9'h0d5);
  assign p2_smul_72184_comb = smul21b_12b_x_9b(p2_clipped__43_comb, 9'h105);
  assign p2_smul_28938_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__59_comb, 8'hb9);
  assign p2_smul_28940_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__75_comb, 8'h47);
  assign p2_smul_72187_comb = smul21b_12b_x_9b(p2_clipped__91_comb, 9'h0fb);
  assign p2_smul_72190_comb = smul21b_12b_x_9b(p2_clipped__123_comb, 9'h12b);
  assign p2_smul_72191_comb = smul21b_12b_x_9b(p2_clipped__12_comb, 9'h0d5);
  assign p2_smul_72194_comb = smul21b_12b_x_9b(p2_clipped__44_comb, 9'h105);
  assign p2_smul_28954_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__60_comb, 8'hb9);
  assign p2_smul_28956_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__76_comb, 8'h47);
  assign p2_smul_72197_comb = smul21b_12b_x_9b(p2_clipped__92_comb, 9'h0fb);
  assign p2_smul_72200_comb = smul21b_12b_x_9b(p2_clipped__124_comb, 9'h12b);
  assign p2_smul_72201_comb = smul21b_12b_x_9b(p2_clipped__13_comb, 9'h0d5);
  assign p2_smul_72204_comb = smul21b_12b_x_9b(p2_clipped__45_comb, 9'h105);
  assign p2_smul_28970_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__61_comb, 8'hb9);
  assign p2_smul_28972_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__77_comb, 8'h47);
  assign p2_smul_72207_comb = smul21b_12b_x_9b(p2_clipped__93_comb, 9'h0fb);
  assign p2_smul_72210_comb = smul21b_12b_x_9b(p2_clipped__125_comb, 9'h12b);
  assign p2_smul_72211_comb = smul21b_12b_x_9b(p2_clipped__14_comb, 9'h0d5);
  assign p2_smul_72214_comb = smul21b_12b_x_9b(p2_clipped__46_comb, 9'h105);
  assign p2_smul_28986_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__62_comb, 8'hb9);
  assign p2_smul_28988_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__78_comb, 8'h47);
  assign p2_smul_72217_comb = smul21b_12b_x_9b(p2_clipped__94_comb, 9'h0fb);
  assign p2_smul_72220_comb = smul21b_12b_x_9b(p2_clipped__126_comb, 9'h12b);
  assign p2_smul_72221_comb = smul21b_12b_x_9b(p2_clipped__15_comb, 9'h0d5);
  assign p2_smul_72224_comb = smul21b_12b_x_9b(p2_clipped__47_comb, 9'h105);
  assign p2_smul_29002_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__63_comb, 8'hb9);
  assign p2_smul_29004_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__79_comb, 8'h47);
  assign p2_smul_72227_comb = smul21b_12b_x_9b(p2_clipped__95_comb, 9'h0fb);
  assign p2_smul_72230_comb = smul21b_12b_x_9b(p2_clipped__127_comb, 9'h12b);
  assign p2_smul_29156_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__9_comb, 8'h47);
  assign p2_smul_72306_comb = smul21b_12b_x_9b(p2_clipped__25_comb, 9'h105);
  assign p2_smul_72309_comb = smul21b_12b_x_9b(p2_clipped__57_comb, 9'h0d5);
  assign p2_smul_72310_comb = smul21b_12b_x_9b(p2_clipped__73_comb, 9'h0d5);
  assign p2_smul_72313_comb = smul21b_12b_x_9b(p2_clipped__105_comb, 9'h105);
  assign p2_smul_29170_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__121_comb, 8'h47);
  assign p2_smul_29172_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__10_comb, 8'h47);
  assign p2_smul_72316_comb = smul21b_12b_x_9b(p2_clipped__26_comb, 9'h105);
  assign p2_smul_72319_comb = smul21b_12b_x_9b(p2_clipped__58_comb, 9'h0d5);
  assign p2_smul_72320_comb = smul21b_12b_x_9b(p2_clipped__74_comb, 9'h0d5);
  assign p2_smul_72323_comb = smul21b_12b_x_9b(p2_clipped__106_comb, 9'h105);
  assign p2_smul_29186_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__122_comb, 8'h47);
  assign p2_smul_29188_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__11_comb, 8'h47);
  assign p2_smul_72326_comb = smul21b_12b_x_9b(p2_clipped__27_comb, 9'h105);
  assign p2_smul_72329_comb = smul21b_12b_x_9b(p2_clipped__59_comb, 9'h0d5);
  assign p2_smul_72330_comb = smul21b_12b_x_9b(p2_clipped__75_comb, 9'h0d5);
  assign p2_smul_72333_comb = smul21b_12b_x_9b(p2_clipped__107_comb, 9'h105);
  assign p2_smul_29202_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__123_comb, 8'h47);
  assign p2_smul_29204_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__12_comb, 8'h47);
  assign p2_smul_72336_comb = smul21b_12b_x_9b(p2_clipped__28_comb, 9'h105);
  assign p2_smul_72339_comb = smul21b_12b_x_9b(p2_clipped__60_comb, 9'h0d5);
  assign p2_smul_72340_comb = smul21b_12b_x_9b(p2_clipped__76_comb, 9'h0d5);
  assign p2_smul_72343_comb = smul21b_12b_x_9b(p2_clipped__108_comb, 9'h105);
  assign p2_smul_29218_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__124_comb, 8'h47);
  assign p2_smul_29220_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__13_comb, 8'h47);
  assign p2_smul_72346_comb = smul21b_12b_x_9b(p2_clipped__29_comb, 9'h105);
  assign p2_smul_72349_comb = smul21b_12b_x_9b(p2_clipped__61_comb, 9'h0d5);
  assign p2_smul_72350_comb = smul21b_12b_x_9b(p2_clipped__77_comb, 9'h0d5);
  assign p2_smul_72353_comb = smul21b_12b_x_9b(p2_clipped__109_comb, 9'h105);
  assign p2_smul_29234_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__125_comb, 8'h47);
  assign p2_smul_29236_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__14_comb, 8'h47);
  assign p2_smul_72356_comb = smul21b_12b_x_9b(p2_clipped__30_comb, 9'h105);
  assign p2_smul_72359_comb = smul21b_12b_x_9b(p2_clipped__62_comb, 9'h0d5);
  assign p2_smul_72360_comb = smul21b_12b_x_9b(p2_clipped__78_comb, 9'h0d5);
  assign p2_smul_72363_comb = smul21b_12b_x_9b(p2_clipped__110_comb, 9'h105);
  assign p2_smul_29250_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__126_comb, 8'h47);
  assign p2_smul_29252_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__15_comb, 8'h47);
  assign p2_smul_72366_comb = smul21b_12b_x_9b(p2_clipped__31_comb, 9'h105);
  assign p2_smul_72369_comb = smul21b_12b_x_9b(p2_clipped__63_comb, 9'h0d5);
  assign p2_smul_72370_comb = smul21b_12b_x_9b(p2_clipped__79_comb, 9'h0d5);
  assign p2_smul_72373_comb = smul21b_12b_x_9b(p2_clipped__111_comb, 9'h105);
  assign p2_smul_29266_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__127_comb, 8'h47);
  assign p2_smul_29286_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__25_comb, 7'h45);
  assign p2_smul_29290_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__57_comb, 7'h3b);
  assign p2_smul_29292_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__73_comb, 7'h3b);
  assign p2_smul_29296_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__105_comb, 7'h45);
  assign p2_smul_29302_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__26_comb, 7'h45);
  assign p2_smul_29306_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__58_comb, 7'h3b);
  assign p2_smul_29308_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__74_comb, 7'h3b);
  assign p2_smul_29312_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__106_comb, 7'h45);
  assign p2_smul_29318_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__27_comb, 7'h45);
  assign p2_smul_29322_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__59_comb, 7'h3b);
  assign p2_smul_29324_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__75_comb, 7'h3b);
  assign p2_smul_29328_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__107_comb, 7'h45);
  assign p2_smul_29334_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__28_comb, 7'h45);
  assign p2_smul_29338_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__60_comb, 7'h3b);
  assign p2_smul_29340_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__76_comb, 7'h3b);
  assign p2_smul_29344_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__108_comb, 7'h45);
  assign p2_smul_29350_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__29_comb, 7'h45);
  assign p2_smul_29354_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__61_comb, 7'h3b);
  assign p2_smul_29356_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__77_comb, 7'h3b);
  assign p2_smul_29360_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__109_comb, 7'h45);
  assign p2_smul_29366_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__30_comb, 7'h45);
  assign p2_smul_29370_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__62_comb, 7'h3b);
  assign p2_smul_29372_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__78_comb, 7'h3b);
  assign p2_smul_29376_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__110_comb, 7'h45);
  assign p2_smul_29382_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__31_comb, 7'h45);
  assign p2_smul_29386_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__63_comb, 7'h3b);
  assign p2_smul_29388_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__79_comb, 7'h3b);
  assign p2_smul_29392_NarrowedMult__comb = smul19b_12b_x_7b(p2_clipped__111_comb, 7'h45);
  assign p2_smul_29414_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__25_comb, 8'hb9);
  assign p2_smul_72484_comb = smul21b_12b_x_9b(p2_clipped__41_comb, 9'h0d5);
  assign p2_smul_72485_comb = smul21b_12b_x_9b(p2_clipped__57_comb, 9'h105);
  assign p2_smul_72486_comb = smul21b_12b_x_9b(p2_clipped__73_comb, 9'h105);
  assign p2_smul_72487_comb = smul21b_12b_x_9b(p2_clipped__89_comb, 9'h0d5);
  assign p2_smul_29424_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__105_comb, 8'hb9);
  assign p2_smul_29430_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__26_comb, 8'hb9);
  assign p2_smul_72494_comb = smul21b_12b_x_9b(p2_clipped__42_comb, 9'h0d5);
  assign p2_smul_72495_comb = smul21b_12b_x_9b(p2_clipped__58_comb, 9'h105);
  assign p2_smul_72496_comb = smul21b_12b_x_9b(p2_clipped__74_comb, 9'h105);
  assign p2_smul_72497_comb = smul21b_12b_x_9b(p2_clipped__90_comb, 9'h0d5);
  assign p2_smul_29440_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__106_comb, 8'hb9);
  assign p2_smul_29446_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__27_comb, 8'hb9);
  assign p2_smul_72504_comb = smul21b_12b_x_9b(p2_clipped__43_comb, 9'h0d5);
  assign p2_smul_72505_comb = smul21b_12b_x_9b(p2_clipped__59_comb, 9'h105);
  assign p2_smul_72506_comb = smul21b_12b_x_9b(p2_clipped__75_comb, 9'h105);
  assign p2_smul_72507_comb = smul21b_12b_x_9b(p2_clipped__91_comb, 9'h0d5);
  assign p2_smul_29456_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__107_comb, 8'hb9);
  assign p2_smul_29462_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__28_comb, 8'hb9);
  assign p2_smul_72514_comb = smul21b_12b_x_9b(p2_clipped__44_comb, 9'h0d5);
  assign p2_smul_72515_comb = smul21b_12b_x_9b(p2_clipped__60_comb, 9'h105);
  assign p2_smul_72516_comb = smul21b_12b_x_9b(p2_clipped__76_comb, 9'h105);
  assign p2_smul_72517_comb = smul21b_12b_x_9b(p2_clipped__92_comb, 9'h0d5);
  assign p2_smul_29472_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__108_comb, 8'hb9);
  assign p2_smul_29478_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__29_comb, 8'hb9);
  assign p2_smul_72524_comb = smul21b_12b_x_9b(p2_clipped__45_comb, 9'h0d5);
  assign p2_smul_72525_comb = smul21b_12b_x_9b(p2_clipped__61_comb, 9'h105);
  assign p2_smul_72526_comb = smul21b_12b_x_9b(p2_clipped__77_comb, 9'h105);
  assign p2_smul_72527_comb = smul21b_12b_x_9b(p2_clipped__93_comb, 9'h0d5);
  assign p2_smul_29488_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__109_comb, 8'hb9);
  assign p2_smul_29494_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__30_comb, 8'hb9);
  assign p2_smul_72534_comb = smul21b_12b_x_9b(p2_clipped__46_comb, 9'h0d5);
  assign p2_smul_72535_comb = smul21b_12b_x_9b(p2_clipped__62_comb, 9'h105);
  assign p2_smul_72536_comb = smul21b_12b_x_9b(p2_clipped__78_comb, 9'h105);
  assign p2_smul_72537_comb = smul21b_12b_x_9b(p2_clipped__94_comb, 9'h0d5);
  assign p2_smul_29504_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__110_comb, 8'hb9);
  assign p2_smul_29510_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__31_comb, 8'hb9);
  assign p2_smul_72544_comb = smul21b_12b_x_9b(p2_clipped__47_comb, 9'h0d5);
  assign p2_smul_72545_comb = smul21b_12b_x_9b(p2_clipped__63_comb, 9'h105);
  assign p2_smul_72546_comb = smul21b_12b_x_9b(p2_clipped__79_comb, 9'h105);
  assign p2_smul_72547_comb = smul21b_12b_x_9b(p2_clipped__95_comb, 9'h0d5);
  assign p2_smul_29520_NarrowedMult__comb = smul20b_12b_x_8b(p2_clipped__111_comb, 8'hb9);
  assign p2_add_73615_comb = p2_smul_72239_comb[20:7] + 14'h0001;
  assign p2_add_73616_comb = p2_smul_72240_comb[20:7] + 14'h0001;
  assign p2_add_73617_comb = p2_smul_72241_comb[20:7] + 14'h0001;
  assign p2_add_73618_comb = p2_smul_72242_comb[20:7] + 14'h0001;
  assign p2_add_73619_comb = p2_smul_72243_comb[20:7] + 14'h0001;
  assign p2_add_73620_comb = p2_smul_72244_comb[20:7] + 14'h0001;
  assign p2_add_73621_comb = p2_smul_72245_comb[20:7] + 14'h0001;
  assign p2_add_73622_comb = p2_smul_72246_comb[20:7] + 14'h0001;
  assign p2_add_73623_comb = p2_smul_72247_comb[20:7] + 14'h0001;
  assign p2_add_73624_comb = p2_smul_72248_comb[20:7] + 14'h0001;
  assign p2_add_73625_comb = p2_smul_72249_comb[20:7] + 14'h0001;
  assign p2_add_73626_comb = p2_smul_72250_comb[20:7] + 14'h0001;
  assign p2_add_73627_comb = p2_smul_72251_comb[20:7] + 14'h0001;
  assign p2_add_73628_comb = p2_smul_72252_comb[20:7] + 14'h0001;
  assign p2_add_73629_comb = p2_smul_72253_comb[20:7] + 14'h0001;
  assign p2_add_73630_comb = p2_smul_72254_comb[20:7] + 14'h0001;
  assign p2_add_73631_comb = p2_smul_72255_comb[20:7] + 14'h0001;
  assign p2_add_73632_comb = p2_smul_72256_comb[20:7] + 14'h0001;
  assign p2_add_73633_comb = p2_smul_72257_comb[20:7] + 14'h0001;
  assign p2_add_73634_comb = p2_smul_72258_comb[20:7] + 14'h0001;
  assign p2_add_73635_comb = p2_smul_72259_comb[20:7] + 14'h0001;
  assign p2_add_73636_comb = p2_smul_72260_comb[20:7] + 14'h0001;
  assign p2_add_73637_comb = p2_smul_72261_comb[20:7] + 14'h0001;
  assign p2_add_73638_comb = p2_smul_72262_comb[20:7] + 14'h0001;
  assign p2_add_73639_comb = p2_smul_72263_comb[20:7] + 14'h0001;
  assign p2_add_73640_comb = p2_smul_72264_comb[20:7] + 14'h0001;
  assign p2_add_73641_comb = p2_smul_72265_comb[20:7] + 14'h0001;
  assign p2_add_73642_comb = p2_smul_72266_comb[20:7] + 14'h0001;
  assign p2_add_73643_comb = p2_smul_72267_comb[20:7] + 14'h0001;
  assign p2_add_73644_comb = p2_smul_72268_comb[20:7] + 14'h0001;
  assign p2_add_73645_comb = p2_smul_72269_comb[20:7] + 14'h0001;
  assign p2_add_73646_comb = p2_smul_72270_comb[20:7] + 14'h0001;
  assign p2_add_73647_comb = p2_smul_72271_comb[20:7] + 14'h0001;
  assign p2_add_73648_comb = p2_smul_72272_comb[20:7] + 14'h0001;
  assign p2_add_73649_comb = p2_smul_72273_comb[20:7] + 14'h0001;
  assign p2_add_73650_comb = p2_smul_72274_comb[20:7] + 14'h0001;
  assign p2_add_73651_comb = p2_smul_72275_comb[20:7] + 14'h0001;
  assign p2_add_73652_comb = p2_smul_72276_comb[20:7] + 14'h0001;
  assign p2_add_73653_comb = p2_smul_72277_comb[20:7] + 14'h0001;
  assign p2_add_73654_comb = p2_smul_72278_comb[20:7] + 14'h0001;
  assign p2_add_73655_comb = p2_smul_72279_comb[20:7] + 14'h0001;
  assign p2_add_73656_comb = p2_smul_72280_comb[20:7] + 14'h0001;
  assign p2_add_73657_comb = p2_smul_72281_comb[20:7] + 14'h0001;
  assign p2_add_73658_comb = p2_smul_72282_comb[20:7] + 14'h0001;
  assign p2_add_73659_comb = p2_smul_72283_comb[20:7] + 14'h0001;
  assign p2_add_73660_comb = p2_smul_72284_comb[20:7] + 14'h0001;
  assign p2_add_73661_comb = p2_smul_72285_comb[20:7] + 14'h0001;
  assign p2_add_73662_comb = p2_smul_72286_comb[20:7] + 14'h0001;
  assign p2_add_73663_comb = p2_smul_72287_comb[20:7] + 14'h0001;
  assign p2_add_73664_comb = p2_smul_72288_comb[20:7] + 14'h0001;
  assign p2_add_73665_comb = p2_smul_72289_comb[20:7] + 14'h0001;
  assign p2_add_73666_comb = p2_smul_72290_comb[20:7] + 14'h0001;
  assign p2_add_73667_comb = p2_smul_72291_comb[20:7] + 14'h0001;
  assign p2_add_73668_comb = p2_smul_72292_comb[20:7] + 14'h0001;
  assign p2_add_73669_comb = p2_smul_72293_comb[20:7] + 14'h0001;
  assign p2_add_73670_comb = p2_smul_72294_comb[20:7] + 14'h0001;
  assign p2_sum__464_comb = {{19{p2_add_73387_comb[12]}}, p2_add_73387_comb};
  assign p2_sum__465_comb = {{19{p2_add_73388_comb[12]}}, p2_add_73388_comb};
  assign p2_sum__466_comb = {{19{p2_add_73389_comb[12]}}, p2_add_73389_comb};
  assign p2_sum__467_comb = {{19{p2_add_73390_comb[12]}}, p2_add_73390_comb};
  assign p2_sum__408_comb = {{19{p2_add_73391_comb[12]}}, p2_add_73391_comb};
  assign p2_sum__409_comb = {{19{p2_add_73392_comb[12]}}, p2_add_73392_comb};
  assign p2_sum__410_comb = {{19{p2_add_73393_comb[12]}}, p2_add_73393_comb};
  assign p2_sum__411_comb = {{19{p2_add_73394_comb[12]}}, p2_add_73394_comb};
  assign p2_sum__352_comb = {{19{p2_add_73395_comb[12]}}, p2_add_73395_comb};
  assign p2_sum__353_comb = {{19{p2_add_73396_comb[12]}}, p2_add_73396_comb};
  assign p2_sum__354_comb = {{19{p2_add_73397_comb[12]}}, p2_add_73397_comb};
  assign p2_sum__355_comb = {{19{p2_add_73398_comb[12]}}, p2_add_73398_comb};
  assign p2_sum__296_comb = {{19{p2_add_73399_comb[12]}}, p2_add_73399_comb};
  assign p2_sum__297_comb = {{19{p2_add_73400_comb[12]}}, p2_add_73400_comb};
  assign p2_sum__298_comb = {{19{p2_add_73401_comb[12]}}, p2_add_73401_comb};
  assign p2_sum__299_comb = {{19{p2_add_73402_comb[12]}}, p2_add_73402_comb};
  assign p2_sum__240_comb = {{19{p2_add_73403_comb[12]}}, p2_add_73403_comb};
  assign p2_sum__241_comb = {{19{p2_add_73404_comb[12]}}, p2_add_73404_comb};
  assign p2_sum__242_comb = {{19{p2_add_73405_comb[12]}}, p2_add_73405_comb};
  assign p2_sum__243_comb = {{19{p2_add_73406_comb[12]}}, p2_add_73406_comb};
  assign p2_sum__184_comb = {{19{p2_add_73407_comb[12]}}, p2_add_73407_comb};
  assign p2_sum__185_comb = {{19{p2_add_73408_comb[12]}}, p2_add_73408_comb};
  assign p2_sum__186_comb = {{19{p2_add_73409_comb[12]}}, p2_add_73409_comb};
  assign p2_sum__187_comb = {{19{p2_add_73410_comb[12]}}, p2_add_73410_comb};
  assign p2_sum__128_comb = {{19{p2_add_73411_comb[12]}}, p2_add_73411_comb};
  assign p2_sum__129_comb = {{19{p2_add_73412_comb[12]}}, p2_add_73412_comb};
  assign p2_sum__130_comb = {{19{p2_add_73413_comb[12]}}, p2_add_73413_comb};
  assign p2_sum__131_comb = {{19{p2_add_73414_comb[12]}}, p2_add_73414_comb};
  assign p2_sum__524_comb = p2_sum__520_comb + p2_sum__521_comb;
  assign p2_sum__525_comb = p2_sum__522_comb + p2_sum__523_comb;
  assign p2_add_74455_comb = p2_add_73607_comb[13:1] + p2_add_73608_comb[13:1];
  assign p2_add_74456_comb = p2_add_73609_comb[13:1] + p2_add_73610_comb[13:1];
  assign p2_add_74457_comb = p2_add_73611_comb[13:1] + p2_add_73612_comb[13:1];
  assign p2_add_74458_comb = p2_add_73613_comb[13:1] + p2_add_73614_comb[13:1];
  assign p2_add_72635_comb = p2_smul_28650_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72636_comb = p2_smul_28652_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72649_comb = p2_smul_28666_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72650_comb = p2_smul_28668_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72663_comb = p2_smul_28682_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72664_comb = p2_smul_28684_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72677_comb = p2_smul_28698_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72678_comb = p2_smul_28700_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72691_comb = p2_smul_28714_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72692_comb = p2_smul_28716_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72705_comb = p2_smul_28730_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72706_comb = p2_smul_28732_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72719_comb = p2_smul_28746_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72720_comb = p2_smul_28748_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72741_comb = p2_smul_28774_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72742_comb = p2_smul_28776_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72747_comb = p2_smul_28782_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72748_comb = p2_smul_28784_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72753_comb = p2_smul_28790_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72754_comb = p2_smul_28792_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72759_comb = p2_smul_28798_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72760_comb = p2_smul_28800_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72765_comb = p2_smul_28806_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72766_comb = p2_smul_28808_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72771_comb = p2_smul_28814_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72772_comb = p2_smul_28816_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72777_comb = p2_smul_28822_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72778_comb = p2_smul_28824_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72783_comb = p2_smul_28830_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72784_comb = p2_smul_28832_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72789_comb = p2_smul_28838_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72790_comb = p2_smul_28840_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72795_comb = p2_smul_28846_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72796_comb = p2_smul_28848_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72801_comb = p2_smul_28854_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72802_comb = p2_smul_28856_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72807_comb = p2_smul_28862_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72808_comb = p2_smul_28864_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72813_comb = p2_smul_28870_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72814_comb = p2_smul_28872_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72819_comb = p2_smul_28878_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72820_comb = p2_smul_28880_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_72839_comb = p2_smul_28902_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72848_comb = p2_smul_28912_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72853_comb = p2_smul_28918_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72862_comb = p2_smul_28928_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72867_comb = p2_smul_28934_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72876_comb = p2_smul_28944_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72881_comb = p2_smul_28950_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72890_comb = p2_smul_28960_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72895_comb = p2_smul_28966_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72904_comb = p2_smul_28976_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72909_comb = p2_smul_28982_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72918_comb = p2_smul_28992_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72923_comb = p2_smul_28998_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_72932_comb = p2_smul_29008_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73081_comb = p2_smul_29160_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73086_comb = p2_smul_29166_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73095_comb = p2_smul_29176_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73100_comb = p2_smul_29182_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73109_comb = p2_smul_29192_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73114_comb = p2_smul_29198_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73123_comb = p2_smul_29208_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73128_comb = p2_smul_29214_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73137_comb = p2_smul_29224_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73142_comb = p2_smul_29230_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73151_comb = p2_smul_29240_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73156_comb = p2_smul_29246_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73165_comb = p2_smul_29256_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73170_comb = p2_smul_29262_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73187_comb = p2_smul_29284_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73190_comb = p2_smul_29288_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73195_comb = p2_smul_29294_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73198_comb = p2_smul_29298_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73199_comb = p2_smul_29300_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73202_comb = p2_smul_29304_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73207_comb = p2_smul_29310_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73210_comb = p2_smul_29314_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73211_comb = p2_smul_29316_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73214_comb = p2_smul_29320_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73219_comb = p2_smul_29326_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73222_comb = p2_smul_29330_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73223_comb = p2_smul_29332_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73226_comb = p2_smul_29336_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73231_comb = p2_smul_29342_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73234_comb = p2_smul_29346_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73235_comb = p2_smul_29348_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73238_comb = p2_smul_29352_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73243_comb = p2_smul_29358_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73246_comb = p2_smul_29362_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73247_comb = p2_smul_29364_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73250_comb = p2_smul_29368_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73255_comb = p2_smul_29374_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73258_comb = p2_smul_29378_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73259_comb = p2_smul_29380_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73262_comb = p2_smul_29384_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73267_comb = p2_smul_29390_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73270_comb = p2_smul_29394_NarrowedMult__comb[18:6] + 13'h0001;
  assign p2_add_73285_comb = p2_smul_29412_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73298_comb = p2_smul_29426_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73299_comb = p2_smul_29428_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73312_comb = p2_smul_29442_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73313_comb = p2_smul_29444_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73326_comb = p2_smul_29458_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73327_comb = p2_smul_29460_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73340_comb = p2_smul_29474_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73341_comb = p2_smul_29476_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73354_comb = p2_smul_29490_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73355_comb = p2_smul_29492_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73368_comb = p2_smul_29506_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73369_comb = p2_smul_29508_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_add_73382_comb = p2_smul_29522_NarrowedMult__comb[17:6] + 12'h001;
  assign p2_sum__468_comb = p2_sum__464_comb + p2_sum__465_comb;
  assign p2_sum__469_comb = p2_sum__466_comb + p2_sum__467_comb;
  assign p2_sum__412_comb = p2_sum__408_comb + p2_sum__409_comb;
  assign p2_sum__413_comb = p2_sum__410_comb + p2_sum__411_comb;
  assign p2_sum__356_comb = p2_sum__352_comb + p2_sum__353_comb;
  assign p2_sum__357_comb = p2_sum__354_comb + p2_sum__355_comb;
  assign p2_sum__300_comb = p2_sum__296_comb + p2_sum__297_comb;
  assign p2_sum__301_comb = p2_sum__298_comb + p2_sum__299_comb;
  assign p2_sum__244_comb = p2_sum__240_comb + p2_sum__241_comb;
  assign p2_sum__245_comb = p2_sum__242_comb + p2_sum__243_comb;
  assign p2_sum__188_comb = p2_sum__184_comb + p2_sum__185_comb;
  assign p2_sum__189_comb = p2_sum__186_comb + p2_sum__187_comb;
  assign p2_sum__132_comb = p2_sum__128_comb + p2_sum__129_comb;
  assign p2_sum__133_comb = p2_sum__130_comb + p2_sum__131_comb;
  assign p2_add_74359_comb = p2_add_73415_comb[13:1] + p2_add_73416_comb[13:1];
  assign p2_add_74360_comb = p2_add_73417_comb[13:1] + {{2{p2_bit_slice_73418_comb[10]}}, p2_bit_slice_73418_comb};
  assign p2_add_74361_comb = {{2{p2_bit_slice_73419_comb[10]}}, p2_bit_slice_73419_comb} + p2_add_73420_comb[13:1];
  assign p2_add_74362_comb = p2_add_73421_comb[13:1] + p2_add_73422_comb[13:1];
  assign p2_add_74391_comb = p2_add_73479_comb[13:1] + {{1{p2_bit_slice_73480_comb[11]}}, p2_bit_slice_73480_comb};
  assign p2_add_74392_comb = {{1{p2_bit_slice_73481_comb[11]}}, p2_bit_slice_73481_comb} + p2_add_73482_comb[13:1];
  assign p2_add_74393_comb = p2_add_73483_comb[13:1] + {{1{p2_bit_slice_73484_comb[11]}}, p2_bit_slice_73484_comb};
  assign p2_add_74394_comb = {{1{p2_bit_slice_73485_comb[11]}}, p2_bit_slice_73485_comb} + p2_add_73486_comb[13:1];
  assign p2_add_74423_comb = p2_add_73543_comb[13:1] + {{2{p2_bit_slice_73544_comb[10]}}, p2_bit_slice_73544_comb};
  assign p2_add_74424_comb = p2_add_73545_comb[13:1] + p2_add_73546_comb[13:1];
  assign p2_add_74425_comb = p2_add_73547_comb[13:1] + p2_add_73548_comb[13:1];
  assign p2_add_74426_comb = {{2{p2_bit_slice_73549_comb[10]}}, p2_bit_slice_73549_comb} + p2_add_73550_comb[13:1];
  assign p2_add_74487_comb = p2_add_73671_comb[13:1] + p2_add_73672_comb[13:1];
  assign p2_add_74488_comb = {{2{p2_bit_slice_73673_comb[10]}}, p2_bit_slice_73673_comb} + p2_add_73674_comb[13:1];
  assign p2_add_74489_comb = p2_add_73675_comb[13:1] + {{2{p2_bit_slice_73676_comb[10]}}, p2_bit_slice_73676_comb};
  assign p2_add_74490_comb = p2_add_73677_comb[13:1] + p2_add_73678_comb[13:1];
  assign p2_add_74519_comb = {{1{p2_bit_slice_73735_comb[11]}}, p2_bit_slice_73735_comb} + p2_add_73736_comb[13:1];
  assign p2_add_74520_comb = {{1{p2_bit_slice_73737_comb[11]}}, p2_bit_slice_73737_comb} + p2_add_73738_comb[13:1];
  assign p2_add_74521_comb = p2_add_73739_comb[13:1] + {{1{p2_bit_slice_73740_comb[11]}}, p2_bit_slice_73740_comb};
  assign p2_add_74522_comb = p2_add_73741_comb[13:1] + {{1{p2_bit_slice_73742_comb[11]}}, p2_bit_slice_73742_comb};
  assign p2_add_74551_comb = {{2{p2_bit_slice_73799_comb[10]}}, p2_bit_slice_73799_comb} + p2_add_73800_comb[13:1];
  assign p2_add_74552_comb = p2_add_73801_comb[13:1] + p2_add_73802_comb[13:1];
  assign p2_add_74553_comb = p2_add_73803_comb[13:1] + p2_add_73804_comb[13:1];
  assign p2_add_74554_comb = p2_add_73805_comb[13:1] + {{2{p2_bit_slice_73806_comb[10]}}, p2_bit_slice_73806_comb};
  assign p2_sum__526_comb = p2_sum__524_comb + p2_sum__525_comb;
  assign p2_sum__1568_comb = {{12{p2_add_74455_comb[12]}}, p2_add_74455_comb};
  assign p2_sum__1569_comb = {{12{p2_add_74456_comb[12]}}, p2_add_74456_comb};
  assign p2_sum__1570_comb = {{12{p2_add_74457_comb[12]}}, p2_add_74457_comb};
  assign p2_sum__1571_comb = {{12{p2_add_74458_comb[12]}}, p2_add_74458_comb};
  assign p2_add_73423_comb = p2_smul_71985_comb[20:7] + 14'h0001;
  assign p2_add_73424_comb = p2_smul_71986_comb[20:7] + 14'h0001;
  assign p2_add_73425_comb = p2_smul_28648_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73426_comb = p2_add_72635_comb[11:1];
  assign p2_bit_slice_73427_comb = p2_add_72636_comb[11:1];
  assign p2_add_73428_comb = p2_smul_28654_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73429_comb = p2_smul_71993_comb[20:7] + 14'h0001;
  assign p2_add_73430_comb = p2_smul_71994_comb[20:7] + 14'h0001;
  assign p2_add_73431_comb = p2_smul_71995_comb[20:7] + 14'h0001;
  assign p2_add_73432_comb = p2_smul_71996_comb[20:7] + 14'h0001;
  assign p2_add_73433_comb = p2_smul_28664_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73434_comb = p2_add_72649_comb[11:1];
  assign p2_bit_slice_73435_comb = p2_add_72650_comb[11:1];
  assign p2_add_73436_comb = p2_smul_28670_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73437_comb = p2_smul_72003_comb[20:7] + 14'h0001;
  assign p2_add_73438_comb = p2_smul_72004_comb[20:7] + 14'h0001;
  assign p2_add_73439_comb = p2_smul_72005_comb[20:7] + 14'h0001;
  assign p2_add_73440_comb = p2_smul_72006_comb[20:7] + 14'h0001;
  assign p2_add_73441_comb = p2_smul_28680_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73442_comb = p2_add_72663_comb[11:1];
  assign p2_bit_slice_73443_comb = p2_add_72664_comb[11:1];
  assign p2_add_73444_comb = p2_smul_28686_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73445_comb = p2_smul_72013_comb[20:7] + 14'h0001;
  assign p2_add_73446_comb = p2_smul_72014_comb[20:7] + 14'h0001;
  assign p2_add_73447_comb = p2_smul_72015_comb[20:7] + 14'h0001;
  assign p2_add_73448_comb = p2_smul_72016_comb[20:7] + 14'h0001;
  assign p2_add_73449_comb = p2_smul_28696_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73450_comb = p2_add_72677_comb[11:1];
  assign p2_bit_slice_73451_comb = p2_add_72678_comb[11:1];
  assign p2_add_73452_comb = p2_smul_28702_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73453_comb = p2_smul_72023_comb[20:7] + 14'h0001;
  assign p2_add_73454_comb = p2_smul_72024_comb[20:7] + 14'h0001;
  assign p2_add_73455_comb = p2_smul_72025_comb[20:7] + 14'h0001;
  assign p2_add_73456_comb = p2_smul_72026_comb[20:7] + 14'h0001;
  assign p2_add_73457_comb = p2_smul_28712_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73458_comb = p2_add_72691_comb[11:1];
  assign p2_bit_slice_73459_comb = p2_add_72692_comb[11:1];
  assign p2_add_73460_comb = p2_smul_28718_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73461_comb = p2_smul_72033_comb[20:7] + 14'h0001;
  assign p2_add_73462_comb = p2_smul_72034_comb[20:7] + 14'h0001;
  assign p2_add_73463_comb = p2_smul_72035_comb[20:7] + 14'h0001;
  assign p2_add_73464_comb = p2_smul_72036_comb[20:7] + 14'h0001;
  assign p2_add_73465_comb = p2_smul_28728_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73466_comb = p2_add_72705_comb[11:1];
  assign p2_bit_slice_73467_comb = p2_add_72706_comb[11:1];
  assign p2_add_73468_comb = p2_smul_28734_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73469_comb = p2_smul_72043_comb[20:7] + 14'h0001;
  assign p2_add_73470_comb = p2_smul_72044_comb[20:7] + 14'h0001;
  assign p2_add_73471_comb = p2_smul_72045_comb[20:7] + 14'h0001;
  assign p2_add_73472_comb = p2_smul_72046_comb[20:7] + 14'h0001;
  assign p2_add_73473_comb = p2_smul_28744_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73474_comb = p2_add_72719_comb[11:1];
  assign p2_bit_slice_73475_comb = p2_add_72720_comb[11:1];
  assign p2_add_73476_comb = p2_smul_28750_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73477_comb = p2_smul_72053_comb[20:7] + 14'h0001;
  assign p2_add_73478_comb = p2_smul_72054_comb[20:7] + 14'h0001;
  assign p2_add_73487_comb = p2_smul_28772_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73488_comb = p2_add_72741_comb[12:1];
  assign p2_bit_slice_73489_comb = p2_add_72742_comb[12:1];
  assign p2_add_73490_comb = p2_smul_28778_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73491_comb = p2_smul_28780_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73492_comb = p2_add_72747_comb[12:1];
  assign p2_bit_slice_73493_comb = p2_add_72748_comb[12:1];
  assign p2_add_73494_comb = p2_smul_28786_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73495_comb = p2_smul_28788_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73496_comb = p2_add_72753_comb[12:1];
  assign p2_bit_slice_73497_comb = p2_add_72754_comb[12:1];
  assign p2_add_73498_comb = p2_smul_28794_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73499_comb = p2_smul_28796_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73500_comb = p2_add_72759_comb[12:1];
  assign p2_bit_slice_73501_comb = p2_add_72760_comb[12:1];
  assign p2_add_73502_comb = p2_smul_28802_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73503_comb = p2_smul_28804_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73504_comb = p2_add_72765_comb[12:1];
  assign p2_bit_slice_73505_comb = p2_add_72766_comb[12:1];
  assign p2_add_73506_comb = p2_smul_28810_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73507_comb = p2_smul_28812_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73508_comb = p2_add_72771_comb[12:1];
  assign p2_bit_slice_73509_comb = p2_add_72772_comb[12:1];
  assign p2_add_73510_comb = p2_smul_28818_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73511_comb = p2_smul_28820_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73512_comb = p2_add_72777_comb[12:1];
  assign p2_bit_slice_73513_comb = p2_add_72778_comb[12:1];
  assign p2_add_73514_comb = p2_smul_28826_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73515_comb = p2_smul_28828_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73516_comb = p2_add_72783_comb[12:1];
  assign p2_bit_slice_73517_comb = p2_add_72784_comb[12:1];
  assign p2_add_73518_comb = p2_smul_28834_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73519_comb = p2_smul_28836_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73520_comb = p2_add_72789_comb[12:1];
  assign p2_bit_slice_73521_comb = p2_add_72790_comb[12:1];
  assign p2_add_73522_comb = p2_smul_28842_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73523_comb = p2_smul_28844_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73524_comb = p2_add_72795_comb[12:1];
  assign p2_bit_slice_73525_comb = p2_add_72796_comb[12:1];
  assign p2_add_73526_comb = p2_smul_28850_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73527_comb = p2_smul_28852_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73528_comb = p2_add_72801_comb[12:1];
  assign p2_bit_slice_73529_comb = p2_add_72802_comb[12:1];
  assign p2_add_73530_comb = p2_smul_28858_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73531_comb = p2_smul_28860_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73532_comb = p2_add_72807_comb[12:1];
  assign p2_bit_slice_73533_comb = p2_add_72808_comb[12:1];
  assign p2_add_73534_comb = p2_smul_28866_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73535_comb = p2_smul_28868_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73536_comb = p2_add_72813_comb[12:1];
  assign p2_bit_slice_73537_comb = p2_add_72814_comb[12:1];
  assign p2_add_73538_comb = p2_smul_28874_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73539_comb = p2_smul_28876_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73540_comb = p2_add_72819_comb[12:1];
  assign p2_bit_slice_73541_comb = p2_add_72820_comb[12:1];
  assign p2_add_73542_comb = p2_smul_28882_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73551_comb = p2_smul_72161_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73552_comb = p2_add_72839_comb[11:1];
  assign p2_add_73553_comb = p2_smul_72164_comb[20:7] + 14'h0001;
  assign p2_add_73554_comb = p2_smul_28906_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73555_comb = p2_smul_28908_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73556_comb = p2_smul_72167_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73557_comb = p2_add_72848_comb[11:1];
  assign p2_add_73558_comb = p2_smul_72170_comb[20:7] + 14'h0001;
  assign p2_add_73559_comb = p2_smul_72171_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73560_comb = p2_add_72853_comb[11:1];
  assign p2_add_73561_comb = p2_smul_72174_comb[20:7] + 14'h0001;
  assign p2_add_73562_comb = p2_smul_28922_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73563_comb = p2_smul_28924_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73564_comb = p2_smul_72177_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73565_comb = p2_add_72862_comb[11:1];
  assign p2_add_73566_comb = p2_smul_72180_comb[20:7] + 14'h0001;
  assign p2_add_73567_comb = p2_smul_72181_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73568_comb = p2_add_72867_comb[11:1];
  assign p2_add_73569_comb = p2_smul_72184_comb[20:7] + 14'h0001;
  assign p2_add_73570_comb = p2_smul_28938_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73571_comb = p2_smul_28940_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73572_comb = p2_smul_72187_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73573_comb = p2_add_72876_comb[11:1];
  assign p2_add_73574_comb = p2_smul_72190_comb[20:7] + 14'h0001;
  assign p2_add_73575_comb = p2_smul_72191_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73576_comb = p2_add_72881_comb[11:1];
  assign p2_add_73577_comb = p2_smul_72194_comb[20:7] + 14'h0001;
  assign p2_add_73578_comb = p2_smul_28954_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73579_comb = p2_smul_28956_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73580_comb = p2_smul_72197_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73581_comb = p2_add_72890_comb[11:1];
  assign p2_add_73582_comb = p2_smul_72200_comb[20:7] + 14'h0001;
  assign p2_add_73583_comb = p2_smul_72201_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73584_comb = p2_add_72895_comb[11:1];
  assign p2_add_73585_comb = p2_smul_72204_comb[20:7] + 14'h0001;
  assign p2_add_73586_comb = p2_smul_28970_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73587_comb = p2_smul_28972_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73588_comb = p2_smul_72207_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73589_comb = p2_add_72904_comb[11:1];
  assign p2_add_73590_comb = p2_smul_72210_comb[20:7] + 14'h0001;
  assign p2_add_73591_comb = p2_smul_72211_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73592_comb = p2_add_72909_comb[11:1];
  assign p2_add_73593_comb = p2_smul_72214_comb[20:7] + 14'h0001;
  assign p2_add_73594_comb = p2_smul_28986_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73595_comb = p2_smul_28988_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73596_comb = p2_smul_72217_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73597_comb = p2_add_72918_comb[11:1];
  assign p2_add_73598_comb = p2_smul_72220_comb[20:7] + 14'h0001;
  assign p2_add_73599_comb = p2_smul_72221_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73600_comb = p2_add_72923_comb[11:1];
  assign p2_add_73601_comb = p2_smul_72224_comb[20:7] + 14'h0001;
  assign p2_add_73602_comb = p2_smul_29002_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73603_comb = p2_smul_29004_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73604_comb = p2_smul_72227_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73605_comb = p2_add_72932_comb[11:1];
  assign p2_add_73606_comb = p2_smul_72230_comb[20:7] + 14'h0001;
  assign p2_add_73679_comb = p2_smul_29156_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73680_comb = p2_smul_72306_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73681_comb = p2_add_73081_comb[11:1];
  assign p2_add_73682_comb = p2_smul_72309_comb[20:7] + 14'h0001;
  assign p2_add_73683_comb = p2_smul_72310_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73684_comb = p2_add_73086_comb[11:1];
  assign p2_add_73685_comb = p2_smul_72313_comb[20:7] + 14'h0001;
  assign p2_add_73686_comb = p2_smul_29170_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73687_comb = p2_smul_29172_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73688_comb = p2_smul_72316_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73689_comb = p2_add_73095_comb[11:1];
  assign p2_add_73690_comb = p2_smul_72319_comb[20:7] + 14'h0001;
  assign p2_add_73691_comb = p2_smul_72320_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73692_comb = p2_add_73100_comb[11:1];
  assign p2_add_73693_comb = p2_smul_72323_comb[20:7] + 14'h0001;
  assign p2_add_73694_comb = p2_smul_29186_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73695_comb = p2_smul_29188_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73696_comb = p2_smul_72326_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73697_comb = p2_add_73109_comb[11:1];
  assign p2_add_73698_comb = p2_smul_72329_comb[20:7] + 14'h0001;
  assign p2_add_73699_comb = p2_smul_72330_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73700_comb = p2_add_73114_comb[11:1];
  assign p2_add_73701_comb = p2_smul_72333_comb[20:7] + 14'h0001;
  assign p2_add_73702_comb = p2_smul_29202_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73703_comb = p2_smul_29204_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73704_comb = p2_smul_72336_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73705_comb = p2_add_73123_comb[11:1];
  assign p2_add_73706_comb = p2_smul_72339_comb[20:7] + 14'h0001;
  assign p2_add_73707_comb = p2_smul_72340_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73708_comb = p2_add_73128_comb[11:1];
  assign p2_add_73709_comb = p2_smul_72343_comb[20:7] + 14'h0001;
  assign p2_add_73710_comb = p2_smul_29218_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73711_comb = p2_smul_29220_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73712_comb = p2_smul_72346_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73713_comb = p2_add_73137_comb[11:1];
  assign p2_add_73714_comb = p2_smul_72349_comb[20:7] + 14'h0001;
  assign p2_add_73715_comb = p2_smul_72350_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73716_comb = p2_add_73142_comb[11:1];
  assign p2_add_73717_comb = p2_smul_72353_comb[20:7] + 14'h0001;
  assign p2_add_73718_comb = p2_smul_29234_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73719_comb = p2_smul_29236_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73720_comb = p2_smul_72356_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73721_comb = p2_add_73151_comb[11:1];
  assign p2_add_73722_comb = p2_smul_72359_comb[20:7] + 14'h0001;
  assign p2_add_73723_comb = p2_smul_72360_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73724_comb = p2_add_73156_comb[11:1];
  assign p2_add_73725_comb = p2_smul_72363_comb[20:7] + 14'h0001;
  assign p2_add_73726_comb = p2_smul_29250_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73727_comb = p2_smul_29252_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73728_comb = p2_smul_72366_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73729_comb = p2_add_73165_comb[11:1];
  assign p2_add_73730_comb = p2_smul_72369_comb[20:7] + 14'h0001;
  assign p2_add_73731_comb = p2_smul_72370_comb[20:7] + 14'h0001;
  assign p2_bit_slice_73732_comb = p2_add_73170_comb[11:1];
  assign p2_add_73733_comb = p2_smul_72373_comb[20:7] + 14'h0001;
  assign p2_add_73734_comb = p2_smul_29266_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73743_comb = p2_add_73187_comb[12:1];
  assign p2_add_73744_comb = p2_smul_29286_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73745_comb = p2_add_73190_comb[12:1];
  assign p2_add_73746_comb = p2_smul_29290_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73747_comb = p2_smul_29292_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73748_comb = p2_add_73195_comb[12:1];
  assign p2_add_73749_comb = p2_smul_29296_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73750_comb = p2_add_73198_comb[12:1];
  assign p2_bit_slice_73751_comb = p2_add_73199_comb[12:1];
  assign p2_add_73752_comb = p2_smul_29302_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73753_comb = p2_add_73202_comb[12:1];
  assign p2_add_73754_comb = p2_smul_29306_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73755_comb = p2_smul_29308_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73756_comb = p2_add_73207_comb[12:1];
  assign p2_add_73757_comb = p2_smul_29312_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73758_comb = p2_add_73210_comb[12:1];
  assign p2_bit_slice_73759_comb = p2_add_73211_comb[12:1];
  assign p2_add_73760_comb = p2_smul_29318_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73761_comb = p2_add_73214_comb[12:1];
  assign p2_add_73762_comb = p2_smul_29322_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73763_comb = p2_smul_29324_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73764_comb = p2_add_73219_comb[12:1];
  assign p2_add_73765_comb = p2_smul_29328_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73766_comb = p2_add_73222_comb[12:1];
  assign p2_bit_slice_73767_comb = p2_add_73223_comb[12:1];
  assign p2_add_73768_comb = p2_smul_29334_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73769_comb = p2_add_73226_comb[12:1];
  assign p2_add_73770_comb = p2_smul_29338_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73771_comb = p2_smul_29340_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73772_comb = p2_add_73231_comb[12:1];
  assign p2_add_73773_comb = p2_smul_29344_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73774_comb = p2_add_73234_comb[12:1];
  assign p2_bit_slice_73775_comb = p2_add_73235_comb[12:1];
  assign p2_add_73776_comb = p2_smul_29350_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73777_comb = p2_add_73238_comb[12:1];
  assign p2_add_73778_comb = p2_smul_29354_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73779_comb = p2_smul_29356_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73780_comb = p2_add_73243_comb[12:1];
  assign p2_add_73781_comb = p2_smul_29360_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73782_comb = p2_add_73246_comb[12:1];
  assign p2_bit_slice_73783_comb = p2_add_73247_comb[12:1];
  assign p2_add_73784_comb = p2_smul_29366_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73785_comb = p2_add_73250_comb[12:1];
  assign p2_add_73786_comb = p2_smul_29370_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73787_comb = p2_smul_29372_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73788_comb = p2_add_73255_comb[12:1];
  assign p2_add_73789_comb = p2_smul_29376_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73790_comb = p2_add_73258_comb[12:1];
  assign p2_bit_slice_73791_comb = p2_add_73259_comb[12:1];
  assign p2_add_73792_comb = p2_smul_29382_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73793_comb = p2_add_73262_comb[12:1];
  assign p2_add_73794_comb = p2_smul_29386_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_add_73795_comb = p2_smul_29388_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73796_comb = p2_add_73267_comb[12:1];
  assign p2_add_73797_comb = p2_smul_29392_NarrowedMult__comb[18:5] + 14'h0001;
  assign p2_bit_slice_73798_comb = p2_add_73270_comb[12:1];
  assign p2_bit_slice_73807_comb = p2_add_73285_comb[11:1];
  assign p2_add_73808_comb = p2_smul_29414_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73809_comb = p2_smul_72484_comb[20:7] + 14'h0001;
  assign p2_add_73810_comb = p2_smul_72485_comb[20:7] + 14'h0001;
  assign p2_add_73811_comb = p2_smul_72486_comb[20:7] + 14'h0001;
  assign p2_add_73812_comb = p2_smul_72487_comb[20:7] + 14'h0001;
  assign p2_add_73813_comb = p2_smul_29424_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73814_comb = p2_add_73298_comb[11:1];
  assign p2_bit_slice_73815_comb = p2_add_73299_comb[11:1];
  assign p2_add_73816_comb = p2_smul_29430_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73817_comb = p2_smul_72494_comb[20:7] + 14'h0001;
  assign p2_add_73818_comb = p2_smul_72495_comb[20:7] + 14'h0001;
  assign p2_add_73819_comb = p2_smul_72496_comb[20:7] + 14'h0001;
  assign p2_add_73820_comb = p2_smul_72497_comb[20:7] + 14'h0001;
  assign p2_add_73821_comb = p2_smul_29440_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73822_comb = p2_add_73312_comb[11:1];
  assign p2_bit_slice_73823_comb = p2_add_73313_comb[11:1];
  assign p2_add_73824_comb = p2_smul_29446_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73825_comb = p2_smul_72504_comb[20:7] + 14'h0001;
  assign p2_add_73826_comb = p2_smul_72505_comb[20:7] + 14'h0001;
  assign p2_add_73827_comb = p2_smul_72506_comb[20:7] + 14'h0001;
  assign p2_add_73828_comb = p2_smul_72507_comb[20:7] + 14'h0001;
  assign p2_add_73829_comb = p2_smul_29456_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73830_comb = p2_add_73326_comb[11:1];
  assign p2_bit_slice_73831_comb = p2_add_73327_comb[11:1];
  assign p2_add_73832_comb = p2_smul_29462_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73833_comb = p2_smul_72514_comb[20:7] + 14'h0001;
  assign p2_add_73834_comb = p2_smul_72515_comb[20:7] + 14'h0001;
  assign p2_add_73835_comb = p2_smul_72516_comb[20:7] + 14'h0001;
  assign p2_add_73836_comb = p2_smul_72517_comb[20:7] + 14'h0001;
  assign p2_add_73837_comb = p2_smul_29472_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73838_comb = p2_add_73340_comb[11:1];
  assign p2_bit_slice_73839_comb = p2_add_73341_comb[11:1];
  assign p2_add_73840_comb = p2_smul_29478_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73841_comb = p2_smul_72524_comb[20:7] + 14'h0001;
  assign p2_add_73842_comb = p2_smul_72525_comb[20:7] + 14'h0001;
  assign p2_add_73843_comb = p2_smul_72526_comb[20:7] + 14'h0001;
  assign p2_add_73844_comb = p2_smul_72527_comb[20:7] + 14'h0001;
  assign p2_add_73845_comb = p2_smul_29488_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73846_comb = p2_add_73354_comb[11:1];
  assign p2_bit_slice_73847_comb = p2_add_73355_comb[11:1];
  assign p2_add_73848_comb = p2_smul_29494_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73849_comb = p2_smul_72534_comb[20:7] + 14'h0001;
  assign p2_add_73850_comb = p2_smul_72535_comb[20:7] + 14'h0001;
  assign p2_add_73851_comb = p2_smul_72536_comb[20:7] + 14'h0001;
  assign p2_add_73852_comb = p2_smul_72537_comb[20:7] + 14'h0001;
  assign p2_add_73853_comb = p2_smul_29504_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73854_comb = p2_add_73368_comb[11:1];
  assign p2_bit_slice_73855_comb = p2_add_73369_comb[11:1];
  assign p2_add_73856_comb = p2_smul_29510_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_add_73857_comb = p2_smul_72544_comb[20:7] + 14'h0001;
  assign p2_add_73858_comb = p2_smul_72545_comb[20:7] + 14'h0001;
  assign p2_add_73859_comb = p2_smul_72546_comb[20:7] + 14'h0001;
  assign p2_add_73860_comb = p2_smul_72547_comb[20:7] + 14'h0001;
  assign p2_add_73861_comb = p2_smul_29520_NarrowedMult__comb[19:6] + 14'h0001;
  assign p2_bit_slice_73862_comb = p2_add_73382_comb[11:1];
  assign p2_add_74459_comb = p2_add_73615_comb[13:1] + p2_add_73616_comb[13:1];
  assign p2_add_74460_comb = p2_add_73617_comb[13:1] + p2_add_73618_comb[13:1];
  assign p2_add_74461_comb = p2_add_73619_comb[13:1] + p2_add_73620_comb[13:1];
  assign p2_add_74462_comb = p2_add_73621_comb[13:1] + p2_add_73622_comb[13:1];
  assign p2_add_74463_comb = p2_add_73623_comb[13:1] + p2_add_73624_comb[13:1];
  assign p2_add_74464_comb = p2_add_73625_comb[13:1] + p2_add_73626_comb[13:1];
  assign p2_add_74465_comb = p2_add_73627_comb[13:1] + p2_add_73628_comb[13:1];
  assign p2_add_74466_comb = p2_add_73629_comb[13:1] + p2_add_73630_comb[13:1];
  assign p2_add_74467_comb = p2_add_73631_comb[13:1] + p2_add_73632_comb[13:1];
  assign p2_add_74468_comb = p2_add_73633_comb[13:1] + p2_add_73634_comb[13:1];
  assign p2_add_74469_comb = p2_add_73635_comb[13:1] + p2_add_73636_comb[13:1];
  assign p2_add_74470_comb = p2_add_73637_comb[13:1] + p2_add_73638_comb[13:1];
  assign p2_add_74471_comb = p2_add_73639_comb[13:1] + p2_add_73640_comb[13:1];
  assign p2_add_74472_comb = p2_add_73641_comb[13:1] + p2_add_73642_comb[13:1];
  assign p2_add_74473_comb = p2_add_73643_comb[13:1] + p2_add_73644_comb[13:1];
  assign p2_add_74474_comb = p2_add_73645_comb[13:1] + p2_add_73646_comb[13:1];
  assign p2_add_74475_comb = p2_add_73647_comb[13:1] + p2_add_73648_comb[13:1];
  assign p2_add_74476_comb = p2_add_73649_comb[13:1] + p2_add_73650_comb[13:1];
  assign p2_add_74477_comb = p2_add_73651_comb[13:1] + p2_add_73652_comb[13:1];
  assign p2_add_74478_comb = p2_add_73653_comb[13:1] + p2_add_73654_comb[13:1];
  assign p2_add_74479_comb = p2_add_73655_comb[13:1] + p2_add_73656_comb[13:1];
  assign p2_add_74480_comb = p2_add_73657_comb[13:1] + p2_add_73658_comb[13:1];
  assign p2_add_74481_comb = p2_add_73659_comb[13:1] + p2_add_73660_comb[13:1];
  assign p2_add_74482_comb = p2_add_73661_comb[13:1] + p2_add_73662_comb[13:1];
  assign p2_add_74483_comb = p2_add_73663_comb[13:1] + p2_add_73664_comb[13:1];
  assign p2_add_74484_comb = p2_add_73665_comb[13:1] + p2_add_73666_comb[13:1];
  assign p2_add_74485_comb = p2_add_73667_comb[13:1] + p2_add_73668_comb[13:1];
  assign p2_add_74486_comb = p2_add_73669_comb[13:1] + p2_add_73670_comb[13:1];
  assign p2_sum__470_comb = p2_sum__468_comb + p2_sum__469_comb;
  assign p2_sum__414_comb = p2_sum__412_comb + p2_sum__413_comb;
  assign p2_sum__358_comb = p2_sum__356_comb + p2_sum__357_comb;
  assign p2_sum__302_comb = p2_sum__300_comb + p2_sum__301_comb;
  assign p2_sum__246_comb = p2_sum__244_comb + p2_sum__245_comb;
  assign p2_sum__190_comb = p2_sum__188_comb + p2_sum__189_comb;
  assign p2_sum__134_comb = p2_sum__132_comb + p2_sum__133_comb;
  assign p2_sum__1580_comb = {{12{p2_add_74359_comb[12]}}, p2_add_74359_comb};
  assign p2_sum__1581_comb = {{12{p2_add_74360_comb[12]}}, p2_add_74360_comb};
  assign p2_sum__1582_comb = {{12{p2_add_74361_comb[12]}}, p2_add_74361_comb};
  assign p2_sum__1583_comb = {{12{p2_add_74362_comb[12]}}, p2_add_74362_comb};
  assign p2_sum__1576_comb = {{12{p2_add_74391_comb[12]}}, p2_add_74391_comb};
  assign p2_sum__1577_comb = {{12{p2_add_74392_comb[12]}}, p2_add_74392_comb};
  assign p2_sum__1578_comb = {{12{p2_add_74393_comb[12]}}, p2_add_74393_comb};
  assign p2_sum__1579_comb = {{12{p2_add_74394_comb[12]}}, p2_add_74394_comb};
  assign p2_sum__1572_comb = {{12{p2_add_74423_comb[12]}}, p2_add_74423_comb};
  assign p2_sum__1573_comb = {{12{p2_add_74424_comb[12]}}, p2_add_74424_comb};
  assign p2_sum__1574_comb = {{12{p2_add_74425_comb[12]}}, p2_add_74425_comb};
  assign p2_sum__1575_comb = {{12{p2_add_74426_comb[12]}}, p2_add_74426_comb};
  assign p2_sum__1564_comb = {{12{p2_add_74487_comb[12]}}, p2_add_74487_comb};
  assign p2_sum__1565_comb = {{12{p2_add_74488_comb[12]}}, p2_add_74488_comb};
  assign p2_sum__1566_comb = {{12{p2_add_74489_comb[12]}}, p2_add_74489_comb};
  assign p2_sum__1567_comb = {{12{p2_add_74490_comb[12]}}, p2_add_74490_comb};
  assign p2_sum__1560_comb = {{12{p2_add_74519_comb[12]}}, p2_add_74519_comb};
  assign p2_sum__1561_comb = {{12{p2_add_74520_comb[12]}}, p2_add_74520_comb};
  assign p2_sum__1562_comb = {{12{p2_add_74521_comb[12]}}, p2_add_74521_comb};
  assign p2_sum__1563_comb = {{12{p2_add_74522_comb[12]}}, p2_add_74522_comb};
  assign p2_sum__1556_comb = {{12{p2_add_74551_comb[12]}}, p2_add_74551_comb};
  assign p2_sum__1557_comb = {{12{p2_add_74552_comb[12]}}, p2_add_74552_comb};
  assign p2_sum__1558_comb = {{12{p2_add_74553_comb[12]}}, p2_add_74553_comb};
  assign p2_sum__1559_comb = {{12{p2_add_74554_comb[12]}}, p2_add_74554_comb};
  assign p2_umul_74655_comb = umul32b_32b_x_7b(p2_sum__526_comb, 7'h5b);
  assign p2_sum__1240_comb = p2_sum__1568_comb + p2_sum__1569_comb;
  assign p2_sum__1241_comb = p2_sum__1570_comb + p2_sum__1571_comb;
  assign p2_sum__1540_comb = {{12{p2_add_74459_comb[12]}}, p2_add_74459_comb};
  assign p2_sum__1541_comb = {{12{p2_add_74460_comb[12]}}, p2_add_74460_comb};
  assign p2_sum__1542_comb = {{12{p2_add_74461_comb[12]}}, p2_add_74461_comb};
  assign p2_sum__1543_comb = {{12{p2_add_74462_comb[12]}}, p2_add_74462_comb};
  assign p2_sum__1512_comb = {{12{p2_add_74463_comb[12]}}, p2_add_74463_comb};
  assign p2_sum__1513_comb = {{12{p2_add_74464_comb[12]}}, p2_add_74464_comb};
  assign p2_sum__1514_comb = {{12{p2_add_74465_comb[12]}}, p2_add_74465_comb};
  assign p2_sum__1515_comb = {{12{p2_add_74466_comb[12]}}, p2_add_74466_comb};
  assign p2_sum__1484_comb = {{12{p2_add_74467_comb[12]}}, p2_add_74467_comb};
  assign p2_sum__1485_comb = {{12{p2_add_74468_comb[12]}}, p2_add_74468_comb};
  assign p2_sum__1486_comb = {{12{p2_add_74469_comb[12]}}, p2_add_74469_comb};
  assign p2_sum__1487_comb = {{12{p2_add_74470_comb[12]}}, p2_add_74470_comb};
  assign p2_sum__1456_comb = {{12{p2_add_74471_comb[12]}}, p2_add_74471_comb};
  assign p2_sum__1457_comb = {{12{p2_add_74472_comb[12]}}, p2_add_74472_comb};
  assign p2_sum__1458_comb = {{12{p2_add_74473_comb[12]}}, p2_add_74473_comb};
  assign p2_sum__1459_comb = {{12{p2_add_74474_comb[12]}}, p2_add_74474_comb};
  assign p2_sum__1428_comb = {{12{p2_add_74475_comb[12]}}, p2_add_74475_comb};
  assign p2_sum__1429_comb = {{12{p2_add_74476_comb[12]}}, p2_add_74476_comb};
  assign p2_sum__1430_comb = {{12{p2_add_74477_comb[12]}}, p2_add_74477_comb};
  assign p2_sum__1431_comb = {{12{p2_add_74478_comb[12]}}, p2_add_74478_comb};
  assign p2_sum__1400_comb = {{12{p2_add_74479_comb[12]}}, p2_add_74479_comb};
  assign p2_sum__1401_comb = {{12{p2_add_74480_comb[12]}}, p2_add_74480_comb};
  assign p2_sum__1402_comb = {{12{p2_add_74481_comb[12]}}, p2_add_74481_comb};
  assign p2_sum__1403_comb = {{12{p2_add_74482_comb[12]}}, p2_add_74482_comb};
  assign p2_sum__1372_comb = {{12{p2_add_74483_comb[12]}}, p2_add_74483_comb};
  assign p2_sum__1373_comb = {{12{p2_add_74484_comb[12]}}, p2_add_74484_comb};
  assign p2_sum__1374_comb = {{12{p2_add_74485_comb[12]}}, p2_add_74485_comb};
  assign p2_sum__1375_comb = {{12{p2_add_74486_comb[12]}}, p2_add_74486_comb};
  assign p2_umul_74656_comb = umul32b_32b_x_7b(p2_sum__470_comb, 7'h5b);
  assign p2_umul_74657_comb = umul32b_32b_x_7b(p2_sum__414_comb, 7'h5b);
  assign p2_umul_74658_comb = umul32b_32b_x_7b(p2_sum__358_comb, 7'h5b);
  assign p2_umul_74659_comb = umul32b_32b_x_7b(p2_sum__302_comb, 7'h5b);
  assign p2_umul_74660_comb = umul32b_32b_x_7b(p2_sum__246_comb, 7'h5b);
  assign p2_umul_74661_comb = umul32b_32b_x_7b(p2_sum__190_comb, 7'h5b);
  assign p2_umul_74662_comb = umul32b_32b_x_7b(p2_sum__134_comb, 7'h5b);
  assign p2_sum__1246_comb = p2_sum__1580_comb + p2_sum__1581_comb;
  assign p2_sum__1247_comb = p2_sum__1582_comb + p2_sum__1583_comb;
  assign p2_sum__1244_comb = p2_sum__1576_comb + p2_sum__1577_comb;
  assign p2_sum__1245_comb = p2_sum__1578_comb + p2_sum__1579_comb;
  assign p2_sum__1242_comb = p2_sum__1572_comb + p2_sum__1573_comb;
  assign p2_sum__1243_comb = p2_sum__1574_comb + p2_sum__1575_comb;
  assign p2_sum__1238_comb = p2_sum__1564_comb + p2_sum__1565_comb;
  assign p2_sum__1239_comb = p2_sum__1566_comb + p2_sum__1567_comb;
  assign p2_sum__1236_comb = p2_sum__1560_comb + p2_sum__1561_comb;
  assign p2_sum__1237_comb = p2_sum__1562_comb + p2_sum__1563_comb;
  assign p2_sum__1234_comb = p2_sum__1556_comb + p2_sum__1557_comb;
  assign p2_sum__1235_comb = p2_sum__1558_comb + p2_sum__1559_comb;
  assign p2_sum__1076_comb = p2_sum__1240_comb + p2_sum__1241_comb;
  assign p2_add_74363_comb = p2_add_73423_comb[13:1] + p2_add_73424_comb[13:1];
  assign p2_add_74364_comb = p2_add_73425_comb[13:1] + {{2{p2_bit_slice_73426_comb[10]}}, p2_bit_slice_73426_comb};
  assign p2_add_74365_comb = {{2{p2_bit_slice_73427_comb[10]}}, p2_bit_slice_73427_comb} + p2_add_73428_comb[13:1];
  assign p2_add_74366_comb = p2_add_73429_comb[13:1] + p2_add_73430_comb[13:1];
  assign p2_add_74367_comb = p2_add_73431_comb[13:1] + p2_add_73432_comb[13:1];
  assign p2_add_74368_comb = p2_add_73433_comb[13:1] + {{2{p2_bit_slice_73434_comb[10]}}, p2_bit_slice_73434_comb};
  assign p2_add_74369_comb = {{2{p2_bit_slice_73435_comb[10]}}, p2_bit_slice_73435_comb} + p2_add_73436_comb[13:1];
  assign p2_add_74370_comb = p2_add_73437_comb[13:1] + p2_add_73438_comb[13:1];
  assign p2_add_74371_comb = p2_add_73439_comb[13:1] + p2_add_73440_comb[13:1];
  assign p2_add_74372_comb = p2_add_73441_comb[13:1] + {{2{p2_bit_slice_73442_comb[10]}}, p2_bit_slice_73442_comb};
  assign p2_add_74373_comb = {{2{p2_bit_slice_73443_comb[10]}}, p2_bit_slice_73443_comb} + p2_add_73444_comb[13:1];
  assign p2_add_74374_comb = p2_add_73445_comb[13:1] + p2_add_73446_comb[13:1];
  assign p2_add_74375_comb = p2_add_73447_comb[13:1] + p2_add_73448_comb[13:1];
  assign p2_add_74376_comb = p2_add_73449_comb[13:1] + {{2{p2_bit_slice_73450_comb[10]}}, p2_bit_slice_73450_comb};
  assign p2_add_74377_comb = {{2{p2_bit_slice_73451_comb[10]}}, p2_bit_slice_73451_comb} + p2_add_73452_comb[13:1];
  assign p2_add_74378_comb = p2_add_73453_comb[13:1] + p2_add_73454_comb[13:1];
  assign p2_add_74379_comb = p2_add_73455_comb[13:1] + p2_add_73456_comb[13:1];
  assign p2_add_74380_comb = p2_add_73457_comb[13:1] + {{2{p2_bit_slice_73458_comb[10]}}, p2_bit_slice_73458_comb};
  assign p2_add_74381_comb = {{2{p2_bit_slice_73459_comb[10]}}, p2_bit_slice_73459_comb} + p2_add_73460_comb[13:1];
  assign p2_add_74382_comb = p2_add_73461_comb[13:1] + p2_add_73462_comb[13:1];
  assign p2_add_74383_comb = p2_add_73463_comb[13:1] + p2_add_73464_comb[13:1];
  assign p2_add_74384_comb = p2_add_73465_comb[13:1] + {{2{p2_bit_slice_73466_comb[10]}}, p2_bit_slice_73466_comb};
  assign p2_add_74385_comb = {{2{p2_bit_slice_73467_comb[10]}}, p2_bit_slice_73467_comb} + p2_add_73468_comb[13:1];
  assign p2_add_74386_comb = p2_add_73469_comb[13:1] + p2_add_73470_comb[13:1];
  assign p2_add_74387_comb = p2_add_73471_comb[13:1] + p2_add_73472_comb[13:1];
  assign p2_add_74388_comb = p2_add_73473_comb[13:1] + {{2{p2_bit_slice_73474_comb[10]}}, p2_bit_slice_73474_comb};
  assign p2_add_74389_comb = {{2{p2_bit_slice_73475_comb[10]}}, p2_bit_slice_73475_comb} + p2_add_73476_comb[13:1];
  assign p2_add_74390_comb = p2_add_73477_comb[13:1] + p2_add_73478_comb[13:1];
  assign p2_add_74395_comb = p2_add_73487_comb[13:1] + {{1{p2_bit_slice_73488_comb[11]}}, p2_bit_slice_73488_comb};
  assign p2_add_74396_comb = {{1{p2_bit_slice_73489_comb[11]}}, p2_bit_slice_73489_comb} + p2_add_73490_comb[13:1];
  assign p2_add_74397_comb = p2_add_73491_comb[13:1] + {{1{p2_bit_slice_73492_comb[11]}}, p2_bit_slice_73492_comb};
  assign p2_add_74398_comb = {{1{p2_bit_slice_73493_comb[11]}}, p2_bit_slice_73493_comb} + p2_add_73494_comb[13:1];
  assign p2_add_74399_comb = p2_add_73495_comb[13:1] + {{1{p2_bit_slice_73496_comb[11]}}, p2_bit_slice_73496_comb};
  assign p2_add_74400_comb = {{1{p2_bit_slice_73497_comb[11]}}, p2_bit_slice_73497_comb} + p2_add_73498_comb[13:1];
  assign p2_add_74401_comb = p2_add_73499_comb[13:1] + {{1{p2_bit_slice_73500_comb[11]}}, p2_bit_slice_73500_comb};
  assign p2_add_74402_comb = {{1{p2_bit_slice_73501_comb[11]}}, p2_bit_slice_73501_comb} + p2_add_73502_comb[13:1];
  assign p2_add_74403_comb = p2_add_73503_comb[13:1] + {{1{p2_bit_slice_73504_comb[11]}}, p2_bit_slice_73504_comb};
  assign p2_add_74404_comb = {{1{p2_bit_slice_73505_comb[11]}}, p2_bit_slice_73505_comb} + p2_add_73506_comb[13:1];
  assign p2_add_74405_comb = p2_add_73507_comb[13:1] + {{1{p2_bit_slice_73508_comb[11]}}, p2_bit_slice_73508_comb};
  assign p2_add_74406_comb = {{1{p2_bit_slice_73509_comb[11]}}, p2_bit_slice_73509_comb} + p2_add_73510_comb[13:1];
  assign p2_add_74407_comb = p2_add_73511_comb[13:1] + {{1{p2_bit_slice_73512_comb[11]}}, p2_bit_slice_73512_comb};
  assign p2_add_74408_comb = {{1{p2_bit_slice_73513_comb[11]}}, p2_bit_slice_73513_comb} + p2_add_73514_comb[13:1];
  assign p2_add_74409_comb = p2_add_73515_comb[13:1] + {{1{p2_bit_slice_73516_comb[11]}}, p2_bit_slice_73516_comb};
  assign p2_add_74410_comb = {{1{p2_bit_slice_73517_comb[11]}}, p2_bit_slice_73517_comb} + p2_add_73518_comb[13:1];
  assign p2_add_74411_comb = p2_add_73519_comb[13:1] + {{1{p2_bit_slice_73520_comb[11]}}, p2_bit_slice_73520_comb};
  assign p2_add_74412_comb = {{1{p2_bit_slice_73521_comb[11]}}, p2_bit_slice_73521_comb} + p2_add_73522_comb[13:1];
  assign p2_add_74413_comb = p2_add_73523_comb[13:1] + {{1{p2_bit_slice_73524_comb[11]}}, p2_bit_slice_73524_comb};
  assign p2_add_74414_comb = {{1{p2_bit_slice_73525_comb[11]}}, p2_bit_slice_73525_comb} + p2_add_73526_comb[13:1];
  assign p2_add_74415_comb = p2_add_73527_comb[13:1] + {{1{p2_bit_slice_73528_comb[11]}}, p2_bit_slice_73528_comb};
  assign p2_add_74416_comb = {{1{p2_bit_slice_73529_comb[11]}}, p2_bit_slice_73529_comb} + p2_add_73530_comb[13:1];
  assign p2_add_74417_comb = p2_add_73531_comb[13:1] + {{1{p2_bit_slice_73532_comb[11]}}, p2_bit_slice_73532_comb};
  assign p2_add_74418_comb = {{1{p2_bit_slice_73533_comb[11]}}, p2_bit_slice_73533_comb} + p2_add_73534_comb[13:1];
  assign p2_add_74419_comb = p2_add_73535_comb[13:1] + {{1{p2_bit_slice_73536_comb[11]}}, p2_bit_slice_73536_comb};
  assign p2_add_74420_comb = {{1{p2_bit_slice_73537_comb[11]}}, p2_bit_slice_73537_comb} + p2_add_73538_comb[13:1];
  assign p2_add_74421_comb = p2_add_73539_comb[13:1] + {{1{p2_bit_slice_73540_comb[11]}}, p2_bit_slice_73540_comb};
  assign p2_add_74422_comb = {{1{p2_bit_slice_73541_comb[11]}}, p2_bit_slice_73541_comb} + p2_add_73542_comb[13:1];
  assign p2_add_74427_comb = p2_add_73551_comb[13:1] + {{2{p2_bit_slice_73552_comb[10]}}, p2_bit_slice_73552_comb};
  assign p2_add_74428_comb = p2_add_73553_comb[13:1] + p2_add_73554_comb[13:1];
  assign p2_add_74429_comb = p2_add_73555_comb[13:1] + p2_add_73556_comb[13:1];
  assign p2_add_74430_comb = {{2{p2_bit_slice_73557_comb[10]}}, p2_bit_slice_73557_comb} + p2_add_73558_comb[13:1];
  assign p2_add_74431_comb = p2_add_73559_comb[13:1] + {{2{p2_bit_slice_73560_comb[10]}}, p2_bit_slice_73560_comb};
  assign p2_add_74432_comb = p2_add_73561_comb[13:1] + p2_add_73562_comb[13:1];
  assign p2_add_74433_comb = p2_add_73563_comb[13:1] + p2_add_73564_comb[13:1];
  assign p2_add_74434_comb = {{2{p2_bit_slice_73565_comb[10]}}, p2_bit_slice_73565_comb} + p2_add_73566_comb[13:1];
  assign p2_add_74435_comb = p2_add_73567_comb[13:1] + {{2{p2_bit_slice_73568_comb[10]}}, p2_bit_slice_73568_comb};
  assign p2_add_74436_comb = p2_add_73569_comb[13:1] + p2_add_73570_comb[13:1];
  assign p2_add_74437_comb = p2_add_73571_comb[13:1] + p2_add_73572_comb[13:1];
  assign p2_add_74438_comb = {{2{p2_bit_slice_73573_comb[10]}}, p2_bit_slice_73573_comb} + p2_add_73574_comb[13:1];
  assign p2_add_74439_comb = p2_add_73575_comb[13:1] + {{2{p2_bit_slice_73576_comb[10]}}, p2_bit_slice_73576_comb};
  assign p2_add_74440_comb = p2_add_73577_comb[13:1] + p2_add_73578_comb[13:1];
  assign p2_add_74441_comb = p2_add_73579_comb[13:1] + p2_add_73580_comb[13:1];
  assign p2_add_74442_comb = {{2{p2_bit_slice_73581_comb[10]}}, p2_bit_slice_73581_comb} + p2_add_73582_comb[13:1];
  assign p2_add_74443_comb = p2_add_73583_comb[13:1] + {{2{p2_bit_slice_73584_comb[10]}}, p2_bit_slice_73584_comb};
  assign p2_add_74444_comb = p2_add_73585_comb[13:1] + p2_add_73586_comb[13:1];
  assign p2_add_74445_comb = p2_add_73587_comb[13:1] + p2_add_73588_comb[13:1];
  assign p2_add_74446_comb = {{2{p2_bit_slice_73589_comb[10]}}, p2_bit_slice_73589_comb} + p2_add_73590_comb[13:1];
  assign p2_add_74447_comb = p2_add_73591_comb[13:1] + {{2{p2_bit_slice_73592_comb[10]}}, p2_bit_slice_73592_comb};
  assign p2_add_74448_comb = p2_add_73593_comb[13:1] + p2_add_73594_comb[13:1];
  assign p2_add_74449_comb = p2_add_73595_comb[13:1] + p2_add_73596_comb[13:1];
  assign p2_add_74450_comb = {{2{p2_bit_slice_73597_comb[10]}}, p2_bit_slice_73597_comb} + p2_add_73598_comb[13:1];
  assign p2_add_74451_comb = p2_add_73599_comb[13:1] + {{2{p2_bit_slice_73600_comb[10]}}, p2_bit_slice_73600_comb};
  assign p2_add_74452_comb = p2_add_73601_comb[13:1] + p2_add_73602_comb[13:1];
  assign p2_add_74453_comb = p2_add_73603_comb[13:1] + p2_add_73604_comb[13:1];
  assign p2_add_74454_comb = {{2{p2_bit_slice_73605_comb[10]}}, p2_bit_slice_73605_comb} + p2_add_73606_comb[13:1];
  assign p2_add_74491_comb = p2_add_73679_comb[13:1] + p2_add_73680_comb[13:1];
  assign p2_add_74492_comb = {{2{p2_bit_slice_73681_comb[10]}}, p2_bit_slice_73681_comb} + p2_add_73682_comb[13:1];
  assign p2_add_74493_comb = p2_add_73683_comb[13:1] + {{2{p2_bit_slice_73684_comb[10]}}, p2_bit_slice_73684_comb};
  assign p2_add_74494_comb = p2_add_73685_comb[13:1] + p2_add_73686_comb[13:1];
  assign p2_add_74495_comb = p2_add_73687_comb[13:1] + p2_add_73688_comb[13:1];
  assign p2_add_74496_comb = {{2{p2_bit_slice_73689_comb[10]}}, p2_bit_slice_73689_comb} + p2_add_73690_comb[13:1];
  assign p2_add_74497_comb = p2_add_73691_comb[13:1] + {{2{p2_bit_slice_73692_comb[10]}}, p2_bit_slice_73692_comb};
  assign p2_add_74498_comb = p2_add_73693_comb[13:1] + p2_add_73694_comb[13:1];
  assign p2_add_74499_comb = p2_add_73695_comb[13:1] + p2_add_73696_comb[13:1];
  assign p2_add_74500_comb = {{2{p2_bit_slice_73697_comb[10]}}, p2_bit_slice_73697_comb} + p2_add_73698_comb[13:1];
  assign p2_add_74501_comb = p2_add_73699_comb[13:1] + {{2{p2_bit_slice_73700_comb[10]}}, p2_bit_slice_73700_comb};
  assign p2_add_74502_comb = p2_add_73701_comb[13:1] + p2_add_73702_comb[13:1];
  assign p2_add_74503_comb = p2_add_73703_comb[13:1] + p2_add_73704_comb[13:1];
  assign p2_add_74504_comb = {{2{p2_bit_slice_73705_comb[10]}}, p2_bit_slice_73705_comb} + p2_add_73706_comb[13:1];
  assign p2_add_74505_comb = p2_add_73707_comb[13:1] + {{2{p2_bit_slice_73708_comb[10]}}, p2_bit_slice_73708_comb};
  assign p2_add_74506_comb = p2_add_73709_comb[13:1] + p2_add_73710_comb[13:1];
  assign p2_add_74507_comb = p2_add_73711_comb[13:1] + p2_add_73712_comb[13:1];
  assign p2_add_74508_comb = {{2{p2_bit_slice_73713_comb[10]}}, p2_bit_slice_73713_comb} + p2_add_73714_comb[13:1];
  assign p2_add_74509_comb = p2_add_73715_comb[13:1] + {{2{p2_bit_slice_73716_comb[10]}}, p2_bit_slice_73716_comb};
  assign p2_add_74510_comb = p2_add_73717_comb[13:1] + p2_add_73718_comb[13:1];
  assign p2_add_74511_comb = p2_add_73719_comb[13:1] + p2_add_73720_comb[13:1];
  assign p2_add_74512_comb = {{2{p2_bit_slice_73721_comb[10]}}, p2_bit_slice_73721_comb} + p2_add_73722_comb[13:1];
  assign p2_add_74513_comb = p2_add_73723_comb[13:1] + {{2{p2_bit_slice_73724_comb[10]}}, p2_bit_slice_73724_comb};
  assign p2_add_74514_comb = p2_add_73725_comb[13:1] + p2_add_73726_comb[13:1];
  assign p2_add_74515_comb = p2_add_73727_comb[13:1] + p2_add_73728_comb[13:1];
  assign p2_add_74516_comb = {{2{p2_bit_slice_73729_comb[10]}}, p2_bit_slice_73729_comb} + p2_add_73730_comb[13:1];
  assign p2_add_74517_comb = p2_add_73731_comb[13:1] + {{2{p2_bit_slice_73732_comb[10]}}, p2_bit_slice_73732_comb};
  assign p2_add_74518_comb = p2_add_73733_comb[13:1] + p2_add_73734_comb[13:1];
  assign p2_add_74523_comb = {{1{p2_bit_slice_73743_comb[11]}}, p2_bit_slice_73743_comb} + p2_add_73744_comb[13:1];
  assign p2_add_74524_comb = {{1{p2_bit_slice_73745_comb[11]}}, p2_bit_slice_73745_comb} + p2_add_73746_comb[13:1];
  assign p2_add_74525_comb = p2_add_73747_comb[13:1] + {{1{p2_bit_slice_73748_comb[11]}}, p2_bit_slice_73748_comb};
  assign p2_add_74526_comb = p2_add_73749_comb[13:1] + {{1{p2_bit_slice_73750_comb[11]}}, p2_bit_slice_73750_comb};
  assign p2_add_74527_comb = {{1{p2_bit_slice_73751_comb[11]}}, p2_bit_slice_73751_comb} + p2_add_73752_comb[13:1];
  assign p2_add_74528_comb = {{1{p2_bit_slice_73753_comb[11]}}, p2_bit_slice_73753_comb} + p2_add_73754_comb[13:1];
  assign p2_add_74529_comb = p2_add_73755_comb[13:1] + {{1{p2_bit_slice_73756_comb[11]}}, p2_bit_slice_73756_comb};
  assign p2_add_74530_comb = p2_add_73757_comb[13:1] + {{1{p2_bit_slice_73758_comb[11]}}, p2_bit_slice_73758_comb};
  assign p2_add_74531_comb = {{1{p2_bit_slice_73759_comb[11]}}, p2_bit_slice_73759_comb} + p2_add_73760_comb[13:1];
  assign p2_add_74532_comb = {{1{p2_bit_slice_73761_comb[11]}}, p2_bit_slice_73761_comb} + p2_add_73762_comb[13:1];
  assign p2_add_74533_comb = p2_add_73763_comb[13:1] + {{1{p2_bit_slice_73764_comb[11]}}, p2_bit_slice_73764_comb};
  assign p2_add_74534_comb = p2_add_73765_comb[13:1] + {{1{p2_bit_slice_73766_comb[11]}}, p2_bit_slice_73766_comb};
  assign p2_add_74535_comb = {{1{p2_bit_slice_73767_comb[11]}}, p2_bit_slice_73767_comb} + p2_add_73768_comb[13:1];
  assign p2_add_74536_comb = {{1{p2_bit_slice_73769_comb[11]}}, p2_bit_slice_73769_comb} + p2_add_73770_comb[13:1];
  assign p2_add_74537_comb = p2_add_73771_comb[13:1] + {{1{p2_bit_slice_73772_comb[11]}}, p2_bit_slice_73772_comb};
  assign p2_add_74538_comb = p2_add_73773_comb[13:1] + {{1{p2_bit_slice_73774_comb[11]}}, p2_bit_slice_73774_comb};
  assign p2_add_74539_comb = {{1{p2_bit_slice_73775_comb[11]}}, p2_bit_slice_73775_comb} + p2_add_73776_comb[13:1];
  assign p2_add_74540_comb = {{1{p2_bit_slice_73777_comb[11]}}, p2_bit_slice_73777_comb} + p2_add_73778_comb[13:1];
  assign p2_add_74541_comb = p2_add_73779_comb[13:1] + {{1{p2_bit_slice_73780_comb[11]}}, p2_bit_slice_73780_comb};
  assign p2_add_74542_comb = p2_add_73781_comb[13:1] + {{1{p2_bit_slice_73782_comb[11]}}, p2_bit_slice_73782_comb};
  assign p2_add_74543_comb = {{1{p2_bit_slice_73783_comb[11]}}, p2_bit_slice_73783_comb} + p2_add_73784_comb[13:1];
  assign p2_add_74544_comb = {{1{p2_bit_slice_73785_comb[11]}}, p2_bit_slice_73785_comb} + p2_add_73786_comb[13:1];
  assign p2_add_74545_comb = p2_add_73787_comb[13:1] + {{1{p2_bit_slice_73788_comb[11]}}, p2_bit_slice_73788_comb};
  assign p2_add_74546_comb = p2_add_73789_comb[13:1] + {{1{p2_bit_slice_73790_comb[11]}}, p2_bit_slice_73790_comb};
  assign p2_add_74547_comb = {{1{p2_bit_slice_73791_comb[11]}}, p2_bit_slice_73791_comb} + p2_add_73792_comb[13:1];
  assign p2_add_74548_comb = {{1{p2_bit_slice_73793_comb[11]}}, p2_bit_slice_73793_comb} + p2_add_73794_comb[13:1];
  assign p2_add_74549_comb = p2_add_73795_comb[13:1] + {{1{p2_bit_slice_73796_comb[11]}}, p2_bit_slice_73796_comb};
  assign p2_add_74550_comb = p2_add_73797_comb[13:1] + {{1{p2_bit_slice_73798_comb[11]}}, p2_bit_slice_73798_comb};
  assign p2_add_74555_comb = {{2{p2_bit_slice_73807_comb[10]}}, p2_bit_slice_73807_comb} + p2_add_73808_comb[13:1];
  assign p2_add_74556_comb = p2_add_73809_comb[13:1] + p2_add_73810_comb[13:1];
  assign p2_add_74557_comb = p2_add_73811_comb[13:1] + p2_add_73812_comb[13:1];
  assign p2_add_74558_comb = p2_add_73813_comb[13:1] + {{2{p2_bit_slice_73814_comb[10]}}, p2_bit_slice_73814_comb};
  assign p2_add_74559_comb = {{2{p2_bit_slice_73815_comb[10]}}, p2_bit_slice_73815_comb} + p2_add_73816_comb[13:1];
  assign p2_add_74560_comb = p2_add_73817_comb[13:1] + p2_add_73818_comb[13:1];
  assign p2_add_74561_comb = p2_add_73819_comb[13:1] + p2_add_73820_comb[13:1];
  assign p2_add_74562_comb = p2_add_73821_comb[13:1] + {{2{p2_bit_slice_73822_comb[10]}}, p2_bit_slice_73822_comb};
  assign p2_add_74563_comb = {{2{p2_bit_slice_73823_comb[10]}}, p2_bit_slice_73823_comb} + p2_add_73824_comb[13:1];
  assign p2_add_74564_comb = p2_add_73825_comb[13:1] + p2_add_73826_comb[13:1];
  assign p2_add_74565_comb = p2_add_73827_comb[13:1] + p2_add_73828_comb[13:1];
  assign p2_add_74566_comb = p2_add_73829_comb[13:1] + {{2{p2_bit_slice_73830_comb[10]}}, p2_bit_slice_73830_comb};
  assign p2_add_74567_comb = {{2{p2_bit_slice_73831_comb[10]}}, p2_bit_slice_73831_comb} + p2_add_73832_comb[13:1];
  assign p2_add_74568_comb = p2_add_73833_comb[13:1] + p2_add_73834_comb[13:1];
  assign p2_add_74569_comb = p2_add_73835_comb[13:1] + p2_add_73836_comb[13:1];
  assign p2_add_74570_comb = p2_add_73837_comb[13:1] + {{2{p2_bit_slice_73838_comb[10]}}, p2_bit_slice_73838_comb};
  assign p2_add_74571_comb = {{2{p2_bit_slice_73839_comb[10]}}, p2_bit_slice_73839_comb} + p2_add_73840_comb[13:1];
  assign p2_add_74572_comb = p2_add_73841_comb[13:1] + p2_add_73842_comb[13:1];
  assign p2_add_74573_comb = p2_add_73843_comb[13:1] + p2_add_73844_comb[13:1];
  assign p2_add_74574_comb = p2_add_73845_comb[13:1] + {{2{p2_bit_slice_73846_comb[10]}}, p2_bit_slice_73846_comb};
  assign p2_add_74575_comb = {{2{p2_bit_slice_73847_comb[10]}}, p2_bit_slice_73847_comb} + p2_add_73848_comb[13:1];
  assign p2_add_74576_comb = p2_add_73849_comb[13:1] + p2_add_73850_comb[13:1];
  assign p2_add_74577_comb = p2_add_73851_comb[13:1] + p2_add_73852_comb[13:1];
  assign p2_add_74578_comb = p2_add_73853_comb[13:1] + {{2{p2_bit_slice_73854_comb[10]}}, p2_bit_slice_73854_comb};
  assign p2_add_74579_comb = {{2{p2_bit_slice_73855_comb[10]}}, p2_bit_slice_73855_comb} + p2_add_73856_comb[13:1];
  assign p2_add_74580_comb = p2_add_73857_comb[13:1] + p2_add_73858_comb[13:1];
  assign p2_add_74581_comb = p2_add_73859_comb[13:1] + p2_add_73860_comb[13:1];
  assign p2_add_74582_comb = p2_add_73861_comb[13:1] + {{2{p2_bit_slice_73862_comb[10]}}, p2_bit_slice_73862_comb};
  assign p2_sum__1226_comb = p2_sum__1540_comb + p2_sum__1541_comb;
  assign p2_sum__1227_comb = p2_sum__1542_comb + p2_sum__1543_comb;
  assign p2_sum__1212_comb = p2_sum__1512_comb + p2_sum__1513_comb;
  assign p2_sum__1213_comb = p2_sum__1514_comb + p2_sum__1515_comb;
  assign p2_sum__1198_comb = p2_sum__1484_comb + p2_sum__1485_comb;
  assign p2_sum__1199_comb = p2_sum__1486_comb + p2_sum__1487_comb;
  assign p2_sum__1184_comb = p2_sum__1456_comb + p2_sum__1457_comb;
  assign p2_sum__1185_comb = p2_sum__1458_comb + p2_sum__1459_comb;
  assign p2_sum__1170_comb = p2_sum__1428_comb + p2_sum__1429_comb;
  assign p2_sum__1171_comb = p2_sum__1430_comb + p2_sum__1431_comb;
  assign p2_sum__1156_comb = p2_sum__1400_comb + p2_sum__1401_comb;
  assign p2_sum__1157_comb = p2_sum__1402_comb + p2_sum__1403_comb;
  assign p2_sum__1142_comb = p2_sum__1372_comb + p2_sum__1373_comb;
  assign p2_sum__1143_comb = p2_sum__1374_comb + p2_sum__1375_comb;
  assign p2_bit_slice_74693_comb = p2_umul_74656_comb[31:7];
  assign p2_bit_slice_74694_comb = p2_umul_74657_comb[31:7];
  assign p2_bit_slice_74695_comb = p2_umul_74658_comb[31:7];
  assign p2_bit_slice_74696_comb = p2_umul_74659_comb[31:7];
  assign p2_bit_slice_74697_comb = p2_umul_74660_comb[31:7];
  assign p2_bit_slice_74698_comb = p2_umul_74661_comb[31:7];
  assign p2_bit_slice_74699_comb = p2_umul_74662_comb[31:7];
  assign p2_sum__1079_comb = p2_sum__1246_comb + p2_sum__1247_comb;
  assign p2_sum__1078_comb = p2_sum__1244_comb + p2_sum__1245_comb;
  assign p2_sum__1077_comb = p2_sum__1242_comb + p2_sum__1243_comb;
  assign p2_sum__1075_comb = p2_sum__1238_comb + p2_sum__1239_comb;
  assign p2_sum__1074_comb = p2_sum__1236_comb + p2_sum__1237_comb;
  assign p2_sum__1073_comb = p2_sum__1234_comb + p2_sum__1235_comb;
  assign p2_add_74708_comb = p2_umul_74655_comb[31:7] + 25'h000_0001;
  assign p2_add_74709_comb = p2_sum__1076_comb + 25'h000_0001;

  // Registers for pipe stage 2:
  reg [12:0] p2_add_74363;
  reg [12:0] p2_add_74364;
  reg [12:0] p2_add_74365;
  reg [12:0] p2_add_74366;
  reg [12:0] p2_add_74367;
  reg [12:0] p2_add_74368;
  reg [12:0] p2_add_74369;
  reg [12:0] p2_add_74370;
  reg [12:0] p2_add_74371;
  reg [12:0] p2_add_74372;
  reg [12:0] p2_add_74373;
  reg [12:0] p2_add_74374;
  reg [12:0] p2_add_74375;
  reg [12:0] p2_add_74376;
  reg [12:0] p2_add_74377;
  reg [12:0] p2_add_74378;
  reg [12:0] p2_add_74379;
  reg [12:0] p2_add_74380;
  reg [12:0] p2_add_74381;
  reg [12:0] p2_add_74382;
  reg [12:0] p2_add_74383;
  reg [12:0] p2_add_74384;
  reg [12:0] p2_add_74385;
  reg [12:0] p2_add_74386;
  reg [12:0] p2_add_74387;
  reg [12:0] p2_add_74388;
  reg [12:0] p2_add_74389;
  reg [12:0] p2_add_74390;
  reg [12:0] p2_add_74395;
  reg [12:0] p2_add_74396;
  reg [12:0] p2_add_74397;
  reg [12:0] p2_add_74398;
  reg [12:0] p2_add_74399;
  reg [12:0] p2_add_74400;
  reg [12:0] p2_add_74401;
  reg [12:0] p2_add_74402;
  reg [12:0] p2_add_74403;
  reg [12:0] p2_add_74404;
  reg [12:0] p2_add_74405;
  reg [12:0] p2_add_74406;
  reg [12:0] p2_add_74407;
  reg [12:0] p2_add_74408;
  reg [12:0] p2_add_74409;
  reg [12:0] p2_add_74410;
  reg [12:0] p2_add_74411;
  reg [12:0] p2_add_74412;
  reg [12:0] p2_add_74413;
  reg [12:0] p2_add_74414;
  reg [12:0] p2_add_74415;
  reg [12:0] p2_add_74416;
  reg [12:0] p2_add_74417;
  reg [12:0] p2_add_74418;
  reg [12:0] p2_add_74419;
  reg [12:0] p2_add_74420;
  reg [12:0] p2_add_74421;
  reg [12:0] p2_add_74422;
  reg [12:0] p2_add_74427;
  reg [12:0] p2_add_74428;
  reg [12:0] p2_add_74429;
  reg [12:0] p2_add_74430;
  reg [12:0] p2_add_74431;
  reg [12:0] p2_add_74432;
  reg [12:0] p2_add_74433;
  reg [12:0] p2_add_74434;
  reg [12:0] p2_add_74435;
  reg [12:0] p2_add_74436;
  reg [12:0] p2_add_74437;
  reg [12:0] p2_add_74438;
  reg [12:0] p2_add_74439;
  reg [12:0] p2_add_74440;
  reg [12:0] p2_add_74441;
  reg [12:0] p2_add_74442;
  reg [12:0] p2_add_74443;
  reg [12:0] p2_add_74444;
  reg [12:0] p2_add_74445;
  reg [12:0] p2_add_74446;
  reg [12:0] p2_add_74447;
  reg [12:0] p2_add_74448;
  reg [12:0] p2_add_74449;
  reg [12:0] p2_add_74450;
  reg [12:0] p2_add_74451;
  reg [12:0] p2_add_74452;
  reg [12:0] p2_add_74453;
  reg [12:0] p2_add_74454;
  reg [12:0] p2_add_74491;
  reg [12:0] p2_add_74492;
  reg [12:0] p2_add_74493;
  reg [12:0] p2_add_74494;
  reg [12:0] p2_add_74495;
  reg [12:0] p2_add_74496;
  reg [12:0] p2_add_74497;
  reg [12:0] p2_add_74498;
  reg [12:0] p2_add_74499;
  reg [12:0] p2_add_74500;
  reg [12:0] p2_add_74501;
  reg [12:0] p2_add_74502;
  reg [12:0] p2_add_74503;
  reg [12:0] p2_add_74504;
  reg [12:0] p2_add_74505;
  reg [12:0] p2_add_74506;
  reg [12:0] p2_add_74507;
  reg [12:0] p2_add_74508;
  reg [12:0] p2_add_74509;
  reg [12:0] p2_add_74510;
  reg [12:0] p2_add_74511;
  reg [12:0] p2_add_74512;
  reg [12:0] p2_add_74513;
  reg [12:0] p2_add_74514;
  reg [12:0] p2_add_74515;
  reg [12:0] p2_add_74516;
  reg [12:0] p2_add_74517;
  reg [12:0] p2_add_74518;
  reg [12:0] p2_add_74523;
  reg [12:0] p2_add_74524;
  reg [12:0] p2_add_74525;
  reg [12:0] p2_add_74526;
  reg [12:0] p2_add_74527;
  reg [12:0] p2_add_74528;
  reg [12:0] p2_add_74529;
  reg [12:0] p2_add_74530;
  reg [12:0] p2_add_74531;
  reg [12:0] p2_add_74532;
  reg [12:0] p2_add_74533;
  reg [12:0] p2_add_74534;
  reg [12:0] p2_add_74535;
  reg [12:0] p2_add_74536;
  reg [12:0] p2_add_74537;
  reg [12:0] p2_add_74538;
  reg [12:0] p2_add_74539;
  reg [12:0] p2_add_74540;
  reg [12:0] p2_add_74541;
  reg [12:0] p2_add_74542;
  reg [12:0] p2_add_74543;
  reg [12:0] p2_add_74544;
  reg [12:0] p2_add_74545;
  reg [12:0] p2_add_74546;
  reg [12:0] p2_add_74547;
  reg [12:0] p2_add_74548;
  reg [12:0] p2_add_74549;
  reg [12:0] p2_add_74550;
  reg [12:0] p2_add_74555;
  reg [12:0] p2_add_74556;
  reg [12:0] p2_add_74557;
  reg [12:0] p2_add_74558;
  reg [12:0] p2_add_74559;
  reg [12:0] p2_add_74560;
  reg [12:0] p2_add_74561;
  reg [12:0] p2_add_74562;
  reg [12:0] p2_add_74563;
  reg [12:0] p2_add_74564;
  reg [12:0] p2_add_74565;
  reg [12:0] p2_add_74566;
  reg [12:0] p2_add_74567;
  reg [12:0] p2_add_74568;
  reg [12:0] p2_add_74569;
  reg [12:0] p2_add_74570;
  reg [12:0] p2_add_74571;
  reg [12:0] p2_add_74572;
  reg [12:0] p2_add_74573;
  reg [12:0] p2_add_74574;
  reg [12:0] p2_add_74575;
  reg [12:0] p2_add_74576;
  reg [12:0] p2_add_74577;
  reg [12:0] p2_add_74578;
  reg [12:0] p2_add_74579;
  reg [12:0] p2_add_74580;
  reg [12:0] p2_add_74581;
  reg [12:0] p2_add_74582;
  reg [24:0] p2_sum__1226;
  reg [24:0] p2_sum__1227;
  reg [24:0] p2_sum__1212;
  reg [24:0] p2_sum__1213;
  reg [24:0] p2_sum__1198;
  reg [24:0] p2_sum__1199;
  reg [24:0] p2_sum__1184;
  reg [24:0] p2_sum__1185;
  reg [24:0] p2_sum__1170;
  reg [24:0] p2_sum__1171;
  reg [24:0] p2_sum__1156;
  reg [24:0] p2_sum__1157;
  reg [24:0] p2_sum__1142;
  reg [24:0] p2_sum__1143;
  reg [24:0] p2_bit_slice_74693;
  reg [24:0] p2_bit_slice_74694;
  reg [24:0] p2_bit_slice_74695;
  reg [24:0] p2_bit_slice_74696;
  reg [24:0] p2_bit_slice_74697;
  reg [24:0] p2_bit_slice_74698;
  reg [24:0] p2_bit_slice_74699;
  reg [24:0] p2_sum__1079;
  reg [24:0] p2_sum__1078;
  reg [24:0] p2_sum__1077;
  reg [24:0] p2_sum__1075;
  reg [24:0] p2_sum__1074;
  reg [24:0] p2_sum__1073;
  reg [24:0] p2_add_74708;
  reg [24:0] p2_add_74709;
  always @ (posedge clk) begin
    p2_add_74363 <= p2_add_74363_comb;
    p2_add_74364 <= p2_add_74364_comb;
    p2_add_74365 <= p2_add_74365_comb;
    p2_add_74366 <= p2_add_74366_comb;
    p2_add_74367 <= p2_add_74367_comb;
    p2_add_74368 <= p2_add_74368_comb;
    p2_add_74369 <= p2_add_74369_comb;
    p2_add_74370 <= p2_add_74370_comb;
    p2_add_74371 <= p2_add_74371_comb;
    p2_add_74372 <= p2_add_74372_comb;
    p2_add_74373 <= p2_add_74373_comb;
    p2_add_74374 <= p2_add_74374_comb;
    p2_add_74375 <= p2_add_74375_comb;
    p2_add_74376 <= p2_add_74376_comb;
    p2_add_74377 <= p2_add_74377_comb;
    p2_add_74378 <= p2_add_74378_comb;
    p2_add_74379 <= p2_add_74379_comb;
    p2_add_74380 <= p2_add_74380_comb;
    p2_add_74381 <= p2_add_74381_comb;
    p2_add_74382 <= p2_add_74382_comb;
    p2_add_74383 <= p2_add_74383_comb;
    p2_add_74384 <= p2_add_74384_comb;
    p2_add_74385 <= p2_add_74385_comb;
    p2_add_74386 <= p2_add_74386_comb;
    p2_add_74387 <= p2_add_74387_comb;
    p2_add_74388 <= p2_add_74388_comb;
    p2_add_74389 <= p2_add_74389_comb;
    p2_add_74390 <= p2_add_74390_comb;
    p2_add_74395 <= p2_add_74395_comb;
    p2_add_74396 <= p2_add_74396_comb;
    p2_add_74397 <= p2_add_74397_comb;
    p2_add_74398 <= p2_add_74398_comb;
    p2_add_74399 <= p2_add_74399_comb;
    p2_add_74400 <= p2_add_74400_comb;
    p2_add_74401 <= p2_add_74401_comb;
    p2_add_74402 <= p2_add_74402_comb;
    p2_add_74403 <= p2_add_74403_comb;
    p2_add_74404 <= p2_add_74404_comb;
    p2_add_74405 <= p2_add_74405_comb;
    p2_add_74406 <= p2_add_74406_comb;
    p2_add_74407 <= p2_add_74407_comb;
    p2_add_74408 <= p2_add_74408_comb;
    p2_add_74409 <= p2_add_74409_comb;
    p2_add_74410 <= p2_add_74410_comb;
    p2_add_74411 <= p2_add_74411_comb;
    p2_add_74412 <= p2_add_74412_comb;
    p2_add_74413 <= p2_add_74413_comb;
    p2_add_74414 <= p2_add_74414_comb;
    p2_add_74415 <= p2_add_74415_comb;
    p2_add_74416 <= p2_add_74416_comb;
    p2_add_74417 <= p2_add_74417_comb;
    p2_add_74418 <= p2_add_74418_comb;
    p2_add_74419 <= p2_add_74419_comb;
    p2_add_74420 <= p2_add_74420_comb;
    p2_add_74421 <= p2_add_74421_comb;
    p2_add_74422 <= p2_add_74422_comb;
    p2_add_74427 <= p2_add_74427_comb;
    p2_add_74428 <= p2_add_74428_comb;
    p2_add_74429 <= p2_add_74429_comb;
    p2_add_74430 <= p2_add_74430_comb;
    p2_add_74431 <= p2_add_74431_comb;
    p2_add_74432 <= p2_add_74432_comb;
    p2_add_74433 <= p2_add_74433_comb;
    p2_add_74434 <= p2_add_74434_comb;
    p2_add_74435 <= p2_add_74435_comb;
    p2_add_74436 <= p2_add_74436_comb;
    p2_add_74437 <= p2_add_74437_comb;
    p2_add_74438 <= p2_add_74438_comb;
    p2_add_74439 <= p2_add_74439_comb;
    p2_add_74440 <= p2_add_74440_comb;
    p2_add_74441 <= p2_add_74441_comb;
    p2_add_74442 <= p2_add_74442_comb;
    p2_add_74443 <= p2_add_74443_comb;
    p2_add_74444 <= p2_add_74444_comb;
    p2_add_74445 <= p2_add_74445_comb;
    p2_add_74446 <= p2_add_74446_comb;
    p2_add_74447 <= p2_add_74447_comb;
    p2_add_74448 <= p2_add_74448_comb;
    p2_add_74449 <= p2_add_74449_comb;
    p2_add_74450 <= p2_add_74450_comb;
    p2_add_74451 <= p2_add_74451_comb;
    p2_add_74452 <= p2_add_74452_comb;
    p2_add_74453 <= p2_add_74453_comb;
    p2_add_74454 <= p2_add_74454_comb;
    p2_add_74491 <= p2_add_74491_comb;
    p2_add_74492 <= p2_add_74492_comb;
    p2_add_74493 <= p2_add_74493_comb;
    p2_add_74494 <= p2_add_74494_comb;
    p2_add_74495 <= p2_add_74495_comb;
    p2_add_74496 <= p2_add_74496_comb;
    p2_add_74497 <= p2_add_74497_comb;
    p2_add_74498 <= p2_add_74498_comb;
    p2_add_74499 <= p2_add_74499_comb;
    p2_add_74500 <= p2_add_74500_comb;
    p2_add_74501 <= p2_add_74501_comb;
    p2_add_74502 <= p2_add_74502_comb;
    p2_add_74503 <= p2_add_74503_comb;
    p2_add_74504 <= p2_add_74504_comb;
    p2_add_74505 <= p2_add_74505_comb;
    p2_add_74506 <= p2_add_74506_comb;
    p2_add_74507 <= p2_add_74507_comb;
    p2_add_74508 <= p2_add_74508_comb;
    p2_add_74509 <= p2_add_74509_comb;
    p2_add_74510 <= p2_add_74510_comb;
    p2_add_74511 <= p2_add_74511_comb;
    p2_add_74512 <= p2_add_74512_comb;
    p2_add_74513 <= p2_add_74513_comb;
    p2_add_74514 <= p2_add_74514_comb;
    p2_add_74515 <= p2_add_74515_comb;
    p2_add_74516 <= p2_add_74516_comb;
    p2_add_74517 <= p2_add_74517_comb;
    p2_add_74518 <= p2_add_74518_comb;
    p2_add_74523 <= p2_add_74523_comb;
    p2_add_74524 <= p2_add_74524_comb;
    p2_add_74525 <= p2_add_74525_comb;
    p2_add_74526 <= p2_add_74526_comb;
    p2_add_74527 <= p2_add_74527_comb;
    p2_add_74528 <= p2_add_74528_comb;
    p2_add_74529 <= p2_add_74529_comb;
    p2_add_74530 <= p2_add_74530_comb;
    p2_add_74531 <= p2_add_74531_comb;
    p2_add_74532 <= p2_add_74532_comb;
    p2_add_74533 <= p2_add_74533_comb;
    p2_add_74534 <= p2_add_74534_comb;
    p2_add_74535 <= p2_add_74535_comb;
    p2_add_74536 <= p2_add_74536_comb;
    p2_add_74537 <= p2_add_74537_comb;
    p2_add_74538 <= p2_add_74538_comb;
    p2_add_74539 <= p2_add_74539_comb;
    p2_add_74540 <= p2_add_74540_comb;
    p2_add_74541 <= p2_add_74541_comb;
    p2_add_74542 <= p2_add_74542_comb;
    p2_add_74543 <= p2_add_74543_comb;
    p2_add_74544 <= p2_add_74544_comb;
    p2_add_74545 <= p2_add_74545_comb;
    p2_add_74546 <= p2_add_74546_comb;
    p2_add_74547 <= p2_add_74547_comb;
    p2_add_74548 <= p2_add_74548_comb;
    p2_add_74549 <= p2_add_74549_comb;
    p2_add_74550 <= p2_add_74550_comb;
    p2_add_74555 <= p2_add_74555_comb;
    p2_add_74556 <= p2_add_74556_comb;
    p2_add_74557 <= p2_add_74557_comb;
    p2_add_74558 <= p2_add_74558_comb;
    p2_add_74559 <= p2_add_74559_comb;
    p2_add_74560 <= p2_add_74560_comb;
    p2_add_74561 <= p2_add_74561_comb;
    p2_add_74562 <= p2_add_74562_comb;
    p2_add_74563 <= p2_add_74563_comb;
    p2_add_74564 <= p2_add_74564_comb;
    p2_add_74565 <= p2_add_74565_comb;
    p2_add_74566 <= p2_add_74566_comb;
    p2_add_74567 <= p2_add_74567_comb;
    p2_add_74568 <= p2_add_74568_comb;
    p2_add_74569 <= p2_add_74569_comb;
    p2_add_74570 <= p2_add_74570_comb;
    p2_add_74571 <= p2_add_74571_comb;
    p2_add_74572 <= p2_add_74572_comb;
    p2_add_74573 <= p2_add_74573_comb;
    p2_add_74574 <= p2_add_74574_comb;
    p2_add_74575 <= p2_add_74575_comb;
    p2_add_74576 <= p2_add_74576_comb;
    p2_add_74577 <= p2_add_74577_comb;
    p2_add_74578 <= p2_add_74578_comb;
    p2_add_74579 <= p2_add_74579_comb;
    p2_add_74580 <= p2_add_74580_comb;
    p2_add_74581 <= p2_add_74581_comb;
    p2_add_74582 <= p2_add_74582_comb;
    p2_sum__1226 <= p2_sum__1226_comb;
    p2_sum__1227 <= p2_sum__1227_comb;
    p2_sum__1212 <= p2_sum__1212_comb;
    p2_sum__1213 <= p2_sum__1213_comb;
    p2_sum__1198 <= p2_sum__1198_comb;
    p2_sum__1199 <= p2_sum__1199_comb;
    p2_sum__1184 <= p2_sum__1184_comb;
    p2_sum__1185 <= p2_sum__1185_comb;
    p2_sum__1170 <= p2_sum__1170_comb;
    p2_sum__1171 <= p2_sum__1171_comb;
    p2_sum__1156 <= p2_sum__1156_comb;
    p2_sum__1157 <= p2_sum__1157_comb;
    p2_sum__1142 <= p2_sum__1142_comb;
    p2_sum__1143 <= p2_sum__1143_comb;
    p2_bit_slice_74693 <= p2_bit_slice_74693_comb;
    p2_bit_slice_74694 <= p2_bit_slice_74694_comb;
    p2_bit_slice_74695 <= p2_bit_slice_74695_comb;
    p2_bit_slice_74696 <= p2_bit_slice_74696_comb;
    p2_bit_slice_74697 <= p2_bit_slice_74697_comb;
    p2_bit_slice_74698 <= p2_bit_slice_74698_comb;
    p2_bit_slice_74699 <= p2_bit_slice_74699_comb;
    p2_sum__1079 <= p2_sum__1079_comb;
    p2_sum__1078 <= p2_sum__1078_comb;
    p2_sum__1077 <= p2_sum__1077_comb;
    p2_sum__1075 <= p2_sum__1075_comb;
    p2_sum__1074 <= p2_sum__1074_comb;
    p2_sum__1073 <= p2_sum__1073_comb;
    p2_add_74708 <= p2_add_74708_comb;
    p2_add_74709 <= p2_add_74709_comb;
  end

  // ===== Pipe stage 3:
  wire [24:0] p3_sum__1552_comb;
  wire [24:0] p3_sum__1553_comb;
  wire [24:0] p3_sum__1554_comb;
  wire [24:0] p3_sum__1555_comb;
  wire [24:0] p3_sum__1524_comb;
  wire [24:0] p3_sum__1525_comb;
  wire [24:0] p3_sum__1526_comb;
  wire [24:0] p3_sum__1527_comb;
  wire [24:0] p3_sum__1496_comb;
  wire [24:0] p3_sum__1497_comb;
  wire [24:0] p3_sum__1498_comb;
  wire [24:0] p3_sum__1499_comb;
  wire [24:0] p3_sum__1468_comb;
  wire [24:0] p3_sum__1469_comb;
  wire [24:0] p3_sum__1470_comb;
  wire [24:0] p3_sum__1471_comb;
  wire [24:0] p3_sum__1440_comb;
  wire [24:0] p3_sum__1441_comb;
  wire [24:0] p3_sum__1442_comb;
  wire [24:0] p3_sum__1443_comb;
  wire [24:0] p3_sum__1412_comb;
  wire [24:0] p3_sum__1413_comb;
  wire [24:0] p3_sum__1414_comb;
  wire [24:0] p3_sum__1415_comb;
  wire [24:0] p3_sum__1384_comb;
  wire [24:0] p3_sum__1385_comb;
  wire [24:0] p3_sum__1386_comb;
  wire [24:0] p3_sum__1387_comb;
  wire [24:0] p3_sum__1548_comb;
  wire [24:0] p3_sum__1549_comb;
  wire [24:0] p3_sum__1550_comb;
  wire [24:0] p3_sum__1551_comb;
  wire [24:0] p3_sum__1520_comb;
  wire [24:0] p3_sum__1521_comb;
  wire [24:0] p3_sum__1522_comb;
  wire [24:0] p3_sum__1523_comb;
  wire [24:0] p3_sum__1492_comb;
  wire [24:0] p3_sum__1493_comb;
  wire [24:0] p3_sum__1494_comb;
  wire [24:0] p3_sum__1495_comb;
  wire [24:0] p3_sum__1464_comb;
  wire [24:0] p3_sum__1465_comb;
  wire [24:0] p3_sum__1466_comb;
  wire [24:0] p3_sum__1467_comb;
  wire [24:0] p3_sum__1436_comb;
  wire [24:0] p3_sum__1437_comb;
  wire [24:0] p3_sum__1438_comb;
  wire [24:0] p3_sum__1439_comb;
  wire [24:0] p3_sum__1408_comb;
  wire [24:0] p3_sum__1409_comb;
  wire [24:0] p3_sum__1410_comb;
  wire [24:0] p3_sum__1411_comb;
  wire [24:0] p3_sum__1380_comb;
  wire [24:0] p3_sum__1381_comb;
  wire [24:0] p3_sum__1382_comb;
  wire [24:0] p3_sum__1383_comb;
  wire [24:0] p3_sum__1544_comb;
  wire [24:0] p3_sum__1545_comb;
  wire [24:0] p3_sum__1546_comb;
  wire [24:0] p3_sum__1547_comb;
  wire [24:0] p3_sum__1516_comb;
  wire [24:0] p3_sum__1517_comb;
  wire [24:0] p3_sum__1518_comb;
  wire [24:0] p3_sum__1519_comb;
  wire [24:0] p3_sum__1488_comb;
  wire [24:0] p3_sum__1489_comb;
  wire [24:0] p3_sum__1490_comb;
  wire [24:0] p3_sum__1491_comb;
  wire [24:0] p3_sum__1460_comb;
  wire [24:0] p3_sum__1461_comb;
  wire [24:0] p3_sum__1462_comb;
  wire [24:0] p3_sum__1463_comb;
  wire [24:0] p3_sum__1432_comb;
  wire [24:0] p3_sum__1433_comb;
  wire [24:0] p3_sum__1434_comb;
  wire [24:0] p3_sum__1435_comb;
  wire [24:0] p3_sum__1404_comb;
  wire [24:0] p3_sum__1405_comb;
  wire [24:0] p3_sum__1406_comb;
  wire [24:0] p3_sum__1407_comb;
  wire [24:0] p3_sum__1376_comb;
  wire [24:0] p3_sum__1377_comb;
  wire [24:0] p3_sum__1378_comb;
  wire [24:0] p3_sum__1379_comb;
  wire [24:0] p3_sum__1536_comb;
  wire [24:0] p3_sum__1537_comb;
  wire [24:0] p3_sum__1538_comb;
  wire [24:0] p3_sum__1539_comb;
  wire [24:0] p3_sum__1508_comb;
  wire [24:0] p3_sum__1509_comb;
  wire [24:0] p3_sum__1510_comb;
  wire [24:0] p3_sum__1511_comb;
  wire [24:0] p3_sum__1480_comb;
  wire [24:0] p3_sum__1481_comb;
  wire [24:0] p3_sum__1482_comb;
  wire [24:0] p3_sum__1483_comb;
  wire [24:0] p3_sum__1452_comb;
  wire [24:0] p3_sum__1453_comb;
  wire [24:0] p3_sum__1454_comb;
  wire [24:0] p3_sum__1455_comb;
  wire [24:0] p3_sum__1424_comb;
  wire [24:0] p3_sum__1425_comb;
  wire [24:0] p3_sum__1426_comb;
  wire [24:0] p3_sum__1427_comb;
  wire [24:0] p3_sum__1396_comb;
  wire [24:0] p3_sum__1397_comb;
  wire [24:0] p3_sum__1398_comb;
  wire [24:0] p3_sum__1399_comb;
  wire [24:0] p3_sum__1368_comb;
  wire [24:0] p3_sum__1369_comb;
  wire [24:0] p3_sum__1370_comb;
  wire [24:0] p3_sum__1371_comb;
  wire [24:0] p3_sum__1532_comb;
  wire [24:0] p3_sum__1533_comb;
  wire [24:0] p3_sum__1534_comb;
  wire [24:0] p3_sum__1535_comb;
  wire [24:0] p3_sum__1504_comb;
  wire [24:0] p3_sum__1505_comb;
  wire [24:0] p3_sum__1506_comb;
  wire [24:0] p3_sum__1507_comb;
  wire [24:0] p3_sum__1476_comb;
  wire [24:0] p3_sum__1477_comb;
  wire [24:0] p3_sum__1478_comb;
  wire [24:0] p3_sum__1479_comb;
  wire [24:0] p3_sum__1448_comb;
  wire [24:0] p3_sum__1449_comb;
  wire [24:0] p3_sum__1450_comb;
  wire [24:0] p3_sum__1451_comb;
  wire [24:0] p3_sum__1420_comb;
  wire [24:0] p3_sum__1421_comb;
  wire [24:0] p3_sum__1422_comb;
  wire [24:0] p3_sum__1423_comb;
  wire [24:0] p3_sum__1392_comb;
  wire [24:0] p3_sum__1393_comb;
  wire [24:0] p3_sum__1394_comb;
  wire [24:0] p3_sum__1395_comb;
  wire [24:0] p3_sum__1364_comb;
  wire [24:0] p3_sum__1365_comb;
  wire [24:0] p3_sum__1366_comb;
  wire [24:0] p3_sum__1367_comb;
  wire [24:0] p3_sum__1528_comb;
  wire [24:0] p3_sum__1529_comb;
  wire [24:0] p3_sum__1530_comb;
  wire [24:0] p3_sum__1531_comb;
  wire [24:0] p3_sum__1500_comb;
  wire [24:0] p3_sum__1501_comb;
  wire [24:0] p3_sum__1502_comb;
  wire [24:0] p3_sum__1503_comb;
  wire [24:0] p3_sum__1472_comb;
  wire [24:0] p3_sum__1473_comb;
  wire [24:0] p3_sum__1474_comb;
  wire [24:0] p3_sum__1475_comb;
  wire [24:0] p3_sum__1444_comb;
  wire [24:0] p3_sum__1445_comb;
  wire [24:0] p3_sum__1446_comb;
  wire [24:0] p3_sum__1447_comb;
  wire [24:0] p3_sum__1416_comb;
  wire [24:0] p3_sum__1417_comb;
  wire [24:0] p3_sum__1418_comb;
  wire [24:0] p3_sum__1419_comb;
  wire [24:0] p3_sum__1388_comb;
  wire [24:0] p3_sum__1389_comb;
  wire [24:0] p3_sum__1390_comb;
  wire [24:0] p3_sum__1391_comb;
  wire [24:0] p3_sum__1360_comb;
  wire [24:0] p3_sum__1361_comb;
  wire [24:0] p3_sum__1362_comb;
  wire [24:0] p3_sum__1363_comb;
  wire [24:0] p3_sum__1232_comb;
  wire [24:0] p3_sum__1233_comb;
  wire [24:0] p3_sum__1218_comb;
  wire [24:0] p3_sum__1219_comb;
  wire [24:0] p3_sum__1204_comb;
  wire [24:0] p3_sum__1205_comb;
  wire [24:0] p3_sum__1190_comb;
  wire [24:0] p3_sum__1191_comb;
  wire [24:0] p3_sum__1176_comb;
  wire [24:0] p3_sum__1177_comb;
  wire [24:0] p3_sum__1162_comb;
  wire [24:0] p3_sum__1163_comb;
  wire [24:0] p3_sum__1148_comb;
  wire [24:0] p3_sum__1149_comb;
  wire [24:0] p3_sum__1230_comb;
  wire [24:0] p3_sum__1231_comb;
  wire [24:0] p3_sum__1216_comb;
  wire [24:0] p3_sum__1217_comb;
  wire [24:0] p3_sum__1202_comb;
  wire [24:0] p3_sum__1203_comb;
  wire [24:0] p3_sum__1188_comb;
  wire [24:0] p3_sum__1189_comb;
  wire [24:0] p3_sum__1174_comb;
  wire [24:0] p3_sum__1175_comb;
  wire [24:0] p3_sum__1160_comb;
  wire [24:0] p3_sum__1161_comb;
  wire [24:0] p3_sum__1146_comb;
  wire [24:0] p3_sum__1147_comb;
  wire [24:0] p3_sum__1228_comb;
  wire [24:0] p3_sum__1229_comb;
  wire [24:0] p3_sum__1214_comb;
  wire [24:0] p3_sum__1215_comb;
  wire [24:0] p3_sum__1200_comb;
  wire [24:0] p3_sum__1201_comb;
  wire [24:0] p3_sum__1186_comb;
  wire [24:0] p3_sum__1187_comb;
  wire [24:0] p3_sum__1172_comb;
  wire [24:0] p3_sum__1173_comb;
  wire [24:0] p3_sum__1158_comb;
  wire [24:0] p3_sum__1159_comb;
  wire [24:0] p3_sum__1144_comb;
  wire [24:0] p3_sum__1145_comb;
  wire [24:0] p3_sum__1224_comb;
  wire [24:0] p3_sum__1225_comb;
  wire [24:0] p3_sum__1210_comb;
  wire [24:0] p3_sum__1211_comb;
  wire [24:0] p3_sum__1196_comb;
  wire [24:0] p3_sum__1197_comb;
  wire [24:0] p3_sum__1182_comb;
  wire [24:0] p3_sum__1183_comb;
  wire [24:0] p3_sum__1168_comb;
  wire [24:0] p3_sum__1169_comb;
  wire [24:0] p3_sum__1154_comb;
  wire [24:0] p3_sum__1155_comb;
  wire [24:0] p3_sum__1140_comb;
  wire [24:0] p3_sum__1141_comb;
  wire [24:0] p3_sum__1222_comb;
  wire [24:0] p3_sum__1223_comb;
  wire [24:0] p3_sum__1208_comb;
  wire [24:0] p3_sum__1209_comb;
  wire [24:0] p3_sum__1194_comb;
  wire [24:0] p3_sum__1195_comb;
  wire [24:0] p3_sum__1180_comb;
  wire [24:0] p3_sum__1181_comb;
  wire [24:0] p3_sum__1166_comb;
  wire [24:0] p3_sum__1167_comb;
  wire [24:0] p3_sum__1152_comb;
  wire [24:0] p3_sum__1153_comb;
  wire [24:0] p3_sum__1138_comb;
  wire [24:0] p3_sum__1139_comb;
  wire [24:0] p3_sum__1220_comb;
  wire [24:0] p3_sum__1221_comb;
  wire [24:0] p3_sum__1206_comb;
  wire [24:0] p3_sum__1207_comb;
  wire [24:0] p3_sum__1192_comb;
  wire [24:0] p3_sum__1193_comb;
  wire [24:0] p3_sum__1178_comb;
  wire [24:0] p3_sum__1179_comb;
  wire [24:0] p3_sum__1164_comb;
  wire [24:0] p3_sum__1165_comb;
  wire [24:0] p3_sum__1150_comb;
  wire [24:0] p3_sum__1151_comb;
  wire [24:0] p3_sum__1136_comb;
  wire [24:0] p3_sum__1137_comb;
  wire [24:0] p3_sum__1072_comb;
  wire [24:0] p3_sum__1065_comb;
  wire [24:0] p3_sum__1058_comb;
  wire [24:0] p3_sum__1051_comb;
  wire [24:0] p3_sum__1044_comb;
  wire [24:0] p3_sum__1037_comb;
  wire [24:0] p3_sum__1030_comb;
  wire [24:0] p3_sum__1071_comb;
  wire [24:0] p3_sum__1064_comb;
  wire [24:0] p3_sum__1057_comb;
  wire [24:0] p3_sum__1050_comb;
  wire [24:0] p3_sum__1043_comb;
  wire [24:0] p3_sum__1036_comb;
  wire [24:0] p3_sum__1029_comb;
  wire [24:0] p3_sum__1070_comb;
  wire [24:0] p3_sum__1063_comb;
  wire [24:0] p3_sum__1056_comb;
  wire [24:0] p3_sum__1049_comb;
  wire [24:0] p3_sum__1042_comb;
  wire [24:0] p3_sum__1035_comb;
  wire [24:0] p3_sum__1028_comb;
  wire [24:0] p3_sum__1069_comb;
  wire [24:0] p3_sum__1062_comb;
  wire [24:0] p3_sum__1055_comb;
  wire [24:0] p3_sum__1048_comb;
  wire [24:0] p3_sum__1041_comb;
  wire [24:0] p3_sum__1034_comb;
  wire [24:0] p3_sum__1027_comb;
  wire [24:0] p3_sum__1068_comb;
  wire [24:0] p3_sum__1061_comb;
  wire [24:0] p3_sum__1054_comb;
  wire [24:0] p3_sum__1047_comb;
  wire [24:0] p3_sum__1040_comb;
  wire [24:0] p3_sum__1033_comb;
  wire [24:0] p3_sum__1026_comb;
  wire [24:0] p3_sum__1067_comb;
  wire [24:0] p3_sum__1060_comb;
  wire [24:0] p3_sum__1053_comb;
  wire [24:0] p3_sum__1046_comb;
  wire [24:0] p3_sum__1039_comb;
  wire [24:0] p3_sum__1032_comb;
  wire [24:0] p3_sum__1025_comb;
  wire [24:0] p3_sum__1066_comb;
  wire [24:0] p3_sum__1059_comb;
  wire [24:0] p3_sum__1052_comb;
  wire [24:0] p3_sum__1045_comb;
  wire [24:0] p3_sum__1038_comb;
  wire [24:0] p3_sum__1031_comb;
  wire [24:0] p3_sum__1024_comb;
  wire [24:0] p3_add_75467_comb;
  wire [24:0] p3_add_75468_comb;
  wire [24:0] p3_add_75469_comb;
  wire [24:0] p3_add_75470_comb;
  wire [24:0] p3_add_75471_comb;
  wire [24:0] p3_add_75472_comb;
  wire [24:0] p3_add_75473_comb;
  wire [24:0] p3_add_75474_comb;
  wire [24:0] p3_add_75475_comb;
  wire [24:0] p3_add_75476_comb;
  wire [24:0] p3_add_75477_comb;
  wire [24:0] p3_add_75478_comb;
  wire [24:0] p3_add_75479_comb;
  wire [24:0] p3_add_75480_comb;
  wire [24:0] p3_add_75481_comb;
  wire [24:0] p3_add_75482_comb;
  wire [24:0] p3_add_75483_comb;
  wire [24:0] p3_add_75484_comb;
  wire [24:0] p3_add_75485_comb;
  wire [24:0] p3_add_75486_comb;
  wire [24:0] p3_add_75487_comb;
  wire [24:0] p3_add_75488_comb;
  wire [24:0] p3_add_75489_comb;
  wire [24:0] p3_add_75490_comb;
  wire [24:0] p3_add_75491_comb;
  wire [24:0] p3_add_75492_comb;
  wire [24:0] p3_add_75493_comb;
  wire [24:0] p3_add_75494_comb;
  wire [24:0] p3_add_75495_comb;
  wire [24:0] p3_add_75496_comb;
  wire [24:0] p3_add_75497_comb;
  wire [24:0] p3_add_75498_comb;
  wire [24:0] p3_add_75499_comb;
  wire [24:0] p3_add_75500_comb;
  wire [24:0] p3_add_75501_comb;
  wire [24:0] p3_add_75502_comb;
  wire [24:0] p3_add_75503_comb;
  wire [24:0] p3_add_75504_comb;
  wire [24:0] p3_add_75505_comb;
  wire [24:0] p3_add_75506_comb;
  wire [24:0] p3_add_75507_comb;
  wire [24:0] p3_add_75508_comb;
  wire [24:0] p3_add_75509_comb;
  wire [24:0] p3_add_75510_comb;
  wire [24:0] p3_add_75511_comb;
  wire [24:0] p3_add_75512_comb;
  wire [24:0] p3_add_75513_comb;
  wire [24:0] p3_add_75514_comb;
  wire [24:0] p3_add_75515_comb;
  wire [24:0] p3_add_75516_comb;
  wire [24:0] p3_add_75517_comb;
  wire [24:0] p3_add_75518_comb;
  wire [24:0] p3_add_75519_comb;
  wire [24:0] p3_add_75520_comb;
  wire [24:0] p3_add_75521_comb;
  wire [24:0] p3_add_75522_comb;
  wire [24:0] p3_add_75523_comb;
  wire [24:0] p3_add_75524_comb;
  wire [24:0] p3_add_75525_comb;
  wire [24:0] p3_add_75526_comb;
  wire [24:0] p3_add_75527_comb;
  wire [24:0] p3_add_75528_comb;
  wire [11:0] p3_clipped__136_comb;
  wire [11:0] p3_clipped__152_comb;
  wire [11:0] p3_clipped__168_comb;
  wire [11:0] p3_clipped__184_comb;
  wire [11:0] p3_clipped__200_comb;
  wire [11:0] p3_clipped__216_comb;
  wire [11:0] p3_clipped__232_comb;
  wire [11:0] p3_clipped__248_comb;
  wire [11:0] p3_clipped__137_comb;
  wire [11:0] p3_clipped__153_comb;
  wire [11:0] p3_clipped__169_comb;
  wire [11:0] p3_clipped__185_comb;
  wire [11:0] p3_clipped__201_comb;
  wire [11:0] p3_clipped__217_comb;
  wire [11:0] p3_clipped__233_comb;
  wire [11:0] p3_clipped__249_comb;
  wire [11:0] p3_clipped__138_comb;
  wire [11:0] p3_clipped__154_comb;
  wire [11:0] p3_clipped__170_comb;
  wire [11:0] p3_clipped__186_comb;
  wire [11:0] p3_clipped__202_comb;
  wire [11:0] p3_clipped__218_comb;
  wire [11:0] p3_clipped__234_comb;
  wire [11:0] p3_clipped__250_comb;
  wire [11:0] p3_clipped__139_comb;
  wire [11:0] p3_clipped__155_comb;
  wire [11:0] p3_clipped__171_comb;
  wire [11:0] p3_clipped__187_comb;
  wire [11:0] p3_clipped__203_comb;
  wire [11:0] p3_clipped__219_comb;
  wire [11:0] p3_clipped__235_comb;
  wire [11:0] p3_clipped__251_comb;
  wire [11:0] p3_clipped__140_comb;
  wire [11:0] p3_clipped__156_comb;
  wire [11:0] p3_clipped__172_comb;
  wire [11:0] p3_clipped__188_comb;
  wire [11:0] p3_clipped__204_comb;
  wire [11:0] p3_clipped__220_comb;
  wire [11:0] p3_clipped__236_comb;
  wire [11:0] p3_clipped__252_comb;
  wire [11:0] p3_clipped__141_comb;
  wire [11:0] p3_clipped__157_comb;
  wire [11:0] p3_clipped__173_comb;
  wire [11:0] p3_clipped__189_comb;
  wire [11:0] p3_clipped__205_comb;
  wire [11:0] p3_clipped__221_comb;
  wire [11:0] p3_clipped__237_comb;
  wire [11:0] p3_clipped__253_comb;
  wire [11:0] p3_clipped__142_comb;
  wire [11:0] p3_clipped__158_comb;
  wire [11:0] p3_clipped__174_comb;
  wire [11:0] p3_clipped__190_comb;
  wire [11:0] p3_clipped__206_comb;
  wire [11:0] p3_clipped__222_comb;
  wire [11:0] p3_clipped__238_comb;
  wire [11:0] p3_clipped__254_comb;
  wire [11:0] p3_clipped__143_comb;
  wire [11:0] p3_clipped__159_comb;
  wire [11:0] p3_clipped__175_comb;
  wire [11:0] p3_clipped__191_comb;
  wire [11:0] p3_clipped__207_comb;
  wire [11:0] p3_clipped__223_comb;
  wire [11:0] p3_clipped__239_comb;
  wire [11:0] p3_clipped__255_comb;
  wire [11:0] p3_array_76169_comb[0:7];
  wire [11:0] p3_array_76170_comb[0:7];
  wire [11:0] p3_array_76171_comb[0:7];
  wire [11:0] p3_array_76172_comb[0:7];
  wire [11:0] p3_array_76173_comb[0:7];
  wire [11:0] p3_array_76174_comb[0:7];
  wire [11:0] p3_array_76175_comb[0:7];
  wire [11:0] p3_array_76176_comb[0:7];
  wire [11:0] p3_col_transformed_comb[0:7][0:7];
  assign p3_sum__1552_comb = {{12{p2_add_74363[12]}}, p2_add_74363};
  assign p3_sum__1553_comb = {{12{p2_add_74364[12]}}, p2_add_74364};
  assign p3_sum__1554_comb = {{12{p2_add_74365[12]}}, p2_add_74365};
  assign p3_sum__1555_comb = {{12{p2_add_74366[12]}}, p2_add_74366};
  assign p3_sum__1524_comb = {{12{p2_add_74367[12]}}, p2_add_74367};
  assign p3_sum__1525_comb = {{12{p2_add_74368[12]}}, p2_add_74368};
  assign p3_sum__1526_comb = {{12{p2_add_74369[12]}}, p2_add_74369};
  assign p3_sum__1527_comb = {{12{p2_add_74370[12]}}, p2_add_74370};
  assign p3_sum__1496_comb = {{12{p2_add_74371[12]}}, p2_add_74371};
  assign p3_sum__1497_comb = {{12{p2_add_74372[12]}}, p2_add_74372};
  assign p3_sum__1498_comb = {{12{p2_add_74373[12]}}, p2_add_74373};
  assign p3_sum__1499_comb = {{12{p2_add_74374[12]}}, p2_add_74374};
  assign p3_sum__1468_comb = {{12{p2_add_74375[12]}}, p2_add_74375};
  assign p3_sum__1469_comb = {{12{p2_add_74376[12]}}, p2_add_74376};
  assign p3_sum__1470_comb = {{12{p2_add_74377[12]}}, p2_add_74377};
  assign p3_sum__1471_comb = {{12{p2_add_74378[12]}}, p2_add_74378};
  assign p3_sum__1440_comb = {{12{p2_add_74379[12]}}, p2_add_74379};
  assign p3_sum__1441_comb = {{12{p2_add_74380[12]}}, p2_add_74380};
  assign p3_sum__1442_comb = {{12{p2_add_74381[12]}}, p2_add_74381};
  assign p3_sum__1443_comb = {{12{p2_add_74382[12]}}, p2_add_74382};
  assign p3_sum__1412_comb = {{12{p2_add_74383[12]}}, p2_add_74383};
  assign p3_sum__1413_comb = {{12{p2_add_74384[12]}}, p2_add_74384};
  assign p3_sum__1414_comb = {{12{p2_add_74385[12]}}, p2_add_74385};
  assign p3_sum__1415_comb = {{12{p2_add_74386[12]}}, p2_add_74386};
  assign p3_sum__1384_comb = {{12{p2_add_74387[12]}}, p2_add_74387};
  assign p3_sum__1385_comb = {{12{p2_add_74388[12]}}, p2_add_74388};
  assign p3_sum__1386_comb = {{12{p2_add_74389[12]}}, p2_add_74389};
  assign p3_sum__1387_comb = {{12{p2_add_74390[12]}}, p2_add_74390};
  assign p3_sum__1548_comb = {{12{p2_add_74395[12]}}, p2_add_74395};
  assign p3_sum__1549_comb = {{12{p2_add_74396[12]}}, p2_add_74396};
  assign p3_sum__1550_comb = {{12{p2_add_74397[12]}}, p2_add_74397};
  assign p3_sum__1551_comb = {{12{p2_add_74398[12]}}, p2_add_74398};
  assign p3_sum__1520_comb = {{12{p2_add_74399[12]}}, p2_add_74399};
  assign p3_sum__1521_comb = {{12{p2_add_74400[12]}}, p2_add_74400};
  assign p3_sum__1522_comb = {{12{p2_add_74401[12]}}, p2_add_74401};
  assign p3_sum__1523_comb = {{12{p2_add_74402[12]}}, p2_add_74402};
  assign p3_sum__1492_comb = {{12{p2_add_74403[12]}}, p2_add_74403};
  assign p3_sum__1493_comb = {{12{p2_add_74404[12]}}, p2_add_74404};
  assign p3_sum__1494_comb = {{12{p2_add_74405[12]}}, p2_add_74405};
  assign p3_sum__1495_comb = {{12{p2_add_74406[12]}}, p2_add_74406};
  assign p3_sum__1464_comb = {{12{p2_add_74407[12]}}, p2_add_74407};
  assign p3_sum__1465_comb = {{12{p2_add_74408[12]}}, p2_add_74408};
  assign p3_sum__1466_comb = {{12{p2_add_74409[12]}}, p2_add_74409};
  assign p3_sum__1467_comb = {{12{p2_add_74410[12]}}, p2_add_74410};
  assign p3_sum__1436_comb = {{12{p2_add_74411[12]}}, p2_add_74411};
  assign p3_sum__1437_comb = {{12{p2_add_74412[12]}}, p2_add_74412};
  assign p3_sum__1438_comb = {{12{p2_add_74413[12]}}, p2_add_74413};
  assign p3_sum__1439_comb = {{12{p2_add_74414[12]}}, p2_add_74414};
  assign p3_sum__1408_comb = {{12{p2_add_74415[12]}}, p2_add_74415};
  assign p3_sum__1409_comb = {{12{p2_add_74416[12]}}, p2_add_74416};
  assign p3_sum__1410_comb = {{12{p2_add_74417[12]}}, p2_add_74417};
  assign p3_sum__1411_comb = {{12{p2_add_74418[12]}}, p2_add_74418};
  assign p3_sum__1380_comb = {{12{p2_add_74419[12]}}, p2_add_74419};
  assign p3_sum__1381_comb = {{12{p2_add_74420[12]}}, p2_add_74420};
  assign p3_sum__1382_comb = {{12{p2_add_74421[12]}}, p2_add_74421};
  assign p3_sum__1383_comb = {{12{p2_add_74422[12]}}, p2_add_74422};
  assign p3_sum__1544_comb = {{12{p2_add_74427[12]}}, p2_add_74427};
  assign p3_sum__1545_comb = {{12{p2_add_74428[12]}}, p2_add_74428};
  assign p3_sum__1546_comb = {{12{p2_add_74429[12]}}, p2_add_74429};
  assign p3_sum__1547_comb = {{12{p2_add_74430[12]}}, p2_add_74430};
  assign p3_sum__1516_comb = {{12{p2_add_74431[12]}}, p2_add_74431};
  assign p3_sum__1517_comb = {{12{p2_add_74432[12]}}, p2_add_74432};
  assign p3_sum__1518_comb = {{12{p2_add_74433[12]}}, p2_add_74433};
  assign p3_sum__1519_comb = {{12{p2_add_74434[12]}}, p2_add_74434};
  assign p3_sum__1488_comb = {{12{p2_add_74435[12]}}, p2_add_74435};
  assign p3_sum__1489_comb = {{12{p2_add_74436[12]}}, p2_add_74436};
  assign p3_sum__1490_comb = {{12{p2_add_74437[12]}}, p2_add_74437};
  assign p3_sum__1491_comb = {{12{p2_add_74438[12]}}, p2_add_74438};
  assign p3_sum__1460_comb = {{12{p2_add_74439[12]}}, p2_add_74439};
  assign p3_sum__1461_comb = {{12{p2_add_74440[12]}}, p2_add_74440};
  assign p3_sum__1462_comb = {{12{p2_add_74441[12]}}, p2_add_74441};
  assign p3_sum__1463_comb = {{12{p2_add_74442[12]}}, p2_add_74442};
  assign p3_sum__1432_comb = {{12{p2_add_74443[12]}}, p2_add_74443};
  assign p3_sum__1433_comb = {{12{p2_add_74444[12]}}, p2_add_74444};
  assign p3_sum__1434_comb = {{12{p2_add_74445[12]}}, p2_add_74445};
  assign p3_sum__1435_comb = {{12{p2_add_74446[12]}}, p2_add_74446};
  assign p3_sum__1404_comb = {{12{p2_add_74447[12]}}, p2_add_74447};
  assign p3_sum__1405_comb = {{12{p2_add_74448[12]}}, p2_add_74448};
  assign p3_sum__1406_comb = {{12{p2_add_74449[12]}}, p2_add_74449};
  assign p3_sum__1407_comb = {{12{p2_add_74450[12]}}, p2_add_74450};
  assign p3_sum__1376_comb = {{12{p2_add_74451[12]}}, p2_add_74451};
  assign p3_sum__1377_comb = {{12{p2_add_74452[12]}}, p2_add_74452};
  assign p3_sum__1378_comb = {{12{p2_add_74453[12]}}, p2_add_74453};
  assign p3_sum__1379_comb = {{12{p2_add_74454[12]}}, p2_add_74454};
  assign p3_sum__1536_comb = {{12{p2_add_74491[12]}}, p2_add_74491};
  assign p3_sum__1537_comb = {{12{p2_add_74492[12]}}, p2_add_74492};
  assign p3_sum__1538_comb = {{12{p2_add_74493[12]}}, p2_add_74493};
  assign p3_sum__1539_comb = {{12{p2_add_74494[12]}}, p2_add_74494};
  assign p3_sum__1508_comb = {{12{p2_add_74495[12]}}, p2_add_74495};
  assign p3_sum__1509_comb = {{12{p2_add_74496[12]}}, p2_add_74496};
  assign p3_sum__1510_comb = {{12{p2_add_74497[12]}}, p2_add_74497};
  assign p3_sum__1511_comb = {{12{p2_add_74498[12]}}, p2_add_74498};
  assign p3_sum__1480_comb = {{12{p2_add_74499[12]}}, p2_add_74499};
  assign p3_sum__1481_comb = {{12{p2_add_74500[12]}}, p2_add_74500};
  assign p3_sum__1482_comb = {{12{p2_add_74501[12]}}, p2_add_74501};
  assign p3_sum__1483_comb = {{12{p2_add_74502[12]}}, p2_add_74502};
  assign p3_sum__1452_comb = {{12{p2_add_74503[12]}}, p2_add_74503};
  assign p3_sum__1453_comb = {{12{p2_add_74504[12]}}, p2_add_74504};
  assign p3_sum__1454_comb = {{12{p2_add_74505[12]}}, p2_add_74505};
  assign p3_sum__1455_comb = {{12{p2_add_74506[12]}}, p2_add_74506};
  assign p3_sum__1424_comb = {{12{p2_add_74507[12]}}, p2_add_74507};
  assign p3_sum__1425_comb = {{12{p2_add_74508[12]}}, p2_add_74508};
  assign p3_sum__1426_comb = {{12{p2_add_74509[12]}}, p2_add_74509};
  assign p3_sum__1427_comb = {{12{p2_add_74510[12]}}, p2_add_74510};
  assign p3_sum__1396_comb = {{12{p2_add_74511[12]}}, p2_add_74511};
  assign p3_sum__1397_comb = {{12{p2_add_74512[12]}}, p2_add_74512};
  assign p3_sum__1398_comb = {{12{p2_add_74513[12]}}, p2_add_74513};
  assign p3_sum__1399_comb = {{12{p2_add_74514[12]}}, p2_add_74514};
  assign p3_sum__1368_comb = {{12{p2_add_74515[12]}}, p2_add_74515};
  assign p3_sum__1369_comb = {{12{p2_add_74516[12]}}, p2_add_74516};
  assign p3_sum__1370_comb = {{12{p2_add_74517[12]}}, p2_add_74517};
  assign p3_sum__1371_comb = {{12{p2_add_74518[12]}}, p2_add_74518};
  assign p3_sum__1532_comb = {{12{p2_add_74523[12]}}, p2_add_74523};
  assign p3_sum__1533_comb = {{12{p2_add_74524[12]}}, p2_add_74524};
  assign p3_sum__1534_comb = {{12{p2_add_74525[12]}}, p2_add_74525};
  assign p3_sum__1535_comb = {{12{p2_add_74526[12]}}, p2_add_74526};
  assign p3_sum__1504_comb = {{12{p2_add_74527[12]}}, p2_add_74527};
  assign p3_sum__1505_comb = {{12{p2_add_74528[12]}}, p2_add_74528};
  assign p3_sum__1506_comb = {{12{p2_add_74529[12]}}, p2_add_74529};
  assign p3_sum__1507_comb = {{12{p2_add_74530[12]}}, p2_add_74530};
  assign p3_sum__1476_comb = {{12{p2_add_74531[12]}}, p2_add_74531};
  assign p3_sum__1477_comb = {{12{p2_add_74532[12]}}, p2_add_74532};
  assign p3_sum__1478_comb = {{12{p2_add_74533[12]}}, p2_add_74533};
  assign p3_sum__1479_comb = {{12{p2_add_74534[12]}}, p2_add_74534};
  assign p3_sum__1448_comb = {{12{p2_add_74535[12]}}, p2_add_74535};
  assign p3_sum__1449_comb = {{12{p2_add_74536[12]}}, p2_add_74536};
  assign p3_sum__1450_comb = {{12{p2_add_74537[12]}}, p2_add_74537};
  assign p3_sum__1451_comb = {{12{p2_add_74538[12]}}, p2_add_74538};
  assign p3_sum__1420_comb = {{12{p2_add_74539[12]}}, p2_add_74539};
  assign p3_sum__1421_comb = {{12{p2_add_74540[12]}}, p2_add_74540};
  assign p3_sum__1422_comb = {{12{p2_add_74541[12]}}, p2_add_74541};
  assign p3_sum__1423_comb = {{12{p2_add_74542[12]}}, p2_add_74542};
  assign p3_sum__1392_comb = {{12{p2_add_74543[12]}}, p2_add_74543};
  assign p3_sum__1393_comb = {{12{p2_add_74544[12]}}, p2_add_74544};
  assign p3_sum__1394_comb = {{12{p2_add_74545[12]}}, p2_add_74545};
  assign p3_sum__1395_comb = {{12{p2_add_74546[12]}}, p2_add_74546};
  assign p3_sum__1364_comb = {{12{p2_add_74547[12]}}, p2_add_74547};
  assign p3_sum__1365_comb = {{12{p2_add_74548[12]}}, p2_add_74548};
  assign p3_sum__1366_comb = {{12{p2_add_74549[12]}}, p2_add_74549};
  assign p3_sum__1367_comb = {{12{p2_add_74550[12]}}, p2_add_74550};
  assign p3_sum__1528_comb = {{12{p2_add_74555[12]}}, p2_add_74555};
  assign p3_sum__1529_comb = {{12{p2_add_74556[12]}}, p2_add_74556};
  assign p3_sum__1530_comb = {{12{p2_add_74557[12]}}, p2_add_74557};
  assign p3_sum__1531_comb = {{12{p2_add_74558[12]}}, p2_add_74558};
  assign p3_sum__1500_comb = {{12{p2_add_74559[12]}}, p2_add_74559};
  assign p3_sum__1501_comb = {{12{p2_add_74560[12]}}, p2_add_74560};
  assign p3_sum__1502_comb = {{12{p2_add_74561[12]}}, p2_add_74561};
  assign p3_sum__1503_comb = {{12{p2_add_74562[12]}}, p2_add_74562};
  assign p3_sum__1472_comb = {{12{p2_add_74563[12]}}, p2_add_74563};
  assign p3_sum__1473_comb = {{12{p2_add_74564[12]}}, p2_add_74564};
  assign p3_sum__1474_comb = {{12{p2_add_74565[12]}}, p2_add_74565};
  assign p3_sum__1475_comb = {{12{p2_add_74566[12]}}, p2_add_74566};
  assign p3_sum__1444_comb = {{12{p2_add_74567[12]}}, p2_add_74567};
  assign p3_sum__1445_comb = {{12{p2_add_74568[12]}}, p2_add_74568};
  assign p3_sum__1446_comb = {{12{p2_add_74569[12]}}, p2_add_74569};
  assign p3_sum__1447_comb = {{12{p2_add_74570[12]}}, p2_add_74570};
  assign p3_sum__1416_comb = {{12{p2_add_74571[12]}}, p2_add_74571};
  assign p3_sum__1417_comb = {{12{p2_add_74572[12]}}, p2_add_74572};
  assign p3_sum__1418_comb = {{12{p2_add_74573[12]}}, p2_add_74573};
  assign p3_sum__1419_comb = {{12{p2_add_74574[12]}}, p2_add_74574};
  assign p3_sum__1388_comb = {{12{p2_add_74575[12]}}, p2_add_74575};
  assign p3_sum__1389_comb = {{12{p2_add_74576[12]}}, p2_add_74576};
  assign p3_sum__1390_comb = {{12{p2_add_74577[12]}}, p2_add_74577};
  assign p3_sum__1391_comb = {{12{p2_add_74578[12]}}, p2_add_74578};
  assign p3_sum__1360_comb = {{12{p2_add_74579[12]}}, p2_add_74579};
  assign p3_sum__1361_comb = {{12{p2_add_74580[12]}}, p2_add_74580};
  assign p3_sum__1362_comb = {{12{p2_add_74581[12]}}, p2_add_74581};
  assign p3_sum__1363_comb = {{12{p2_add_74582[12]}}, p2_add_74582};
  assign p3_sum__1232_comb = p3_sum__1552_comb + p3_sum__1553_comb;
  assign p3_sum__1233_comb = p3_sum__1554_comb + p3_sum__1555_comb;
  assign p3_sum__1218_comb = p3_sum__1524_comb + p3_sum__1525_comb;
  assign p3_sum__1219_comb = p3_sum__1526_comb + p3_sum__1527_comb;
  assign p3_sum__1204_comb = p3_sum__1496_comb + p3_sum__1497_comb;
  assign p3_sum__1205_comb = p3_sum__1498_comb + p3_sum__1499_comb;
  assign p3_sum__1190_comb = p3_sum__1468_comb + p3_sum__1469_comb;
  assign p3_sum__1191_comb = p3_sum__1470_comb + p3_sum__1471_comb;
  assign p3_sum__1176_comb = p3_sum__1440_comb + p3_sum__1441_comb;
  assign p3_sum__1177_comb = p3_sum__1442_comb + p3_sum__1443_comb;
  assign p3_sum__1162_comb = p3_sum__1412_comb + p3_sum__1413_comb;
  assign p3_sum__1163_comb = p3_sum__1414_comb + p3_sum__1415_comb;
  assign p3_sum__1148_comb = p3_sum__1384_comb + p3_sum__1385_comb;
  assign p3_sum__1149_comb = p3_sum__1386_comb + p3_sum__1387_comb;
  assign p3_sum__1230_comb = p3_sum__1548_comb + p3_sum__1549_comb;
  assign p3_sum__1231_comb = p3_sum__1550_comb + p3_sum__1551_comb;
  assign p3_sum__1216_comb = p3_sum__1520_comb + p3_sum__1521_comb;
  assign p3_sum__1217_comb = p3_sum__1522_comb + p3_sum__1523_comb;
  assign p3_sum__1202_comb = p3_sum__1492_comb + p3_sum__1493_comb;
  assign p3_sum__1203_comb = p3_sum__1494_comb + p3_sum__1495_comb;
  assign p3_sum__1188_comb = p3_sum__1464_comb + p3_sum__1465_comb;
  assign p3_sum__1189_comb = p3_sum__1466_comb + p3_sum__1467_comb;
  assign p3_sum__1174_comb = p3_sum__1436_comb + p3_sum__1437_comb;
  assign p3_sum__1175_comb = p3_sum__1438_comb + p3_sum__1439_comb;
  assign p3_sum__1160_comb = p3_sum__1408_comb + p3_sum__1409_comb;
  assign p3_sum__1161_comb = p3_sum__1410_comb + p3_sum__1411_comb;
  assign p3_sum__1146_comb = p3_sum__1380_comb + p3_sum__1381_comb;
  assign p3_sum__1147_comb = p3_sum__1382_comb + p3_sum__1383_comb;
  assign p3_sum__1228_comb = p3_sum__1544_comb + p3_sum__1545_comb;
  assign p3_sum__1229_comb = p3_sum__1546_comb + p3_sum__1547_comb;
  assign p3_sum__1214_comb = p3_sum__1516_comb + p3_sum__1517_comb;
  assign p3_sum__1215_comb = p3_sum__1518_comb + p3_sum__1519_comb;
  assign p3_sum__1200_comb = p3_sum__1488_comb + p3_sum__1489_comb;
  assign p3_sum__1201_comb = p3_sum__1490_comb + p3_sum__1491_comb;
  assign p3_sum__1186_comb = p3_sum__1460_comb + p3_sum__1461_comb;
  assign p3_sum__1187_comb = p3_sum__1462_comb + p3_sum__1463_comb;
  assign p3_sum__1172_comb = p3_sum__1432_comb + p3_sum__1433_comb;
  assign p3_sum__1173_comb = p3_sum__1434_comb + p3_sum__1435_comb;
  assign p3_sum__1158_comb = p3_sum__1404_comb + p3_sum__1405_comb;
  assign p3_sum__1159_comb = p3_sum__1406_comb + p3_sum__1407_comb;
  assign p3_sum__1144_comb = p3_sum__1376_comb + p3_sum__1377_comb;
  assign p3_sum__1145_comb = p3_sum__1378_comb + p3_sum__1379_comb;
  assign p3_sum__1224_comb = p3_sum__1536_comb + p3_sum__1537_comb;
  assign p3_sum__1225_comb = p3_sum__1538_comb + p3_sum__1539_comb;
  assign p3_sum__1210_comb = p3_sum__1508_comb + p3_sum__1509_comb;
  assign p3_sum__1211_comb = p3_sum__1510_comb + p3_sum__1511_comb;
  assign p3_sum__1196_comb = p3_sum__1480_comb + p3_sum__1481_comb;
  assign p3_sum__1197_comb = p3_sum__1482_comb + p3_sum__1483_comb;
  assign p3_sum__1182_comb = p3_sum__1452_comb + p3_sum__1453_comb;
  assign p3_sum__1183_comb = p3_sum__1454_comb + p3_sum__1455_comb;
  assign p3_sum__1168_comb = p3_sum__1424_comb + p3_sum__1425_comb;
  assign p3_sum__1169_comb = p3_sum__1426_comb + p3_sum__1427_comb;
  assign p3_sum__1154_comb = p3_sum__1396_comb + p3_sum__1397_comb;
  assign p3_sum__1155_comb = p3_sum__1398_comb + p3_sum__1399_comb;
  assign p3_sum__1140_comb = p3_sum__1368_comb + p3_sum__1369_comb;
  assign p3_sum__1141_comb = p3_sum__1370_comb + p3_sum__1371_comb;
  assign p3_sum__1222_comb = p3_sum__1532_comb + p3_sum__1533_comb;
  assign p3_sum__1223_comb = p3_sum__1534_comb + p3_sum__1535_comb;
  assign p3_sum__1208_comb = p3_sum__1504_comb + p3_sum__1505_comb;
  assign p3_sum__1209_comb = p3_sum__1506_comb + p3_sum__1507_comb;
  assign p3_sum__1194_comb = p3_sum__1476_comb + p3_sum__1477_comb;
  assign p3_sum__1195_comb = p3_sum__1478_comb + p3_sum__1479_comb;
  assign p3_sum__1180_comb = p3_sum__1448_comb + p3_sum__1449_comb;
  assign p3_sum__1181_comb = p3_sum__1450_comb + p3_sum__1451_comb;
  assign p3_sum__1166_comb = p3_sum__1420_comb + p3_sum__1421_comb;
  assign p3_sum__1167_comb = p3_sum__1422_comb + p3_sum__1423_comb;
  assign p3_sum__1152_comb = p3_sum__1392_comb + p3_sum__1393_comb;
  assign p3_sum__1153_comb = p3_sum__1394_comb + p3_sum__1395_comb;
  assign p3_sum__1138_comb = p3_sum__1364_comb + p3_sum__1365_comb;
  assign p3_sum__1139_comb = p3_sum__1366_comb + p3_sum__1367_comb;
  assign p3_sum__1220_comb = p3_sum__1528_comb + p3_sum__1529_comb;
  assign p3_sum__1221_comb = p3_sum__1530_comb + p3_sum__1531_comb;
  assign p3_sum__1206_comb = p3_sum__1500_comb + p3_sum__1501_comb;
  assign p3_sum__1207_comb = p3_sum__1502_comb + p3_sum__1503_comb;
  assign p3_sum__1192_comb = p3_sum__1472_comb + p3_sum__1473_comb;
  assign p3_sum__1193_comb = p3_sum__1474_comb + p3_sum__1475_comb;
  assign p3_sum__1178_comb = p3_sum__1444_comb + p3_sum__1445_comb;
  assign p3_sum__1179_comb = p3_sum__1446_comb + p3_sum__1447_comb;
  assign p3_sum__1164_comb = p3_sum__1416_comb + p3_sum__1417_comb;
  assign p3_sum__1165_comb = p3_sum__1418_comb + p3_sum__1419_comb;
  assign p3_sum__1150_comb = p3_sum__1388_comb + p3_sum__1389_comb;
  assign p3_sum__1151_comb = p3_sum__1390_comb + p3_sum__1391_comb;
  assign p3_sum__1136_comb = p3_sum__1360_comb + p3_sum__1361_comb;
  assign p3_sum__1137_comb = p3_sum__1362_comb + p3_sum__1363_comb;
  assign p3_sum__1072_comb = p3_sum__1232_comb + p3_sum__1233_comb;
  assign p3_sum__1065_comb = p3_sum__1218_comb + p3_sum__1219_comb;
  assign p3_sum__1058_comb = p3_sum__1204_comb + p3_sum__1205_comb;
  assign p3_sum__1051_comb = p3_sum__1190_comb + p3_sum__1191_comb;
  assign p3_sum__1044_comb = p3_sum__1176_comb + p3_sum__1177_comb;
  assign p3_sum__1037_comb = p3_sum__1162_comb + p3_sum__1163_comb;
  assign p3_sum__1030_comb = p3_sum__1148_comb + p3_sum__1149_comb;
  assign p3_sum__1071_comb = p3_sum__1230_comb + p3_sum__1231_comb;
  assign p3_sum__1064_comb = p3_sum__1216_comb + p3_sum__1217_comb;
  assign p3_sum__1057_comb = p3_sum__1202_comb + p3_sum__1203_comb;
  assign p3_sum__1050_comb = p3_sum__1188_comb + p3_sum__1189_comb;
  assign p3_sum__1043_comb = p3_sum__1174_comb + p3_sum__1175_comb;
  assign p3_sum__1036_comb = p3_sum__1160_comb + p3_sum__1161_comb;
  assign p3_sum__1029_comb = p3_sum__1146_comb + p3_sum__1147_comb;
  assign p3_sum__1070_comb = p3_sum__1228_comb + p3_sum__1229_comb;
  assign p3_sum__1063_comb = p3_sum__1214_comb + p3_sum__1215_comb;
  assign p3_sum__1056_comb = p3_sum__1200_comb + p3_sum__1201_comb;
  assign p3_sum__1049_comb = p3_sum__1186_comb + p3_sum__1187_comb;
  assign p3_sum__1042_comb = p3_sum__1172_comb + p3_sum__1173_comb;
  assign p3_sum__1035_comb = p3_sum__1158_comb + p3_sum__1159_comb;
  assign p3_sum__1028_comb = p3_sum__1144_comb + p3_sum__1145_comb;
  assign p3_sum__1069_comb = p2_sum__1226 + p2_sum__1227;
  assign p3_sum__1062_comb = p2_sum__1212 + p2_sum__1213;
  assign p3_sum__1055_comb = p2_sum__1198 + p2_sum__1199;
  assign p3_sum__1048_comb = p2_sum__1184 + p2_sum__1185;
  assign p3_sum__1041_comb = p2_sum__1170 + p2_sum__1171;
  assign p3_sum__1034_comb = p2_sum__1156 + p2_sum__1157;
  assign p3_sum__1027_comb = p2_sum__1142 + p2_sum__1143;
  assign p3_sum__1068_comb = p3_sum__1224_comb + p3_sum__1225_comb;
  assign p3_sum__1061_comb = p3_sum__1210_comb + p3_sum__1211_comb;
  assign p3_sum__1054_comb = p3_sum__1196_comb + p3_sum__1197_comb;
  assign p3_sum__1047_comb = p3_sum__1182_comb + p3_sum__1183_comb;
  assign p3_sum__1040_comb = p3_sum__1168_comb + p3_sum__1169_comb;
  assign p3_sum__1033_comb = p3_sum__1154_comb + p3_sum__1155_comb;
  assign p3_sum__1026_comb = p3_sum__1140_comb + p3_sum__1141_comb;
  assign p3_sum__1067_comb = p3_sum__1222_comb + p3_sum__1223_comb;
  assign p3_sum__1060_comb = p3_sum__1208_comb + p3_sum__1209_comb;
  assign p3_sum__1053_comb = p3_sum__1194_comb + p3_sum__1195_comb;
  assign p3_sum__1046_comb = p3_sum__1180_comb + p3_sum__1181_comb;
  assign p3_sum__1039_comb = p3_sum__1166_comb + p3_sum__1167_comb;
  assign p3_sum__1032_comb = p3_sum__1152_comb + p3_sum__1153_comb;
  assign p3_sum__1025_comb = p3_sum__1138_comb + p3_sum__1139_comb;
  assign p3_sum__1066_comb = p3_sum__1220_comb + p3_sum__1221_comb;
  assign p3_sum__1059_comb = p3_sum__1206_comb + p3_sum__1207_comb;
  assign p3_sum__1052_comb = p3_sum__1192_comb + p3_sum__1193_comb;
  assign p3_sum__1045_comb = p3_sum__1178_comb + p3_sum__1179_comb;
  assign p3_sum__1038_comb = p3_sum__1164_comb + p3_sum__1165_comb;
  assign p3_sum__1031_comb = p3_sum__1150_comb + p3_sum__1151_comb;
  assign p3_sum__1024_comb = p3_sum__1136_comb + p3_sum__1137_comb;
  assign p3_add_75467_comb = p2_bit_slice_74693 + 25'h000_0001;
  assign p3_add_75468_comb = p2_bit_slice_74694 + 25'h000_0001;
  assign p3_add_75469_comb = p2_bit_slice_74695 + 25'h000_0001;
  assign p3_add_75470_comb = p2_bit_slice_74696 + 25'h000_0001;
  assign p3_add_75471_comb = p2_bit_slice_74697 + 25'h000_0001;
  assign p3_add_75472_comb = p2_bit_slice_74698 + 25'h000_0001;
  assign p3_add_75473_comb = p2_bit_slice_74699 + 25'h000_0001;
  assign p3_add_75474_comb = p2_sum__1079 + 25'h000_0001;
  assign p3_add_75475_comb = p3_sum__1072_comb + 25'h000_0001;
  assign p3_add_75476_comb = p3_sum__1065_comb + 25'h000_0001;
  assign p3_add_75477_comb = p3_sum__1058_comb + 25'h000_0001;
  assign p3_add_75478_comb = p3_sum__1051_comb + 25'h000_0001;
  assign p3_add_75479_comb = p3_sum__1044_comb + 25'h000_0001;
  assign p3_add_75480_comb = p3_sum__1037_comb + 25'h000_0001;
  assign p3_add_75481_comb = p3_sum__1030_comb + 25'h000_0001;
  assign p3_add_75482_comb = p2_sum__1078 + 25'h000_0001;
  assign p3_add_75483_comb = p3_sum__1071_comb + 25'h000_0001;
  assign p3_add_75484_comb = p3_sum__1064_comb + 25'h000_0001;
  assign p3_add_75485_comb = p3_sum__1057_comb + 25'h000_0001;
  assign p3_add_75486_comb = p3_sum__1050_comb + 25'h000_0001;
  assign p3_add_75487_comb = p3_sum__1043_comb + 25'h000_0001;
  assign p3_add_75488_comb = p3_sum__1036_comb + 25'h000_0001;
  assign p3_add_75489_comb = p3_sum__1029_comb + 25'h000_0001;
  assign p3_add_75490_comb = p2_sum__1077 + 25'h000_0001;
  assign p3_add_75491_comb = p3_sum__1070_comb + 25'h000_0001;
  assign p3_add_75492_comb = p3_sum__1063_comb + 25'h000_0001;
  assign p3_add_75493_comb = p3_sum__1056_comb + 25'h000_0001;
  assign p3_add_75494_comb = p3_sum__1049_comb + 25'h000_0001;
  assign p3_add_75495_comb = p3_sum__1042_comb + 25'h000_0001;
  assign p3_add_75496_comb = p3_sum__1035_comb + 25'h000_0001;
  assign p3_add_75497_comb = p3_sum__1028_comb + 25'h000_0001;
  assign p3_add_75498_comb = p3_sum__1069_comb + 25'h000_0001;
  assign p3_add_75499_comb = p3_sum__1062_comb + 25'h000_0001;
  assign p3_add_75500_comb = p3_sum__1055_comb + 25'h000_0001;
  assign p3_add_75501_comb = p3_sum__1048_comb + 25'h000_0001;
  assign p3_add_75502_comb = p3_sum__1041_comb + 25'h000_0001;
  assign p3_add_75503_comb = p3_sum__1034_comb + 25'h000_0001;
  assign p3_add_75504_comb = p3_sum__1027_comb + 25'h000_0001;
  assign p3_add_75505_comb = p2_sum__1075 + 25'h000_0001;
  assign p3_add_75506_comb = p3_sum__1068_comb + 25'h000_0001;
  assign p3_add_75507_comb = p3_sum__1061_comb + 25'h000_0001;
  assign p3_add_75508_comb = p3_sum__1054_comb + 25'h000_0001;
  assign p3_add_75509_comb = p3_sum__1047_comb + 25'h000_0001;
  assign p3_add_75510_comb = p3_sum__1040_comb + 25'h000_0001;
  assign p3_add_75511_comb = p3_sum__1033_comb + 25'h000_0001;
  assign p3_add_75512_comb = p3_sum__1026_comb + 25'h000_0001;
  assign p3_add_75513_comb = p2_sum__1074 + 25'h000_0001;
  assign p3_add_75514_comb = p3_sum__1067_comb + 25'h000_0001;
  assign p3_add_75515_comb = p3_sum__1060_comb + 25'h000_0001;
  assign p3_add_75516_comb = p3_sum__1053_comb + 25'h000_0001;
  assign p3_add_75517_comb = p3_sum__1046_comb + 25'h000_0001;
  assign p3_add_75518_comb = p3_sum__1039_comb + 25'h000_0001;
  assign p3_add_75519_comb = p3_sum__1032_comb + 25'h000_0001;
  assign p3_add_75520_comb = p3_sum__1025_comb + 25'h000_0001;
  assign p3_add_75521_comb = p2_sum__1073 + 25'h000_0001;
  assign p3_add_75522_comb = p3_sum__1066_comb + 25'h000_0001;
  assign p3_add_75523_comb = p3_sum__1059_comb + 25'h000_0001;
  assign p3_add_75524_comb = p3_sum__1052_comb + 25'h000_0001;
  assign p3_add_75525_comb = p3_sum__1045_comb + 25'h000_0001;
  assign p3_add_75526_comb = p3_sum__1038_comb + 25'h000_0001;
  assign p3_add_75527_comb = p3_sum__1031_comb + 25'h000_0001;
  assign p3_add_75528_comb = p3_sum__1024_comb + 25'h000_0001;
  assign p3_clipped__136_comb = $signed(p2_add_74708[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p2_add_74708[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p2_add_74708[12:1]);
  assign p3_clipped__152_comb = $signed(p3_add_75467_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75467_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75467_comb[12:1]);
  assign p3_clipped__168_comb = $signed(p3_add_75468_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75468_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75468_comb[12:1]);
  assign p3_clipped__184_comb = $signed(p3_add_75469_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75469_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75469_comb[12:1]);
  assign p3_clipped__200_comb = $signed(p3_add_75470_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75470_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75470_comb[12:1]);
  assign p3_clipped__216_comb = $signed(p3_add_75471_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75471_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75471_comb[12:1]);
  assign p3_clipped__232_comb = $signed(p3_add_75472_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75472_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75472_comb[12:1]);
  assign p3_clipped__248_comb = $signed(p3_add_75473_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75473_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75473_comb[12:1]);
  assign p3_clipped__137_comb = $signed(p3_add_75474_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75474_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75474_comb[12:1]);
  assign p3_clipped__153_comb = $signed(p3_add_75475_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75475_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75475_comb[12:1]);
  assign p3_clipped__169_comb = $signed(p3_add_75476_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75476_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75476_comb[12:1]);
  assign p3_clipped__185_comb = $signed(p3_add_75477_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75477_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75477_comb[12:1]);
  assign p3_clipped__201_comb = $signed(p3_add_75478_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75478_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75478_comb[12:1]);
  assign p3_clipped__217_comb = $signed(p3_add_75479_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75479_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75479_comb[12:1]);
  assign p3_clipped__233_comb = $signed(p3_add_75480_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75480_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75480_comb[12:1]);
  assign p3_clipped__249_comb = $signed(p3_add_75481_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75481_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75481_comb[12:1]);
  assign p3_clipped__138_comb = $signed(p3_add_75482_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75482_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75482_comb[12:1]);
  assign p3_clipped__154_comb = $signed(p3_add_75483_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75483_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75483_comb[12:1]);
  assign p3_clipped__170_comb = $signed(p3_add_75484_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75484_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75484_comb[12:1]);
  assign p3_clipped__186_comb = $signed(p3_add_75485_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75485_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75485_comb[12:1]);
  assign p3_clipped__202_comb = $signed(p3_add_75486_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75486_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75486_comb[12:1]);
  assign p3_clipped__218_comb = $signed(p3_add_75487_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75487_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75487_comb[12:1]);
  assign p3_clipped__234_comb = $signed(p3_add_75488_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75488_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75488_comb[12:1]);
  assign p3_clipped__250_comb = $signed(p3_add_75489_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75489_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75489_comb[12:1]);
  assign p3_clipped__139_comb = $signed(p3_add_75490_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75490_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75490_comb[12:1]);
  assign p3_clipped__155_comb = $signed(p3_add_75491_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75491_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75491_comb[12:1]);
  assign p3_clipped__171_comb = $signed(p3_add_75492_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75492_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75492_comb[12:1]);
  assign p3_clipped__187_comb = $signed(p3_add_75493_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75493_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75493_comb[12:1]);
  assign p3_clipped__203_comb = $signed(p3_add_75494_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75494_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75494_comb[12:1]);
  assign p3_clipped__219_comb = $signed(p3_add_75495_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75495_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75495_comb[12:1]);
  assign p3_clipped__235_comb = $signed(p3_add_75496_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75496_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75496_comb[12:1]);
  assign p3_clipped__251_comb = $signed(p3_add_75497_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75497_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75497_comb[12:1]);
  assign p3_clipped__140_comb = $signed(p2_add_74709[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p2_add_74709[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p2_add_74709[12:1]);
  assign p3_clipped__156_comb = $signed(p3_add_75498_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75498_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75498_comb[12:1]);
  assign p3_clipped__172_comb = $signed(p3_add_75499_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75499_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75499_comb[12:1]);
  assign p3_clipped__188_comb = $signed(p3_add_75500_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75500_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75500_comb[12:1]);
  assign p3_clipped__204_comb = $signed(p3_add_75501_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75501_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75501_comb[12:1]);
  assign p3_clipped__220_comb = $signed(p3_add_75502_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75502_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75502_comb[12:1]);
  assign p3_clipped__236_comb = $signed(p3_add_75503_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75503_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75503_comb[12:1]);
  assign p3_clipped__252_comb = $signed(p3_add_75504_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75504_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75504_comb[12:1]);
  assign p3_clipped__141_comb = $signed(p3_add_75505_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75505_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75505_comb[12:1]);
  assign p3_clipped__157_comb = $signed(p3_add_75506_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75506_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75506_comb[12:1]);
  assign p3_clipped__173_comb = $signed(p3_add_75507_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75507_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75507_comb[12:1]);
  assign p3_clipped__189_comb = $signed(p3_add_75508_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75508_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75508_comb[12:1]);
  assign p3_clipped__205_comb = $signed(p3_add_75509_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75509_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75509_comb[12:1]);
  assign p3_clipped__221_comb = $signed(p3_add_75510_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75510_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75510_comb[12:1]);
  assign p3_clipped__237_comb = $signed(p3_add_75511_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75511_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75511_comb[12:1]);
  assign p3_clipped__253_comb = $signed(p3_add_75512_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75512_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75512_comb[12:1]);
  assign p3_clipped__142_comb = $signed(p3_add_75513_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75513_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75513_comb[12:1]);
  assign p3_clipped__158_comb = $signed(p3_add_75514_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75514_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75514_comb[12:1]);
  assign p3_clipped__174_comb = $signed(p3_add_75515_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75515_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75515_comb[12:1]);
  assign p3_clipped__190_comb = $signed(p3_add_75516_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75516_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75516_comb[12:1]);
  assign p3_clipped__206_comb = $signed(p3_add_75517_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75517_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75517_comb[12:1]);
  assign p3_clipped__222_comb = $signed(p3_add_75518_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75518_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75518_comb[12:1]);
  assign p3_clipped__238_comb = $signed(p3_add_75519_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75519_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75519_comb[12:1]);
  assign p3_clipped__254_comb = $signed(p3_add_75520_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75520_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75520_comb[12:1]);
  assign p3_clipped__143_comb = $signed(p3_add_75521_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75521_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75521_comb[12:1]);
  assign p3_clipped__159_comb = $signed(p3_add_75522_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75522_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75522_comb[12:1]);
  assign p3_clipped__175_comb = $signed(p3_add_75523_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75523_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75523_comb[12:1]);
  assign p3_clipped__191_comb = $signed(p3_add_75524_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75524_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75524_comb[12:1]);
  assign p3_clipped__207_comb = $signed(p3_add_75525_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75525_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75525_comb[12:1]);
  assign p3_clipped__223_comb = $signed(p3_add_75526_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75526_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75526_comb[12:1]);
  assign p3_clipped__239_comb = $signed(p3_add_75527_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75527_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75527_comb[12:1]);
  assign p3_clipped__255_comb = $signed(p3_add_75528_comb[24:1]) < $signed(24'hff_f800) ? 12'h800 : ($signed(p3_add_75528_comb[24:1]) > $signed(24'h00_07ff) ? 12'h7ff : p3_add_75528_comb[12:1]);
  assign p3_array_76169_comb[0] = p3_clipped__136_comb;
  assign p3_array_76169_comb[1] = p3_clipped__152_comb;
  assign p3_array_76169_comb[2] = p3_clipped__168_comb;
  assign p3_array_76169_comb[3] = p3_clipped__184_comb;
  assign p3_array_76169_comb[4] = p3_clipped__200_comb;
  assign p3_array_76169_comb[5] = p3_clipped__216_comb;
  assign p3_array_76169_comb[6] = p3_clipped__232_comb;
  assign p3_array_76169_comb[7] = p3_clipped__248_comb;
  assign p3_array_76170_comb[0] = p3_clipped__137_comb;
  assign p3_array_76170_comb[1] = p3_clipped__153_comb;
  assign p3_array_76170_comb[2] = p3_clipped__169_comb;
  assign p3_array_76170_comb[3] = p3_clipped__185_comb;
  assign p3_array_76170_comb[4] = p3_clipped__201_comb;
  assign p3_array_76170_comb[5] = p3_clipped__217_comb;
  assign p3_array_76170_comb[6] = p3_clipped__233_comb;
  assign p3_array_76170_comb[7] = p3_clipped__249_comb;
  assign p3_array_76171_comb[0] = p3_clipped__138_comb;
  assign p3_array_76171_comb[1] = p3_clipped__154_comb;
  assign p3_array_76171_comb[2] = p3_clipped__170_comb;
  assign p3_array_76171_comb[3] = p3_clipped__186_comb;
  assign p3_array_76171_comb[4] = p3_clipped__202_comb;
  assign p3_array_76171_comb[5] = p3_clipped__218_comb;
  assign p3_array_76171_comb[6] = p3_clipped__234_comb;
  assign p3_array_76171_comb[7] = p3_clipped__250_comb;
  assign p3_array_76172_comb[0] = p3_clipped__139_comb;
  assign p3_array_76172_comb[1] = p3_clipped__155_comb;
  assign p3_array_76172_comb[2] = p3_clipped__171_comb;
  assign p3_array_76172_comb[3] = p3_clipped__187_comb;
  assign p3_array_76172_comb[4] = p3_clipped__203_comb;
  assign p3_array_76172_comb[5] = p3_clipped__219_comb;
  assign p3_array_76172_comb[6] = p3_clipped__235_comb;
  assign p3_array_76172_comb[7] = p3_clipped__251_comb;
  assign p3_array_76173_comb[0] = p3_clipped__140_comb;
  assign p3_array_76173_comb[1] = p3_clipped__156_comb;
  assign p3_array_76173_comb[2] = p3_clipped__172_comb;
  assign p3_array_76173_comb[3] = p3_clipped__188_comb;
  assign p3_array_76173_comb[4] = p3_clipped__204_comb;
  assign p3_array_76173_comb[5] = p3_clipped__220_comb;
  assign p3_array_76173_comb[6] = p3_clipped__236_comb;
  assign p3_array_76173_comb[7] = p3_clipped__252_comb;
  assign p3_array_76174_comb[0] = p3_clipped__141_comb;
  assign p3_array_76174_comb[1] = p3_clipped__157_comb;
  assign p3_array_76174_comb[2] = p3_clipped__173_comb;
  assign p3_array_76174_comb[3] = p3_clipped__189_comb;
  assign p3_array_76174_comb[4] = p3_clipped__205_comb;
  assign p3_array_76174_comb[5] = p3_clipped__221_comb;
  assign p3_array_76174_comb[6] = p3_clipped__237_comb;
  assign p3_array_76174_comb[7] = p3_clipped__253_comb;
  assign p3_array_76175_comb[0] = p3_clipped__142_comb;
  assign p3_array_76175_comb[1] = p3_clipped__158_comb;
  assign p3_array_76175_comb[2] = p3_clipped__174_comb;
  assign p3_array_76175_comb[3] = p3_clipped__190_comb;
  assign p3_array_76175_comb[4] = p3_clipped__206_comb;
  assign p3_array_76175_comb[5] = p3_clipped__222_comb;
  assign p3_array_76175_comb[6] = p3_clipped__238_comb;
  assign p3_array_76175_comb[7] = p3_clipped__254_comb;
  assign p3_array_76176_comb[0] = p3_clipped__143_comb;
  assign p3_array_76176_comb[1] = p3_clipped__159_comb;
  assign p3_array_76176_comb[2] = p3_clipped__175_comb;
  assign p3_array_76176_comb[3] = p3_clipped__191_comb;
  assign p3_array_76176_comb[4] = p3_clipped__207_comb;
  assign p3_array_76176_comb[5] = p3_clipped__223_comb;
  assign p3_array_76176_comb[6] = p3_clipped__239_comb;
  assign p3_array_76176_comb[7] = p3_clipped__255_comb;
  assign p3_col_transformed_comb[0][0] = p3_array_76169_comb[0];
  assign p3_col_transformed_comb[0][1] = p3_array_76169_comb[1];
  assign p3_col_transformed_comb[0][2] = p3_array_76169_comb[2];
  assign p3_col_transformed_comb[0][3] = p3_array_76169_comb[3];
  assign p3_col_transformed_comb[0][4] = p3_array_76169_comb[4];
  assign p3_col_transformed_comb[0][5] = p3_array_76169_comb[5];
  assign p3_col_transformed_comb[0][6] = p3_array_76169_comb[6];
  assign p3_col_transformed_comb[0][7] = p3_array_76169_comb[7];
  assign p3_col_transformed_comb[1][0] = p3_array_76170_comb[0];
  assign p3_col_transformed_comb[1][1] = p3_array_76170_comb[1];
  assign p3_col_transformed_comb[1][2] = p3_array_76170_comb[2];
  assign p3_col_transformed_comb[1][3] = p3_array_76170_comb[3];
  assign p3_col_transformed_comb[1][4] = p3_array_76170_comb[4];
  assign p3_col_transformed_comb[1][5] = p3_array_76170_comb[5];
  assign p3_col_transformed_comb[1][6] = p3_array_76170_comb[6];
  assign p3_col_transformed_comb[1][7] = p3_array_76170_comb[7];
  assign p3_col_transformed_comb[2][0] = p3_array_76171_comb[0];
  assign p3_col_transformed_comb[2][1] = p3_array_76171_comb[1];
  assign p3_col_transformed_comb[2][2] = p3_array_76171_comb[2];
  assign p3_col_transformed_comb[2][3] = p3_array_76171_comb[3];
  assign p3_col_transformed_comb[2][4] = p3_array_76171_comb[4];
  assign p3_col_transformed_comb[2][5] = p3_array_76171_comb[5];
  assign p3_col_transformed_comb[2][6] = p3_array_76171_comb[6];
  assign p3_col_transformed_comb[2][7] = p3_array_76171_comb[7];
  assign p3_col_transformed_comb[3][0] = p3_array_76172_comb[0];
  assign p3_col_transformed_comb[3][1] = p3_array_76172_comb[1];
  assign p3_col_transformed_comb[3][2] = p3_array_76172_comb[2];
  assign p3_col_transformed_comb[3][3] = p3_array_76172_comb[3];
  assign p3_col_transformed_comb[3][4] = p3_array_76172_comb[4];
  assign p3_col_transformed_comb[3][5] = p3_array_76172_comb[5];
  assign p3_col_transformed_comb[3][6] = p3_array_76172_comb[6];
  assign p3_col_transformed_comb[3][7] = p3_array_76172_comb[7];
  assign p3_col_transformed_comb[4][0] = p3_array_76173_comb[0];
  assign p3_col_transformed_comb[4][1] = p3_array_76173_comb[1];
  assign p3_col_transformed_comb[4][2] = p3_array_76173_comb[2];
  assign p3_col_transformed_comb[4][3] = p3_array_76173_comb[3];
  assign p3_col_transformed_comb[4][4] = p3_array_76173_comb[4];
  assign p3_col_transformed_comb[4][5] = p3_array_76173_comb[5];
  assign p3_col_transformed_comb[4][6] = p3_array_76173_comb[6];
  assign p3_col_transformed_comb[4][7] = p3_array_76173_comb[7];
  assign p3_col_transformed_comb[5][0] = p3_array_76174_comb[0];
  assign p3_col_transformed_comb[5][1] = p3_array_76174_comb[1];
  assign p3_col_transformed_comb[5][2] = p3_array_76174_comb[2];
  assign p3_col_transformed_comb[5][3] = p3_array_76174_comb[3];
  assign p3_col_transformed_comb[5][4] = p3_array_76174_comb[4];
  assign p3_col_transformed_comb[5][5] = p3_array_76174_comb[5];
  assign p3_col_transformed_comb[5][6] = p3_array_76174_comb[6];
  assign p3_col_transformed_comb[5][7] = p3_array_76174_comb[7];
  assign p3_col_transformed_comb[6][0] = p3_array_76175_comb[0];
  assign p3_col_transformed_comb[6][1] = p3_array_76175_comb[1];
  assign p3_col_transformed_comb[6][2] = p3_array_76175_comb[2];
  assign p3_col_transformed_comb[6][3] = p3_array_76175_comb[3];
  assign p3_col_transformed_comb[6][4] = p3_array_76175_comb[4];
  assign p3_col_transformed_comb[6][5] = p3_array_76175_comb[5];
  assign p3_col_transformed_comb[6][6] = p3_array_76175_comb[6];
  assign p3_col_transformed_comb[6][7] = p3_array_76175_comb[7];
  assign p3_col_transformed_comb[7][0] = p3_array_76176_comb[0];
  assign p3_col_transformed_comb[7][1] = p3_array_76176_comb[1];
  assign p3_col_transformed_comb[7][2] = p3_array_76176_comb[2];
  assign p3_col_transformed_comb[7][3] = p3_array_76176_comb[3];
  assign p3_col_transformed_comb[7][4] = p3_array_76176_comb[4];
  assign p3_col_transformed_comb[7][5] = p3_array_76176_comb[5];
  assign p3_col_transformed_comb[7][6] = p3_array_76176_comb[6];
  assign p3_col_transformed_comb[7][7] = p3_array_76176_comb[7];

  // Registers for pipe stage 3:
  reg [11:0] p3_col_transformed[0:7][0:7];
  always @ (posedge clk) begin
    p3_col_transformed[0][0] <= p3_col_transformed_comb[0][0];
    p3_col_transformed[0][1] <= p3_col_transformed_comb[0][1];
    p3_col_transformed[0][2] <= p3_col_transformed_comb[0][2];
    p3_col_transformed[0][3] <= p3_col_transformed_comb[0][3];
    p3_col_transformed[0][4] <= p3_col_transformed_comb[0][4];
    p3_col_transformed[0][5] <= p3_col_transformed_comb[0][5];
    p3_col_transformed[0][6] <= p3_col_transformed_comb[0][6];
    p3_col_transformed[0][7] <= p3_col_transformed_comb[0][7];
    p3_col_transformed[1][0] <= p3_col_transformed_comb[1][0];
    p3_col_transformed[1][1] <= p3_col_transformed_comb[1][1];
    p3_col_transformed[1][2] <= p3_col_transformed_comb[1][2];
    p3_col_transformed[1][3] <= p3_col_transformed_comb[1][3];
    p3_col_transformed[1][4] <= p3_col_transformed_comb[1][4];
    p3_col_transformed[1][5] <= p3_col_transformed_comb[1][5];
    p3_col_transformed[1][6] <= p3_col_transformed_comb[1][6];
    p3_col_transformed[1][7] <= p3_col_transformed_comb[1][7];
    p3_col_transformed[2][0] <= p3_col_transformed_comb[2][0];
    p3_col_transformed[2][1] <= p3_col_transformed_comb[2][1];
    p3_col_transformed[2][2] <= p3_col_transformed_comb[2][2];
    p3_col_transformed[2][3] <= p3_col_transformed_comb[2][3];
    p3_col_transformed[2][4] <= p3_col_transformed_comb[2][4];
    p3_col_transformed[2][5] <= p3_col_transformed_comb[2][5];
    p3_col_transformed[2][6] <= p3_col_transformed_comb[2][6];
    p3_col_transformed[2][7] <= p3_col_transformed_comb[2][7];
    p3_col_transformed[3][0] <= p3_col_transformed_comb[3][0];
    p3_col_transformed[3][1] <= p3_col_transformed_comb[3][1];
    p3_col_transformed[3][2] <= p3_col_transformed_comb[3][2];
    p3_col_transformed[3][3] <= p3_col_transformed_comb[3][3];
    p3_col_transformed[3][4] <= p3_col_transformed_comb[3][4];
    p3_col_transformed[3][5] <= p3_col_transformed_comb[3][5];
    p3_col_transformed[3][6] <= p3_col_transformed_comb[3][6];
    p3_col_transformed[3][7] <= p3_col_transformed_comb[3][7];
    p3_col_transformed[4][0] <= p3_col_transformed_comb[4][0];
    p3_col_transformed[4][1] <= p3_col_transformed_comb[4][1];
    p3_col_transformed[4][2] <= p3_col_transformed_comb[4][2];
    p3_col_transformed[4][3] <= p3_col_transformed_comb[4][3];
    p3_col_transformed[4][4] <= p3_col_transformed_comb[4][4];
    p3_col_transformed[4][5] <= p3_col_transformed_comb[4][5];
    p3_col_transformed[4][6] <= p3_col_transformed_comb[4][6];
    p3_col_transformed[4][7] <= p3_col_transformed_comb[4][7];
    p3_col_transformed[5][0] <= p3_col_transformed_comb[5][0];
    p3_col_transformed[5][1] <= p3_col_transformed_comb[5][1];
    p3_col_transformed[5][2] <= p3_col_transformed_comb[5][2];
    p3_col_transformed[5][3] <= p3_col_transformed_comb[5][3];
    p3_col_transformed[5][4] <= p3_col_transformed_comb[5][4];
    p3_col_transformed[5][5] <= p3_col_transformed_comb[5][5];
    p3_col_transformed[5][6] <= p3_col_transformed_comb[5][6];
    p3_col_transformed[5][7] <= p3_col_transformed_comb[5][7];
    p3_col_transformed[6][0] <= p3_col_transformed_comb[6][0];
    p3_col_transformed[6][1] <= p3_col_transformed_comb[6][1];
    p3_col_transformed[6][2] <= p3_col_transformed_comb[6][2];
    p3_col_transformed[6][3] <= p3_col_transformed_comb[6][3];
    p3_col_transformed[6][4] <= p3_col_transformed_comb[6][4];
    p3_col_transformed[6][5] <= p3_col_transformed_comb[6][5];
    p3_col_transformed[6][6] <= p3_col_transformed_comb[6][6];
    p3_col_transformed[6][7] <= p3_col_transformed_comb[6][7];
    p3_col_transformed[7][0] <= p3_col_transformed_comb[7][0];
    p3_col_transformed[7][1] <= p3_col_transformed_comb[7][1];
    p3_col_transformed[7][2] <= p3_col_transformed_comb[7][2];
    p3_col_transformed[7][3] <= p3_col_transformed_comb[7][3];
    p3_col_transformed[7][4] <= p3_col_transformed_comb[7][4];
    p3_col_transformed[7][5] <= p3_col_transformed_comb[7][5];
    p3_col_transformed[7][6] <= p3_col_transformed_comb[7][6];
    p3_col_transformed[7][7] <= p3_col_transformed_comb[7][7];
  end
  assign out = {{p3_col_transformed[7][7], p3_col_transformed[7][6], p3_col_transformed[7][5], p3_col_transformed[7][4], p3_col_transformed[7][3], p3_col_transformed[7][2], p3_col_transformed[7][1], p3_col_transformed[7][0]}, {p3_col_transformed[6][7], p3_col_transformed[6][6], p3_col_transformed[6][5], p3_col_transformed[6][4], p3_col_transformed[6][3], p3_col_transformed[6][2], p3_col_transformed[6][1], p3_col_transformed[6][0]}, {p3_col_transformed[5][7], p3_col_transformed[5][6], p3_col_transformed[5][5], p3_col_transformed[5][4], p3_col_transformed[5][3], p3_col_transformed[5][2], p3_col_transformed[5][1], p3_col_transformed[5][0]}, {p3_col_transformed[4][7], p3_col_transformed[4][6], p3_col_transformed[4][5], p3_col_transformed[4][4], p3_col_transformed[4][3], p3_col_transformed[4][2], p3_col_transformed[4][1], p3_col_transformed[4][0]}, {p3_col_transformed[3][7], p3_col_transformed[3][6], p3_col_transformed[3][5], p3_col_transformed[3][4], p3_col_transformed[3][3], p3_col_transformed[3][2], p3_col_transformed[3][1], p3_col_transformed[3][0]}, {p3_col_transformed[2][7], p3_col_transformed[2][6], p3_col_transformed[2][5], p3_col_transformed[2][4], p3_col_transformed[2][3], p3_col_transformed[2][2], p3_col_transformed[2][1], p3_col_transformed[2][0]}, {p3_col_transformed[1][7], p3_col_transformed[1][6], p3_col_transformed[1][5], p3_col_transformed[1][4], p3_col_transformed[1][3], p3_col_transformed[1][2], p3_col_transformed[1][1], p3_col_transformed[1][0]}, {p3_col_transformed[0][7], p3_col_transformed[0][6], p3_col_transformed[0][5], p3_col_transformed[0][4], p3_col_transformed[0][3], p3_col_transformed[0][2], p3_col_transformed[0][1], p3_col_transformed[0][0]}};
endmodule
