module dct_2d_s10(
  input wire clk,
  input wire [639:0] x,
  output wire [639:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [18:0] smul19b_11b_x_9b (input reg [10:0] lhs, input reg [8:0] rhs);
    reg signed [10:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [18:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul19b_11b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [19:0] smul20b_11b_x_9b (input reg [10:0] lhs, input reg [8:0] rhs);
    reg signed [10:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [19:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul20b_11b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [17:0] smul18b_18b_x_8b (input reg [17:0] lhs, input reg [7:0] rhs);
    reg signed [17:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [17:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul18b_18b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [17:0] smul18b_18b_x_6b (input reg [17:0] lhs, input reg [5:0] rhs);
    reg signed [17:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [17:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul18b_18b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [18:0] smul19b_19b_x_7b (input reg [18:0] lhs, input reg [6:0] rhs);
    reg signed [18:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [18:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul19b_19b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [18:0] smul19b_19b_x_6b (input reg [18:0] lhs, input reg [5:0] rhs);
    reg signed [18:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [18:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul19b_19b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [18:0] smul19b_19b_x_8b (input reg [18:0] lhs, input reg [7:0] rhs);
    reg signed [18:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [18:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul19b_19b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [17:0] smul18b_18b_x_7b (input reg [17:0] lhs, input reg [6:0] rhs);
    reg signed [17:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [17:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul18b_18b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [23:0] umul24b_24b_x_7b (input reg [23:0] lhs, input reg [6:0] rhs);
    begin
      umul24b_24b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [9:0] x_unflattened[0:7][0:7];
  assign x_unflattened[0][0] = x[9:0];
  assign x_unflattened[0][1] = x[19:10];
  assign x_unflattened[0][2] = x[29:20];
  assign x_unflattened[0][3] = x[39:30];
  assign x_unflattened[0][4] = x[49:40];
  assign x_unflattened[0][5] = x[59:50];
  assign x_unflattened[0][6] = x[69:60];
  assign x_unflattened[0][7] = x[79:70];
  assign x_unflattened[1][0] = x[89:80];
  assign x_unflattened[1][1] = x[99:90];
  assign x_unflattened[1][2] = x[109:100];
  assign x_unflattened[1][3] = x[119:110];
  assign x_unflattened[1][4] = x[129:120];
  assign x_unflattened[1][5] = x[139:130];
  assign x_unflattened[1][6] = x[149:140];
  assign x_unflattened[1][7] = x[159:150];
  assign x_unflattened[2][0] = x[169:160];
  assign x_unflattened[2][1] = x[179:170];
  assign x_unflattened[2][2] = x[189:180];
  assign x_unflattened[2][3] = x[199:190];
  assign x_unflattened[2][4] = x[209:200];
  assign x_unflattened[2][5] = x[219:210];
  assign x_unflattened[2][6] = x[229:220];
  assign x_unflattened[2][7] = x[239:230];
  assign x_unflattened[3][0] = x[249:240];
  assign x_unflattened[3][1] = x[259:250];
  assign x_unflattened[3][2] = x[269:260];
  assign x_unflattened[3][3] = x[279:270];
  assign x_unflattened[3][4] = x[289:280];
  assign x_unflattened[3][5] = x[299:290];
  assign x_unflattened[3][6] = x[309:300];
  assign x_unflattened[3][7] = x[319:310];
  assign x_unflattened[4][0] = x[329:320];
  assign x_unflattened[4][1] = x[339:330];
  assign x_unflattened[4][2] = x[349:340];
  assign x_unflattened[4][3] = x[359:350];
  assign x_unflattened[4][4] = x[369:360];
  assign x_unflattened[4][5] = x[379:370];
  assign x_unflattened[4][6] = x[389:380];
  assign x_unflattened[4][7] = x[399:390];
  assign x_unflattened[5][0] = x[409:400];
  assign x_unflattened[5][1] = x[419:410];
  assign x_unflattened[5][2] = x[429:420];
  assign x_unflattened[5][3] = x[439:430];
  assign x_unflattened[5][4] = x[449:440];
  assign x_unflattened[5][5] = x[459:450];
  assign x_unflattened[5][6] = x[469:460];
  assign x_unflattened[5][7] = x[479:470];
  assign x_unflattened[6][0] = x[489:480];
  assign x_unflattened[6][1] = x[499:490];
  assign x_unflattened[6][2] = x[509:500];
  assign x_unflattened[6][3] = x[519:510];
  assign x_unflattened[6][4] = x[529:520];
  assign x_unflattened[6][5] = x[539:530];
  assign x_unflattened[6][6] = x[549:540];
  assign x_unflattened[6][7] = x[559:550];
  assign x_unflattened[7][0] = x[569:560];
  assign x_unflattened[7][1] = x[579:570];
  assign x_unflattened[7][2] = x[589:580];
  assign x_unflattened[7][3] = x[599:590];
  assign x_unflattened[7][4] = x[609:600];
  assign x_unflattened[7][5] = x[619:610];
  assign x_unflattened[7][6] = x[629:620];
  assign x_unflattened[7][7] = x[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_x[0:7][0:7];
  always @ (posedge clk) begin
    p0_x[0][0] <= x_unflattened[0][0];
    p0_x[0][1] <= x_unflattened[0][1];
    p0_x[0][2] <= x_unflattened[0][2];
    p0_x[0][3] <= x_unflattened[0][3];
    p0_x[0][4] <= x_unflattened[0][4];
    p0_x[0][5] <= x_unflattened[0][5];
    p0_x[0][6] <= x_unflattened[0][6];
    p0_x[0][7] <= x_unflattened[0][7];
    p0_x[1][0] <= x_unflattened[1][0];
    p0_x[1][1] <= x_unflattened[1][1];
    p0_x[1][2] <= x_unflattened[1][2];
    p0_x[1][3] <= x_unflattened[1][3];
    p0_x[1][4] <= x_unflattened[1][4];
    p0_x[1][5] <= x_unflattened[1][5];
    p0_x[1][6] <= x_unflattened[1][6];
    p0_x[1][7] <= x_unflattened[1][7];
    p0_x[2][0] <= x_unflattened[2][0];
    p0_x[2][1] <= x_unflattened[2][1];
    p0_x[2][2] <= x_unflattened[2][2];
    p0_x[2][3] <= x_unflattened[2][3];
    p0_x[2][4] <= x_unflattened[2][4];
    p0_x[2][5] <= x_unflattened[2][5];
    p0_x[2][6] <= x_unflattened[2][6];
    p0_x[2][7] <= x_unflattened[2][7];
    p0_x[3][0] <= x_unflattened[3][0];
    p0_x[3][1] <= x_unflattened[3][1];
    p0_x[3][2] <= x_unflattened[3][2];
    p0_x[3][3] <= x_unflattened[3][3];
    p0_x[3][4] <= x_unflattened[3][4];
    p0_x[3][5] <= x_unflattened[3][5];
    p0_x[3][6] <= x_unflattened[3][6];
    p0_x[3][7] <= x_unflattened[3][7];
    p0_x[4][0] <= x_unflattened[4][0];
    p0_x[4][1] <= x_unflattened[4][1];
    p0_x[4][2] <= x_unflattened[4][2];
    p0_x[4][3] <= x_unflattened[4][3];
    p0_x[4][4] <= x_unflattened[4][4];
    p0_x[4][5] <= x_unflattened[4][5];
    p0_x[4][6] <= x_unflattened[4][6];
    p0_x[4][7] <= x_unflattened[4][7];
    p0_x[5][0] <= x_unflattened[5][0];
    p0_x[5][1] <= x_unflattened[5][1];
    p0_x[5][2] <= x_unflattened[5][2];
    p0_x[5][3] <= x_unflattened[5][3];
    p0_x[5][4] <= x_unflattened[5][4];
    p0_x[5][5] <= x_unflattened[5][5];
    p0_x[5][6] <= x_unflattened[5][6];
    p0_x[5][7] <= x_unflattened[5][7];
    p0_x[6][0] <= x_unflattened[6][0];
    p0_x[6][1] <= x_unflattened[6][1];
    p0_x[6][2] <= x_unflattened[6][2];
    p0_x[6][3] <= x_unflattened[6][3];
    p0_x[6][4] <= x_unflattened[6][4];
    p0_x[6][5] <= x_unflattened[6][5];
    p0_x[6][6] <= x_unflattened[6][6];
    p0_x[6][7] <= x_unflattened[6][7];
    p0_x[7][0] <= x_unflattened[7][0];
    p0_x[7][1] <= x_unflattened[7][1];
    p0_x[7][2] <= x_unflattened[7][2];
    p0_x[7][3] <= x_unflattened[7][3];
    p0_x[7][4] <= x_unflattened[7][4];
    p0_x[7][5] <= x_unflattened[7][5];
    p0_x[7][6] <= x_unflattened[7][6];
    p0_x[7][7] <= x_unflattened[7][7];
  end

  // ===== Pipe stage 1:
  wire [9:0] p1_array_index_79763_comb;
  wire [9:0] p1_array_index_79764_comb;
  wire [9:0] p1_array_index_79765_comb;
  wire [9:0] p1_array_index_79766_comb;
  wire [9:0] p1_array_index_79767_comb;
  wire [9:0] p1_array_index_79768_comb;
  wire [9:0] p1_array_index_79769_comb;
  wire [9:0] p1_array_index_79770_comb;
  wire [9:0] p1_array_index_79771_comb;
  wire [9:0] p1_array_index_79772_comb;
  wire [9:0] p1_array_index_79773_comb;
  wire [9:0] p1_array_index_79774_comb;
  wire [9:0] p1_array_index_79775_comb;
  wire [9:0] p1_array_index_79776_comb;
  wire [9:0] p1_array_index_79777_comb;
  wire [9:0] p1_array_index_79778_comb;
  wire [9:0] p1_array_index_79779_comb;
  wire [9:0] p1_array_index_79780_comb;
  wire [9:0] p1_array_index_79781_comb;
  wire [9:0] p1_array_index_79782_comb;
  wire [9:0] p1_array_index_79783_comb;
  wire [9:0] p1_array_index_79784_comb;
  wire [9:0] p1_array_index_79785_comb;
  wire [9:0] p1_array_index_79786_comb;
  wire [9:0] p1_array_index_79787_comb;
  wire [9:0] p1_array_index_79788_comb;
  wire [9:0] p1_array_index_79789_comb;
  wire [9:0] p1_array_index_79790_comb;
  wire [9:0] p1_array_index_79791_comb;
  wire [9:0] p1_array_index_79792_comb;
  wire [9:0] p1_array_index_79793_comb;
  wire [9:0] p1_array_index_79794_comb;
  wire [9:0] p1_array_index_79795_comb;
  wire [9:0] p1_array_index_79796_comb;
  wire [9:0] p1_array_index_79797_comb;
  wire [9:0] p1_array_index_79798_comb;
  wire [9:0] p1_array_index_79799_comb;
  wire [9:0] p1_array_index_79800_comb;
  wire [9:0] p1_array_index_79801_comb;
  wire [9:0] p1_array_index_79802_comb;
  wire [9:0] p1_array_index_79803_comb;
  wire [9:0] p1_array_index_79804_comb;
  wire [9:0] p1_array_index_79805_comb;
  wire [9:0] p1_array_index_79806_comb;
  wire [9:0] p1_array_index_79807_comb;
  wire [9:0] p1_array_index_79808_comb;
  wire [9:0] p1_array_index_79809_comb;
  wire [9:0] p1_array_index_79810_comb;
  wire [9:0] p1_array_index_79811_comb;
  wire [9:0] p1_array_index_79812_comb;
  wire [9:0] p1_array_index_79813_comb;
  wire [9:0] p1_array_index_79814_comb;
  wire [9:0] p1_array_index_79815_comb;
  wire [9:0] p1_array_index_79816_comb;
  wire [9:0] p1_array_index_79817_comb;
  wire [9:0] p1_array_index_79818_comb;
  wire [9:0] p1_array_index_79819_comb;
  wire [9:0] p1_array_index_79820_comb;
  wire [9:0] p1_array_index_79821_comb;
  wire [9:0] p1_array_index_79822_comb;
  wire [9:0] p1_array_index_79823_comb;
  wire [9:0] p1_array_index_79824_comb;
  wire [9:0] p1_array_index_79825_comb;
  wire [9:0] p1_array_index_79826_comb;
  wire [2:0] p1_bit_slice_79827_comb;
  wire [2:0] p1_bit_slice_79828_comb;
  wire [2:0] p1_bit_slice_79829_comb;
  wire [2:0] p1_bit_slice_79830_comb;
  wire [2:0] p1_bit_slice_79831_comb;
  wire [2:0] p1_bit_slice_79832_comb;
  wire [2:0] p1_bit_slice_79833_comb;
  wire [2:0] p1_bit_slice_79834_comb;
  wire [2:0] p1_bit_slice_79835_comb;
  wire [2:0] p1_bit_slice_79836_comb;
  wire [2:0] p1_bit_slice_79837_comb;
  wire [2:0] p1_bit_slice_79838_comb;
  wire [2:0] p1_bit_slice_79839_comb;
  wire [2:0] p1_bit_slice_79840_comb;
  wire [2:0] p1_bit_slice_79841_comb;
  wire [2:0] p1_bit_slice_79842_comb;
  wire [2:0] p1_bit_slice_79843_comb;
  wire [2:0] p1_bit_slice_79844_comb;
  wire [2:0] p1_bit_slice_79845_comb;
  wire [2:0] p1_bit_slice_79846_comb;
  wire [2:0] p1_bit_slice_79847_comb;
  wire [2:0] p1_bit_slice_79848_comb;
  wire [2:0] p1_bit_slice_79849_comb;
  wire [2:0] p1_bit_slice_79850_comb;
  wire [2:0] p1_bit_slice_79851_comb;
  wire [2:0] p1_bit_slice_79852_comb;
  wire [2:0] p1_bit_slice_79853_comb;
  wire [2:0] p1_bit_slice_79854_comb;
  wire [2:0] p1_bit_slice_79855_comb;
  wire [2:0] p1_bit_slice_79856_comb;
  wire [2:0] p1_bit_slice_79857_comb;
  wire [2:0] p1_bit_slice_79858_comb;
  wire [2:0] p1_bit_slice_79859_comb;
  wire [2:0] p1_bit_slice_79860_comb;
  wire [2:0] p1_bit_slice_79861_comb;
  wire [2:0] p1_bit_slice_79862_comb;
  wire [2:0] p1_bit_slice_79863_comb;
  wire [2:0] p1_bit_slice_79864_comb;
  wire [2:0] p1_bit_slice_79865_comb;
  wire [2:0] p1_bit_slice_79866_comb;
  wire [2:0] p1_bit_slice_79867_comb;
  wire [2:0] p1_bit_slice_79868_comb;
  wire [2:0] p1_bit_slice_79869_comb;
  wire [2:0] p1_bit_slice_79870_comb;
  wire [2:0] p1_bit_slice_79871_comb;
  wire [2:0] p1_bit_slice_79872_comb;
  wire [2:0] p1_bit_slice_79873_comb;
  wire [2:0] p1_bit_slice_79874_comb;
  wire [2:0] p1_bit_slice_79875_comb;
  wire [2:0] p1_bit_slice_79876_comb;
  wire [2:0] p1_bit_slice_79877_comb;
  wire [2:0] p1_bit_slice_79878_comb;
  wire [2:0] p1_bit_slice_79879_comb;
  wire [2:0] p1_bit_slice_79880_comb;
  wire [2:0] p1_bit_slice_79881_comb;
  wire [2:0] p1_bit_slice_79882_comb;
  wire [2:0] p1_bit_slice_79883_comb;
  wire [2:0] p1_bit_slice_79884_comb;
  wire [2:0] p1_bit_slice_79885_comb;
  wire [2:0] p1_bit_slice_79886_comb;
  wire [2:0] p1_bit_slice_79887_comb;
  wire [2:0] p1_bit_slice_79888_comb;
  wire [2:0] p1_bit_slice_79889_comb;
  wire [2:0] p1_bit_slice_79890_comb;
  wire [3:0] p1_add_80019_comb;
  wire [3:0] p1_add_80021_comb;
  wire [3:0] p1_add_80023_comb;
  wire [3:0] p1_add_80025_comb;
  wire [3:0] p1_add_80027_comb;
  wire [3:0] p1_add_80029_comb;
  wire [3:0] p1_add_80031_comb;
  wire [3:0] p1_add_80033_comb;
  wire [3:0] p1_add_80035_comb;
  wire [3:0] p1_add_80037_comb;
  wire [3:0] p1_add_80039_comb;
  wire [3:0] p1_add_80041_comb;
  wire [3:0] p1_add_80043_comb;
  wire [3:0] p1_add_80045_comb;
  wire [3:0] p1_add_80047_comb;
  wire [3:0] p1_add_80049_comb;
  wire [3:0] p1_add_80051_comb;
  wire [3:0] p1_add_80053_comb;
  wire [3:0] p1_add_80055_comb;
  wire [3:0] p1_add_80057_comb;
  wire [3:0] p1_add_80059_comb;
  wire [3:0] p1_add_80061_comb;
  wire [3:0] p1_add_80063_comb;
  wire [3:0] p1_add_80065_comb;
  wire [3:0] p1_add_80067_comb;
  wire [3:0] p1_add_80069_comb;
  wire [3:0] p1_add_80071_comb;
  wire [3:0] p1_add_80073_comb;
  wire [3:0] p1_add_80075_comb;
  wire [3:0] p1_add_80077_comb;
  wire [3:0] p1_add_80079_comb;
  wire [3:0] p1_add_80081_comb;
  wire [3:0] p1_add_80083_comb;
  wire [3:0] p1_add_80085_comb;
  wire [3:0] p1_add_80087_comb;
  wire [3:0] p1_add_80089_comb;
  wire [3:0] p1_add_80091_comb;
  wire [3:0] p1_add_80093_comb;
  wire [3:0] p1_add_80095_comb;
  wire [3:0] p1_add_80097_comb;
  wire [3:0] p1_add_80099_comb;
  wire [3:0] p1_add_80101_comb;
  wire [3:0] p1_add_80103_comb;
  wire [3:0] p1_add_80105_comb;
  wire [3:0] p1_add_80107_comb;
  wire [3:0] p1_add_80109_comb;
  wire [3:0] p1_add_80111_comb;
  wire [3:0] p1_add_80113_comb;
  wire [3:0] p1_add_80115_comb;
  wire [3:0] p1_add_80117_comb;
  wire [3:0] p1_add_80119_comb;
  wire [3:0] p1_add_80121_comb;
  wire [3:0] p1_add_80123_comb;
  wire [3:0] p1_add_80125_comb;
  wire [3:0] p1_add_80127_comb;
  wire [3:0] p1_add_80129_comb;
  wire [3:0] p1_add_80131_comb;
  wire [3:0] p1_add_80133_comb;
  wire [3:0] p1_add_80135_comb;
  wire [3:0] p1_add_80137_comb;
  wire [3:0] p1_add_80139_comb;
  wire [3:0] p1_add_80141_comb;
  wire [3:0] p1_add_80143_comb;
  wire [3:0] p1_add_80145_comb;
  wire [10:0] p1_concat_80147_comb;
  wire [10:0] p1_concat_80148_comb;
  wire [10:0] p1_concat_80149_comb;
  wire [10:0] p1_concat_80150_comb;
  wire [10:0] p1_concat_80151_comb;
  wire [10:0] p1_concat_80152_comb;
  wire [10:0] p1_concat_80153_comb;
  wire [10:0] p1_concat_80154_comb;
  wire [10:0] p1_concat_80155_comb;
  wire [10:0] p1_concat_80156_comb;
  wire [10:0] p1_concat_80157_comb;
  wire [10:0] p1_concat_80158_comb;
  wire [10:0] p1_concat_80159_comb;
  wire [10:0] p1_concat_80160_comb;
  wire [10:0] p1_concat_80161_comb;
  wire [10:0] p1_concat_80162_comb;
  wire [10:0] p1_concat_80163_comb;
  wire [10:0] p1_concat_80164_comb;
  wire [10:0] p1_concat_80165_comb;
  wire [10:0] p1_concat_80166_comb;
  wire [10:0] p1_concat_80167_comb;
  wire [10:0] p1_concat_80168_comb;
  wire [10:0] p1_concat_80169_comb;
  wire [10:0] p1_concat_80170_comb;
  wire [10:0] p1_concat_80171_comb;
  wire [10:0] p1_concat_80172_comb;
  wire [10:0] p1_concat_80173_comb;
  wire [10:0] p1_concat_80174_comb;
  wire [10:0] p1_concat_80175_comb;
  wire [10:0] p1_concat_80176_comb;
  wire [10:0] p1_concat_80177_comb;
  wire [10:0] p1_concat_80178_comb;
  wire [10:0] p1_concat_80179_comb;
  wire [10:0] p1_concat_80180_comb;
  wire [10:0] p1_concat_80181_comb;
  wire [10:0] p1_concat_80182_comb;
  wire [10:0] p1_concat_80183_comb;
  wire [10:0] p1_concat_80184_comb;
  wire [10:0] p1_concat_80185_comb;
  wire [10:0] p1_concat_80186_comb;
  wire [10:0] p1_concat_80187_comb;
  wire [10:0] p1_concat_80188_comb;
  wire [10:0] p1_concat_80189_comb;
  wire [10:0] p1_concat_80190_comb;
  wire [10:0] p1_concat_80191_comb;
  wire [10:0] p1_concat_80192_comb;
  wire [10:0] p1_concat_80193_comb;
  wire [10:0] p1_concat_80194_comb;
  wire [10:0] p1_concat_80195_comb;
  wire [10:0] p1_concat_80196_comb;
  wire [10:0] p1_concat_80197_comb;
  wire [10:0] p1_concat_80198_comb;
  wire [10:0] p1_concat_80199_comb;
  wire [10:0] p1_concat_80200_comb;
  wire [10:0] p1_concat_80201_comb;
  wire [10:0] p1_concat_80202_comb;
  wire [10:0] p1_concat_80203_comb;
  wire [10:0] p1_concat_80204_comb;
  wire [10:0] p1_concat_80205_comb;
  wire [10:0] p1_concat_80206_comb;
  wire [10:0] p1_concat_80207_comb;
  wire [10:0] p1_concat_80208_comb;
  wire [10:0] p1_concat_80209_comb;
  wire [10:0] p1_concat_80210_comb;
  wire [23:0] p1_sign_ext_80213_comb;
  wire [23:0] p1_sign_ext_80214_comb;
  wire [23:0] p1_sign_ext_80215_comb;
  wire [23:0] p1_sign_ext_80216_comb;
  wire [23:0] p1_sign_ext_80221_comb;
  wire [23:0] p1_sign_ext_80222_comb;
  wire [23:0] p1_sign_ext_80223_comb;
  wire [23:0] p1_sign_ext_80224_comb;
  wire [23:0] p1_sign_ext_80229_comb;
  wire [23:0] p1_sign_ext_80230_comb;
  wire [23:0] p1_sign_ext_80231_comb;
  wire [23:0] p1_sign_ext_80232_comb;
  wire [23:0] p1_sign_ext_80237_comb;
  wire [23:0] p1_sign_ext_80238_comb;
  wire [23:0] p1_sign_ext_80239_comb;
  wire [23:0] p1_sign_ext_80240_comb;
  wire [23:0] p1_sign_ext_80243_comb;
  wire [23:0] p1_sign_ext_80244_comb;
  wire [23:0] p1_sign_ext_80245_comb;
  wire [23:0] p1_sign_ext_80246_comb;
  wire [23:0] p1_sign_ext_80247_comb;
  wire [23:0] p1_sign_ext_80248_comb;
  wire [23:0] p1_sign_ext_80249_comb;
  wire [23:0] p1_sign_ext_80250_comb;
  wire [23:0] p1_sign_ext_80267_comb;
  wire [23:0] p1_sign_ext_80272_comb;
  wire [23:0] p1_sign_ext_80273_comb;
  wire [23:0] p1_sign_ext_80278_comb;
  wire [23:0] p1_sign_ext_80279_comb;
  wire [23:0] p1_sign_ext_80284_comb;
  wire [23:0] p1_sign_ext_80285_comb;
  wire [23:0] p1_sign_ext_80290_comb;
  wire [23:0] p1_sign_ext_80309_comb;
  wire [23:0] p1_sign_ext_80310_comb;
  wire [23:0] p1_sign_ext_80311_comb;
  wire [23:0] p1_sign_ext_80312_comb;
  wire [23:0] p1_sign_ext_80317_comb;
  wire [23:0] p1_sign_ext_80318_comb;
  wire [23:0] p1_sign_ext_80319_comb;
  wire [23:0] p1_sign_ext_80320_comb;
  wire [23:0] p1_sign_ext_80323_comb;
  wire [23:0] p1_sign_ext_80324_comb;
  wire [23:0] p1_sign_ext_80325_comb;
  wire [23:0] p1_sign_ext_80326_comb;
  wire [23:0] p1_sign_ext_80335_comb;
  wire [23:0] p1_sign_ext_80340_comb;
  wire [23:0] p1_sign_ext_80341_comb;
  wire [23:0] p1_sign_ext_80346_comb;
  wire [23:0] p1_sign_ext_80357_comb;
  wire [23:0] p1_sign_ext_80358_comb;
  wire [23:0] p1_sign_ext_80359_comb;
  wire [23:0] p1_sign_ext_80360_comb;
  wire [23:0] p1_sign_ext_80365_comb;
  wire [23:0] p1_sign_ext_80366_comb;
  wire [23:0] p1_sign_ext_80367_comb;
  wire [23:0] p1_sign_ext_80368_comb;
  wire [23:0] p1_sign_ext_80371_comb;
  wire [23:0] p1_sign_ext_80372_comb;
  wire [23:0] p1_sign_ext_80373_comb;
  wire [23:0] p1_sign_ext_80374_comb;
  wire [23:0] p1_sign_ext_80383_comb;
  wire [23:0] p1_sign_ext_80388_comb;
  wire [23:0] p1_sign_ext_80389_comb;
  wire [23:0] p1_sign_ext_80394_comb;
  wire [18:0] p1_smul_81379_comb;
  wire [18:0] p1_smul_81380_comb;
  wire [18:0] p1_smul_81381_comb;
  wire [18:0] p1_smul_81382_comb;
  wire [18:0] p1_smul_81383_comb;
  wire [18:0] p1_smul_81384_comb;
  wire [18:0] p1_smul_81385_comb;
  wire [18:0] p1_smul_81386_comb;
  wire [18:0] p1_smul_81387_comb;
  wire [18:0] p1_smul_81388_comb;
  wire [18:0] p1_smul_81389_comb;
  wire [18:0] p1_smul_81390_comb;
  wire [18:0] p1_smul_81391_comb;
  wire [18:0] p1_smul_81392_comb;
  wire [18:0] p1_smul_81393_comb;
  wire [18:0] p1_smul_81394_comb;
  wire [18:0] p1_smul_81395_comb;
  wire [18:0] p1_smul_81396_comb;
  wire [18:0] p1_smul_81397_comb;
  wire [18:0] p1_smul_81398_comb;
  wire [18:0] p1_smul_81399_comb;
  wire [18:0] p1_smul_81400_comb;
  wire [18:0] p1_smul_81401_comb;
  wire [18:0] p1_smul_81402_comb;
  wire [18:0] p1_smul_81403_comb;
  wire [18:0] p1_smul_81404_comb;
  wire [18:0] p1_smul_81405_comb;
  wire [18:0] p1_smul_81406_comb;
  wire [18:0] p1_smul_81407_comb;
  wire [18:0] p1_smul_81408_comb;
  wire [18:0] p1_smul_81409_comb;
  wire [18:0] p1_smul_81410_comb;
  wire [18:0] p1_smul_81547_comb;
  wire [18:0] p1_smul_81548_comb;
  wire [18:0] p1_smul_81549_comb;
  wire [18:0] p1_smul_81550_comb;
  wire [18:0] p1_smul_81551_comb;
  wire [18:0] p1_smul_81552_comb;
  wire [18:0] p1_smul_81553_comb;
  wire [18:0] p1_smul_81554_comb;
  wire [18:0] p1_smul_81555_comb;
  wire [18:0] p1_smul_81556_comb;
  wire [18:0] p1_smul_81557_comb;
  wire [18:0] p1_smul_81558_comb;
  wire [18:0] p1_smul_81559_comb;
  wire [18:0] p1_smul_81560_comb;
  wire [18:0] p1_smul_81561_comb;
  wire [18:0] p1_smul_81562_comb;
  wire [18:0] p1_smul_81659_comb;
  wire [18:0] p1_smul_81660_comb;
  wire [18:0] p1_smul_81661_comb;
  wire [18:0] p1_smul_81662_comb;
  wire [18:0] p1_smul_81663_comb;
  wire [18:0] p1_smul_81664_comb;
  wire [18:0] p1_smul_81665_comb;
  wire [18:0] p1_smul_81666_comb;
  wire [18:0] p1_smul_81667_comb;
  wire [18:0] p1_smul_81668_comb;
  wire [18:0] p1_smul_81669_comb;
  wire [18:0] p1_smul_81670_comb;
  wire [18:0] p1_smul_81671_comb;
  wire [18:0] p1_smul_81672_comb;
  wire [18:0] p1_smul_81673_comb;
  wire [18:0] p1_smul_81674_comb;
  wire [19:0] p1_smul_80403_comb;
  wire [19:0] p1_smul_80404_comb;
  wire [19:0] p1_smul_80413_comb;
  wire [19:0] p1_smul_80414_comb;
  wire [19:0] p1_smul_80415_comb;
  wire [19:0] p1_smul_80416_comb;
  wire [19:0] p1_smul_80425_comb;
  wire [19:0] p1_smul_80426_comb;
  wire [19:0] p1_smul_80427_comb;
  wire [19:0] p1_smul_80428_comb;
  wire [19:0] p1_smul_80437_comb;
  wire [19:0] p1_smul_80438_comb;
  wire [19:0] p1_smul_80439_comb;
  wire [19:0] p1_smul_80440_comb;
  wire [19:0] p1_smul_80449_comb;
  wire [19:0] p1_smul_80450_comb;
  wire [19:0] p1_smul_80483_comb;
  wire [19:0] p1_smul_80485_comb;
  wire [19:0] p1_smul_80490_comb;
  wire [19:0] p1_smul_80492_comb;
  wire [19:0] p1_smul_80493_comb;
  wire [19:0] p1_smul_80495_comb;
  wire [19:0] p1_smul_80500_comb;
  wire [19:0] p1_smul_80502_comb;
  wire [19:0] p1_smul_80503_comb;
  wire [19:0] p1_smul_80505_comb;
  wire [19:0] p1_smul_80510_comb;
  wire [19:0] p1_smul_80512_comb;
  wire [19:0] p1_smul_80513_comb;
  wire [19:0] p1_smul_80515_comb;
  wire [19:0] p1_smul_80520_comb;
  wire [19:0] p1_smul_80522_comb;
  wire [19:0] p1_smul_80525_comb;
  wire [19:0] p1_smul_80527_comb;
  wire [19:0] p1_smul_80528_comb;
  wire [19:0] p1_smul_80530_comb;
  wire [19:0] p1_smul_80535_comb;
  wire [19:0] p1_smul_80537_comb;
  wire [19:0] p1_smul_80538_comb;
  wire [19:0] p1_smul_80540_comb;
  wire [19:0] p1_smul_80545_comb;
  wire [19:0] p1_smul_80547_comb;
  wire [19:0] p1_smul_80548_comb;
  wire [19:0] p1_smul_80550_comb;
  wire [19:0] p1_smul_80555_comb;
  wire [19:0] p1_smul_80557_comb;
  wire [19:0] p1_smul_80558_comb;
  wire [19:0] p1_smul_80560_comb;
  wire [19:0] p1_smul_80583_comb;
  wire [19:0] p1_smul_80584_comb;
  wire [19:0] p1_smul_80585_comb;
  wire [19:0] p1_smul_80586_comb;
  wire [19:0] p1_smul_80595_comb;
  wire [19:0] p1_smul_80596_comb;
  wire [19:0] p1_smul_80597_comb;
  wire [19:0] p1_smul_80598_comb;
  wire [19:0] p1_smul_80607_comb;
  wire [19:0] p1_smul_80608_comb;
  wire [19:0] p1_smul_80609_comb;
  wire [19:0] p1_smul_80610_comb;
  wire [19:0] p1_smul_80619_comb;
  wire [19:0] p1_smul_80620_comb;
  wire [19:0] p1_smul_80621_comb;
  wire [19:0] p1_smul_80622_comb;
  wire [19:0] p1_smul_80627_comb;
  wire [19:0] p1_smul_80628_comb;
  wire [19:0] p1_smul_80637_comb;
  wire [19:0] p1_smul_80638_comb;
  wire [19:0] p1_smul_80639_comb;
  wire [19:0] p1_smul_80640_comb;
  wire [19:0] p1_smul_80649_comb;
  wire [19:0] p1_smul_80650_comb;
  wire [19:0] p1_smul_80667_comb;
  wire [19:0] p1_smul_80669_comb;
  wire [19:0] p1_smul_80674_comb;
  wire [19:0] p1_smul_80676_comb;
  wire [19:0] p1_smul_80677_comb;
  wire [19:0] p1_smul_80679_comb;
  wire [19:0] p1_smul_80684_comb;
  wire [19:0] p1_smul_80686_comb;
  wire [19:0] p1_smul_80689_comb;
  wire [19:0] p1_smul_80691_comb;
  wire [19:0] p1_smul_80692_comb;
  wire [19:0] p1_smul_80694_comb;
  wire [19:0] p1_smul_80699_comb;
  wire [19:0] p1_smul_80701_comb;
  wire [19:0] p1_smul_80702_comb;
  wire [19:0] p1_smul_80704_comb;
  wire [19:0] p1_smul_80719_comb;
  wire [19:0] p1_smul_80720_comb;
  wire [19:0] p1_smul_80721_comb;
  wire [19:0] p1_smul_80722_comb;
  wire [19:0] p1_smul_80731_comb;
  wire [19:0] p1_smul_80732_comb;
  wire [19:0] p1_smul_80733_comb;
  wire [19:0] p1_smul_80734_comb;
  wire [19:0] p1_smul_80739_comb;
  wire [19:0] p1_smul_80740_comb;
  wire [19:0] p1_smul_80749_comb;
  wire [19:0] p1_smul_80750_comb;
  wire [19:0] p1_smul_80751_comb;
  wire [19:0] p1_smul_80752_comb;
  wire [19:0] p1_smul_80761_comb;
  wire [19:0] p1_smul_80762_comb;
  wire [19:0] p1_smul_80779_comb;
  wire [19:0] p1_smul_80781_comb;
  wire [19:0] p1_smul_80786_comb;
  wire [19:0] p1_smul_80788_comb;
  wire [19:0] p1_smul_80789_comb;
  wire [19:0] p1_smul_80791_comb;
  wire [19:0] p1_smul_80796_comb;
  wire [19:0] p1_smul_80798_comb;
  wire [19:0] p1_smul_80801_comb;
  wire [19:0] p1_smul_80803_comb;
  wire [19:0] p1_smul_80804_comb;
  wire [19:0] p1_smul_80806_comb;
  wire [19:0] p1_smul_80811_comb;
  wire [19:0] p1_smul_80813_comb;
  wire [19:0] p1_smul_80814_comb;
  wire [19:0] p1_smul_80816_comb;
  wire [19:0] p1_smul_80831_comb;
  wire [19:0] p1_smul_80832_comb;
  wire [19:0] p1_smul_80833_comb;
  wire [19:0] p1_smul_80834_comb;
  wire [19:0] p1_smul_80843_comb;
  wire [19:0] p1_smul_80844_comb;
  wire [19:0] p1_smul_80845_comb;
  wire [19:0] p1_smul_80846_comb;
  wire [18:0] p1_add_81795_comb;
  wire [18:0] p1_add_81796_comb;
  wire [18:0] p1_add_81797_comb;
  wire [18:0] p1_add_81798_comb;
  wire [18:0] p1_add_81799_comb;
  wire [18:0] p1_add_81800_comb;
  wire [18:0] p1_add_81801_comb;
  wire [18:0] p1_add_81802_comb;
  wire [18:0] p1_add_81803_comb;
  wire [18:0] p1_add_81804_comb;
  wire [18:0] p1_add_81805_comb;
  wire [18:0] p1_add_81806_comb;
  wire [18:0] p1_add_81807_comb;
  wire [18:0] p1_add_81808_comb;
  wire [18:0] p1_add_81809_comb;
  wire [18:0] p1_add_81810_comb;
  wire [18:0] p1_add_81915_comb;
  wire [18:0] p1_add_81916_comb;
  wire [18:0] p1_add_81917_comb;
  wire [18:0] p1_add_81918_comb;
  wire [18:0] p1_add_81919_comb;
  wire [18:0] p1_add_81920_comb;
  wire [18:0] p1_add_81921_comb;
  wire [18:0] p1_add_81922_comb;
  wire [18:0] p1_add_81995_comb;
  wire [18:0] p1_add_81996_comb;
  wire [18:0] p1_add_81997_comb;
  wire [18:0] p1_add_81998_comb;
  wire [18:0] p1_add_81999_comb;
  wire [18:0] p1_add_82000_comb;
  wire [18:0] p1_add_82001_comb;
  wire [18:0] p1_add_82002_comb;
  wire [19:0] p1_add_80851_comb;
  wire [17:0] p1_smul_80852_comb;
  wire [17:0] p1_smul_80853_comb;
  wire [17:0] p1_smul_80854_comb;
  wire [17:0] p1_smul_80855_comb;
  wire [19:0] p1_add_80856_comb;
  wire [19:0] p1_add_80857_comb;
  wire [17:0] p1_smul_80858_comb;
  wire [17:0] p1_smul_80859_comb;
  wire [17:0] p1_smul_80860_comb;
  wire [17:0] p1_smul_80861_comb;
  wire [19:0] p1_add_80862_comb;
  wire [19:0] p1_add_80863_comb;
  wire [17:0] p1_smul_80864_comb;
  wire [17:0] p1_smul_80865_comb;
  wire [17:0] p1_smul_80866_comb;
  wire [17:0] p1_smul_80867_comb;
  wire [19:0] p1_add_80868_comb;
  wire [19:0] p1_add_80869_comb;
  wire [17:0] p1_smul_80870_comb;
  wire [17:0] p1_smul_80871_comb;
  wire [17:0] p1_smul_80872_comb;
  wire [17:0] p1_smul_80873_comb;
  wire [19:0] p1_add_80874_comb;
  wire [18:0] p1_smul_80876_comb;
  wire [18:0] p1_smul_80877_comb;
  wire [18:0] p1_smul_80880_comb;
  wire [18:0] p1_smul_80881_comb;
  wire [18:0] p1_smul_80884_comb;
  wire [18:0] p1_smul_80885_comb;
  wire [18:0] p1_smul_80888_comb;
  wire [18:0] p1_smul_80889_comb;
  wire [18:0] p1_smul_80892_comb;
  wire [18:0] p1_smul_80893_comb;
  wire [18:0] p1_smul_80896_comb;
  wire [18:0] p1_smul_80897_comb;
  wire [18:0] p1_smul_80900_comb;
  wire [18:0] p1_smul_80901_comb;
  wire [18:0] p1_smul_80904_comb;
  wire [18:0] p1_smul_80905_comb;
  wire [18:0] p1_smul_80908_comb;
  wire [18:0] p1_smul_80910_comb;
  wire [18:0] p1_smul_80911_comb;
  wire [18:0] p1_smul_80913_comb;
  wire [18:0] p1_smul_80916_comb;
  wire [18:0] p1_smul_80918_comb;
  wire [18:0] p1_smul_80919_comb;
  wire [18:0] p1_smul_80921_comb;
  wire [18:0] p1_smul_80924_comb;
  wire [18:0] p1_smul_80926_comb;
  wire [18:0] p1_smul_80927_comb;
  wire [18:0] p1_smul_80929_comb;
  wire [18:0] p1_smul_80932_comb;
  wire [18:0] p1_smul_80934_comb;
  wire [18:0] p1_smul_80935_comb;
  wire [18:0] p1_smul_80937_comb;
  wire [18:0] p1_smul_80971_comb;
  wire [18:0] p1_smul_80973_comb;
  wire [18:0] p1_smul_80976_comb;
  wire [18:0] p1_smul_80978_comb;
  wire [18:0] p1_smul_80979_comb;
  wire [18:0] p1_smul_80981_comb;
  wire [18:0] p1_smul_80984_comb;
  wire [18:0] p1_smul_80986_comb;
  wire [18:0] p1_smul_80987_comb;
  wire [18:0] p1_smul_80989_comb;
  wire [18:0] p1_smul_80992_comb;
  wire [18:0] p1_smul_80994_comb;
  wire [18:0] p1_smul_80995_comb;
  wire [18:0] p1_smul_80997_comb;
  wire [18:0] p1_smul_81000_comb;
  wire [18:0] p1_smul_81002_comb;
  wire [18:0] p1_smul_81003_comb;
  wire [18:0] p1_smul_81005_comb;
  wire [18:0] p1_smul_81008_comb;
  wire [18:0] p1_smul_81010_comb;
  wire [18:0] p1_smul_81011_comb;
  wire [18:0] p1_smul_81013_comb;
  wire [18:0] p1_smul_81016_comb;
  wire [18:0] p1_smul_81018_comb;
  wire [18:0] p1_smul_81019_comb;
  wire [18:0] p1_smul_81021_comb;
  wire [18:0] p1_smul_81024_comb;
  wire [18:0] p1_smul_81026_comb;
  wire [18:0] p1_smul_81027_comb;
  wire [18:0] p1_smul_81029_comb;
  wire [18:0] p1_smul_81032_comb;
  wire [18:0] p1_smul_81034_comb;
  wire [17:0] p1_smul_81035_comb;
  wire [17:0] p1_smul_81036_comb;
  wire [19:0] p1_add_81037_comb;
  wire [19:0] p1_add_81038_comb;
  wire [17:0] p1_smul_81039_comb;
  wire [17:0] p1_smul_81040_comb;
  wire [17:0] p1_smul_81041_comb;
  wire [17:0] p1_smul_81042_comb;
  wire [19:0] p1_add_81043_comb;
  wire [19:0] p1_add_81044_comb;
  wire [17:0] p1_smul_81045_comb;
  wire [17:0] p1_smul_81046_comb;
  wire [17:0] p1_smul_81047_comb;
  wire [17:0] p1_smul_81048_comb;
  wire [19:0] p1_add_81049_comb;
  wire [19:0] p1_add_81050_comb;
  wire [17:0] p1_smul_81051_comb;
  wire [17:0] p1_smul_81052_comb;
  wire [17:0] p1_smul_81053_comb;
  wire [17:0] p1_smul_81054_comb;
  wire [19:0] p1_add_81055_comb;
  wire [19:0] p1_add_81056_comb;
  wire [17:0] p1_smul_81057_comb;
  wire [17:0] p1_smul_81058_comb;
  wire [19:0] p1_add_81059_comb;
  wire [17:0] p1_smul_81060_comb;
  wire [17:0] p1_smul_81061_comb;
  wire [17:0] p1_smul_81062_comb;
  wire [17:0] p1_smul_81063_comb;
  wire [19:0] p1_add_81064_comb;
  wire [19:0] p1_add_81065_comb;
  wire [17:0] p1_smul_81066_comb;
  wire [17:0] p1_smul_81067_comb;
  wire [17:0] p1_smul_81068_comb;
  wire [17:0] p1_smul_81069_comb;
  wire [19:0] p1_add_81070_comb;
  wire [18:0] p1_smul_81072_comb;
  wire [18:0] p1_smul_81073_comb;
  wire [18:0] p1_smul_81076_comb;
  wire [18:0] p1_smul_81077_comb;
  wire [18:0] p1_smul_81080_comb;
  wire [18:0] p1_smul_81081_comb;
  wire [18:0] p1_smul_81084_comb;
  wire [18:0] p1_smul_81085_comb;
  wire [18:0] p1_smul_81088_comb;
  wire [18:0] p1_smul_81090_comb;
  wire [18:0] p1_smul_81091_comb;
  wire [18:0] p1_smul_81093_comb;
  wire [18:0] p1_smul_81096_comb;
  wire [18:0] p1_smul_81098_comb;
  wire [18:0] p1_smul_81099_comb;
  wire [18:0] p1_smul_81101_comb;
  wire [18:0] p1_smul_81119_comb;
  wire [18:0] p1_smul_81121_comb;
  wire [18:0] p1_smul_81124_comb;
  wire [18:0] p1_smul_81126_comb;
  wire [18:0] p1_smul_81127_comb;
  wire [18:0] p1_smul_81129_comb;
  wire [18:0] p1_smul_81132_comb;
  wire [18:0] p1_smul_81134_comb;
  wire [18:0] p1_smul_81135_comb;
  wire [18:0] p1_smul_81137_comb;
  wire [18:0] p1_smul_81140_comb;
  wire [18:0] p1_smul_81142_comb;
  wire [18:0] p1_smul_81143_comb;
  wire [18:0] p1_smul_81145_comb;
  wire [18:0] p1_smul_81148_comb;
  wire [18:0] p1_smul_81150_comb;
  wire [17:0] p1_smul_81151_comb;
  wire [17:0] p1_smul_81152_comb;
  wire [19:0] p1_add_81153_comb;
  wire [19:0] p1_add_81154_comb;
  wire [17:0] p1_smul_81155_comb;
  wire [17:0] p1_smul_81156_comb;
  wire [17:0] p1_smul_81157_comb;
  wire [17:0] p1_smul_81158_comb;
  wire [19:0] p1_add_81159_comb;
  wire [19:0] p1_add_81160_comb;
  wire [17:0] p1_smul_81161_comb;
  wire [17:0] p1_smul_81162_comb;
  wire [19:0] p1_add_81163_comb;
  wire [17:0] p1_smul_81164_comb;
  wire [17:0] p1_smul_81165_comb;
  wire [17:0] p1_smul_81166_comb;
  wire [17:0] p1_smul_81167_comb;
  wire [19:0] p1_add_81168_comb;
  wire [19:0] p1_add_81169_comb;
  wire [17:0] p1_smul_81170_comb;
  wire [17:0] p1_smul_81171_comb;
  wire [17:0] p1_smul_81172_comb;
  wire [17:0] p1_smul_81173_comb;
  wire [19:0] p1_add_81174_comb;
  wire [18:0] p1_smul_81176_comb;
  wire [18:0] p1_smul_81177_comb;
  wire [18:0] p1_smul_81180_comb;
  wire [18:0] p1_smul_81181_comb;
  wire [18:0] p1_smul_81184_comb;
  wire [18:0] p1_smul_81185_comb;
  wire [18:0] p1_smul_81188_comb;
  wire [18:0] p1_smul_81189_comb;
  wire [18:0] p1_smul_81192_comb;
  wire [18:0] p1_smul_81194_comb;
  wire [18:0] p1_smul_81195_comb;
  wire [18:0] p1_smul_81197_comb;
  wire [18:0] p1_smul_81200_comb;
  wire [18:0] p1_smul_81202_comb;
  wire [18:0] p1_smul_81203_comb;
  wire [18:0] p1_smul_81205_comb;
  wire [18:0] p1_smul_81223_comb;
  wire [18:0] p1_smul_81225_comb;
  wire [18:0] p1_smul_81228_comb;
  wire [18:0] p1_smul_81230_comb;
  wire [18:0] p1_smul_81231_comb;
  wire [18:0] p1_smul_81233_comb;
  wire [18:0] p1_smul_81236_comb;
  wire [18:0] p1_smul_81238_comb;
  wire [18:0] p1_smul_81239_comb;
  wire [18:0] p1_smul_81241_comb;
  wire [18:0] p1_smul_81244_comb;
  wire [18:0] p1_smul_81246_comb;
  wire [18:0] p1_smul_81247_comb;
  wire [18:0] p1_smul_81249_comb;
  wire [18:0] p1_smul_81252_comb;
  wire [18:0] p1_smul_81254_comb;
  wire [17:0] p1_smul_81255_comb;
  wire [17:0] p1_smul_81256_comb;
  wire [19:0] p1_add_81257_comb;
  wire [19:0] p1_add_81258_comb;
  wire [17:0] p1_smul_81259_comb;
  wire [17:0] p1_smul_81260_comb;
  wire [17:0] p1_smul_81261_comb;
  wire [17:0] p1_smul_81262_comb;
  wire [19:0] p1_add_81263_comb;
  wire [19:0] p1_add_81264_comb;
  wire [17:0] p1_smul_81265_comb;
  wire [17:0] p1_smul_81266_comb;
  wire [11:0] p1_add_81715_comb;
  wire [11:0] p1_add_81716_comb;
  wire [11:0] p1_add_81717_comb;
  wire [11:0] p1_add_81718_comb;
  wire [11:0] p1_add_81719_comb;
  wire [11:0] p1_add_81720_comb;
  wire [11:0] p1_add_81721_comb;
  wire [11:0] p1_add_81722_comb;
  wire [11:0] p1_add_81723_comb;
  wire [11:0] p1_add_81724_comb;
  wire [11:0] p1_add_81725_comb;
  wire [11:0] p1_add_81726_comb;
  wire [11:0] p1_add_81727_comb;
  wire [11:0] p1_add_81728_comb;
  wire [11:0] p1_add_81729_comb;
  wire [11:0] p1_add_81730_comb;
  wire [11:0] p1_add_81875_comb;
  wire [11:0] p1_add_81876_comb;
  wire [11:0] p1_add_81877_comb;
  wire [11:0] p1_add_81878_comb;
  wire [11:0] p1_add_81879_comb;
  wire [11:0] p1_add_81880_comb;
  wire [11:0] p1_add_81881_comb;
  wire [11:0] p1_add_81882_comb;
  wire [11:0] p1_add_81955_comb;
  wire [11:0] p1_add_81956_comb;
  wire [11:0] p1_add_81957_comb;
  wire [11:0] p1_add_81958_comb;
  wire [11:0] p1_add_81959_comb;
  wire [11:0] p1_add_81960_comb;
  wire [11:0] p1_add_81961_comb;
  wire [11:0] p1_add_81962_comb;
  wire [24:0] p1_sum__1736_comb;
  wire [24:0] p1_sum__1737_comb;
  wire [24:0] p1_sum__1738_comb;
  wire [24:0] p1_sum__1739_comb;
  wire [24:0] p1_sum__1708_comb;
  wire [24:0] p1_sum__1709_comb;
  wire [24:0] p1_sum__1710_comb;
  wire [24:0] p1_sum__1711_comb;
  wire [24:0] p1_sum__1680_comb;
  wire [24:0] p1_sum__1681_comb;
  wire [24:0] p1_sum__1682_comb;
  wire [24:0] p1_sum__1683_comb;
  wire [24:0] p1_sum__1652_comb;
  wire [24:0] p1_sum__1653_comb;
  wire [24:0] p1_sum__1654_comb;
  wire [24:0] p1_sum__1655_comb;
  wire [24:0] p1_sum__1760_comb;
  wire [24:0] p1_sum__1761_comb;
  wire [24:0] p1_sum__1762_comb;
  wire [24:0] p1_sum__1763_comb;
  wire [24:0] p1_sum__1628_comb;
  wire [24:0] p1_sum__1629_comb;
  wire [24:0] p1_sum__1630_comb;
  wire [24:0] p1_sum__1631_comb;
  wire [24:0] p1_sum__1780_comb;
  wire [24:0] p1_sum__1781_comb;
  wire [24:0] p1_sum__1782_comb;
  wire [24:0] p1_sum__1783_comb;
  wire [24:0] p1_sum__1608_comb;
  wire [24:0] p1_sum__1609_comb;
  wire [24:0] p1_sum__1610_comb;
  wire [24:0] p1_sum__1611_comb;
  wire [18:0] p1_bit_slice_81299_comb;
  wire [17:0] p1_add_81300_comb;
  wire [17:0] p1_add_81301_comb;
  wire [18:0] p1_bit_slice_81302_comb;
  wire [18:0] p1_bit_slice_81303_comb;
  wire [17:0] p1_add_81304_comb;
  wire [17:0] p1_add_81305_comb;
  wire [18:0] p1_bit_slice_81306_comb;
  wire [18:0] p1_bit_slice_81307_comb;
  wire [17:0] p1_add_81308_comb;
  wire [17:0] p1_add_81309_comb;
  wire [18:0] p1_bit_slice_81310_comb;
  wire [18:0] p1_bit_slice_81311_comb;
  wire [17:0] p1_add_81312_comb;
  wire [17:0] p1_add_81313_comb;
  wire [18:0] p1_bit_slice_81314_comb;
  wire [17:0] p1_smul_81315_comb;
  wire [17:0] p1_smul_81318_comb;
  wire [17:0] p1_smul_81319_comb;
  wire [17:0] p1_smul_81322_comb;
  wire [17:0] p1_smul_81323_comb;
  wire [17:0] p1_smul_81326_comb;
  wire [17:0] p1_smul_81327_comb;
  wire [17:0] p1_smul_81330_comb;
  wire [17:0] p1_smul_81331_comb;
  wire [17:0] p1_smul_81334_comb;
  wire [17:0] p1_smul_81335_comb;
  wire [17:0] p1_smul_81338_comb;
  wire [17:0] p1_smul_81339_comb;
  wire [17:0] p1_smul_81342_comb;
  wire [17:0] p1_smul_81343_comb;
  wire [17:0] p1_smul_81346_comb;
  wire [18:0] p1_add_81347_comb;
  wire [18:0] p1_add_81349_comb;
  wire [18:0] p1_add_81351_comb;
  wire [18:0] p1_add_81353_comb;
  wire [18:0] p1_add_81355_comb;
  wire [18:0] p1_add_81357_comb;
  wire [18:0] p1_add_81359_comb;
  wire [18:0] p1_add_81361_comb;
  wire [18:0] p1_add_81363_comb;
  wire [18:0] p1_add_81365_comb;
  wire [18:0] p1_add_81367_comb;
  wire [18:0] p1_add_81369_comb;
  wire [18:0] p1_add_81371_comb;
  wire [18:0] p1_add_81373_comb;
  wire [18:0] p1_add_81375_comb;
  wire [18:0] p1_add_81377_comb;
  wire [18:0] p1_add_81411_comb;
  wire [18:0] p1_add_81413_comb;
  wire [18:0] p1_add_81415_comb;
  wire [18:0] p1_add_81417_comb;
  wire [18:0] p1_add_81419_comb;
  wire [18:0] p1_add_81421_comb;
  wire [18:0] p1_add_81423_comb;
  wire [18:0] p1_add_81425_comb;
  wire [18:0] p1_add_81427_comb;
  wire [18:0] p1_add_81429_comb;
  wire [18:0] p1_add_81431_comb;
  wire [18:0] p1_add_81433_comb;
  wire [18:0] p1_add_81435_comb;
  wire [18:0] p1_add_81437_comb;
  wire [18:0] p1_add_81439_comb;
  wire [18:0] p1_add_81441_comb;
  wire [17:0] p1_smul_81444_comb;
  wire [17:0] p1_smul_81446_comb;
  wire [17:0] p1_smul_81447_comb;
  wire [17:0] p1_smul_81449_comb;
  wire [17:0] p1_smul_81452_comb;
  wire [17:0] p1_smul_81454_comb;
  wire [17:0] p1_smul_81455_comb;
  wire [17:0] p1_smul_81457_comb;
  wire [17:0] p1_smul_81460_comb;
  wire [17:0] p1_smul_81462_comb;
  wire [17:0] p1_smul_81463_comb;
  wire [17:0] p1_smul_81465_comb;
  wire [17:0] p1_smul_81468_comb;
  wire [17:0] p1_smul_81470_comb;
  wire [17:0] p1_smul_81471_comb;
  wire [17:0] p1_smul_81473_comb;
  wire [17:0] p1_add_81475_comb;
  wire [18:0] p1_bit_slice_81476_comb;
  wire [18:0] p1_bit_slice_81477_comb;
  wire [17:0] p1_add_81478_comb;
  wire [17:0] p1_add_81479_comb;
  wire [18:0] p1_bit_slice_81480_comb;
  wire [18:0] p1_bit_slice_81481_comb;
  wire [17:0] p1_add_81482_comb;
  wire [17:0] p1_add_81483_comb;
  wire [18:0] p1_bit_slice_81484_comb;
  wire [18:0] p1_bit_slice_81485_comb;
  wire [17:0] p1_add_81486_comb;
  wire [17:0] p1_add_81487_comb;
  wire [18:0] p1_bit_slice_81488_comb;
  wire [18:0] p1_bit_slice_81489_comb;
  wire [17:0] p1_add_81490_comb;
  wire [18:0] p1_bit_slice_81507_comb;
  wire [17:0] p1_add_81508_comb;
  wire [17:0] p1_add_81509_comb;
  wire [18:0] p1_bit_slice_81510_comb;
  wire [18:0] p1_bit_slice_81511_comb;
  wire [17:0] p1_add_81512_comb;
  wire [17:0] p1_add_81513_comb;
  wire [18:0] p1_bit_slice_81514_comb;
  wire [17:0] p1_smul_81515_comb;
  wire [17:0] p1_smul_81518_comb;
  wire [17:0] p1_smul_81519_comb;
  wire [17:0] p1_smul_81522_comb;
  wire [17:0] p1_smul_81523_comb;
  wire [17:0] p1_smul_81526_comb;
  wire [17:0] p1_smul_81527_comb;
  wire [17:0] p1_smul_81530_comb;
  wire [18:0] p1_add_81531_comb;
  wire [18:0] p1_add_81533_comb;
  wire [18:0] p1_add_81535_comb;
  wire [18:0] p1_add_81537_comb;
  wire [18:0] p1_add_81539_comb;
  wire [18:0] p1_add_81541_comb;
  wire [18:0] p1_add_81543_comb;
  wire [18:0] p1_add_81545_comb;
  wire [18:0] p1_add_81563_comb;
  wire [18:0] p1_add_81565_comb;
  wire [18:0] p1_add_81567_comb;
  wire [18:0] p1_add_81569_comb;
  wire [18:0] p1_add_81571_comb;
  wire [18:0] p1_add_81573_comb;
  wire [18:0] p1_add_81575_comb;
  wire [18:0] p1_add_81577_comb;
  wire [17:0] p1_smul_81580_comb;
  wire [17:0] p1_smul_81582_comb;
  wire [17:0] p1_smul_81583_comb;
  wire [17:0] p1_smul_81585_comb;
  wire [17:0] p1_smul_81588_comb;
  wire [17:0] p1_smul_81590_comb;
  wire [17:0] p1_smul_81591_comb;
  wire [17:0] p1_smul_81593_comb;
  wire [17:0] p1_add_81595_comb;
  wire [18:0] p1_bit_slice_81596_comb;
  wire [18:0] p1_bit_slice_81597_comb;
  wire [17:0] p1_add_81598_comb;
  wire [17:0] p1_add_81599_comb;
  wire [18:0] p1_bit_slice_81600_comb;
  wire [18:0] p1_bit_slice_81601_comb;
  wire [17:0] p1_add_81602_comb;
  wire [18:0] p1_bit_slice_81619_comb;
  wire [17:0] p1_add_81620_comb;
  wire [17:0] p1_add_81621_comb;
  wire [18:0] p1_bit_slice_81622_comb;
  wire [18:0] p1_bit_slice_81623_comb;
  wire [17:0] p1_add_81624_comb;
  wire [17:0] p1_add_81625_comb;
  wire [18:0] p1_bit_slice_81626_comb;
  wire [17:0] p1_smul_81627_comb;
  wire [17:0] p1_smul_81630_comb;
  wire [17:0] p1_smul_81631_comb;
  wire [17:0] p1_smul_81634_comb;
  wire [17:0] p1_smul_81635_comb;
  wire [17:0] p1_smul_81638_comb;
  wire [17:0] p1_smul_81639_comb;
  wire [17:0] p1_smul_81642_comb;
  wire [18:0] p1_add_81643_comb;
  wire [18:0] p1_add_81645_comb;
  wire [18:0] p1_add_81647_comb;
  wire [18:0] p1_add_81649_comb;
  wire [18:0] p1_add_81651_comb;
  wire [18:0] p1_add_81653_comb;
  wire [18:0] p1_add_81655_comb;
  wire [18:0] p1_add_81657_comb;
  wire [18:0] p1_add_81675_comb;
  wire [18:0] p1_add_81677_comb;
  wire [18:0] p1_add_81679_comb;
  wire [18:0] p1_add_81681_comb;
  wire [18:0] p1_add_81683_comb;
  wire [18:0] p1_add_81685_comb;
  wire [18:0] p1_add_81687_comb;
  wire [18:0] p1_add_81689_comb;
  wire [17:0] p1_smul_81692_comb;
  wire [17:0] p1_smul_81694_comb;
  wire [17:0] p1_smul_81695_comb;
  wire [17:0] p1_smul_81697_comb;
  wire [17:0] p1_smul_81700_comb;
  wire [17:0] p1_smul_81702_comb;
  wire [17:0] p1_smul_81703_comb;
  wire [17:0] p1_smul_81705_comb;
  wire [17:0] p1_add_81707_comb;
  wire [18:0] p1_bit_slice_81708_comb;
  wire [18:0] p1_bit_slice_81709_comb;
  wire [17:0] p1_add_81710_comb;
  wire [17:0] p1_add_81711_comb;
  wire [18:0] p1_bit_slice_81712_comb;
  wire [18:0] p1_bit_slice_81713_comb;
  wire [17:0] p1_add_81714_comb;
  wire [24:0] p1_sum__1324_comb;
  wire [24:0] p1_sum__1325_comb;
  wire [24:0] p1_sum__1310_comb;
  wire [24:0] p1_sum__1311_comb;
  wire [24:0] p1_sum__1296_comb;
  wire [24:0] p1_sum__1297_comb;
  wire [24:0] p1_sum__1282_comb;
  wire [24:0] p1_sum__1283_comb;
  wire [24:0] p1_sum__1336_comb;
  wire [24:0] p1_sum__1337_comb;
  wire [24:0] p1_sum__1270_comb;
  wire [24:0] p1_sum__1271_comb;
  wire [24:0] p1_sum__1346_comb;
  wire [24:0] p1_sum__1347_comb;
  wire [24:0] p1_sum__1260_comb;
  wire [24:0] p1_sum__1261_comb;
  wire [17:0] p1_add_81747_comb;
  wire [17:0] p1_add_81749_comb;
  wire [17:0] p1_add_81751_comb;
  wire [17:0] p1_add_81753_comb;
  wire [17:0] p1_add_81755_comb;
  wire [17:0] p1_add_81757_comb;
  wire [17:0] p1_add_81759_comb;
  wire [17:0] p1_add_81761_comb;
  wire [17:0] p1_add_81763_comb;
  wire [17:0] p1_add_81765_comb;
  wire [17:0] p1_add_81767_comb;
  wire [17:0] p1_add_81769_comb;
  wire [17:0] p1_add_81771_comb;
  wire [17:0] p1_add_81773_comb;
  wire [17:0] p1_add_81775_comb;
  wire [17:0] p1_add_81777_comb;
  wire [19:0] p1_concat_81779_comb;
  wire [19:0] p1_concat_81780_comb;
  wire [19:0] p1_concat_81781_comb;
  wire [19:0] p1_concat_81782_comb;
  wire [19:0] p1_concat_81783_comb;
  wire [19:0] p1_concat_81784_comb;
  wire [19:0] p1_concat_81785_comb;
  wire [19:0] p1_concat_81786_comb;
  wire [19:0] p1_concat_81787_comb;
  wire [19:0] p1_concat_81788_comb;
  wire [19:0] p1_concat_81789_comb;
  wire [19:0] p1_concat_81790_comb;
  wire [19:0] p1_concat_81791_comb;
  wire [19:0] p1_concat_81792_comb;
  wire [19:0] p1_concat_81793_comb;
  wire [19:0] p1_concat_81794_comb;
  wire [19:0] p1_concat_81811_comb;
  wire [19:0] p1_concat_81812_comb;
  wire [19:0] p1_concat_81813_comb;
  wire [19:0] p1_concat_81814_comb;
  wire [19:0] p1_concat_81815_comb;
  wire [19:0] p1_concat_81816_comb;
  wire [19:0] p1_concat_81817_comb;
  wire [19:0] p1_concat_81818_comb;
  wire [19:0] p1_concat_81819_comb;
  wire [19:0] p1_concat_81820_comb;
  wire [19:0] p1_concat_81821_comb;
  wire [19:0] p1_concat_81822_comb;
  wire [19:0] p1_concat_81823_comb;
  wire [19:0] p1_concat_81824_comb;
  wire [19:0] p1_concat_81825_comb;
  wire [19:0] p1_concat_81826_comb;
  wire [17:0] p1_add_81827_comb;
  wire [17:0] p1_add_81829_comb;
  wire [17:0] p1_add_81831_comb;
  wire [17:0] p1_add_81833_comb;
  wire [17:0] p1_add_81835_comb;
  wire [17:0] p1_add_81837_comb;
  wire [17:0] p1_add_81839_comb;
  wire [17:0] p1_add_81841_comb;
  wire [17:0] p1_add_81843_comb;
  wire [17:0] p1_add_81845_comb;
  wire [17:0] p1_add_81847_comb;
  wire [17:0] p1_add_81849_comb;
  wire [17:0] p1_add_81851_comb;
  wire [17:0] p1_add_81853_comb;
  wire [17:0] p1_add_81855_comb;
  wire [17:0] p1_add_81857_comb;
  wire [17:0] p1_add_81891_comb;
  wire [17:0] p1_add_81893_comb;
  wire [17:0] p1_add_81895_comb;
  wire [17:0] p1_add_81897_comb;
  wire [17:0] p1_add_81899_comb;
  wire [17:0] p1_add_81901_comb;
  wire [17:0] p1_add_81903_comb;
  wire [17:0] p1_add_81905_comb;
  wire [19:0] p1_concat_81907_comb;
  wire [19:0] p1_concat_81908_comb;
  wire [19:0] p1_concat_81909_comb;
  wire [19:0] p1_concat_81910_comb;
  wire [19:0] p1_concat_81911_comb;
  wire [19:0] p1_concat_81912_comb;
  wire [19:0] p1_concat_81913_comb;
  wire [19:0] p1_concat_81914_comb;
  wire [19:0] p1_concat_81923_comb;
  wire [19:0] p1_concat_81924_comb;
  wire [19:0] p1_concat_81925_comb;
  wire [19:0] p1_concat_81926_comb;
  wire [19:0] p1_concat_81927_comb;
  wire [19:0] p1_concat_81928_comb;
  wire [19:0] p1_concat_81929_comb;
  wire [19:0] p1_concat_81930_comb;
  wire [17:0] p1_add_81931_comb;
  wire [17:0] p1_add_81933_comb;
  wire [17:0] p1_add_81935_comb;
  wire [17:0] p1_add_81937_comb;
  wire [17:0] p1_add_81939_comb;
  wire [17:0] p1_add_81941_comb;
  wire [17:0] p1_add_81943_comb;
  wire [17:0] p1_add_81945_comb;
  wire [17:0] p1_add_81971_comb;
  wire [17:0] p1_add_81973_comb;
  wire [17:0] p1_add_81975_comb;
  wire [17:0] p1_add_81977_comb;
  wire [17:0] p1_add_81979_comb;
  wire [17:0] p1_add_81981_comb;
  wire [17:0] p1_add_81983_comb;
  wire [17:0] p1_add_81985_comb;
  wire [19:0] p1_concat_81987_comb;
  wire [19:0] p1_concat_81988_comb;
  wire [19:0] p1_concat_81989_comb;
  wire [19:0] p1_concat_81990_comb;
  wire [19:0] p1_concat_81991_comb;
  wire [19:0] p1_concat_81992_comb;
  wire [19:0] p1_concat_81993_comb;
  wire [19:0] p1_concat_81994_comb;
  wire [19:0] p1_concat_82003_comb;
  wire [19:0] p1_concat_82004_comb;
  wire [19:0] p1_concat_82005_comb;
  wire [19:0] p1_concat_82006_comb;
  wire [19:0] p1_concat_82007_comb;
  wire [19:0] p1_concat_82008_comb;
  wire [19:0] p1_concat_82009_comb;
  wire [19:0] p1_concat_82010_comb;
  wire [17:0] p1_add_82011_comb;
  wire [17:0] p1_add_82013_comb;
  wire [17:0] p1_add_82015_comb;
  wire [17:0] p1_add_82017_comb;
  wire [17:0] p1_add_82019_comb;
  wire [17:0] p1_add_82021_comb;
  wire [17:0] p1_add_82023_comb;
  wire [17:0] p1_add_82025_comb;
  wire [23:0] p1_add_82291_comb;
  wire [23:0] p1_add_82292_comb;
  wire [23:0] p1_add_82293_comb;
  wire [23:0] p1_add_82294_comb;
  wire [23:0] p1_add_82295_comb;
  wire [23:0] p1_add_82296_comb;
  wire [23:0] p1_add_82297_comb;
  wire [23:0] p1_add_82298_comb;
  wire [23:0] p1_add_82371_comb;
  wire [23:0] p1_add_82372_comb;
  wire [23:0] p1_add_82373_comb;
  wire [23:0] p1_add_82374_comb;
  wire [23:0] p1_add_82411_comb;
  wire [23:0] p1_add_82412_comb;
  wire [23:0] p1_add_82413_comb;
  wire [23:0] p1_add_82414_comb;
  wire [24:0] p1_sum__1118_comb;
  wire [24:0] p1_sum__1111_comb;
  wire [24:0] p1_sum__1104_comb;
  wire [24:0] p1_sum__1097_comb;
  wire [24:0] p1_sum__1124_comb;
  wire [24:0] p1_sum__1091_comb;
  wire [24:0] p1_sum__1129_comb;
  wire [24:0] p1_sum__1086_comb;
  wire [23:0] p1_add_82051_comb;
  wire [23:0] p1_add_82053_comb;
  wire [23:0] p1_add_82055_comb;
  wire [23:0] p1_add_82057_comb;
  wire [23:0] p1_add_82059_comb;
  wire [23:0] p1_add_82061_comb;
  wire [23:0] p1_add_82063_comb;
  wire [23:0] p1_add_82065_comb;
  wire [18:0] p1_concat_82067_comb;
  wire [18:0] p1_concat_82068_comb;
  wire [18:0] p1_concat_82069_comb;
  wire [18:0] p1_concat_82070_comb;
  wire [18:0] p1_concat_82071_comb;
  wire [18:0] p1_concat_82072_comb;
  wire [18:0] p1_concat_82073_comb;
  wire [18:0] p1_concat_82074_comb;
  wire [18:0] p1_concat_82075_comb;
  wire [18:0] p1_concat_82076_comb;
  wire [18:0] p1_concat_82077_comb;
  wire [18:0] p1_concat_82078_comb;
  wire [18:0] p1_concat_82079_comb;
  wire [18:0] p1_concat_82080_comb;
  wire [18:0] p1_concat_82081_comb;
  wire [18:0] p1_concat_82082_comb;
  wire [24:0] p1_sum__1756_comb;
  wire [24:0] p1_sum__1757_comb;
  wire [24:0] p1_sum__1758_comb;
  wire [24:0] p1_sum__1759_comb;
  wire [24:0] p1_sum__1732_comb;
  wire [24:0] p1_sum__1733_comb;
  wire [24:0] p1_sum__1734_comb;
  wire [24:0] p1_sum__1735_comb;
  wire [24:0] p1_sum__1704_comb;
  wire [24:0] p1_sum__1705_comb;
  wire [24:0] p1_sum__1706_comb;
  wire [24:0] p1_sum__1707_comb;
  wire [24:0] p1_sum__1676_comb;
  wire [24:0] p1_sum__1677_comb;
  wire [24:0] p1_sum__1678_comb;
  wire [24:0] p1_sum__1679_comb;
  wire [24:0] p1_sum__1712_comb;
  wire [24:0] p1_sum__1713_comb;
  wire [24:0] p1_sum__1714_comb;
  wire [24:0] p1_sum__1715_comb;
  wire [24:0] p1_sum__1684_comb;
  wire [24:0] p1_sum__1685_comb;
  wire [24:0] p1_sum__1686_comb;
  wire [24:0] p1_sum__1687_comb;
  wire [24:0] p1_sum__1656_comb;
  wire [24:0] p1_sum__1657_comb;
  wire [24:0] p1_sum__1658_comb;
  wire [24:0] p1_sum__1659_comb;
  wire [24:0] p1_sum__1632_comb;
  wire [24:0] p1_sum__1633_comb;
  wire [24:0] p1_sum__1634_comb;
  wire [24:0] p1_sum__1635_comb;
  wire [18:0] p1_concat_82131_comb;
  wire [18:0] p1_concat_82132_comb;
  wire [18:0] p1_concat_82133_comb;
  wire [18:0] p1_concat_82134_comb;
  wire [18:0] p1_concat_82135_comb;
  wire [18:0] p1_concat_82136_comb;
  wire [18:0] p1_concat_82137_comb;
  wire [18:0] p1_concat_82138_comb;
  wire [18:0] p1_concat_82139_comb;
  wire [18:0] p1_concat_82140_comb;
  wire [18:0] p1_concat_82141_comb;
  wire [18:0] p1_concat_82142_comb;
  wire [18:0] p1_concat_82143_comb;
  wire [18:0] p1_concat_82144_comb;
  wire [18:0] p1_concat_82145_comb;
  wire [18:0] p1_concat_82146_comb;
  wire [23:0] p1_add_82147_comb;
  wire [23:0] p1_add_82149_comb;
  wire [23:0] p1_add_82151_comb;
  wire [23:0] p1_add_82153_comb;
  wire [23:0] p1_add_82155_comb;
  wire [23:0] p1_add_82157_comb;
  wire [23:0] p1_add_82159_comb;
  wire [23:0] p1_add_82161_comb;
  wire [23:0] p1_add_82171_comb;
  wire [23:0] p1_add_82173_comb;
  wire [23:0] p1_add_82175_comb;
  wire [23:0] p1_add_82177_comb;
  wire [18:0] p1_concat_82179_comb;
  wire [18:0] p1_concat_82180_comb;
  wire [18:0] p1_concat_82181_comb;
  wire [18:0] p1_concat_82182_comb;
  wire [18:0] p1_concat_82183_comb;
  wire [18:0] p1_concat_82184_comb;
  wire [18:0] p1_concat_82185_comb;
  wire [18:0] p1_concat_82186_comb;
  wire [24:0] p1_sum__1776_comb;
  wire [24:0] p1_sum__1777_comb;
  wire [24:0] p1_sum__1778_comb;
  wire [24:0] p1_sum__1779_comb;
  wire [24:0] p1_sum__1648_comb;
  wire [24:0] p1_sum__1649_comb;
  wire [24:0] p1_sum__1650_comb;
  wire [24:0] p1_sum__1651_comb;
  wire [24:0] p1_sum__1740_comb;
  wire [24:0] p1_sum__1741_comb;
  wire [24:0] p1_sum__1742_comb;
  wire [24:0] p1_sum__1743_comb;
  wire [24:0] p1_sum__1612_comb;
  wire [24:0] p1_sum__1613_comb;
  wire [24:0] p1_sum__1614_comb;
  wire [24:0] p1_sum__1615_comb;
  wire [18:0] p1_concat_82211_comb;
  wire [18:0] p1_concat_82212_comb;
  wire [18:0] p1_concat_82213_comb;
  wire [18:0] p1_concat_82214_comb;
  wire [18:0] p1_concat_82215_comb;
  wire [18:0] p1_concat_82216_comb;
  wire [18:0] p1_concat_82217_comb;
  wire [18:0] p1_concat_82218_comb;
  wire [23:0] p1_add_82219_comb;
  wire [23:0] p1_add_82221_comb;
  wire [23:0] p1_add_82223_comb;
  wire [23:0] p1_add_82225_comb;
  wire [23:0] p1_add_82235_comb;
  wire [23:0] p1_add_82237_comb;
  wire [23:0] p1_add_82239_comb;
  wire [23:0] p1_add_82241_comb;
  wire [18:0] p1_concat_82243_comb;
  wire [18:0] p1_concat_82244_comb;
  wire [18:0] p1_concat_82245_comb;
  wire [18:0] p1_concat_82246_comb;
  wire [18:0] p1_concat_82247_comb;
  wire [18:0] p1_concat_82248_comb;
  wire [18:0] p1_concat_82249_comb;
  wire [18:0] p1_concat_82250_comb;
  wire [24:0] p1_sum__1792_comb;
  wire [24:0] p1_sum__1793_comb;
  wire [24:0] p1_sum__1794_comb;
  wire [24:0] p1_sum__1795_comb;
  wire [24:0] p1_sum__1624_comb;
  wire [24:0] p1_sum__1625_comb;
  wire [24:0] p1_sum__1626_comb;
  wire [24:0] p1_sum__1627_comb;
  wire [24:0] p1_sum__1764_comb;
  wire [24:0] p1_sum__1765_comb;
  wire [24:0] p1_sum__1766_comb;
  wire [24:0] p1_sum__1767_comb;
  wire [24:0] p1_sum__1596_comb;
  wire [24:0] p1_sum__1597_comb;
  wire [24:0] p1_sum__1598_comb;
  wire [24:0] p1_sum__1599_comb;
  wire [18:0] p1_concat_82275_comb;
  wire [18:0] p1_concat_82276_comb;
  wire [18:0] p1_concat_82277_comb;
  wire [18:0] p1_concat_82278_comb;
  wire [18:0] p1_concat_82279_comb;
  wire [18:0] p1_concat_82280_comb;
  wire [18:0] p1_concat_82281_comb;
  wire [18:0] p1_concat_82282_comb;
  wire [23:0] p1_add_82283_comb;
  wire [23:0] p1_add_82285_comb;
  wire [23:0] p1_add_82287_comb;
  wire [23:0] p1_add_82289_comb;
  wire [23:0] p1_add_82451_comb;
  wire [23:0] p1_add_82453_comb;
  wire [23:0] p1_add_82455_comb;
  wire [23:0] p1_add_82457_comb;
  wire [23:0] p1_add_82515_comb;
  wire [23:0] p1_add_82517_comb;
  wire [23:0] p1_add_82547_comb;
  wire [23:0] p1_add_82549_comb;
  wire [24:0] p1_add_82595_comb;
  wire [24:0] p1_add_82596_comb;
  wire [24:0] p1_add_82597_comb;
  wire [24:0] p1_add_82598_comb;
  wire [24:0] p1_add_82619_comb;
  wire [24:0] p1_add_82620_comb;
  wire [24:0] p1_add_82635_comb;
  wire [24:0] p1_add_82636_comb;
  wire [24:0] p1_sum__1348_comb;
  wire [24:0] p1_sum__1349_comb;
  wire [24:0] p1_sum__1340_comb;
  wire [24:0] p1_sum__1341_comb;
  wire [24:0] p1_sum__1330_comb;
  wire [24:0] p1_sum__1331_comb;
  wire [24:0] p1_sum__1318_comb;
  wire [24:0] p1_sum__1319_comb;
  wire [24:0] p1_sum__1334_comb;
  wire [24:0] p1_sum__1335_comb;
  wire [24:0] p1_sum__1322_comb;
  wire [24:0] p1_sum__1323_comb;
  wire [24:0] p1_sum__1308_comb;
  wire [24:0] p1_sum__1309_comb;
  wire [24:0] p1_sum__1294_comb;
  wire [24:0] p1_sum__1295_comb;
  wire [24:0] p1_sum__1312_comb;
  wire [24:0] p1_sum__1313_comb;
  wire [24:0] p1_sum__1298_comb;
  wire [24:0] p1_sum__1299_comb;
  wire [24:0] p1_sum__1284_comb;
  wire [24:0] p1_sum__1285_comb;
  wire [24:0] p1_sum__1272_comb;
  wire [24:0] p1_sum__1273_comb;
  wire [24:0] p1_sum__1288_comb;
  wire [24:0] p1_sum__1289_comb;
  wire [24:0] p1_sum__1276_comb;
  wire [24:0] p1_sum__1277_comb;
  wire [24:0] p1_sum__1266_comb;
  wire [24:0] p1_sum__1267_comb;
  wire [24:0] p1_sum__1258_comb;
  wire [24:0] p1_sum__1259_comb;
  wire [24:0] p1_sum__1354_comb;
  wire [24:0] p1_sum__1355_comb;
  wire [24:0] p1_sum__1304_comb;
  wire [24:0] p1_sum__1305_comb;
  wire [24:0] p1_sum__1344_comb;
  wire [24:0] p1_sum__1345_comb;
  wire [24:0] p1_sum__1280_comb;
  wire [24:0] p1_sum__1281_comb;
  wire [24:0] p1_sum__1326_comb;
  wire [24:0] p1_sum__1327_comb;
  wire [24:0] p1_sum__1262_comb;
  wire [24:0] p1_sum__1263_comb;
  wire [24:0] p1_sum__1302_comb;
  wire [24:0] p1_sum__1303_comb;
  wire [24:0] p1_sum__1252_comb;
  wire [24:0] p1_sum__1253_comb;
  wire [24:0] p1_sum__1358_comb;
  wire [24:0] p1_sum__1359_comb;
  wire [24:0] p1_sum__1290_comb;
  wire [24:0] p1_sum__1291_comb;
  wire [24:0] p1_sum__1352_comb;
  wire [24:0] p1_sum__1353_comb;
  wire [24:0] p1_sum__1268_comb;
  wire [24:0] p1_sum__1269_comb;
  wire [24:0] p1_sum__1338_comb;
  wire [24:0] p1_sum__1339_comb;
  wire [24:0] p1_sum__1254_comb;
  wire [24:0] p1_sum__1255_comb;
  wire [24:0] p1_sum__1316_comb;
  wire [24:0] p1_sum__1317_comb;
  wire [24:0] p1_sum__1248_comb;
  wire [24:0] p1_sum__1249_comb;
  wire [23:0] p1_umul_28108_NarrowedMult__comb;
  wire [23:0] p1_umul_28110_NarrowedMult__comb;
  wire [23:0] p1_umul_28112_NarrowedMult__comb;
  wire [23:0] p1_umul_28114_NarrowedMult__comb;
  wire [23:0] p1_umul_28106_NarrowedMult__comb;
  wire [23:0] p1_umul_28116_NarrowedMult__comb;
  wire [23:0] p1_umul_28104_NarrowedMult__comb;
  wire [23:0] p1_umul_28118_NarrowedMult__comb;
  wire [16:0] p1_bit_slice_82659_comb;
  wire [16:0] p1_bit_slice_82660_comb;
  wire [16:0] p1_bit_slice_82661_comb;
  wire [16:0] p1_bit_slice_82662_comb;
  wire [16:0] p1_bit_slice_82683_comb;
  wire [16:0] p1_bit_slice_82684_comb;
  wire [16:0] p1_bit_slice_82699_comb;
  wire [16:0] p1_bit_slice_82700_comb;
  wire [24:0] p1_sum__1130_comb;
  wire [24:0] p1_sum__1126_comb;
  wire [24:0] p1_sum__1121_comb;
  wire [24:0] p1_sum__1115_comb;
  wire [23:0] p1_add_82467_comb;
  wire [23:0] p1_add_82468_comb;
  wire [23:0] p1_add_82469_comb;
  wire [23:0] p1_add_82470_comb;
  wire [23:0] p1_add_82471_comb;
  wire [23:0] p1_add_82472_comb;
  wire [23:0] p1_add_82473_comb;
  wire [23:0] p1_add_82474_comb;
  wire [24:0] p1_sum__1123_comb;
  wire [24:0] p1_sum__1117_comb;
  wire [24:0] p1_sum__1110_comb;
  wire [24:0] p1_sum__1103_comb;
  wire [24:0] p1_sum__1112_comb;
  wire [24:0] p1_sum__1105_comb;
  wire [24:0] p1_sum__1098_comb;
  wire [24:0] p1_sum__1092_comb;
  wire [23:0] p1_add_82499_comb;
  wire [23:0] p1_add_82500_comb;
  wire [23:0] p1_add_82501_comb;
  wire [23:0] p1_add_82502_comb;
  wire [23:0] p1_add_82503_comb;
  wire [23:0] p1_add_82504_comb;
  wire [23:0] p1_add_82505_comb;
  wire [23:0] p1_add_82506_comb;
  wire [24:0] p1_sum__1100_comb;
  wire [24:0] p1_sum__1094_comb;
  wire [24:0] p1_sum__1089_comb;
  wire [24:0] p1_sum__1085_comb;
  wire [24:0] p1_sum__1133_comb;
  wire [24:0] p1_sum__1108_comb;
  wire [23:0] p1_add_82523_comb;
  wire [23:0] p1_add_82524_comb;
  wire [23:0] p1_add_82525_comb;
  wire [23:0] p1_add_82526_comb;
  wire [24:0] p1_sum__1128_comb;
  wire [24:0] p1_sum__1096_comb;
  wire [24:0] p1_sum__1119_comb;
  wire [24:0] p1_sum__1087_comb;
  wire [23:0] p1_add_82539_comb;
  wire [23:0] p1_add_82540_comb;
  wire [23:0] p1_add_82541_comb;
  wire [23:0] p1_add_82542_comb;
  wire [24:0] p1_sum__1107_comb;
  wire [24:0] p1_sum__1082_comb;
  wire [24:0] p1_sum__1135_comb;
  wire [24:0] p1_sum__1101_comb;
  wire [23:0] p1_add_82555_comb;
  wire [23:0] p1_add_82556_comb;
  wire [23:0] p1_add_82557_comb;
  wire [23:0] p1_add_82558_comb;
  wire [24:0] p1_sum__1132_comb;
  wire [24:0] p1_sum__1090_comb;
  wire [24:0] p1_sum__1125_comb;
  wire [24:0] p1_sum__1083_comb;
  wire [23:0] p1_add_82571_comb;
  wire [23:0] p1_add_82572_comb;
  wire [23:0] p1_add_82573_comb;
  wire [23:0] p1_add_82574_comb;
  wire [24:0] p1_sum__1114_comb;
  wire [24:0] p1_sum__1080_comb;
  wire [16:0] p1_bit_slice_82643_comb;
  wire [16:0] p1_bit_slice_82644_comb;
  wire [16:0] p1_bit_slice_82645_comb;
  wire [16:0] p1_bit_slice_82646_comb;
  wire [16:0] p1_bit_slice_82675_comb;
  wire [16:0] p1_bit_slice_82676_comb;
  wire [16:0] p1_bit_slice_82691_comb;
  wire [16:0] p1_bit_slice_82692_comb;
  wire [24:0] p1_add_82583_comb;
  wire [24:0] p1_add_82584_comb;
  wire [24:0] p1_add_82585_comb;
  wire [24:0] p1_add_82586_comb;
  wire [23:0] p1_add_82587_comb;
  wire [23:0] p1_add_82588_comb;
  wire [23:0] p1_add_82589_comb;
  wire [23:0] p1_add_82590_comb;
  wire [24:0] p1_add_82591_comb;
  wire [24:0] p1_add_82592_comb;
  wire [24:0] p1_add_82593_comb;
  wire [24:0] p1_add_82594_comb;
  wire [24:0] p1_add_82599_comb;
  wire [24:0] p1_add_82600_comb;
  wire [24:0] p1_add_82601_comb;
  wire [24:0] p1_add_82602_comb;
  wire [23:0] p1_add_82603_comb;
  wire [23:0] p1_add_82604_comb;
  wire [23:0] p1_add_82605_comb;
  wire [23:0] p1_add_82606_comb;
  wire [24:0] p1_add_82607_comb;
  wire [24:0] p1_add_82608_comb;
  wire [24:0] p1_add_82609_comb;
  wire [24:0] p1_add_82610_comb;
  wire [24:0] p1_add_82613_comb;
  wire [24:0] p1_add_82614_comb;
  wire [23:0] p1_add_82615_comb;
  wire [23:0] p1_add_82616_comb;
  wire [24:0] p1_add_82617_comb;
  wire [24:0] p1_add_82618_comb;
  wire [24:0] p1_add_82621_comb;
  wire [24:0] p1_add_82622_comb;
  wire [23:0] p1_add_82623_comb;
  wire [23:0] p1_add_82624_comb;
  wire [24:0] p1_add_82625_comb;
  wire [24:0] p1_add_82626_comb;
  wire [24:0] p1_add_82629_comb;
  wire [24:0] p1_add_82630_comb;
  wire [23:0] p1_add_82631_comb;
  wire [23:0] p1_add_82632_comb;
  wire [24:0] p1_add_82633_comb;
  wire [24:0] p1_add_82634_comb;
  wire [24:0] p1_add_82637_comb;
  wire [24:0] p1_add_82638_comb;
  wire [23:0] p1_add_82639_comb;
  wire [23:0] p1_add_82640_comb;
  wire [24:0] p1_add_82641_comb;
  wire [24:0] p1_add_82642_comb;
  wire [17:0] p1_add_82851_comb;
  wire [17:0] p1_add_82852_comb;
  wire [17:0] p1_add_82853_comb;
  wire [17:0] p1_add_82854_comb;
  wire [17:0] p1_add_82875_comb;
  wire [17:0] p1_add_82876_comb;
  wire [17:0] p1_add_82891_comb;
  wire [17:0] p1_add_82892_comb;
  wire [16:0] p1_bit_slice_82647_comb;
  wire [16:0] p1_bit_slice_82648_comb;
  wire [16:0] p1_bit_slice_82649_comb;
  wire [16:0] p1_bit_slice_82650_comb;
  wire [16:0] p1_bit_slice_82651_comb;
  wire [16:0] p1_bit_slice_82652_comb;
  wire [16:0] p1_bit_slice_82653_comb;
  wire [16:0] p1_bit_slice_82654_comb;
  wire [16:0] p1_bit_slice_82655_comb;
  wire [16:0] p1_bit_slice_82656_comb;
  wire [16:0] p1_bit_slice_82657_comb;
  wire [16:0] p1_bit_slice_82658_comb;
  wire [16:0] p1_bit_slice_82663_comb;
  wire [16:0] p1_bit_slice_82664_comb;
  wire [16:0] p1_bit_slice_82665_comb;
  wire [16:0] p1_bit_slice_82666_comb;
  wire [16:0] p1_bit_slice_82667_comb;
  wire [16:0] p1_bit_slice_82668_comb;
  wire [16:0] p1_bit_slice_82669_comb;
  wire [16:0] p1_bit_slice_82670_comb;
  wire [16:0] p1_bit_slice_82671_comb;
  wire [16:0] p1_bit_slice_82672_comb;
  wire [16:0] p1_bit_slice_82673_comb;
  wire [16:0] p1_bit_slice_82674_comb;
  wire [16:0] p1_bit_slice_82677_comb;
  wire [16:0] p1_bit_slice_82678_comb;
  wire [16:0] p1_bit_slice_82679_comb;
  wire [16:0] p1_bit_slice_82680_comb;
  wire [16:0] p1_bit_slice_82681_comb;
  wire [16:0] p1_bit_slice_82682_comb;
  wire [16:0] p1_bit_slice_82685_comb;
  wire [16:0] p1_bit_slice_82686_comb;
  wire [16:0] p1_bit_slice_82687_comb;
  wire [16:0] p1_bit_slice_82688_comb;
  wire [16:0] p1_bit_slice_82689_comb;
  wire [16:0] p1_bit_slice_82690_comb;
  wire [16:0] p1_bit_slice_82693_comb;
  wire [16:0] p1_bit_slice_82694_comb;
  wire [16:0] p1_bit_slice_82695_comb;
  wire [16:0] p1_bit_slice_82696_comb;
  wire [16:0] p1_bit_slice_82697_comb;
  wire [16:0] p1_bit_slice_82698_comb;
  wire [16:0] p1_bit_slice_82701_comb;
  wire [16:0] p1_bit_slice_82702_comb;
  wire [16:0] p1_bit_slice_82703_comb;
  wire [16:0] p1_bit_slice_82704_comb;
  wire [16:0] p1_bit_slice_82705_comb;
  wire [16:0] p1_bit_slice_82706_comb;
  wire [17:0] p1_add_82835_comb;
  wire [17:0] p1_add_82836_comb;
  wire [17:0] p1_add_82837_comb;
  wire [17:0] p1_add_82838_comb;
  wire [17:0] p1_add_82867_comb;
  wire [17:0] p1_add_82868_comb;
  wire [17:0] p1_add_82883_comb;
  wire [17:0] p1_add_82884_comb;
  wire [9:0] p1_bit_slice_82903_comb;
  wire [9:0] p1_bit_slice_82904_comb;
  wire [9:0] p1_bit_slice_82905_comb;
  wire [9:0] p1_bit_slice_82906_comb;
  wire [9:0] p1_bit_slice_82909_comb;
  wire [9:0] p1_bit_slice_82910_comb;
  wire [9:0] p1_bit_slice_82913_comb;
  wire [9:0] p1_bit_slice_82914_comb;
  wire [9:0] p1_bit_slice_82899_comb;
  wire [9:0] p1_bit_slice_82900_comb;
  wire [9:0] p1_bit_slice_82901_comb;
  wire [9:0] p1_bit_slice_82902_comb;
  wire [9:0] p1_bit_slice_82907_comb;
  wire [9:0] p1_bit_slice_82908_comb;
  wire [9:0] p1_bit_slice_82911_comb;
  wire [9:0] p1_bit_slice_82912_comb;
  wire [17:0] p1_add_82839_comb;
  wire [17:0] p1_add_82840_comb;
  wire [17:0] p1_add_82841_comb;
  wire [17:0] p1_add_82842_comb;
  wire [17:0] p1_add_82843_comb;
  wire [17:0] p1_add_82844_comb;
  wire [17:0] p1_add_82845_comb;
  wire [17:0] p1_add_82846_comb;
  wire [17:0] p1_add_82847_comb;
  wire [17:0] p1_add_82848_comb;
  wire [17:0] p1_add_82849_comb;
  wire [17:0] p1_add_82850_comb;
  wire [17:0] p1_add_82855_comb;
  wire [17:0] p1_add_82856_comb;
  wire [17:0] p1_add_82857_comb;
  wire [17:0] p1_add_82858_comb;
  wire [17:0] p1_add_82859_comb;
  wire [17:0] p1_add_82860_comb;
  wire [17:0] p1_add_82861_comb;
  wire [17:0] p1_add_82862_comb;
  wire [17:0] p1_add_82863_comb;
  wire [17:0] p1_add_82864_comb;
  wire [17:0] p1_add_82865_comb;
  wire [17:0] p1_add_82866_comb;
  wire [17:0] p1_add_82869_comb;
  wire [17:0] p1_add_82870_comb;
  wire [17:0] p1_add_82871_comb;
  wire [17:0] p1_add_82872_comb;
  wire [17:0] p1_add_82873_comb;
  wire [17:0] p1_add_82874_comb;
  wire [17:0] p1_add_82877_comb;
  wire [17:0] p1_add_82878_comb;
  wire [17:0] p1_add_82879_comb;
  wire [17:0] p1_add_82880_comb;
  wire [17:0] p1_add_82881_comb;
  wire [17:0] p1_add_82882_comb;
  wire [17:0] p1_add_82885_comb;
  wire [17:0] p1_add_82886_comb;
  wire [17:0] p1_add_82887_comb;
  wire [17:0] p1_add_82888_comb;
  wire [17:0] p1_add_82889_comb;
  wire [17:0] p1_add_82890_comb;
  wire [17:0] p1_add_82893_comb;
  wire [17:0] p1_add_82894_comb;
  wire [17:0] p1_add_82895_comb;
  wire [17:0] p1_add_82896_comb;
  wire [17:0] p1_add_82897_comb;
  wire [17:0] p1_add_82898_comb;
  wire [10:0] p1_sign_ext_82915_comb;
  wire [10:0] p1_sign_ext_82916_comb;
  wire [10:0] p1_sign_ext_82917_comb;
  wire [10:0] p1_sign_ext_82918_comb;
  wire [10:0] p1_sign_ext_82927_comb;
  wire [10:0] p1_sign_ext_82928_comb;
  wire [10:0] p1_sign_ext_82933_comb;
  wire [10:0] p1_sign_ext_82934_comb;
  wire [6:0] p1_bit_slice_82939_comb;
  wire [6:0] p1_bit_slice_82940_comb;
  wire [6:0] p1_bit_slice_82941_comb;
  wire [6:0] p1_bit_slice_82942_comb;
  wire [10:0] p1_add_82943_comb;
  wire [6:0] p1_bit_slice_82944_comb;
  wire [10:0] p1_add_82945_comb;
  wire [6:0] p1_bit_slice_82946_comb;
  wire [10:0] p1_add_82947_comb;
  wire [6:0] p1_bit_slice_82948_comb;
  wire [10:0] p1_add_82949_comb;
  wire [6:0] p1_bit_slice_82950_comb;
  wire [6:0] p1_bit_slice_82951_comb;
  wire [6:0] p1_bit_slice_82952_comb;
  wire [10:0] p1_add_82953_comb;
  wire [6:0] p1_bit_slice_82954_comb;
  wire [10:0] p1_add_82955_comb;
  wire [6:0] p1_bit_slice_82956_comb;
  wire [6:0] p1_bit_slice_82957_comb;
  wire [6:0] p1_bit_slice_82958_comb;
  wire [10:0] p1_add_82959_comb;
  wire [6:0] p1_bit_slice_82960_comb;
  wire [10:0] p1_add_82961_comb;
  wire [6:0] p1_bit_slice_82962_comb;
  assign p1_array_index_79763_comb = p0_x[3'h2][3'h2];
  assign p1_array_index_79764_comb = p0_x[3'h2][3'h3];
  assign p1_array_index_79765_comb = p0_x[3'h2][3'h4];
  assign p1_array_index_79766_comb = p0_x[3'h2][3'h5];
  assign p1_array_index_79767_comb = p0_x[3'h3][3'h2];
  assign p1_array_index_79768_comb = p0_x[3'h3][3'h3];
  assign p1_array_index_79769_comb = p0_x[3'h3][3'h4];
  assign p1_array_index_79770_comb = p0_x[3'h3][3'h5];
  assign p1_array_index_79771_comb = p0_x[3'h4][3'h2];
  assign p1_array_index_79772_comb = p0_x[3'h4][3'h3];
  assign p1_array_index_79773_comb = p0_x[3'h4][3'h4];
  assign p1_array_index_79774_comb = p0_x[3'h4][3'h5];
  assign p1_array_index_79775_comb = p0_x[3'h5][3'h2];
  assign p1_array_index_79776_comb = p0_x[3'h5][3'h3];
  assign p1_array_index_79777_comb = p0_x[3'h5][3'h4];
  assign p1_array_index_79778_comb = p0_x[3'h5][3'h5];
  assign p1_array_index_79779_comb = p0_x[3'h2][3'h1];
  assign p1_array_index_79780_comb = p0_x[3'h2][3'h6];
  assign p1_array_index_79781_comb = p0_x[3'h3][3'h1];
  assign p1_array_index_79782_comb = p0_x[3'h3][3'h6];
  assign p1_array_index_79783_comb = p0_x[3'h4][3'h1];
  assign p1_array_index_79784_comb = p0_x[3'h4][3'h6];
  assign p1_array_index_79785_comb = p0_x[3'h5][3'h1];
  assign p1_array_index_79786_comb = p0_x[3'h5][3'h6];
  assign p1_array_index_79787_comb = p0_x[3'h2][3'h0];
  assign p1_array_index_79788_comb = p0_x[3'h2][3'h7];
  assign p1_array_index_79789_comb = p0_x[3'h3][3'h0];
  assign p1_array_index_79790_comb = p0_x[3'h3][3'h7];
  assign p1_array_index_79791_comb = p0_x[3'h4][3'h0];
  assign p1_array_index_79792_comb = p0_x[3'h4][3'h7];
  assign p1_array_index_79793_comb = p0_x[3'h5][3'h0];
  assign p1_array_index_79794_comb = p0_x[3'h5][3'h7];
  assign p1_array_index_79795_comb = p0_x[3'h1][3'h2];
  assign p1_array_index_79796_comb = p0_x[3'h1][3'h3];
  assign p1_array_index_79797_comb = p0_x[3'h1][3'h4];
  assign p1_array_index_79798_comb = p0_x[3'h1][3'h5];
  assign p1_array_index_79799_comb = p0_x[3'h6][3'h2];
  assign p1_array_index_79800_comb = p0_x[3'h6][3'h3];
  assign p1_array_index_79801_comb = p0_x[3'h6][3'h4];
  assign p1_array_index_79802_comb = p0_x[3'h6][3'h5];
  assign p1_array_index_79803_comb = p0_x[3'h1][3'h1];
  assign p1_array_index_79804_comb = p0_x[3'h1][3'h6];
  assign p1_array_index_79805_comb = p0_x[3'h6][3'h1];
  assign p1_array_index_79806_comb = p0_x[3'h6][3'h6];
  assign p1_array_index_79807_comb = p0_x[3'h1][3'h0];
  assign p1_array_index_79808_comb = p0_x[3'h1][3'h7];
  assign p1_array_index_79809_comb = p0_x[3'h6][3'h0];
  assign p1_array_index_79810_comb = p0_x[3'h6][3'h7];
  assign p1_array_index_79811_comb = p0_x[3'h0][3'h2];
  assign p1_array_index_79812_comb = p0_x[3'h0][3'h3];
  assign p1_array_index_79813_comb = p0_x[3'h0][3'h4];
  assign p1_array_index_79814_comb = p0_x[3'h0][3'h5];
  assign p1_array_index_79815_comb = p0_x[3'h7][3'h2];
  assign p1_array_index_79816_comb = p0_x[3'h7][3'h3];
  assign p1_array_index_79817_comb = p0_x[3'h7][3'h4];
  assign p1_array_index_79818_comb = p0_x[3'h7][3'h5];
  assign p1_array_index_79819_comb = p0_x[3'h0][3'h1];
  assign p1_array_index_79820_comb = p0_x[3'h0][3'h6];
  assign p1_array_index_79821_comb = p0_x[3'h7][3'h1];
  assign p1_array_index_79822_comb = p0_x[3'h7][3'h6];
  assign p1_array_index_79823_comb = p0_x[3'h0][3'h0];
  assign p1_array_index_79824_comb = p0_x[3'h0][3'h7];
  assign p1_array_index_79825_comb = p0_x[3'h7][3'h0];
  assign p1_array_index_79826_comb = p0_x[3'h7][3'h7];
  assign p1_bit_slice_79827_comb = p1_array_index_79763_comb[9:7];
  assign p1_bit_slice_79828_comb = p1_array_index_79764_comb[9:7];
  assign p1_bit_slice_79829_comb = p1_array_index_79765_comb[9:7];
  assign p1_bit_slice_79830_comb = p1_array_index_79766_comb[9:7];
  assign p1_bit_slice_79831_comb = p1_array_index_79767_comb[9:7];
  assign p1_bit_slice_79832_comb = p1_array_index_79768_comb[9:7];
  assign p1_bit_slice_79833_comb = p1_array_index_79769_comb[9:7];
  assign p1_bit_slice_79834_comb = p1_array_index_79770_comb[9:7];
  assign p1_bit_slice_79835_comb = p1_array_index_79771_comb[9:7];
  assign p1_bit_slice_79836_comb = p1_array_index_79772_comb[9:7];
  assign p1_bit_slice_79837_comb = p1_array_index_79773_comb[9:7];
  assign p1_bit_slice_79838_comb = p1_array_index_79774_comb[9:7];
  assign p1_bit_slice_79839_comb = p1_array_index_79775_comb[9:7];
  assign p1_bit_slice_79840_comb = p1_array_index_79776_comb[9:7];
  assign p1_bit_slice_79841_comb = p1_array_index_79777_comb[9:7];
  assign p1_bit_slice_79842_comb = p1_array_index_79778_comb[9:7];
  assign p1_bit_slice_79843_comb = p1_array_index_79779_comb[9:7];
  assign p1_bit_slice_79844_comb = p1_array_index_79780_comb[9:7];
  assign p1_bit_slice_79845_comb = p1_array_index_79781_comb[9:7];
  assign p1_bit_slice_79846_comb = p1_array_index_79782_comb[9:7];
  assign p1_bit_slice_79847_comb = p1_array_index_79783_comb[9:7];
  assign p1_bit_slice_79848_comb = p1_array_index_79784_comb[9:7];
  assign p1_bit_slice_79849_comb = p1_array_index_79785_comb[9:7];
  assign p1_bit_slice_79850_comb = p1_array_index_79786_comb[9:7];
  assign p1_bit_slice_79851_comb = p1_array_index_79787_comb[9:7];
  assign p1_bit_slice_79852_comb = p1_array_index_79788_comb[9:7];
  assign p1_bit_slice_79853_comb = p1_array_index_79789_comb[9:7];
  assign p1_bit_slice_79854_comb = p1_array_index_79790_comb[9:7];
  assign p1_bit_slice_79855_comb = p1_array_index_79791_comb[9:7];
  assign p1_bit_slice_79856_comb = p1_array_index_79792_comb[9:7];
  assign p1_bit_slice_79857_comb = p1_array_index_79793_comb[9:7];
  assign p1_bit_slice_79858_comb = p1_array_index_79794_comb[9:7];
  assign p1_bit_slice_79859_comb = p1_array_index_79795_comb[9:7];
  assign p1_bit_slice_79860_comb = p1_array_index_79796_comb[9:7];
  assign p1_bit_slice_79861_comb = p1_array_index_79797_comb[9:7];
  assign p1_bit_slice_79862_comb = p1_array_index_79798_comb[9:7];
  assign p1_bit_slice_79863_comb = p1_array_index_79799_comb[9:7];
  assign p1_bit_slice_79864_comb = p1_array_index_79800_comb[9:7];
  assign p1_bit_slice_79865_comb = p1_array_index_79801_comb[9:7];
  assign p1_bit_slice_79866_comb = p1_array_index_79802_comb[9:7];
  assign p1_bit_slice_79867_comb = p1_array_index_79803_comb[9:7];
  assign p1_bit_slice_79868_comb = p1_array_index_79804_comb[9:7];
  assign p1_bit_slice_79869_comb = p1_array_index_79805_comb[9:7];
  assign p1_bit_slice_79870_comb = p1_array_index_79806_comb[9:7];
  assign p1_bit_slice_79871_comb = p1_array_index_79807_comb[9:7];
  assign p1_bit_slice_79872_comb = p1_array_index_79808_comb[9:7];
  assign p1_bit_slice_79873_comb = p1_array_index_79809_comb[9:7];
  assign p1_bit_slice_79874_comb = p1_array_index_79810_comb[9:7];
  assign p1_bit_slice_79875_comb = p1_array_index_79811_comb[9:7];
  assign p1_bit_slice_79876_comb = p1_array_index_79812_comb[9:7];
  assign p1_bit_slice_79877_comb = p1_array_index_79813_comb[9:7];
  assign p1_bit_slice_79878_comb = p1_array_index_79814_comb[9:7];
  assign p1_bit_slice_79879_comb = p1_array_index_79815_comb[9:7];
  assign p1_bit_slice_79880_comb = p1_array_index_79816_comb[9:7];
  assign p1_bit_slice_79881_comb = p1_array_index_79817_comb[9:7];
  assign p1_bit_slice_79882_comb = p1_array_index_79818_comb[9:7];
  assign p1_bit_slice_79883_comb = p1_array_index_79819_comb[9:7];
  assign p1_bit_slice_79884_comb = p1_array_index_79820_comb[9:7];
  assign p1_bit_slice_79885_comb = p1_array_index_79821_comb[9:7];
  assign p1_bit_slice_79886_comb = p1_array_index_79822_comb[9:7];
  assign p1_bit_slice_79887_comb = p1_array_index_79823_comb[9:7];
  assign p1_bit_slice_79888_comb = p1_array_index_79824_comb[9:7];
  assign p1_bit_slice_79889_comb = p1_array_index_79825_comb[9:7];
  assign p1_bit_slice_79890_comb = p1_array_index_79826_comb[9:7];
  assign p1_add_80019_comb = {{1{p1_bit_slice_79827_comb[2]}}, p1_bit_slice_79827_comb} + 4'hf;
  assign p1_add_80021_comb = {{1{p1_bit_slice_79828_comb[2]}}, p1_bit_slice_79828_comb} + 4'hf;
  assign p1_add_80023_comb = {{1{p1_bit_slice_79829_comb[2]}}, p1_bit_slice_79829_comb} + 4'hf;
  assign p1_add_80025_comb = {{1{p1_bit_slice_79830_comb[2]}}, p1_bit_slice_79830_comb} + 4'hf;
  assign p1_add_80027_comb = {{1{p1_bit_slice_79831_comb[2]}}, p1_bit_slice_79831_comb} + 4'hf;
  assign p1_add_80029_comb = {{1{p1_bit_slice_79832_comb[2]}}, p1_bit_slice_79832_comb} + 4'hf;
  assign p1_add_80031_comb = {{1{p1_bit_slice_79833_comb[2]}}, p1_bit_slice_79833_comb} + 4'hf;
  assign p1_add_80033_comb = {{1{p1_bit_slice_79834_comb[2]}}, p1_bit_slice_79834_comb} + 4'hf;
  assign p1_add_80035_comb = {{1{p1_bit_slice_79835_comb[2]}}, p1_bit_slice_79835_comb} + 4'hf;
  assign p1_add_80037_comb = {{1{p1_bit_slice_79836_comb[2]}}, p1_bit_slice_79836_comb} + 4'hf;
  assign p1_add_80039_comb = {{1{p1_bit_slice_79837_comb[2]}}, p1_bit_slice_79837_comb} + 4'hf;
  assign p1_add_80041_comb = {{1{p1_bit_slice_79838_comb[2]}}, p1_bit_slice_79838_comb} + 4'hf;
  assign p1_add_80043_comb = {{1{p1_bit_slice_79839_comb[2]}}, p1_bit_slice_79839_comb} + 4'hf;
  assign p1_add_80045_comb = {{1{p1_bit_slice_79840_comb[2]}}, p1_bit_slice_79840_comb} + 4'hf;
  assign p1_add_80047_comb = {{1{p1_bit_slice_79841_comb[2]}}, p1_bit_slice_79841_comb} + 4'hf;
  assign p1_add_80049_comb = {{1{p1_bit_slice_79842_comb[2]}}, p1_bit_slice_79842_comb} + 4'hf;
  assign p1_add_80051_comb = {{1{p1_bit_slice_79843_comb[2]}}, p1_bit_slice_79843_comb} + 4'hf;
  assign p1_add_80053_comb = {{1{p1_bit_slice_79844_comb[2]}}, p1_bit_slice_79844_comb} + 4'hf;
  assign p1_add_80055_comb = {{1{p1_bit_slice_79845_comb[2]}}, p1_bit_slice_79845_comb} + 4'hf;
  assign p1_add_80057_comb = {{1{p1_bit_slice_79846_comb[2]}}, p1_bit_slice_79846_comb} + 4'hf;
  assign p1_add_80059_comb = {{1{p1_bit_slice_79847_comb[2]}}, p1_bit_slice_79847_comb} + 4'hf;
  assign p1_add_80061_comb = {{1{p1_bit_slice_79848_comb[2]}}, p1_bit_slice_79848_comb} + 4'hf;
  assign p1_add_80063_comb = {{1{p1_bit_slice_79849_comb[2]}}, p1_bit_slice_79849_comb} + 4'hf;
  assign p1_add_80065_comb = {{1{p1_bit_slice_79850_comb[2]}}, p1_bit_slice_79850_comb} + 4'hf;
  assign p1_add_80067_comb = {{1{p1_bit_slice_79851_comb[2]}}, p1_bit_slice_79851_comb} + 4'hf;
  assign p1_add_80069_comb = {{1{p1_bit_slice_79852_comb[2]}}, p1_bit_slice_79852_comb} + 4'hf;
  assign p1_add_80071_comb = {{1{p1_bit_slice_79853_comb[2]}}, p1_bit_slice_79853_comb} + 4'hf;
  assign p1_add_80073_comb = {{1{p1_bit_slice_79854_comb[2]}}, p1_bit_slice_79854_comb} + 4'hf;
  assign p1_add_80075_comb = {{1{p1_bit_slice_79855_comb[2]}}, p1_bit_slice_79855_comb} + 4'hf;
  assign p1_add_80077_comb = {{1{p1_bit_slice_79856_comb[2]}}, p1_bit_slice_79856_comb} + 4'hf;
  assign p1_add_80079_comb = {{1{p1_bit_slice_79857_comb[2]}}, p1_bit_slice_79857_comb} + 4'hf;
  assign p1_add_80081_comb = {{1{p1_bit_slice_79858_comb[2]}}, p1_bit_slice_79858_comb} + 4'hf;
  assign p1_add_80083_comb = {{1{p1_bit_slice_79859_comb[2]}}, p1_bit_slice_79859_comb} + 4'hf;
  assign p1_add_80085_comb = {{1{p1_bit_slice_79860_comb[2]}}, p1_bit_slice_79860_comb} + 4'hf;
  assign p1_add_80087_comb = {{1{p1_bit_slice_79861_comb[2]}}, p1_bit_slice_79861_comb} + 4'hf;
  assign p1_add_80089_comb = {{1{p1_bit_slice_79862_comb[2]}}, p1_bit_slice_79862_comb} + 4'hf;
  assign p1_add_80091_comb = {{1{p1_bit_slice_79863_comb[2]}}, p1_bit_slice_79863_comb} + 4'hf;
  assign p1_add_80093_comb = {{1{p1_bit_slice_79864_comb[2]}}, p1_bit_slice_79864_comb} + 4'hf;
  assign p1_add_80095_comb = {{1{p1_bit_slice_79865_comb[2]}}, p1_bit_slice_79865_comb} + 4'hf;
  assign p1_add_80097_comb = {{1{p1_bit_slice_79866_comb[2]}}, p1_bit_slice_79866_comb} + 4'hf;
  assign p1_add_80099_comb = {{1{p1_bit_slice_79867_comb[2]}}, p1_bit_slice_79867_comb} + 4'hf;
  assign p1_add_80101_comb = {{1{p1_bit_slice_79868_comb[2]}}, p1_bit_slice_79868_comb} + 4'hf;
  assign p1_add_80103_comb = {{1{p1_bit_slice_79869_comb[2]}}, p1_bit_slice_79869_comb} + 4'hf;
  assign p1_add_80105_comb = {{1{p1_bit_slice_79870_comb[2]}}, p1_bit_slice_79870_comb} + 4'hf;
  assign p1_add_80107_comb = {{1{p1_bit_slice_79871_comb[2]}}, p1_bit_slice_79871_comb} + 4'hf;
  assign p1_add_80109_comb = {{1{p1_bit_slice_79872_comb[2]}}, p1_bit_slice_79872_comb} + 4'hf;
  assign p1_add_80111_comb = {{1{p1_bit_slice_79873_comb[2]}}, p1_bit_slice_79873_comb} + 4'hf;
  assign p1_add_80113_comb = {{1{p1_bit_slice_79874_comb[2]}}, p1_bit_slice_79874_comb} + 4'hf;
  assign p1_add_80115_comb = {{1{p1_bit_slice_79875_comb[2]}}, p1_bit_slice_79875_comb} + 4'hf;
  assign p1_add_80117_comb = {{1{p1_bit_slice_79876_comb[2]}}, p1_bit_slice_79876_comb} + 4'hf;
  assign p1_add_80119_comb = {{1{p1_bit_slice_79877_comb[2]}}, p1_bit_slice_79877_comb} + 4'hf;
  assign p1_add_80121_comb = {{1{p1_bit_slice_79878_comb[2]}}, p1_bit_slice_79878_comb} + 4'hf;
  assign p1_add_80123_comb = {{1{p1_bit_slice_79879_comb[2]}}, p1_bit_slice_79879_comb} + 4'hf;
  assign p1_add_80125_comb = {{1{p1_bit_slice_79880_comb[2]}}, p1_bit_slice_79880_comb} + 4'hf;
  assign p1_add_80127_comb = {{1{p1_bit_slice_79881_comb[2]}}, p1_bit_slice_79881_comb} + 4'hf;
  assign p1_add_80129_comb = {{1{p1_bit_slice_79882_comb[2]}}, p1_bit_slice_79882_comb} + 4'hf;
  assign p1_add_80131_comb = {{1{p1_bit_slice_79883_comb[2]}}, p1_bit_slice_79883_comb} + 4'hf;
  assign p1_add_80133_comb = {{1{p1_bit_slice_79884_comb[2]}}, p1_bit_slice_79884_comb} + 4'hf;
  assign p1_add_80135_comb = {{1{p1_bit_slice_79885_comb[2]}}, p1_bit_slice_79885_comb} + 4'hf;
  assign p1_add_80137_comb = {{1{p1_bit_slice_79886_comb[2]}}, p1_bit_slice_79886_comb} + 4'hf;
  assign p1_add_80139_comb = {{1{p1_bit_slice_79887_comb[2]}}, p1_bit_slice_79887_comb} + 4'hf;
  assign p1_add_80141_comb = {{1{p1_bit_slice_79888_comb[2]}}, p1_bit_slice_79888_comb} + 4'hf;
  assign p1_add_80143_comb = {{1{p1_bit_slice_79889_comb[2]}}, p1_bit_slice_79889_comb} + 4'hf;
  assign p1_add_80145_comb = {{1{p1_bit_slice_79890_comb[2]}}, p1_bit_slice_79890_comb} + 4'hf;
  assign p1_concat_80147_comb = {p1_add_80019_comb, p1_array_index_79763_comb[6:0]};
  assign p1_concat_80148_comb = {p1_add_80021_comb, p1_array_index_79764_comb[6:0]};
  assign p1_concat_80149_comb = {p1_add_80023_comb, p1_array_index_79765_comb[6:0]};
  assign p1_concat_80150_comb = {p1_add_80025_comb, p1_array_index_79766_comb[6:0]};
  assign p1_concat_80151_comb = {p1_add_80027_comb, p1_array_index_79767_comb[6:0]};
  assign p1_concat_80152_comb = {p1_add_80029_comb, p1_array_index_79768_comb[6:0]};
  assign p1_concat_80153_comb = {p1_add_80031_comb, p1_array_index_79769_comb[6:0]};
  assign p1_concat_80154_comb = {p1_add_80033_comb, p1_array_index_79770_comb[6:0]};
  assign p1_concat_80155_comb = {p1_add_80035_comb, p1_array_index_79771_comb[6:0]};
  assign p1_concat_80156_comb = {p1_add_80037_comb, p1_array_index_79772_comb[6:0]};
  assign p1_concat_80157_comb = {p1_add_80039_comb, p1_array_index_79773_comb[6:0]};
  assign p1_concat_80158_comb = {p1_add_80041_comb, p1_array_index_79774_comb[6:0]};
  assign p1_concat_80159_comb = {p1_add_80043_comb, p1_array_index_79775_comb[6:0]};
  assign p1_concat_80160_comb = {p1_add_80045_comb, p1_array_index_79776_comb[6:0]};
  assign p1_concat_80161_comb = {p1_add_80047_comb, p1_array_index_79777_comb[6:0]};
  assign p1_concat_80162_comb = {p1_add_80049_comb, p1_array_index_79778_comb[6:0]};
  assign p1_concat_80163_comb = {p1_add_80051_comb, p1_array_index_79779_comb[6:0]};
  assign p1_concat_80164_comb = {p1_add_80053_comb, p1_array_index_79780_comb[6:0]};
  assign p1_concat_80165_comb = {p1_add_80055_comb, p1_array_index_79781_comb[6:0]};
  assign p1_concat_80166_comb = {p1_add_80057_comb, p1_array_index_79782_comb[6:0]};
  assign p1_concat_80167_comb = {p1_add_80059_comb, p1_array_index_79783_comb[6:0]};
  assign p1_concat_80168_comb = {p1_add_80061_comb, p1_array_index_79784_comb[6:0]};
  assign p1_concat_80169_comb = {p1_add_80063_comb, p1_array_index_79785_comb[6:0]};
  assign p1_concat_80170_comb = {p1_add_80065_comb, p1_array_index_79786_comb[6:0]};
  assign p1_concat_80171_comb = {p1_add_80067_comb, p1_array_index_79787_comb[6:0]};
  assign p1_concat_80172_comb = {p1_add_80069_comb, p1_array_index_79788_comb[6:0]};
  assign p1_concat_80173_comb = {p1_add_80071_comb, p1_array_index_79789_comb[6:0]};
  assign p1_concat_80174_comb = {p1_add_80073_comb, p1_array_index_79790_comb[6:0]};
  assign p1_concat_80175_comb = {p1_add_80075_comb, p1_array_index_79791_comb[6:0]};
  assign p1_concat_80176_comb = {p1_add_80077_comb, p1_array_index_79792_comb[6:0]};
  assign p1_concat_80177_comb = {p1_add_80079_comb, p1_array_index_79793_comb[6:0]};
  assign p1_concat_80178_comb = {p1_add_80081_comb, p1_array_index_79794_comb[6:0]};
  assign p1_concat_80179_comb = {p1_add_80083_comb, p1_array_index_79795_comb[6:0]};
  assign p1_concat_80180_comb = {p1_add_80085_comb, p1_array_index_79796_comb[6:0]};
  assign p1_concat_80181_comb = {p1_add_80087_comb, p1_array_index_79797_comb[6:0]};
  assign p1_concat_80182_comb = {p1_add_80089_comb, p1_array_index_79798_comb[6:0]};
  assign p1_concat_80183_comb = {p1_add_80091_comb, p1_array_index_79799_comb[6:0]};
  assign p1_concat_80184_comb = {p1_add_80093_comb, p1_array_index_79800_comb[6:0]};
  assign p1_concat_80185_comb = {p1_add_80095_comb, p1_array_index_79801_comb[6:0]};
  assign p1_concat_80186_comb = {p1_add_80097_comb, p1_array_index_79802_comb[6:0]};
  assign p1_concat_80187_comb = {p1_add_80099_comb, p1_array_index_79803_comb[6:0]};
  assign p1_concat_80188_comb = {p1_add_80101_comb, p1_array_index_79804_comb[6:0]};
  assign p1_concat_80189_comb = {p1_add_80103_comb, p1_array_index_79805_comb[6:0]};
  assign p1_concat_80190_comb = {p1_add_80105_comb, p1_array_index_79806_comb[6:0]};
  assign p1_concat_80191_comb = {p1_add_80107_comb, p1_array_index_79807_comb[6:0]};
  assign p1_concat_80192_comb = {p1_add_80109_comb, p1_array_index_79808_comb[6:0]};
  assign p1_concat_80193_comb = {p1_add_80111_comb, p1_array_index_79809_comb[6:0]};
  assign p1_concat_80194_comb = {p1_add_80113_comb, p1_array_index_79810_comb[6:0]};
  assign p1_concat_80195_comb = {p1_add_80115_comb, p1_array_index_79811_comb[6:0]};
  assign p1_concat_80196_comb = {p1_add_80117_comb, p1_array_index_79812_comb[6:0]};
  assign p1_concat_80197_comb = {p1_add_80119_comb, p1_array_index_79813_comb[6:0]};
  assign p1_concat_80198_comb = {p1_add_80121_comb, p1_array_index_79814_comb[6:0]};
  assign p1_concat_80199_comb = {p1_add_80123_comb, p1_array_index_79815_comb[6:0]};
  assign p1_concat_80200_comb = {p1_add_80125_comb, p1_array_index_79816_comb[6:0]};
  assign p1_concat_80201_comb = {p1_add_80127_comb, p1_array_index_79817_comb[6:0]};
  assign p1_concat_80202_comb = {p1_add_80129_comb, p1_array_index_79818_comb[6:0]};
  assign p1_concat_80203_comb = {p1_add_80131_comb, p1_array_index_79819_comb[6:0]};
  assign p1_concat_80204_comb = {p1_add_80133_comb, p1_array_index_79820_comb[6:0]};
  assign p1_concat_80205_comb = {p1_add_80135_comb, p1_array_index_79821_comb[6:0]};
  assign p1_concat_80206_comb = {p1_add_80137_comb, p1_array_index_79822_comb[6:0]};
  assign p1_concat_80207_comb = {p1_add_80139_comb, p1_array_index_79823_comb[6:0]};
  assign p1_concat_80208_comb = {p1_add_80141_comb, p1_array_index_79824_comb[6:0]};
  assign p1_concat_80209_comb = {p1_add_80143_comb, p1_array_index_79825_comb[6:0]};
  assign p1_concat_80210_comb = {p1_add_80145_comb, p1_array_index_79826_comb[6:0]};
  assign p1_sign_ext_80213_comb = {{13{p1_concat_80147_comb[10]}}, p1_concat_80147_comb};
  assign p1_sign_ext_80214_comb = {{13{p1_concat_80148_comb[10]}}, p1_concat_80148_comb};
  assign p1_sign_ext_80215_comb = {{13{p1_concat_80149_comb[10]}}, p1_concat_80149_comb};
  assign p1_sign_ext_80216_comb = {{13{p1_concat_80150_comb[10]}}, p1_concat_80150_comb};
  assign p1_sign_ext_80221_comb = {{13{p1_concat_80151_comb[10]}}, p1_concat_80151_comb};
  assign p1_sign_ext_80222_comb = {{13{p1_concat_80152_comb[10]}}, p1_concat_80152_comb};
  assign p1_sign_ext_80223_comb = {{13{p1_concat_80153_comb[10]}}, p1_concat_80153_comb};
  assign p1_sign_ext_80224_comb = {{13{p1_concat_80154_comb[10]}}, p1_concat_80154_comb};
  assign p1_sign_ext_80229_comb = {{13{p1_concat_80155_comb[10]}}, p1_concat_80155_comb};
  assign p1_sign_ext_80230_comb = {{13{p1_concat_80156_comb[10]}}, p1_concat_80156_comb};
  assign p1_sign_ext_80231_comb = {{13{p1_concat_80157_comb[10]}}, p1_concat_80157_comb};
  assign p1_sign_ext_80232_comb = {{13{p1_concat_80158_comb[10]}}, p1_concat_80158_comb};
  assign p1_sign_ext_80237_comb = {{13{p1_concat_80159_comb[10]}}, p1_concat_80159_comb};
  assign p1_sign_ext_80238_comb = {{13{p1_concat_80160_comb[10]}}, p1_concat_80160_comb};
  assign p1_sign_ext_80239_comb = {{13{p1_concat_80161_comb[10]}}, p1_concat_80161_comb};
  assign p1_sign_ext_80240_comb = {{13{p1_concat_80162_comb[10]}}, p1_concat_80162_comb};
  assign p1_sign_ext_80243_comb = {{13{p1_concat_80163_comb[10]}}, p1_concat_80163_comb};
  assign p1_sign_ext_80244_comb = {{13{p1_concat_80164_comb[10]}}, p1_concat_80164_comb};
  assign p1_sign_ext_80245_comb = {{13{p1_concat_80165_comb[10]}}, p1_concat_80165_comb};
  assign p1_sign_ext_80246_comb = {{13{p1_concat_80166_comb[10]}}, p1_concat_80166_comb};
  assign p1_sign_ext_80247_comb = {{13{p1_concat_80167_comb[10]}}, p1_concat_80167_comb};
  assign p1_sign_ext_80248_comb = {{13{p1_concat_80168_comb[10]}}, p1_concat_80168_comb};
  assign p1_sign_ext_80249_comb = {{13{p1_concat_80169_comb[10]}}, p1_concat_80169_comb};
  assign p1_sign_ext_80250_comb = {{13{p1_concat_80170_comb[10]}}, p1_concat_80170_comb};
  assign p1_sign_ext_80267_comb = {{13{p1_concat_80171_comb[10]}}, p1_concat_80171_comb};
  assign p1_sign_ext_80272_comb = {{13{p1_concat_80172_comb[10]}}, p1_concat_80172_comb};
  assign p1_sign_ext_80273_comb = {{13{p1_concat_80173_comb[10]}}, p1_concat_80173_comb};
  assign p1_sign_ext_80278_comb = {{13{p1_concat_80174_comb[10]}}, p1_concat_80174_comb};
  assign p1_sign_ext_80279_comb = {{13{p1_concat_80175_comb[10]}}, p1_concat_80175_comb};
  assign p1_sign_ext_80284_comb = {{13{p1_concat_80176_comb[10]}}, p1_concat_80176_comb};
  assign p1_sign_ext_80285_comb = {{13{p1_concat_80177_comb[10]}}, p1_concat_80177_comb};
  assign p1_sign_ext_80290_comb = {{13{p1_concat_80178_comb[10]}}, p1_concat_80178_comb};
  assign p1_sign_ext_80309_comb = {{13{p1_concat_80179_comb[10]}}, p1_concat_80179_comb};
  assign p1_sign_ext_80310_comb = {{13{p1_concat_80180_comb[10]}}, p1_concat_80180_comb};
  assign p1_sign_ext_80311_comb = {{13{p1_concat_80181_comb[10]}}, p1_concat_80181_comb};
  assign p1_sign_ext_80312_comb = {{13{p1_concat_80182_comb[10]}}, p1_concat_80182_comb};
  assign p1_sign_ext_80317_comb = {{13{p1_concat_80183_comb[10]}}, p1_concat_80183_comb};
  assign p1_sign_ext_80318_comb = {{13{p1_concat_80184_comb[10]}}, p1_concat_80184_comb};
  assign p1_sign_ext_80319_comb = {{13{p1_concat_80185_comb[10]}}, p1_concat_80185_comb};
  assign p1_sign_ext_80320_comb = {{13{p1_concat_80186_comb[10]}}, p1_concat_80186_comb};
  assign p1_sign_ext_80323_comb = {{13{p1_concat_80187_comb[10]}}, p1_concat_80187_comb};
  assign p1_sign_ext_80324_comb = {{13{p1_concat_80188_comb[10]}}, p1_concat_80188_comb};
  assign p1_sign_ext_80325_comb = {{13{p1_concat_80189_comb[10]}}, p1_concat_80189_comb};
  assign p1_sign_ext_80326_comb = {{13{p1_concat_80190_comb[10]}}, p1_concat_80190_comb};
  assign p1_sign_ext_80335_comb = {{13{p1_concat_80191_comb[10]}}, p1_concat_80191_comb};
  assign p1_sign_ext_80340_comb = {{13{p1_concat_80192_comb[10]}}, p1_concat_80192_comb};
  assign p1_sign_ext_80341_comb = {{13{p1_concat_80193_comb[10]}}, p1_concat_80193_comb};
  assign p1_sign_ext_80346_comb = {{13{p1_concat_80194_comb[10]}}, p1_concat_80194_comb};
  assign p1_sign_ext_80357_comb = {{13{p1_concat_80195_comb[10]}}, p1_concat_80195_comb};
  assign p1_sign_ext_80358_comb = {{13{p1_concat_80196_comb[10]}}, p1_concat_80196_comb};
  assign p1_sign_ext_80359_comb = {{13{p1_concat_80197_comb[10]}}, p1_concat_80197_comb};
  assign p1_sign_ext_80360_comb = {{13{p1_concat_80198_comb[10]}}, p1_concat_80198_comb};
  assign p1_sign_ext_80365_comb = {{13{p1_concat_80199_comb[10]}}, p1_concat_80199_comb};
  assign p1_sign_ext_80366_comb = {{13{p1_concat_80200_comb[10]}}, p1_concat_80200_comb};
  assign p1_sign_ext_80367_comb = {{13{p1_concat_80201_comb[10]}}, p1_concat_80201_comb};
  assign p1_sign_ext_80368_comb = {{13{p1_concat_80202_comb[10]}}, p1_concat_80202_comb};
  assign p1_sign_ext_80371_comb = {{13{p1_concat_80203_comb[10]}}, p1_concat_80203_comb};
  assign p1_sign_ext_80372_comb = {{13{p1_concat_80204_comb[10]}}, p1_concat_80204_comb};
  assign p1_sign_ext_80373_comb = {{13{p1_concat_80205_comb[10]}}, p1_concat_80205_comb};
  assign p1_sign_ext_80374_comb = {{13{p1_concat_80206_comb[10]}}, p1_concat_80206_comb};
  assign p1_sign_ext_80383_comb = {{13{p1_concat_80207_comb[10]}}, p1_concat_80207_comb};
  assign p1_sign_ext_80388_comb = {{13{p1_concat_80208_comb[10]}}, p1_concat_80208_comb};
  assign p1_sign_ext_80389_comb = {{13{p1_concat_80209_comb[10]}}, p1_concat_80209_comb};
  assign p1_sign_ext_80394_comb = {{13{p1_concat_80210_comb[10]}}, p1_concat_80210_comb};
  assign p1_smul_81379_comb = smul19b_11b_x_9b(p1_concat_80171_comb, 9'h0b5);
  assign p1_smul_81380_comb = smul19b_11b_x_9b(p1_concat_80163_comb, 9'h14b);
  assign p1_smul_81381_comb = smul19b_11b_x_9b(p1_concat_80147_comb, 9'h14b);
  assign p1_smul_81382_comb = smul19b_11b_x_9b(p1_concat_80148_comb, 9'h0b5);
  assign p1_smul_81383_comb = smul19b_11b_x_9b(p1_concat_80149_comb, 9'h0b5);
  assign p1_smul_81384_comb = smul19b_11b_x_9b(p1_concat_80150_comb, 9'h14b);
  assign p1_smul_81385_comb = smul19b_11b_x_9b(p1_concat_80164_comb, 9'h14b);
  assign p1_smul_81386_comb = smul19b_11b_x_9b(p1_concat_80172_comb, 9'h0b5);
  assign p1_smul_81387_comb = smul19b_11b_x_9b(p1_concat_80173_comb, 9'h0b5);
  assign p1_smul_81388_comb = smul19b_11b_x_9b(p1_concat_80165_comb, 9'h14b);
  assign p1_smul_81389_comb = smul19b_11b_x_9b(p1_concat_80151_comb, 9'h14b);
  assign p1_smul_81390_comb = smul19b_11b_x_9b(p1_concat_80152_comb, 9'h0b5);
  assign p1_smul_81391_comb = smul19b_11b_x_9b(p1_concat_80153_comb, 9'h0b5);
  assign p1_smul_81392_comb = smul19b_11b_x_9b(p1_concat_80154_comb, 9'h14b);
  assign p1_smul_81393_comb = smul19b_11b_x_9b(p1_concat_80166_comb, 9'h14b);
  assign p1_smul_81394_comb = smul19b_11b_x_9b(p1_concat_80174_comb, 9'h0b5);
  assign p1_smul_81395_comb = smul19b_11b_x_9b(p1_concat_80175_comb, 9'h0b5);
  assign p1_smul_81396_comb = smul19b_11b_x_9b(p1_concat_80167_comb, 9'h14b);
  assign p1_smul_81397_comb = smul19b_11b_x_9b(p1_concat_80155_comb, 9'h14b);
  assign p1_smul_81398_comb = smul19b_11b_x_9b(p1_concat_80156_comb, 9'h0b5);
  assign p1_smul_81399_comb = smul19b_11b_x_9b(p1_concat_80157_comb, 9'h0b5);
  assign p1_smul_81400_comb = smul19b_11b_x_9b(p1_concat_80158_comb, 9'h14b);
  assign p1_smul_81401_comb = smul19b_11b_x_9b(p1_concat_80168_comb, 9'h14b);
  assign p1_smul_81402_comb = smul19b_11b_x_9b(p1_concat_80176_comb, 9'h0b5);
  assign p1_smul_81403_comb = smul19b_11b_x_9b(p1_concat_80177_comb, 9'h0b5);
  assign p1_smul_81404_comb = smul19b_11b_x_9b(p1_concat_80169_comb, 9'h14b);
  assign p1_smul_81405_comb = smul19b_11b_x_9b(p1_concat_80159_comb, 9'h14b);
  assign p1_smul_81406_comb = smul19b_11b_x_9b(p1_concat_80160_comb, 9'h0b5);
  assign p1_smul_81407_comb = smul19b_11b_x_9b(p1_concat_80161_comb, 9'h0b5);
  assign p1_smul_81408_comb = smul19b_11b_x_9b(p1_concat_80162_comb, 9'h14b);
  assign p1_smul_81409_comb = smul19b_11b_x_9b(p1_concat_80170_comb, 9'h14b);
  assign p1_smul_81410_comb = smul19b_11b_x_9b(p1_concat_80178_comb, 9'h0b5);
  assign p1_smul_81547_comb = smul19b_11b_x_9b(p1_concat_80191_comb, 9'h0b5);
  assign p1_smul_81548_comb = smul19b_11b_x_9b(p1_concat_80187_comb, 9'h14b);
  assign p1_smul_81549_comb = smul19b_11b_x_9b(p1_concat_80179_comb, 9'h14b);
  assign p1_smul_81550_comb = smul19b_11b_x_9b(p1_concat_80180_comb, 9'h0b5);
  assign p1_smul_81551_comb = smul19b_11b_x_9b(p1_concat_80181_comb, 9'h0b5);
  assign p1_smul_81552_comb = smul19b_11b_x_9b(p1_concat_80182_comb, 9'h14b);
  assign p1_smul_81553_comb = smul19b_11b_x_9b(p1_concat_80188_comb, 9'h14b);
  assign p1_smul_81554_comb = smul19b_11b_x_9b(p1_concat_80192_comb, 9'h0b5);
  assign p1_smul_81555_comb = smul19b_11b_x_9b(p1_concat_80193_comb, 9'h0b5);
  assign p1_smul_81556_comb = smul19b_11b_x_9b(p1_concat_80189_comb, 9'h14b);
  assign p1_smul_81557_comb = smul19b_11b_x_9b(p1_concat_80183_comb, 9'h14b);
  assign p1_smul_81558_comb = smul19b_11b_x_9b(p1_concat_80184_comb, 9'h0b5);
  assign p1_smul_81559_comb = smul19b_11b_x_9b(p1_concat_80185_comb, 9'h0b5);
  assign p1_smul_81560_comb = smul19b_11b_x_9b(p1_concat_80186_comb, 9'h14b);
  assign p1_smul_81561_comb = smul19b_11b_x_9b(p1_concat_80190_comb, 9'h14b);
  assign p1_smul_81562_comb = smul19b_11b_x_9b(p1_concat_80194_comb, 9'h0b5);
  assign p1_smul_81659_comb = smul19b_11b_x_9b(p1_concat_80207_comb, 9'h0b5);
  assign p1_smul_81660_comb = smul19b_11b_x_9b(p1_concat_80203_comb, 9'h14b);
  assign p1_smul_81661_comb = smul19b_11b_x_9b(p1_concat_80195_comb, 9'h14b);
  assign p1_smul_81662_comb = smul19b_11b_x_9b(p1_concat_80196_comb, 9'h0b5);
  assign p1_smul_81663_comb = smul19b_11b_x_9b(p1_concat_80197_comb, 9'h0b5);
  assign p1_smul_81664_comb = smul19b_11b_x_9b(p1_concat_80198_comb, 9'h14b);
  assign p1_smul_81665_comb = smul19b_11b_x_9b(p1_concat_80204_comb, 9'h14b);
  assign p1_smul_81666_comb = smul19b_11b_x_9b(p1_concat_80208_comb, 9'h0b5);
  assign p1_smul_81667_comb = smul19b_11b_x_9b(p1_concat_80209_comb, 9'h0b5);
  assign p1_smul_81668_comb = smul19b_11b_x_9b(p1_concat_80205_comb, 9'h14b);
  assign p1_smul_81669_comb = smul19b_11b_x_9b(p1_concat_80199_comb, 9'h14b);
  assign p1_smul_81670_comb = smul19b_11b_x_9b(p1_concat_80200_comb, 9'h0b5);
  assign p1_smul_81671_comb = smul19b_11b_x_9b(p1_concat_80201_comb, 9'h0b5);
  assign p1_smul_81672_comb = smul19b_11b_x_9b(p1_concat_80202_comb, 9'h14b);
  assign p1_smul_81673_comb = smul19b_11b_x_9b(p1_concat_80206_comb, 9'h14b);
  assign p1_smul_81674_comb = smul19b_11b_x_9b(p1_concat_80210_comb, 9'h0b5);
  assign p1_smul_80403_comb = smul20b_11b_x_9b(p1_concat_80171_comb, 9'h0fb);
  assign p1_smul_80404_comb = smul20b_11b_x_9b(p1_concat_80163_comb, 9'h0d5);
  assign p1_smul_80413_comb = smul20b_11b_x_9b(p1_concat_80164_comb, 9'h12b);
  assign p1_smul_80414_comb = smul20b_11b_x_9b(p1_concat_80172_comb, 9'h105);
  assign p1_smul_80415_comb = smul20b_11b_x_9b(p1_concat_80173_comb, 9'h0fb);
  assign p1_smul_80416_comb = smul20b_11b_x_9b(p1_concat_80165_comb, 9'h0d5);
  assign p1_smul_80425_comb = smul20b_11b_x_9b(p1_concat_80166_comb, 9'h12b);
  assign p1_smul_80426_comb = smul20b_11b_x_9b(p1_concat_80174_comb, 9'h105);
  assign p1_smul_80427_comb = smul20b_11b_x_9b(p1_concat_80175_comb, 9'h0fb);
  assign p1_smul_80428_comb = smul20b_11b_x_9b(p1_concat_80167_comb, 9'h0d5);
  assign p1_smul_80437_comb = smul20b_11b_x_9b(p1_concat_80168_comb, 9'h12b);
  assign p1_smul_80438_comb = smul20b_11b_x_9b(p1_concat_80176_comb, 9'h105);
  assign p1_smul_80439_comb = smul20b_11b_x_9b(p1_concat_80177_comb, 9'h0fb);
  assign p1_smul_80440_comb = smul20b_11b_x_9b(p1_concat_80169_comb, 9'h0d5);
  assign p1_smul_80449_comb = smul20b_11b_x_9b(p1_concat_80170_comb, 9'h12b);
  assign p1_smul_80450_comb = smul20b_11b_x_9b(p1_concat_80178_comb, 9'h105);
  assign p1_smul_80483_comb = smul20b_11b_x_9b(p1_concat_80171_comb, 9'h0d5);
  assign p1_smul_80485_comb = smul20b_11b_x_9b(p1_concat_80147_comb, 9'h105);
  assign p1_smul_80490_comb = smul20b_11b_x_9b(p1_concat_80150_comb, 9'h0fb);
  assign p1_smul_80492_comb = smul20b_11b_x_9b(p1_concat_80172_comb, 9'h12b);
  assign p1_smul_80493_comb = smul20b_11b_x_9b(p1_concat_80173_comb, 9'h0d5);
  assign p1_smul_80495_comb = smul20b_11b_x_9b(p1_concat_80151_comb, 9'h105);
  assign p1_smul_80500_comb = smul20b_11b_x_9b(p1_concat_80154_comb, 9'h0fb);
  assign p1_smul_80502_comb = smul20b_11b_x_9b(p1_concat_80174_comb, 9'h12b);
  assign p1_smul_80503_comb = smul20b_11b_x_9b(p1_concat_80175_comb, 9'h0d5);
  assign p1_smul_80505_comb = smul20b_11b_x_9b(p1_concat_80155_comb, 9'h105);
  assign p1_smul_80510_comb = smul20b_11b_x_9b(p1_concat_80158_comb, 9'h0fb);
  assign p1_smul_80512_comb = smul20b_11b_x_9b(p1_concat_80176_comb, 9'h12b);
  assign p1_smul_80513_comb = smul20b_11b_x_9b(p1_concat_80177_comb, 9'h0d5);
  assign p1_smul_80515_comb = smul20b_11b_x_9b(p1_concat_80159_comb, 9'h105);
  assign p1_smul_80520_comb = smul20b_11b_x_9b(p1_concat_80162_comb, 9'h0fb);
  assign p1_smul_80522_comb = smul20b_11b_x_9b(p1_concat_80178_comb, 9'h12b);
  assign p1_smul_80525_comb = smul20b_11b_x_9b(p1_concat_80163_comb, 9'h105);
  assign p1_smul_80527_comb = smul20b_11b_x_9b(p1_concat_80148_comb, 9'h0d5);
  assign p1_smul_80528_comb = smul20b_11b_x_9b(p1_concat_80149_comb, 9'h0d5);
  assign p1_smul_80530_comb = smul20b_11b_x_9b(p1_concat_80164_comb, 9'h105);
  assign p1_smul_80535_comb = smul20b_11b_x_9b(p1_concat_80165_comb, 9'h105);
  assign p1_smul_80537_comb = smul20b_11b_x_9b(p1_concat_80152_comb, 9'h0d5);
  assign p1_smul_80538_comb = smul20b_11b_x_9b(p1_concat_80153_comb, 9'h0d5);
  assign p1_smul_80540_comb = smul20b_11b_x_9b(p1_concat_80166_comb, 9'h105);
  assign p1_smul_80545_comb = smul20b_11b_x_9b(p1_concat_80167_comb, 9'h105);
  assign p1_smul_80547_comb = smul20b_11b_x_9b(p1_concat_80156_comb, 9'h0d5);
  assign p1_smul_80548_comb = smul20b_11b_x_9b(p1_concat_80157_comb, 9'h0d5);
  assign p1_smul_80550_comb = smul20b_11b_x_9b(p1_concat_80168_comb, 9'h105);
  assign p1_smul_80555_comb = smul20b_11b_x_9b(p1_concat_80169_comb, 9'h105);
  assign p1_smul_80557_comb = smul20b_11b_x_9b(p1_concat_80160_comb, 9'h0d5);
  assign p1_smul_80558_comb = smul20b_11b_x_9b(p1_concat_80161_comb, 9'h0d5);
  assign p1_smul_80560_comb = smul20b_11b_x_9b(p1_concat_80170_comb, 9'h105);
  assign p1_smul_80583_comb = smul20b_11b_x_9b(p1_concat_80147_comb, 9'h0d5);
  assign p1_smul_80584_comb = smul20b_11b_x_9b(p1_concat_80148_comb, 9'h105);
  assign p1_smul_80585_comb = smul20b_11b_x_9b(p1_concat_80149_comb, 9'h105);
  assign p1_smul_80586_comb = smul20b_11b_x_9b(p1_concat_80150_comb, 9'h0d5);
  assign p1_smul_80595_comb = smul20b_11b_x_9b(p1_concat_80151_comb, 9'h0d5);
  assign p1_smul_80596_comb = smul20b_11b_x_9b(p1_concat_80152_comb, 9'h105);
  assign p1_smul_80597_comb = smul20b_11b_x_9b(p1_concat_80153_comb, 9'h105);
  assign p1_smul_80598_comb = smul20b_11b_x_9b(p1_concat_80154_comb, 9'h0d5);
  assign p1_smul_80607_comb = smul20b_11b_x_9b(p1_concat_80155_comb, 9'h0d5);
  assign p1_smul_80608_comb = smul20b_11b_x_9b(p1_concat_80156_comb, 9'h105);
  assign p1_smul_80609_comb = smul20b_11b_x_9b(p1_concat_80157_comb, 9'h105);
  assign p1_smul_80610_comb = smul20b_11b_x_9b(p1_concat_80158_comb, 9'h0d5);
  assign p1_smul_80619_comb = smul20b_11b_x_9b(p1_concat_80159_comb, 9'h0d5);
  assign p1_smul_80620_comb = smul20b_11b_x_9b(p1_concat_80160_comb, 9'h105);
  assign p1_smul_80621_comb = smul20b_11b_x_9b(p1_concat_80161_comb, 9'h105);
  assign p1_smul_80622_comb = smul20b_11b_x_9b(p1_concat_80162_comb, 9'h0d5);
  assign p1_smul_80627_comb = smul20b_11b_x_9b(p1_concat_80191_comb, 9'h0fb);
  assign p1_smul_80628_comb = smul20b_11b_x_9b(p1_concat_80187_comb, 9'h0d5);
  assign p1_smul_80637_comb = smul20b_11b_x_9b(p1_concat_80188_comb, 9'h12b);
  assign p1_smul_80638_comb = smul20b_11b_x_9b(p1_concat_80192_comb, 9'h105);
  assign p1_smul_80639_comb = smul20b_11b_x_9b(p1_concat_80193_comb, 9'h0fb);
  assign p1_smul_80640_comb = smul20b_11b_x_9b(p1_concat_80189_comb, 9'h0d5);
  assign p1_smul_80649_comb = smul20b_11b_x_9b(p1_concat_80190_comb, 9'h12b);
  assign p1_smul_80650_comb = smul20b_11b_x_9b(p1_concat_80194_comb, 9'h105);
  assign p1_smul_80667_comb = smul20b_11b_x_9b(p1_concat_80191_comb, 9'h0d5);
  assign p1_smul_80669_comb = smul20b_11b_x_9b(p1_concat_80179_comb, 9'h105);
  assign p1_smul_80674_comb = smul20b_11b_x_9b(p1_concat_80182_comb, 9'h0fb);
  assign p1_smul_80676_comb = smul20b_11b_x_9b(p1_concat_80192_comb, 9'h12b);
  assign p1_smul_80677_comb = smul20b_11b_x_9b(p1_concat_80193_comb, 9'h0d5);
  assign p1_smul_80679_comb = smul20b_11b_x_9b(p1_concat_80183_comb, 9'h105);
  assign p1_smul_80684_comb = smul20b_11b_x_9b(p1_concat_80186_comb, 9'h0fb);
  assign p1_smul_80686_comb = smul20b_11b_x_9b(p1_concat_80194_comb, 9'h12b);
  assign p1_smul_80689_comb = smul20b_11b_x_9b(p1_concat_80187_comb, 9'h105);
  assign p1_smul_80691_comb = smul20b_11b_x_9b(p1_concat_80180_comb, 9'h0d5);
  assign p1_smul_80692_comb = smul20b_11b_x_9b(p1_concat_80181_comb, 9'h0d5);
  assign p1_smul_80694_comb = smul20b_11b_x_9b(p1_concat_80188_comb, 9'h105);
  assign p1_smul_80699_comb = smul20b_11b_x_9b(p1_concat_80189_comb, 9'h105);
  assign p1_smul_80701_comb = smul20b_11b_x_9b(p1_concat_80184_comb, 9'h0d5);
  assign p1_smul_80702_comb = smul20b_11b_x_9b(p1_concat_80185_comb, 9'h0d5);
  assign p1_smul_80704_comb = smul20b_11b_x_9b(p1_concat_80190_comb, 9'h105);
  assign p1_smul_80719_comb = smul20b_11b_x_9b(p1_concat_80179_comb, 9'h0d5);
  assign p1_smul_80720_comb = smul20b_11b_x_9b(p1_concat_80180_comb, 9'h105);
  assign p1_smul_80721_comb = smul20b_11b_x_9b(p1_concat_80181_comb, 9'h105);
  assign p1_smul_80722_comb = smul20b_11b_x_9b(p1_concat_80182_comb, 9'h0d5);
  assign p1_smul_80731_comb = smul20b_11b_x_9b(p1_concat_80183_comb, 9'h0d5);
  assign p1_smul_80732_comb = smul20b_11b_x_9b(p1_concat_80184_comb, 9'h105);
  assign p1_smul_80733_comb = smul20b_11b_x_9b(p1_concat_80185_comb, 9'h105);
  assign p1_smul_80734_comb = smul20b_11b_x_9b(p1_concat_80186_comb, 9'h0d5);
  assign p1_smul_80739_comb = smul20b_11b_x_9b(p1_concat_80207_comb, 9'h0fb);
  assign p1_smul_80740_comb = smul20b_11b_x_9b(p1_concat_80203_comb, 9'h0d5);
  assign p1_smul_80749_comb = smul20b_11b_x_9b(p1_concat_80204_comb, 9'h12b);
  assign p1_smul_80750_comb = smul20b_11b_x_9b(p1_concat_80208_comb, 9'h105);
  assign p1_smul_80751_comb = smul20b_11b_x_9b(p1_concat_80209_comb, 9'h0fb);
  assign p1_smul_80752_comb = smul20b_11b_x_9b(p1_concat_80205_comb, 9'h0d5);
  assign p1_smul_80761_comb = smul20b_11b_x_9b(p1_concat_80206_comb, 9'h12b);
  assign p1_smul_80762_comb = smul20b_11b_x_9b(p1_concat_80210_comb, 9'h105);
  assign p1_smul_80779_comb = smul20b_11b_x_9b(p1_concat_80207_comb, 9'h0d5);
  assign p1_smul_80781_comb = smul20b_11b_x_9b(p1_concat_80195_comb, 9'h105);
  assign p1_smul_80786_comb = smul20b_11b_x_9b(p1_concat_80198_comb, 9'h0fb);
  assign p1_smul_80788_comb = smul20b_11b_x_9b(p1_concat_80208_comb, 9'h12b);
  assign p1_smul_80789_comb = smul20b_11b_x_9b(p1_concat_80209_comb, 9'h0d5);
  assign p1_smul_80791_comb = smul20b_11b_x_9b(p1_concat_80199_comb, 9'h105);
  assign p1_smul_80796_comb = smul20b_11b_x_9b(p1_concat_80202_comb, 9'h0fb);
  assign p1_smul_80798_comb = smul20b_11b_x_9b(p1_concat_80210_comb, 9'h12b);
  assign p1_smul_80801_comb = smul20b_11b_x_9b(p1_concat_80203_comb, 9'h105);
  assign p1_smul_80803_comb = smul20b_11b_x_9b(p1_concat_80196_comb, 9'h0d5);
  assign p1_smul_80804_comb = smul20b_11b_x_9b(p1_concat_80197_comb, 9'h0d5);
  assign p1_smul_80806_comb = smul20b_11b_x_9b(p1_concat_80204_comb, 9'h105);
  assign p1_smul_80811_comb = smul20b_11b_x_9b(p1_concat_80205_comb, 9'h105);
  assign p1_smul_80813_comb = smul20b_11b_x_9b(p1_concat_80200_comb, 9'h0d5);
  assign p1_smul_80814_comb = smul20b_11b_x_9b(p1_concat_80201_comb, 9'h0d5);
  assign p1_smul_80816_comb = smul20b_11b_x_9b(p1_concat_80206_comb, 9'h105);
  assign p1_smul_80831_comb = smul20b_11b_x_9b(p1_concat_80195_comb, 9'h0d5);
  assign p1_smul_80832_comb = smul20b_11b_x_9b(p1_concat_80196_comb, 9'h105);
  assign p1_smul_80833_comb = smul20b_11b_x_9b(p1_concat_80197_comb, 9'h105);
  assign p1_smul_80834_comb = smul20b_11b_x_9b(p1_concat_80198_comb, 9'h0d5);
  assign p1_smul_80843_comb = smul20b_11b_x_9b(p1_concat_80199_comb, 9'h0d5);
  assign p1_smul_80844_comb = smul20b_11b_x_9b(p1_concat_80200_comb, 9'h105);
  assign p1_smul_80845_comb = smul20b_11b_x_9b(p1_concat_80201_comb, 9'h105);
  assign p1_smul_80846_comb = smul20b_11b_x_9b(p1_concat_80202_comb, 9'h0d5);
  assign p1_add_81795_comb = p1_smul_81379_comb + p1_smul_81380_comb;
  assign p1_add_81796_comb = p1_smul_81381_comb + p1_smul_81382_comb;
  assign p1_add_81797_comb = p1_smul_81383_comb + p1_smul_81384_comb;
  assign p1_add_81798_comb = p1_smul_81385_comb + p1_smul_81386_comb;
  assign p1_add_81799_comb = p1_smul_81387_comb + p1_smul_81388_comb;
  assign p1_add_81800_comb = p1_smul_81389_comb + p1_smul_81390_comb;
  assign p1_add_81801_comb = p1_smul_81391_comb + p1_smul_81392_comb;
  assign p1_add_81802_comb = p1_smul_81393_comb + p1_smul_81394_comb;
  assign p1_add_81803_comb = p1_smul_81395_comb + p1_smul_81396_comb;
  assign p1_add_81804_comb = p1_smul_81397_comb + p1_smul_81398_comb;
  assign p1_add_81805_comb = p1_smul_81399_comb + p1_smul_81400_comb;
  assign p1_add_81806_comb = p1_smul_81401_comb + p1_smul_81402_comb;
  assign p1_add_81807_comb = p1_smul_81403_comb + p1_smul_81404_comb;
  assign p1_add_81808_comb = p1_smul_81405_comb + p1_smul_81406_comb;
  assign p1_add_81809_comb = p1_smul_81407_comb + p1_smul_81408_comb;
  assign p1_add_81810_comb = p1_smul_81409_comb + p1_smul_81410_comb;
  assign p1_add_81915_comb = p1_smul_81547_comb + p1_smul_81548_comb;
  assign p1_add_81916_comb = p1_smul_81549_comb + p1_smul_81550_comb;
  assign p1_add_81917_comb = p1_smul_81551_comb + p1_smul_81552_comb;
  assign p1_add_81918_comb = p1_smul_81553_comb + p1_smul_81554_comb;
  assign p1_add_81919_comb = p1_smul_81555_comb + p1_smul_81556_comb;
  assign p1_add_81920_comb = p1_smul_81557_comb + p1_smul_81558_comb;
  assign p1_add_81921_comb = p1_smul_81559_comb + p1_smul_81560_comb;
  assign p1_add_81922_comb = p1_smul_81561_comb + p1_smul_81562_comb;
  assign p1_add_81995_comb = p1_smul_81659_comb + p1_smul_81660_comb;
  assign p1_add_81996_comb = p1_smul_81661_comb + p1_smul_81662_comb;
  assign p1_add_81997_comb = p1_smul_81663_comb + p1_smul_81664_comb;
  assign p1_add_81998_comb = p1_smul_81665_comb + p1_smul_81666_comb;
  assign p1_add_81999_comb = p1_smul_81667_comb + p1_smul_81668_comb;
  assign p1_add_82000_comb = p1_smul_81669_comb + p1_smul_81670_comb;
  assign p1_add_82001_comb = p1_smul_81671_comb + p1_smul_81672_comb;
  assign p1_add_82002_comb = p1_smul_81673_comb + p1_smul_81674_comb;
  assign p1_add_80851_comb = p1_smul_80403_comb + p1_smul_80404_comb;
  assign p1_smul_80852_comb = smul18b_18b_x_8b(p1_sign_ext_80213_comb[17:0], 8'h47);
  assign p1_smul_80853_comb = smul18b_18b_x_6b(p1_sign_ext_80214_comb[17:0], 6'h19);
  assign p1_smul_80854_comb = smul18b_18b_x_6b(p1_sign_ext_80215_comb[17:0], 6'h27);
  assign p1_smul_80855_comb = smul18b_18b_x_8b(p1_sign_ext_80216_comb[17:0], 8'hb9);
  assign p1_add_80856_comb = p1_smul_80413_comb + p1_smul_80414_comb;
  assign p1_add_80857_comb = p1_smul_80415_comb + p1_smul_80416_comb;
  assign p1_smul_80858_comb = smul18b_18b_x_8b(p1_sign_ext_80221_comb[17:0], 8'h47);
  assign p1_smul_80859_comb = smul18b_18b_x_6b(p1_sign_ext_80222_comb[17:0], 6'h19);
  assign p1_smul_80860_comb = smul18b_18b_x_6b(p1_sign_ext_80223_comb[17:0], 6'h27);
  assign p1_smul_80861_comb = smul18b_18b_x_8b(p1_sign_ext_80224_comb[17:0], 8'hb9);
  assign p1_add_80862_comb = p1_smul_80425_comb + p1_smul_80426_comb;
  assign p1_add_80863_comb = p1_smul_80427_comb + p1_smul_80428_comb;
  assign p1_smul_80864_comb = smul18b_18b_x_8b(p1_sign_ext_80229_comb[17:0], 8'h47);
  assign p1_smul_80865_comb = smul18b_18b_x_6b(p1_sign_ext_80230_comb[17:0], 6'h19);
  assign p1_smul_80866_comb = smul18b_18b_x_6b(p1_sign_ext_80231_comb[17:0], 6'h27);
  assign p1_smul_80867_comb = smul18b_18b_x_8b(p1_sign_ext_80232_comb[17:0], 8'hb9);
  assign p1_add_80868_comb = p1_smul_80437_comb + p1_smul_80438_comb;
  assign p1_add_80869_comb = p1_smul_80439_comb + p1_smul_80440_comb;
  assign p1_smul_80870_comb = smul18b_18b_x_8b(p1_sign_ext_80237_comb[17:0], 8'h47);
  assign p1_smul_80871_comb = smul18b_18b_x_6b(p1_sign_ext_80238_comb[17:0], 6'h19);
  assign p1_smul_80872_comb = smul18b_18b_x_6b(p1_sign_ext_80239_comb[17:0], 6'h27);
  assign p1_smul_80873_comb = smul18b_18b_x_8b(p1_sign_ext_80240_comb[17:0], 8'hb9);
  assign p1_add_80874_comb = p1_smul_80449_comb + p1_smul_80450_comb;
  assign p1_smul_80876_comb = smul19b_19b_x_7b(p1_sign_ext_80243_comb[18:0], 7'h31);
  assign p1_smul_80877_comb = smul19b_19b_x_7b(p1_sign_ext_80213_comb[18:0], 7'h4f);
  assign p1_smul_80880_comb = smul19b_19b_x_7b(p1_sign_ext_80216_comb[18:0], 7'h4f);
  assign p1_smul_80881_comb = smul19b_19b_x_7b(p1_sign_ext_80244_comb[18:0], 7'h31);
  assign p1_smul_80884_comb = smul19b_19b_x_7b(p1_sign_ext_80245_comb[18:0], 7'h31);
  assign p1_smul_80885_comb = smul19b_19b_x_7b(p1_sign_ext_80221_comb[18:0], 7'h4f);
  assign p1_smul_80888_comb = smul19b_19b_x_7b(p1_sign_ext_80224_comb[18:0], 7'h4f);
  assign p1_smul_80889_comb = smul19b_19b_x_7b(p1_sign_ext_80246_comb[18:0], 7'h31);
  assign p1_smul_80892_comb = smul19b_19b_x_7b(p1_sign_ext_80247_comb[18:0], 7'h31);
  assign p1_smul_80893_comb = smul19b_19b_x_7b(p1_sign_ext_80229_comb[18:0], 7'h4f);
  assign p1_smul_80896_comb = smul19b_19b_x_7b(p1_sign_ext_80232_comb[18:0], 7'h4f);
  assign p1_smul_80897_comb = smul19b_19b_x_7b(p1_sign_ext_80248_comb[18:0], 7'h31);
  assign p1_smul_80900_comb = smul19b_19b_x_7b(p1_sign_ext_80249_comb[18:0], 7'h31);
  assign p1_smul_80901_comb = smul19b_19b_x_7b(p1_sign_ext_80237_comb[18:0], 7'h4f);
  assign p1_smul_80904_comb = smul19b_19b_x_7b(p1_sign_ext_80240_comb[18:0], 7'h4f);
  assign p1_smul_80905_comb = smul19b_19b_x_7b(p1_sign_ext_80250_comb[18:0], 7'h31);
  assign p1_smul_80908_comb = smul19b_19b_x_6b(p1_sign_ext_80243_comb[18:0], 6'h27);
  assign p1_smul_80910_comb = smul19b_19b_x_8b(p1_sign_ext_80214_comb[18:0], 8'hb9);
  assign p1_smul_80911_comb = smul19b_19b_x_8b(p1_sign_ext_80215_comb[18:0], 8'h47);
  assign p1_smul_80913_comb = smul19b_19b_x_6b(p1_sign_ext_80244_comb[18:0], 6'h19);
  assign p1_smul_80916_comb = smul19b_19b_x_6b(p1_sign_ext_80245_comb[18:0], 6'h27);
  assign p1_smul_80918_comb = smul19b_19b_x_8b(p1_sign_ext_80222_comb[18:0], 8'hb9);
  assign p1_smul_80919_comb = smul19b_19b_x_8b(p1_sign_ext_80223_comb[18:0], 8'h47);
  assign p1_smul_80921_comb = smul19b_19b_x_6b(p1_sign_ext_80246_comb[18:0], 6'h19);
  assign p1_smul_80924_comb = smul19b_19b_x_6b(p1_sign_ext_80247_comb[18:0], 6'h27);
  assign p1_smul_80926_comb = smul19b_19b_x_8b(p1_sign_ext_80230_comb[18:0], 8'hb9);
  assign p1_smul_80927_comb = smul19b_19b_x_8b(p1_sign_ext_80231_comb[18:0], 8'h47);
  assign p1_smul_80929_comb = smul19b_19b_x_6b(p1_sign_ext_80248_comb[18:0], 6'h19);
  assign p1_smul_80932_comb = smul19b_19b_x_6b(p1_sign_ext_80249_comb[18:0], 6'h27);
  assign p1_smul_80934_comb = smul19b_19b_x_8b(p1_sign_ext_80238_comb[18:0], 8'hb9);
  assign p1_smul_80935_comb = smul19b_19b_x_8b(p1_sign_ext_80239_comb[18:0], 8'h47);
  assign p1_smul_80937_comb = smul19b_19b_x_6b(p1_sign_ext_80250_comb[18:0], 6'h19);
  assign p1_smul_80971_comb = smul19b_19b_x_8b(p1_sign_ext_80267_comb[18:0], 8'h47);
  assign p1_smul_80973_comb = smul19b_19b_x_6b(p1_sign_ext_80213_comb[18:0], 6'h27);
  assign p1_smul_80976_comb = smul19b_19b_x_6b(p1_sign_ext_80216_comb[18:0], 6'h27);
  assign p1_smul_80978_comb = smul19b_19b_x_8b(p1_sign_ext_80272_comb[18:0], 8'h47);
  assign p1_smul_80979_comb = smul19b_19b_x_8b(p1_sign_ext_80273_comb[18:0], 8'h47);
  assign p1_smul_80981_comb = smul19b_19b_x_6b(p1_sign_ext_80221_comb[18:0], 6'h27);
  assign p1_smul_80984_comb = smul19b_19b_x_6b(p1_sign_ext_80224_comb[18:0], 6'h27);
  assign p1_smul_80986_comb = smul19b_19b_x_8b(p1_sign_ext_80278_comb[18:0], 8'h47);
  assign p1_smul_80987_comb = smul19b_19b_x_8b(p1_sign_ext_80279_comb[18:0], 8'h47);
  assign p1_smul_80989_comb = smul19b_19b_x_6b(p1_sign_ext_80229_comb[18:0], 6'h27);
  assign p1_smul_80992_comb = smul19b_19b_x_6b(p1_sign_ext_80232_comb[18:0], 6'h27);
  assign p1_smul_80994_comb = smul19b_19b_x_8b(p1_sign_ext_80284_comb[18:0], 8'h47);
  assign p1_smul_80995_comb = smul19b_19b_x_8b(p1_sign_ext_80285_comb[18:0], 8'h47);
  assign p1_smul_80997_comb = smul19b_19b_x_6b(p1_sign_ext_80237_comb[18:0], 6'h27);
  assign p1_smul_81000_comb = smul19b_19b_x_6b(p1_sign_ext_80240_comb[18:0], 6'h27);
  assign p1_smul_81002_comb = smul19b_19b_x_8b(p1_sign_ext_80290_comb[18:0], 8'h47);
  assign p1_smul_81003_comb = smul19b_19b_x_7b(p1_sign_ext_80267_comb[18:0], 7'h31);
  assign p1_smul_81005_comb = smul19b_19b_x_7b(p1_sign_ext_80213_comb[18:0], 7'h31);
  assign p1_smul_81008_comb = smul19b_19b_x_7b(p1_sign_ext_80216_comb[18:0], 7'h31);
  assign p1_smul_81010_comb = smul19b_19b_x_7b(p1_sign_ext_80272_comb[18:0], 7'h31);
  assign p1_smul_81011_comb = smul19b_19b_x_7b(p1_sign_ext_80273_comb[18:0], 7'h31);
  assign p1_smul_81013_comb = smul19b_19b_x_7b(p1_sign_ext_80221_comb[18:0], 7'h31);
  assign p1_smul_81016_comb = smul19b_19b_x_7b(p1_sign_ext_80224_comb[18:0], 7'h31);
  assign p1_smul_81018_comb = smul19b_19b_x_7b(p1_sign_ext_80278_comb[18:0], 7'h31);
  assign p1_smul_81019_comb = smul19b_19b_x_7b(p1_sign_ext_80279_comb[18:0], 7'h31);
  assign p1_smul_81021_comb = smul19b_19b_x_7b(p1_sign_ext_80229_comb[18:0], 7'h31);
  assign p1_smul_81024_comb = smul19b_19b_x_7b(p1_sign_ext_80232_comb[18:0], 7'h31);
  assign p1_smul_81026_comb = smul19b_19b_x_7b(p1_sign_ext_80284_comb[18:0], 7'h31);
  assign p1_smul_81027_comb = smul19b_19b_x_7b(p1_sign_ext_80285_comb[18:0], 7'h31);
  assign p1_smul_81029_comb = smul19b_19b_x_7b(p1_sign_ext_80237_comb[18:0], 7'h31);
  assign p1_smul_81032_comb = smul19b_19b_x_7b(p1_sign_ext_80240_comb[18:0], 7'h31);
  assign p1_smul_81034_comb = smul19b_19b_x_7b(p1_sign_ext_80290_comb[18:0], 7'h31);
  assign p1_smul_81035_comb = smul18b_18b_x_6b(p1_sign_ext_80267_comb[17:0], 6'h19);
  assign p1_smul_81036_comb = smul18b_18b_x_8b(p1_sign_ext_80243_comb[17:0], 8'hb9);
  assign p1_add_81037_comb = p1_smul_80583_comb + p1_smul_80584_comb;
  assign p1_add_81038_comb = p1_smul_80585_comb + p1_smul_80586_comb;
  assign p1_smul_81039_comb = smul18b_18b_x_8b(p1_sign_ext_80244_comb[17:0], 8'hb9);
  assign p1_smul_81040_comb = smul18b_18b_x_6b(p1_sign_ext_80272_comb[17:0], 6'h19);
  assign p1_smul_81041_comb = smul18b_18b_x_6b(p1_sign_ext_80273_comb[17:0], 6'h19);
  assign p1_smul_81042_comb = smul18b_18b_x_8b(p1_sign_ext_80245_comb[17:0], 8'hb9);
  assign p1_add_81043_comb = p1_smul_80595_comb + p1_smul_80596_comb;
  assign p1_add_81044_comb = p1_smul_80597_comb + p1_smul_80598_comb;
  assign p1_smul_81045_comb = smul18b_18b_x_8b(p1_sign_ext_80246_comb[17:0], 8'hb9);
  assign p1_smul_81046_comb = smul18b_18b_x_6b(p1_sign_ext_80278_comb[17:0], 6'h19);
  assign p1_smul_81047_comb = smul18b_18b_x_6b(p1_sign_ext_80279_comb[17:0], 6'h19);
  assign p1_smul_81048_comb = smul18b_18b_x_8b(p1_sign_ext_80247_comb[17:0], 8'hb9);
  assign p1_add_81049_comb = p1_smul_80607_comb + p1_smul_80608_comb;
  assign p1_add_81050_comb = p1_smul_80609_comb + p1_smul_80610_comb;
  assign p1_smul_81051_comb = smul18b_18b_x_8b(p1_sign_ext_80248_comb[17:0], 8'hb9);
  assign p1_smul_81052_comb = smul18b_18b_x_6b(p1_sign_ext_80284_comb[17:0], 6'h19);
  assign p1_smul_81053_comb = smul18b_18b_x_6b(p1_sign_ext_80285_comb[17:0], 6'h19);
  assign p1_smul_81054_comb = smul18b_18b_x_8b(p1_sign_ext_80249_comb[17:0], 8'hb9);
  assign p1_add_81055_comb = p1_smul_80619_comb + p1_smul_80620_comb;
  assign p1_add_81056_comb = p1_smul_80621_comb + p1_smul_80622_comb;
  assign p1_smul_81057_comb = smul18b_18b_x_8b(p1_sign_ext_80250_comb[17:0], 8'hb9);
  assign p1_smul_81058_comb = smul18b_18b_x_6b(p1_sign_ext_80290_comb[17:0], 6'h19);
  assign p1_add_81059_comb = p1_smul_80627_comb + p1_smul_80628_comb;
  assign p1_smul_81060_comb = smul18b_18b_x_8b(p1_sign_ext_80309_comb[17:0], 8'h47);
  assign p1_smul_81061_comb = smul18b_18b_x_6b(p1_sign_ext_80310_comb[17:0], 6'h19);
  assign p1_smul_81062_comb = smul18b_18b_x_6b(p1_sign_ext_80311_comb[17:0], 6'h27);
  assign p1_smul_81063_comb = smul18b_18b_x_8b(p1_sign_ext_80312_comb[17:0], 8'hb9);
  assign p1_add_81064_comb = p1_smul_80637_comb + p1_smul_80638_comb;
  assign p1_add_81065_comb = p1_smul_80639_comb + p1_smul_80640_comb;
  assign p1_smul_81066_comb = smul18b_18b_x_8b(p1_sign_ext_80317_comb[17:0], 8'h47);
  assign p1_smul_81067_comb = smul18b_18b_x_6b(p1_sign_ext_80318_comb[17:0], 6'h19);
  assign p1_smul_81068_comb = smul18b_18b_x_6b(p1_sign_ext_80319_comb[17:0], 6'h27);
  assign p1_smul_81069_comb = smul18b_18b_x_8b(p1_sign_ext_80320_comb[17:0], 8'hb9);
  assign p1_add_81070_comb = p1_smul_80649_comb + p1_smul_80650_comb;
  assign p1_smul_81072_comb = smul19b_19b_x_7b(p1_sign_ext_80323_comb[18:0], 7'h31);
  assign p1_smul_81073_comb = smul19b_19b_x_7b(p1_sign_ext_80309_comb[18:0], 7'h4f);
  assign p1_smul_81076_comb = smul19b_19b_x_7b(p1_sign_ext_80312_comb[18:0], 7'h4f);
  assign p1_smul_81077_comb = smul19b_19b_x_7b(p1_sign_ext_80324_comb[18:0], 7'h31);
  assign p1_smul_81080_comb = smul19b_19b_x_7b(p1_sign_ext_80325_comb[18:0], 7'h31);
  assign p1_smul_81081_comb = smul19b_19b_x_7b(p1_sign_ext_80317_comb[18:0], 7'h4f);
  assign p1_smul_81084_comb = smul19b_19b_x_7b(p1_sign_ext_80320_comb[18:0], 7'h4f);
  assign p1_smul_81085_comb = smul19b_19b_x_7b(p1_sign_ext_80326_comb[18:0], 7'h31);
  assign p1_smul_81088_comb = smul19b_19b_x_6b(p1_sign_ext_80323_comb[18:0], 6'h27);
  assign p1_smul_81090_comb = smul19b_19b_x_8b(p1_sign_ext_80310_comb[18:0], 8'hb9);
  assign p1_smul_81091_comb = smul19b_19b_x_8b(p1_sign_ext_80311_comb[18:0], 8'h47);
  assign p1_smul_81093_comb = smul19b_19b_x_6b(p1_sign_ext_80324_comb[18:0], 6'h19);
  assign p1_smul_81096_comb = smul19b_19b_x_6b(p1_sign_ext_80325_comb[18:0], 6'h27);
  assign p1_smul_81098_comb = smul19b_19b_x_8b(p1_sign_ext_80318_comb[18:0], 8'hb9);
  assign p1_smul_81099_comb = smul19b_19b_x_8b(p1_sign_ext_80319_comb[18:0], 8'h47);
  assign p1_smul_81101_comb = smul19b_19b_x_6b(p1_sign_ext_80326_comb[18:0], 6'h19);
  assign p1_smul_81119_comb = smul19b_19b_x_8b(p1_sign_ext_80335_comb[18:0], 8'h47);
  assign p1_smul_81121_comb = smul19b_19b_x_6b(p1_sign_ext_80309_comb[18:0], 6'h27);
  assign p1_smul_81124_comb = smul19b_19b_x_6b(p1_sign_ext_80312_comb[18:0], 6'h27);
  assign p1_smul_81126_comb = smul19b_19b_x_8b(p1_sign_ext_80340_comb[18:0], 8'h47);
  assign p1_smul_81127_comb = smul19b_19b_x_8b(p1_sign_ext_80341_comb[18:0], 8'h47);
  assign p1_smul_81129_comb = smul19b_19b_x_6b(p1_sign_ext_80317_comb[18:0], 6'h27);
  assign p1_smul_81132_comb = smul19b_19b_x_6b(p1_sign_ext_80320_comb[18:0], 6'h27);
  assign p1_smul_81134_comb = smul19b_19b_x_8b(p1_sign_ext_80346_comb[18:0], 8'h47);
  assign p1_smul_81135_comb = smul19b_19b_x_7b(p1_sign_ext_80335_comb[18:0], 7'h31);
  assign p1_smul_81137_comb = smul19b_19b_x_7b(p1_sign_ext_80309_comb[18:0], 7'h31);
  assign p1_smul_81140_comb = smul19b_19b_x_7b(p1_sign_ext_80312_comb[18:0], 7'h31);
  assign p1_smul_81142_comb = smul19b_19b_x_7b(p1_sign_ext_80340_comb[18:0], 7'h31);
  assign p1_smul_81143_comb = smul19b_19b_x_7b(p1_sign_ext_80341_comb[18:0], 7'h31);
  assign p1_smul_81145_comb = smul19b_19b_x_7b(p1_sign_ext_80317_comb[18:0], 7'h31);
  assign p1_smul_81148_comb = smul19b_19b_x_7b(p1_sign_ext_80320_comb[18:0], 7'h31);
  assign p1_smul_81150_comb = smul19b_19b_x_7b(p1_sign_ext_80346_comb[18:0], 7'h31);
  assign p1_smul_81151_comb = smul18b_18b_x_6b(p1_sign_ext_80335_comb[17:0], 6'h19);
  assign p1_smul_81152_comb = smul18b_18b_x_8b(p1_sign_ext_80323_comb[17:0], 8'hb9);
  assign p1_add_81153_comb = p1_smul_80719_comb + p1_smul_80720_comb;
  assign p1_add_81154_comb = p1_smul_80721_comb + p1_smul_80722_comb;
  assign p1_smul_81155_comb = smul18b_18b_x_8b(p1_sign_ext_80324_comb[17:0], 8'hb9);
  assign p1_smul_81156_comb = smul18b_18b_x_6b(p1_sign_ext_80340_comb[17:0], 6'h19);
  assign p1_smul_81157_comb = smul18b_18b_x_6b(p1_sign_ext_80341_comb[17:0], 6'h19);
  assign p1_smul_81158_comb = smul18b_18b_x_8b(p1_sign_ext_80325_comb[17:0], 8'hb9);
  assign p1_add_81159_comb = p1_smul_80731_comb + p1_smul_80732_comb;
  assign p1_add_81160_comb = p1_smul_80733_comb + p1_smul_80734_comb;
  assign p1_smul_81161_comb = smul18b_18b_x_8b(p1_sign_ext_80326_comb[17:0], 8'hb9);
  assign p1_smul_81162_comb = smul18b_18b_x_6b(p1_sign_ext_80346_comb[17:0], 6'h19);
  assign p1_add_81163_comb = p1_smul_80739_comb + p1_smul_80740_comb;
  assign p1_smul_81164_comb = smul18b_18b_x_8b(p1_sign_ext_80357_comb[17:0], 8'h47);
  assign p1_smul_81165_comb = smul18b_18b_x_6b(p1_sign_ext_80358_comb[17:0], 6'h19);
  assign p1_smul_81166_comb = smul18b_18b_x_6b(p1_sign_ext_80359_comb[17:0], 6'h27);
  assign p1_smul_81167_comb = smul18b_18b_x_8b(p1_sign_ext_80360_comb[17:0], 8'hb9);
  assign p1_add_81168_comb = p1_smul_80749_comb + p1_smul_80750_comb;
  assign p1_add_81169_comb = p1_smul_80751_comb + p1_smul_80752_comb;
  assign p1_smul_81170_comb = smul18b_18b_x_8b(p1_sign_ext_80365_comb[17:0], 8'h47);
  assign p1_smul_81171_comb = smul18b_18b_x_6b(p1_sign_ext_80366_comb[17:0], 6'h19);
  assign p1_smul_81172_comb = smul18b_18b_x_6b(p1_sign_ext_80367_comb[17:0], 6'h27);
  assign p1_smul_81173_comb = smul18b_18b_x_8b(p1_sign_ext_80368_comb[17:0], 8'hb9);
  assign p1_add_81174_comb = p1_smul_80761_comb + p1_smul_80762_comb;
  assign p1_smul_81176_comb = smul19b_19b_x_7b(p1_sign_ext_80371_comb[18:0], 7'h31);
  assign p1_smul_81177_comb = smul19b_19b_x_7b(p1_sign_ext_80357_comb[18:0], 7'h4f);
  assign p1_smul_81180_comb = smul19b_19b_x_7b(p1_sign_ext_80360_comb[18:0], 7'h4f);
  assign p1_smul_81181_comb = smul19b_19b_x_7b(p1_sign_ext_80372_comb[18:0], 7'h31);
  assign p1_smul_81184_comb = smul19b_19b_x_7b(p1_sign_ext_80373_comb[18:0], 7'h31);
  assign p1_smul_81185_comb = smul19b_19b_x_7b(p1_sign_ext_80365_comb[18:0], 7'h4f);
  assign p1_smul_81188_comb = smul19b_19b_x_7b(p1_sign_ext_80368_comb[18:0], 7'h4f);
  assign p1_smul_81189_comb = smul19b_19b_x_7b(p1_sign_ext_80374_comb[18:0], 7'h31);
  assign p1_smul_81192_comb = smul19b_19b_x_6b(p1_sign_ext_80371_comb[18:0], 6'h27);
  assign p1_smul_81194_comb = smul19b_19b_x_8b(p1_sign_ext_80358_comb[18:0], 8'hb9);
  assign p1_smul_81195_comb = smul19b_19b_x_8b(p1_sign_ext_80359_comb[18:0], 8'h47);
  assign p1_smul_81197_comb = smul19b_19b_x_6b(p1_sign_ext_80372_comb[18:0], 6'h19);
  assign p1_smul_81200_comb = smul19b_19b_x_6b(p1_sign_ext_80373_comb[18:0], 6'h27);
  assign p1_smul_81202_comb = smul19b_19b_x_8b(p1_sign_ext_80366_comb[18:0], 8'hb9);
  assign p1_smul_81203_comb = smul19b_19b_x_8b(p1_sign_ext_80367_comb[18:0], 8'h47);
  assign p1_smul_81205_comb = smul19b_19b_x_6b(p1_sign_ext_80374_comb[18:0], 6'h19);
  assign p1_smul_81223_comb = smul19b_19b_x_8b(p1_sign_ext_80383_comb[18:0], 8'h47);
  assign p1_smul_81225_comb = smul19b_19b_x_6b(p1_sign_ext_80357_comb[18:0], 6'h27);
  assign p1_smul_81228_comb = smul19b_19b_x_6b(p1_sign_ext_80360_comb[18:0], 6'h27);
  assign p1_smul_81230_comb = smul19b_19b_x_8b(p1_sign_ext_80388_comb[18:0], 8'h47);
  assign p1_smul_81231_comb = smul19b_19b_x_8b(p1_sign_ext_80389_comb[18:0], 8'h47);
  assign p1_smul_81233_comb = smul19b_19b_x_6b(p1_sign_ext_80365_comb[18:0], 6'h27);
  assign p1_smul_81236_comb = smul19b_19b_x_6b(p1_sign_ext_80368_comb[18:0], 6'h27);
  assign p1_smul_81238_comb = smul19b_19b_x_8b(p1_sign_ext_80394_comb[18:0], 8'h47);
  assign p1_smul_81239_comb = smul19b_19b_x_7b(p1_sign_ext_80383_comb[18:0], 7'h31);
  assign p1_smul_81241_comb = smul19b_19b_x_7b(p1_sign_ext_80357_comb[18:0], 7'h31);
  assign p1_smul_81244_comb = smul19b_19b_x_7b(p1_sign_ext_80360_comb[18:0], 7'h31);
  assign p1_smul_81246_comb = smul19b_19b_x_7b(p1_sign_ext_80388_comb[18:0], 7'h31);
  assign p1_smul_81247_comb = smul19b_19b_x_7b(p1_sign_ext_80389_comb[18:0], 7'h31);
  assign p1_smul_81249_comb = smul19b_19b_x_7b(p1_sign_ext_80365_comb[18:0], 7'h31);
  assign p1_smul_81252_comb = smul19b_19b_x_7b(p1_sign_ext_80368_comb[18:0], 7'h31);
  assign p1_smul_81254_comb = smul19b_19b_x_7b(p1_sign_ext_80394_comb[18:0], 7'h31);
  assign p1_smul_81255_comb = smul18b_18b_x_6b(p1_sign_ext_80383_comb[17:0], 6'h19);
  assign p1_smul_81256_comb = smul18b_18b_x_8b(p1_sign_ext_80371_comb[17:0], 8'hb9);
  assign p1_add_81257_comb = p1_smul_80831_comb + p1_smul_80832_comb;
  assign p1_add_81258_comb = p1_smul_80833_comb + p1_smul_80834_comb;
  assign p1_smul_81259_comb = smul18b_18b_x_8b(p1_sign_ext_80372_comb[17:0], 8'hb9);
  assign p1_smul_81260_comb = smul18b_18b_x_6b(p1_sign_ext_80388_comb[17:0], 6'h19);
  assign p1_smul_81261_comb = smul18b_18b_x_6b(p1_sign_ext_80389_comb[17:0], 6'h19);
  assign p1_smul_81262_comb = smul18b_18b_x_8b(p1_sign_ext_80373_comb[17:0], 8'hb9);
  assign p1_add_81263_comb = p1_smul_80843_comb + p1_smul_80844_comb;
  assign p1_add_81264_comb = p1_smul_80845_comb + p1_smul_80846_comb;
  assign p1_smul_81265_comb = smul18b_18b_x_8b(p1_sign_ext_80374_comb[17:0], 8'hb9);
  assign p1_smul_81266_comb = smul18b_18b_x_6b(p1_sign_ext_80394_comb[17:0], 6'h19);
  assign p1_add_81715_comb = p1_sign_ext_80267_comb[11:0] + p1_sign_ext_80243_comb[11:0];
  assign p1_add_81716_comb = p1_sign_ext_80213_comb[11:0] + p1_sign_ext_80214_comb[11:0];
  assign p1_add_81717_comb = p1_sign_ext_80215_comb[11:0] + p1_sign_ext_80216_comb[11:0];
  assign p1_add_81718_comb = p1_sign_ext_80244_comb[11:0] + p1_sign_ext_80272_comb[11:0];
  assign p1_add_81719_comb = p1_sign_ext_80273_comb[11:0] + p1_sign_ext_80245_comb[11:0];
  assign p1_add_81720_comb = p1_sign_ext_80221_comb[11:0] + p1_sign_ext_80222_comb[11:0];
  assign p1_add_81721_comb = p1_sign_ext_80223_comb[11:0] + p1_sign_ext_80224_comb[11:0];
  assign p1_add_81722_comb = p1_sign_ext_80246_comb[11:0] + p1_sign_ext_80278_comb[11:0];
  assign p1_add_81723_comb = p1_sign_ext_80279_comb[11:0] + p1_sign_ext_80247_comb[11:0];
  assign p1_add_81724_comb = p1_sign_ext_80229_comb[11:0] + p1_sign_ext_80230_comb[11:0];
  assign p1_add_81725_comb = p1_sign_ext_80231_comb[11:0] + p1_sign_ext_80232_comb[11:0];
  assign p1_add_81726_comb = p1_sign_ext_80248_comb[11:0] + p1_sign_ext_80284_comb[11:0];
  assign p1_add_81727_comb = p1_sign_ext_80285_comb[11:0] + p1_sign_ext_80249_comb[11:0];
  assign p1_add_81728_comb = p1_sign_ext_80237_comb[11:0] + p1_sign_ext_80238_comb[11:0];
  assign p1_add_81729_comb = p1_sign_ext_80239_comb[11:0] + p1_sign_ext_80240_comb[11:0];
  assign p1_add_81730_comb = p1_sign_ext_80250_comb[11:0] + p1_sign_ext_80290_comb[11:0];
  assign p1_add_81875_comb = p1_sign_ext_80335_comb[11:0] + p1_sign_ext_80323_comb[11:0];
  assign p1_add_81876_comb = p1_sign_ext_80309_comb[11:0] + p1_sign_ext_80310_comb[11:0];
  assign p1_add_81877_comb = p1_sign_ext_80311_comb[11:0] + p1_sign_ext_80312_comb[11:0];
  assign p1_add_81878_comb = p1_sign_ext_80324_comb[11:0] + p1_sign_ext_80340_comb[11:0];
  assign p1_add_81879_comb = p1_sign_ext_80341_comb[11:0] + p1_sign_ext_80325_comb[11:0];
  assign p1_add_81880_comb = p1_sign_ext_80317_comb[11:0] + p1_sign_ext_80318_comb[11:0];
  assign p1_add_81881_comb = p1_sign_ext_80319_comb[11:0] + p1_sign_ext_80320_comb[11:0];
  assign p1_add_81882_comb = p1_sign_ext_80326_comb[11:0] + p1_sign_ext_80346_comb[11:0];
  assign p1_add_81955_comb = p1_sign_ext_80383_comb[11:0] + p1_sign_ext_80371_comb[11:0];
  assign p1_add_81956_comb = p1_sign_ext_80357_comb[11:0] + p1_sign_ext_80358_comb[11:0];
  assign p1_add_81957_comb = p1_sign_ext_80359_comb[11:0] + p1_sign_ext_80360_comb[11:0];
  assign p1_add_81958_comb = p1_sign_ext_80372_comb[11:0] + p1_sign_ext_80388_comb[11:0];
  assign p1_add_81959_comb = p1_sign_ext_80389_comb[11:0] + p1_sign_ext_80373_comb[11:0];
  assign p1_add_81960_comb = p1_sign_ext_80365_comb[11:0] + p1_sign_ext_80366_comb[11:0];
  assign p1_add_81961_comb = p1_sign_ext_80367_comb[11:0] + p1_sign_ext_80368_comb[11:0];
  assign p1_add_81962_comb = p1_sign_ext_80374_comb[11:0] + p1_sign_ext_80394_comb[11:0];
  assign p1_sum__1736_comb = {{6{p1_add_81795_comb[18]}}, p1_add_81795_comb};
  assign p1_sum__1737_comb = {{6{p1_add_81796_comb[18]}}, p1_add_81796_comb};
  assign p1_sum__1738_comb = {{6{p1_add_81797_comb[18]}}, p1_add_81797_comb};
  assign p1_sum__1739_comb = {{6{p1_add_81798_comb[18]}}, p1_add_81798_comb};
  assign p1_sum__1708_comb = {{6{p1_add_81799_comb[18]}}, p1_add_81799_comb};
  assign p1_sum__1709_comb = {{6{p1_add_81800_comb[18]}}, p1_add_81800_comb};
  assign p1_sum__1710_comb = {{6{p1_add_81801_comb[18]}}, p1_add_81801_comb};
  assign p1_sum__1711_comb = {{6{p1_add_81802_comb[18]}}, p1_add_81802_comb};
  assign p1_sum__1680_comb = {{6{p1_add_81803_comb[18]}}, p1_add_81803_comb};
  assign p1_sum__1681_comb = {{6{p1_add_81804_comb[18]}}, p1_add_81804_comb};
  assign p1_sum__1682_comb = {{6{p1_add_81805_comb[18]}}, p1_add_81805_comb};
  assign p1_sum__1683_comb = {{6{p1_add_81806_comb[18]}}, p1_add_81806_comb};
  assign p1_sum__1652_comb = {{6{p1_add_81807_comb[18]}}, p1_add_81807_comb};
  assign p1_sum__1653_comb = {{6{p1_add_81808_comb[18]}}, p1_add_81808_comb};
  assign p1_sum__1654_comb = {{6{p1_add_81809_comb[18]}}, p1_add_81809_comb};
  assign p1_sum__1655_comb = {{6{p1_add_81810_comb[18]}}, p1_add_81810_comb};
  assign p1_sum__1760_comb = {{6{p1_add_81915_comb[18]}}, p1_add_81915_comb};
  assign p1_sum__1761_comb = {{6{p1_add_81916_comb[18]}}, p1_add_81916_comb};
  assign p1_sum__1762_comb = {{6{p1_add_81917_comb[18]}}, p1_add_81917_comb};
  assign p1_sum__1763_comb = {{6{p1_add_81918_comb[18]}}, p1_add_81918_comb};
  assign p1_sum__1628_comb = {{6{p1_add_81919_comb[18]}}, p1_add_81919_comb};
  assign p1_sum__1629_comb = {{6{p1_add_81920_comb[18]}}, p1_add_81920_comb};
  assign p1_sum__1630_comb = {{6{p1_add_81921_comb[18]}}, p1_add_81921_comb};
  assign p1_sum__1631_comb = {{6{p1_add_81922_comb[18]}}, p1_add_81922_comb};
  assign p1_sum__1780_comb = {{6{p1_add_81995_comb[18]}}, p1_add_81995_comb};
  assign p1_sum__1781_comb = {{6{p1_add_81996_comb[18]}}, p1_add_81996_comb};
  assign p1_sum__1782_comb = {{6{p1_add_81997_comb[18]}}, p1_add_81997_comb};
  assign p1_sum__1783_comb = {{6{p1_add_81998_comb[18]}}, p1_add_81998_comb};
  assign p1_sum__1608_comb = {{6{p1_add_81999_comb[18]}}, p1_add_81999_comb};
  assign p1_sum__1609_comb = {{6{p1_add_82000_comb[18]}}, p1_add_82000_comb};
  assign p1_sum__1610_comb = {{6{p1_add_82001_comb[18]}}, p1_add_82001_comb};
  assign p1_sum__1611_comb = {{6{p1_add_82002_comb[18]}}, p1_add_82002_comb};
  assign p1_bit_slice_81299_comb = p1_add_80851_comb[19:1];
  assign p1_add_81300_comb = p1_smul_80852_comb + p1_smul_80853_comb;
  assign p1_add_81301_comb = p1_smul_80854_comb + p1_smul_80855_comb;
  assign p1_bit_slice_81302_comb = p1_add_80856_comb[19:1];
  assign p1_bit_slice_81303_comb = p1_add_80857_comb[19:1];
  assign p1_add_81304_comb = p1_smul_80858_comb + p1_smul_80859_comb;
  assign p1_add_81305_comb = p1_smul_80860_comb + p1_smul_80861_comb;
  assign p1_bit_slice_81306_comb = p1_add_80862_comb[19:1];
  assign p1_bit_slice_81307_comb = p1_add_80863_comb[19:1];
  assign p1_add_81308_comb = p1_smul_80864_comb + p1_smul_80865_comb;
  assign p1_add_81309_comb = p1_smul_80866_comb + p1_smul_80867_comb;
  assign p1_bit_slice_81310_comb = p1_add_80868_comb[19:1];
  assign p1_bit_slice_81311_comb = p1_add_80869_comb[19:1];
  assign p1_add_81312_comb = p1_smul_80870_comb + p1_smul_80871_comb;
  assign p1_add_81313_comb = p1_smul_80872_comb + p1_smul_80873_comb;
  assign p1_bit_slice_81314_comb = p1_add_80874_comb[19:1];
  assign p1_smul_81315_comb = smul18b_18b_x_7b(p1_sign_ext_80267_comb[17:0], 7'h3b);
  assign p1_smul_81318_comb = smul18b_18b_x_7b(p1_sign_ext_80214_comb[17:0], 7'h45);
  assign p1_smul_81319_comb = smul18b_18b_x_7b(p1_sign_ext_80215_comb[17:0], 7'h45);
  assign p1_smul_81322_comb = smul18b_18b_x_7b(p1_sign_ext_80272_comb[17:0], 7'h3b);
  assign p1_smul_81323_comb = smul18b_18b_x_7b(p1_sign_ext_80273_comb[17:0], 7'h3b);
  assign p1_smul_81326_comb = smul18b_18b_x_7b(p1_sign_ext_80222_comb[17:0], 7'h45);
  assign p1_smul_81327_comb = smul18b_18b_x_7b(p1_sign_ext_80223_comb[17:0], 7'h45);
  assign p1_smul_81330_comb = smul18b_18b_x_7b(p1_sign_ext_80278_comb[17:0], 7'h3b);
  assign p1_smul_81331_comb = smul18b_18b_x_7b(p1_sign_ext_80279_comb[17:0], 7'h3b);
  assign p1_smul_81334_comb = smul18b_18b_x_7b(p1_sign_ext_80230_comb[17:0], 7'h45);
  assign p1_smul_81335_comb = smul18b_18b_x_7b(p1_sign_ext_80231_comb[17:0], 7'h45);
  assign p1_smul_81338_comb = smul18b_18b_x_7b(p1_sign_ext_80284_comb[17:0], 7'h3b);
  assign p1_smul_81339_comb = smul18b_18b_x_7b(p1_sign_ext_80285_comb[17:0], 7'h3b);
  assign p1_smul_81342_comb = smul18b_18b_x_7b(p1_sign_ext_80238_comb[17:0], 7'h45);
  assign p1_smul_81343_comb = smul18b_18b_x_7b(p1_sign_ext_80239_comb[17:0], 7'h45);
  assign p1_smul_81346_comb = smul18b_18b_x_7b(p1_sign_ext_80290_comb[17:0], 7'h3b);
  assign p1_add_81347_comb = p1_smul_80483_comb[19:1] + p1_smul_80908_comb;
  assign p1_add_81349_comb = p1_smul_80485_comb[19:1] + p1_smul_80910_comb;
  assign p1_add_81351_comb = p1_smul_80911_comb + p1_smul_80490_comb[19:1];
  assign p1_add_81353_comb = p1_smul_80913_comb + p1_smul_80492_comb[19:1];
  assign p1_add_81355_comb = p1_smul_80493_comb[19:1] + p1_smul_80916_comb;
  assign p1_add_81357_comb = p1_smul_80495_comb[19:1] + p1_smul_80918_comb;
  assign p1_add_81359_comb = p1_smul_80919_comb + p1_smul_80500_comb[19:1];
  assign p1_add_81361_comb = p1_smul_80921_comb + p1_smul_80502_comb[19:1];
  assign p1_add_81363_comb = p1_smul_80503_comb[19:1] + p1_smul_80924_comb;
  assign p1_add_81365_comb = p1_smul_80505_comb[19:1] + p1_smul_80926_comb;
  assign p1_add_81367_comb = p1_smul_80927_comb + p1_smul_80510_comb[19:1];
  assign p1_add_81369_comb = p1_smul_80929_comb + p1_smul_80512_comb[19:1];
  assign p1_add_81371_comb = p1_smul_80513_comb[19:1] + p1_smul_80932_comb;
  assign p1_add_81373_comb = p1_smul_80515_comb[19:1] + p1_smul_80934_comb;
  assign p1_add_81375_comb = p1_smul_80935_comb + p1_smul_80520_comb[19:1];
  assign p1_add_81377_comb = p1_smul_80937_comb + p1_smul_80522_comb[19:1];
  assign p1_add_81411_comb = p1_smul_80971_comb + p1_smul_80525_comb[19:1];
  assign p1_add_81413_comb = p1_smul_80973_comb + p1_smul_80527_comb[19:1];
  assign p1_add_81415_comb = p1_smul_80528_comb[19:1] + p1_smul_80976_comb;
  assign p1_add_81417_comb = p1_smul_80530_comb[19:1] + p1_smul_80978_comb;
  assign p1_add_81419_comb = p1_smul_80979_comb + p1_smul_80535_comb[19:1];
  assign p1_add_81421_comb = p1_smul_80981_comb + p1_smul_80537_comb[19:1];
  assign p1_add_81423_comb = p1_smul_80538_comb[19:1] + p1_smul_80984_comb;
  assign p1_add_81425_comb = p1_smul_80540_comb[19:1] + p1_smul_80986_comb;
  assign p1_add_81427_comb = p1_smul_80987_comb + p1_smul_80545_comb[19:1];
  assign p1_add_81429_comb = p1_smul_80989_comb + p1_smul_80547_comb[19:1];
  assign p1_add_81431_comb = p1_smul_80548_comb[19:1] + p1_smul_80992_comb;
  assign p1_add_81433_comb = p1_smul_80550_comb[19:1] + p1_smul_80994_comb;
  assign p1_add_81435_comb = p1_smul_80995_comb + p1_smul_80555_comb[19:1];
  assign p1_add_81437_comb = p1_smul_80997_comb + p1_smul_80557_comb[19:1];
  assign p1_add_81439_comb = p1_smul_80558_comb[19:1] + p1_smul_81000_comb;
  assign p1_add_81441_comb = p1_smul_80560_comb[19:1] + p1_smul_81002_comb;
  assign p1_smul_81444_comb = smul18b_18b_x_7b(p1_sign_ext_80243_comb[17:0], 7'h45);
  assign p1_smul_81446_comb = smul18b_18b_x_7b(p1_sign_ext_80214_comb[17:0], 7'h3b);
  assign p1_smul_81447_comb = smul18b_18b_x_7b(p1_sign_ext_80215_comb[17:0], 7'h3b);
  assign p1_smul_81449_comb = smul18b_18b_x_7b(p1_sign_ext_80244_comb[17:0], 7'h45);
  assign p1_smul_81452_comb = smul18b_18b_x_7b(p1_sign_ext_80245_comb[17:0], 7'h45);
  assign p1_smul_81454_comb = smul18b_18b_x_7b(p1_sign_ext_80222_comb[17:0], 7'h3b);
  assign p1_smul_81455_comb = smul18b_18b_x_7b(p1_sign_ext_80223_comb[17:0], 7'h3b);
  assign p1_smul_81457_comb = smul18b_18b_x_7b(p1_sign_ext_80246_comb[17:0], 7'h45);
  assign p1_smul_81460_comb = smul18b_18b_x_7b(p1_sign_ext_80247_comb[17:0], 7'h45);
  assign p1_smul_81462_comb = smul18b_18b_x_7b(p1_sign_ext_80230_comb[17:0], 7'h3b);
  assign p1_smul_81463_comb = smul18b_18b_x_7b(p1_sign_ext_80231_comb[17:0], 7'h3b);
  assign p1_smul_81465_comb = smul18b_18b_x_7b(p1_sign_ext_80248_comb[17:0], 7'h45);
  assign p1_smul_81468_comb = smul18b_18b_x_7b(p1_sign_ext_80249_comb[17:0], 7'h45);
  assign p1_smul_81470_comb = smul18b_18b_x_7b(p1_sign_ext_80238_comb[17:0], 7'h3b);
  assign p1_smul_81471_comb = smul18b_18b_x_7b(p1_sign_ext_80239_comb[17:0], 7'h3b);
  assign p1_smul_81473_comb = smul18b_18b_x_7b(p1_sign_ext_80250_comb[17:0], 7'h45);
  assign p1_add_81475_comb = p1_smul_81035_comb + p1_smul_81036_comb;
  assign p1_bit_slice_81476_comb = p1_add_81037_comb[19:1];
  assign p1_bit_slice_81477_comb = p1_add_81038_comb[19:1];
  assign p1_add_81478_comb = p1_smul_81039_comb + p1_smul_81040_comb;
  assign p1_add_81479_comb = p1_smul_81041_comb + p1_smul_81042_comb;
  assign p1_bit_slice_81480_comb = p1_add_81043_comb[19:1];
  assign p1_bit_slice_81481_comb = p1_add_81044_comb[19:1];
  assign p1_add_81482_comb = p1_smul_81045_comb + p1_smul_81046_comb;
  assign p1_add_81483_comb = p1_smul_81047_comb + p1_smul_81048_comb;
  assign p1_bit_slice_81484_comb = p1_add_81049_comb[19:1];
  assign p1_bit_slice_81485_comb = p1_add_81050_comb[19:1];
  assign p1_add_81486_comb = p1_smul_81051_comb + p1_smul_81052_comb;
  assign p1_add_81487_comb = p1_smul_81053_comb + p1_smul_81054_comb;
  assign p1_bit_slice_81488_comb = p1_add_81055_comb[19:1];
  assign p1_bit_slice_81489_comb = p1_add_81056_comb[19:1];
  assign p1_add_81490_comb = p1_smul_81057_comb + p1_smul_81058_comb;
  assign p1_bit_slice_81507_comb = p1_add_81059_comb[19:1];
  assign p1_add_81508_comb = p1_smul_81060_comb + p1_smul_81061_comb;
  assign p1_add_81509_comb = p1_smul_81062_comb + p1_smul_81063_comb;
  assign p1_bit_slice_81510_comb = p1_add_81064_comb[19:1];
  assign p1_bit_slice_81511_comb = p1_add_81065_comb[19:1];
  assign p1_add_81512_comb = p1_smul_81066_comb + p1_smul_81067_comb;
  assign p1_add_81513_comb = p1_smul_81068_comb + p1_smul_81069_comb;
  assign p1_bit_slice_81514_comb = p1_add_81070_comb[19:1];
  assign p1_smul_81515_comb = smul18b_18b_x_7b(p1_sign_ext_80335_comb[17:0], 7'h3b);
  assign p1_smul_81518_comb = smul18b_18b_x_7b(p1_sign_ext_80310_comb[17:0], 7'h45);
  assign p1_smul_81519_comb = smul18b_18b_x_7b(p1_sign_ext_80311_comb[17:0], 7'h45);
  assign p1_smul_81522_comb = smul18b_18b_x_7b(p1_sign_ext_80340_comb[17:0], 7'h3b);
  assign p1_smul_81523_comb = smul18b_18b_x_7b(p1_sign_ext_80341_comb[17:0], 7'h3b);
  assign p1_smul_81526_comb = smul18b_18b_x_7b(p1_sign_ext_80318_comb[17:0], 7'h45);
  assign p1_smul_81527_comb = smul18b_18b_x_7b(p1_sign_ext_80319_comb[17:0], 7'h45);
  assign p1_smul_81530_comb = smul18b_18b_x_7b(p1_sign_ext_80346_comb[17:0], 7'h3b);
  assign p1_add_81531_comb = p1_smul_80667_comb[19:1] + p1_smul_81088_comb;
  assign p1_add_81533_comb = p1_smul_80669_comb[19:1] + p1_smul_81090_comb;
  assign p1_add_81535_comb = p1_smul_81091_comb + p1_smul_80674_comb[19:1];
  assign p1_add_81537_comb = p1_smul_81093_comb + p1_smul_80676_comb[19:1];
  assign p1_add_81539_comb = p1_smul_80677_comb[19:1] + p1_smul_81096_comb;
  assign p1_add_81541_comb = p1_smul_80679_comb[19:1] + p1_smul_81098_comb;
  assign p1_add_81543_comb = p1_smul_81099_comb + p1_smul_80684_comb[19:1];
  assign p1_add_81545_comb = p1_smul_81101_comb + p1_smul_80686_comb[19:1];
  assign p1_add_81563_comb = p1_smul_81119_comb + p1_smul_80689_comb[19:1];
  assign p1_add_81565_comb = p1_smul_81121_comb + p1_smul_80691_comb[19:1];
  assign p1_add_81567_comb = p1_smul_80692_comb[19:1] + p1_smul_81124_comb;
  assign p1_add_81569_comb = p1_smul_80694_comb[19:1] + p1_smul_81126_comb;
  assign p1_add_81571_comb = p1_smul_81127_comb + p1_smul_80699_comb[19:1];
  assign p1_add_81573_comb = p1_smul_81129_comb + p1_smul_80701_comb[19:1];
  assign p1_add_81575_comb = p1_smul_80702_comb[19:1] + p1_smul_81132_comb;
  assign p1_add_81577_comb = p1_smul_80704_comb[19:1] + p1_smul_81134_comb;
  assign p1_smul_81580_comb = smul18b_18b_x_7b(p1_sign_ext_80323_comb[17:0], 7'h45);
  assign p1_smul_81582_comb = smul18b_18b_x_7b(p1_sign_ext_80310_comb[17:0], 7'h3b);
  assign p1_smul_81583_comb = smul18b_18b_x_7b(p1_sign_ext_80311_comb[17:0], 7'h3b);
  assign p1_smul_81585_comb = smul18b_18b_x_7b(p1_sign_ext_80324_comb[17:0], 7'h45);
  assign p1_smul_81588_comb = smul18b_18b_x_7b(p1_sign_ext_80325_comb[17:0], 7'h45);
  assign p1_smul_81590_comb = smul18b_18b_x_7b(p1_sign_ext_80318_comb[17:0], 7'h3b);
  assign p1_smul_81591_comb = smul18b_18b_x_7b(p1_sign_ext_80319_comb[17:0], 7'h3b);
  assign p1_smul_81593_comb = smul18b_18b_x_7b(p1_sign_ext_80326_comb[17:0], 7'h45);
  assign p1_add_81595_comb = p1_smul_81151_comb + p1_smul_81152_comb;
  assign p1_bit_slice_81596_comb = p1_add_81153_comb[19:1];
  assign p1_bit_slice_81597_comb = p1_add_81154_comb[19:1];
  assign p1_add_81598_comb = p1_smul_81155_comb + p1_smul_81156_comb;
  assign p1_add_81599_comb = p1_smul_81157_comb + p1_smul_81158_comb;
  assign p1_bit_slice_81600_comb = p1_add_81159_comb[19:1];
  assign p1_bit_slice_81601_comb = p1_add_81160_comb[19:1];
  assign p1_add_81602_comb = p1_smul_81161_comb + p1_smul_81162_comb;
  assign p1_bit_slice_81619_comb = p1_add_81163_comb[19:1];
  assign p1_add_81620_comb = p1_smul_81164_comb + p1_smul_81165_comb;
  assign p1_add_81621_comb = p1_smul_81166_comb + p1_smul_81167_comb;
  assign p1_bit_slice_81622_comb = p1_add_81168_comb[19:1];
  assign p1_bit_slice_81623_comb = p1_add_81169_comb[19:1];
  assign p1_add_81624_comb = p1_smul_81170_comb + p1_smul_81171_comb;
  assign p1_add_81625_comb = p1_smul_81172_comb + p1_smul_81173_comb;
  assign p1_bit_slice_81626_comb = p1_add_81174_comb[19:1];
  assign p1_smul_81627_comb = smul18b_18b_x_7b(p1_sign_ext_80383_comb[17:0], 7'h3b);
  assign p1_smul_81630_comb = smul18b_18b_x_7b(p1_sign_ext_80358_comb[17:0], 7'h45);
  assign p1_smul_81631_comb = smul18b_18b_x_7b(p1_sign_ext_80359_comb[17:0], 7'h45);
  assign p1_smul_81634_comb = smul18b_18b_x_7b(p1_sign_ext_80388_comb[17:0], 7'h3b);
  assign p1_smul_81635_comb = smul18b_18b_x_7b(p1_sign_ext_80389_comb[17:0], 7'h3b);
  assign p1_smul_81638_comb = smul18b_18b_x_7b(p1_sign_ext_80366_comb[17:0], 7'h45);
  assign p1_smul_81639_comb = smul18b_18b_x_7b(p1_sign_ext_80367_comb[17:0], 7'h45);
  assign p1_smul_81642_comb = smul18b_18b_x_7b(p1_sign_ext_80394_comb[17:0], 7'h3b);
  assign p1_add_81643_comb = p1_smul_80779_comb[19:1] + p1_smul_81192_comb;
  assign p1_add_81645_comb = p1_smul_80781_comb[19:1] + p1_smul_81194_comb;
  assign p1_add_81647_comb = p1_smul_81195_comb + p1_smul_80786_comb[19:1];
  assign p1_add_81649_comb = p1_smul_81197_comb + p1_smul_80788_comb[19:1];
  assign p1_add_81651_comb = p1_smul_80789_comb[19:1] + p1_smul_81200_comb;
  assign p1_add_81653_comb = p1_smul_80791_comb[19:1] + p1_smul_81202_comb;
  assign p1_add_81655_comb = p1_smul_81203_comb + p1_smul_80796_comb[19:1];
  assign p1_add_81657_comb = p1_smul_81205_comb + p1_smul_80798_comb[19:1];
  assign p1_add_81675_comb = p1_smul_81223_comb + p1_smul_80801_comb[19:1];
  assign p1_add_81677_comb = p1_smul_81225_comb + p1_smul_80803_comb[19:1];
  assign p1_add_81679_comb = p1_smul_80804_comb[19:1] + p1_smul_81228_comb;
  assign p1_add_81681_comb = p1_smul_80806_comb[19:1] + p1_smul_81230_comb;
  assign p1_add_81683_comb = p1_smul_81231_comb + p1_smul_80811_comb[19:1];
  assign p1_add_81685_comb = p1_smul_81233_comb + p1_smul_80813_comb[19:1];
  assign p1_add_81687_comb = p1_smul_80814_comb[19:1] + p1_smul_81236_comb;
  assign p1_add_81689_comb = p1_smul_80816_comb[19:1] + p1_smul_81238_comb;
  assign p1_smul_81692_comb = smul18b_18b_x_7b(p1_sign_ext_80371_comb[17:0], 7'h45);
  assign p1_smul_81694_comb = smul18b_18b_x_7b(p1_sign_ext_80358_comb[17:0], 7'h3b);
  assign p1_smul_81695_comb = smul18b_18b_x_7b(p1_sign_ext_80359_comb[17:0], 7'h3b);
  assign p1_smul_81697_comb = smul18b_18b_x_7b(p1_sign_ext_80372_comb[17:0], 7'h45);
  assign p1_smul_81700_comb = smul18b_18b_x_7b(p1_sign_ext_80373_comb[17:0], 7'h45);
  assign p1_smul_81702_comb = smul18b_18b_x_7b(p1_sign_ext_80366_comb[17:0], 7'h3b);
  assign p1_smul_81703_comb = smul18b_18b_x_7b(p1_sign_ext_80367_comb[17:0], 7'h3b);
  assign p1_smul_81705_comb = smul18b_18b_x_7b(p1_sign_ext_80374_comb[17:0], 7'h45);
  assign p1_add_81707_comb = p1_smul_81255_comb + p1_smul_81256_comb;
  assign p1_bit_slice_81708_comb = p1_add_81257_comb[19:1];
  assign p1_bit_slice_81709_comb = p1_add_81258_comb[19:1];
  assign p1_add_81710_comb = p1_smul_81259_comb + p1_smul_81260_comb;
  assign p1_add_81711_comb = p1_smul_81261_comb + p1_smul_81262_comb;
  assign p1_bit_slice_81712_comb = p1_add_81263_comb[19:1];
  assign p1_bit_slice_81713_comb = p1_add_81264_comb[19:1];
  assign p1_add_81714_comb = p1_smul_81265_comb + p1_smul_81266_comb;
  assign p1_sum__1324_comb = p1_sum__1736_comb + p1_sum__1737_comb;
  assign p1_sum__1325_comb = p1_sum__1738_comb + p1_sum__1739_comb;
  assign p1_sum__1310_comb = p1_sum__1708_comb + p1_sum__1709_comb;
  assign p1_sum__1311_comb = p1_sum__1710_comb + p1_sum__1711_comb;
  assign p1_sum__1296_comb = p1_sum__1680_comb + p1_sum__1681_comb;
  assign p1_sum__1297_comb = p1_sum__1682_comb + p1_sum__1683_comb;
  assign p1_sum__1282_comb = p1_sum__1652_comb + p1_sum__1653_comb;
  assign p1_sum__1283_comb = p1_sum__1654_comb + p1_sum__1655_comb;
  assign p1_sum__1336_comb = p1_sum__1760_comb + p1_sum__1761_comb;
  assign p1_sum__1337_comb = p1_sum__1762_comb + p1_sum__1763_comb;
  assign p1_sum__1270_comb = p1_sum__1628_comb + p1_sum__1629_comb;
  assign p1_sum__1271_comb = p1_sum__1630_comb + p1_sum__1631_comb;
  assign p1_sum__1346_comb = p1_sum__1780_comb + p1_sum__1781_comb;
  assign p1_sum__1347_comb = p1_sum__1782_comb + p1_sum__1783_comb;
  assign p1_sum__1260_comb = p1_sum__1608_comb + p1_sum__1609_comb;
  assign p1_sum__1261_comb = p1_sum__1610_comb + p1_sum__1611_comb;
  assign p1_add_81747_comb = p1_smul_81315_comb + p1_smul_80876_comb[18:1];
  assign p1_add_81749_comb = p1_smul_80877_comb[18:1] + p1_smul_81318_comb;
  assign p1_add_81751_comb = p1_smul_81319_comb + p1_smul_80880_comb[18:1];
  assign p1_add_81753_comb = p1_smul_80881_comb[18:1] + p1_smul_81322_comb;
  assign p1_add_81755_comb = p1_smul_81323_comb + p1_smul_80884_comb[18:1];
  assign p1_add_81757_comb = p1_smul_80885_comb[18:1] + p1_smul_81326_comb;
  assign p1_add_81759_comb = p1_smul_81327_comb + p1_smul_80888_comb[18:1];
  assign p1_add_81761_comb = p1_smul_80889_comb[18:1] + p1_smul_81330_comb;
  assign p1_add_81763_comb = p1_smul_81331_comb + p1_smul_80892_comb[18:1];
  assign p1_add_81765_comb = p1_smul_80893_comb[18:1] + p1_smul_81334_comb;
  assign p1_add_81767_comb = p1_smul_81335_comb + p1_smul_80896_comb[18:1];
  assign p1_add_81769_comb = p1_smul_80897_comb[18:1] + p1_smul_81338_comb;
  assign p1_add_81771_comb = p1_smul_81339_comb + p1_smul_80900_comb[18:1];
  assign p1_add_81773_comb = p1_smul_80901_comb[18:1] + p1_smul_81342_comb;
  assign p1_add_81775_comb = p1_smul_81343_comb + p1_smul_80904_comb[18:1];
  assign p1_add_81777_comb = p1_smul_80905_comb[18:1] + p1_smul_81346_comb;
  assign p1_concat_81779_comb = {p1_add_81347_comb, p1_smul_80483_comb[0]};
  assign p1_concat_81780_comb = {p1_add_81349_comb, p1_smul_80485_comb[0]};
  assign p1_concat_81781_comb = {p1_add_81351_comb, p1_smul_80490_comb[0]};
  assign p1_concat_81782_comb = {p1_add_81353_comb, p1_smul_80492_comb[0]};
  assign p1_concat_81783_comb = {p1_add_81355_comb, p1_smul_80493_comb[0]};
  assign p1_concat_81784_comb = {p1_add_81357_comb, p1_smul_80495_comb[0]};
  assign p1_concat_81785_comb = {p1_add_81359_comb, p1_smul_80500_comb[0]};
  assign p1_concat_81786_comb = {p1_add_81361_comb, p1_smul_80502_comb[0]};
  assign p1_concat_81787_comb = {p1_add_81363_comb, p1_smul_80503_comb[0]};
  assign p1_concat_81788_comb = {p1_add_81365_comb, p1_smul_80505_comb[0]};
  assign p1_concat_81789_comb = {p1_add_81367_comb, p1_smul_80510_comb[0]};
  assign p1_concat_81790_comb = {p1_add_81369_comb, p1_smul_80512_comb[0]};
  assign p1_concat_81791_comb = {p1_add_81371_comb, p1_smul_80513_comb[0]};
  assign p1_concat_81792_comb = {p1_add_81373_comb, p1_smul_80515_comb[0]};
  assign p1_concat_81793_comb = {p1_add_81375_comb, p1_smul_80520_comb[0]};
  assign p1_concat_81794_comb = {p1_add_81377_comb, p1_smul_80522_comb[0]};
  assign p1_concat_81811_comb = {p1_add_81411_comb, p1_smul_80525_comb[0]};
  assign p1_concat_81812_comb = {p1_add_81413_comb, p1_smul_80527_comb[0]};
  assign p1_concat_81813_comb = {p1_add_81415_comb, p1_smul_80528_comb[0]};
  assign p1_concat_81814_comb = {p1_add_81417_comb, p1_smul_80530_comb[0]};
  assign p1_concat_81815_comb = {p1_add_81419_comb, p1_smul_80535_comb[0]};
  assign p1_concat_81816_comb = {p1_add_81421_comb, p1_smul_80537_comb[0]};
  assign p1_concat_81817_comb = {p1_add_81423_comb, p1_smul_80538_comb[0]};
  assign p1_concat_81818_comb = {p1_add_81425_comb, p1_smul_80540_comb[0]};
  assign p1_concat_81819_comb = {p1_add_81427_comb, p1_smul_80545_comb[0]};
  assign p1_concat_81820_comb = {p1_add_81429_comb, p1_smul_80547_comb[0]};
  assign p1_concat_81821_comb = {p1_add_81431_comb, p1_smul_80548_comb[0]};
  assign p1_concat_81822_comb = {p1_add_81433_comb, p1_smul_80550_comb[0]};
  assign p1_concat_81823_comb = {p1_add_81435_comb, p1_smul_80555_comb[0]};
  assign p1_concat_81824_comb = {p1_add_81437_comb, p1_smul_80557_comb[0]};
  assign p1_concat_81825_comb = {p1_add_81439_comb, p1_smul_80558_comb[0]};
  assign p1_concat_81826_comb = {p1_add_81441_comb, p1_smul_80560_comb[0]};
  assign p1_add_81827_comb = p1_smul_81003_comb[18:1] + p1_smul_81444_comb;
  assign p1_add_81829_comb = p1_smul_81005_comb[18:1] + p1_smul_81446_comb;
  assign p1_add_81831_comb = p1_smul_81447_comb + p1_smul_81008_comb[18:1];
  assign p1_add_81833_comb = p1_smul_81449_comb + p1_smul_81010_comb[18:1];
  assign p1_add_81835_comb = p1_smul_81011_comb[18:1] + p1_smul_81452_comb;
  assign p1_add_81837_comb = p1_smul_81013_comb[18:1] + p1_smul_81454_comb;
  assign p1_add_81839_comb = p1_smul_81455_comb + p1_smul_81016_comb[18:1];
  assign p1_add_81841_comb = p1_smul_81457_comb + p1_smul_81018_comb[18:1];
  assign p1_add_81843_comb = p1_smul_81019_comb[18:1] + p1_smul_81460_comb;
  assign p1_add_81845_comb = p1_smul_81021_comb[18:1] + p1_smul_81462_comb;
  assign p1_add_81847_comb = p1_smul_81463_comb + p1_smul_81024_comb[18:1];
  assign p1_add_81849_comb = p1_smul_81465_comb + p1_smul_81026_comb[18:1];
  assign p1_add_81851_comb = p1_smul_81027_comb[18:1] + p1_smul_81468_comb;
  assign p1_add_81853_comb = p1_smul_81029_comb[18:1] + p1_smul_81470_comb;
  assign p1_add_81855_comb = p1_smul_81471_comb + p1_smul_81032_comb[18:1];
  assign p1_add_81857_comb = p1_smul_81473_comb + p1_smul_81034_comb[18:1];
  assign p1_add_81891_comb = p1_smul_81515_comb + p1_smul_81072_comb[18:1];
  assign p1_add_81893_comb = p1_smul_81073_comb[18:1] + p1_smul_81518_comb;
  assign p1_add_81895_comb = p1_smul_81519_comb + p1_smul_81076_comb[18:1];
  assign p1_add_81897_comb = p1_smul_81077_comb[18:1] + p1_smul_81522_comb;
  assign p1_add_81899_comb = p1_smul_81523_comb + p1_smul_81080_comb[18:1];
  assign p1_add_81901_comb = p1_smul_81081_comb[18:1] + p1_smul_81526_comb;
  assign p1_add_81903_comb = p1_smul_81527_comb + p1_smul_81084_comb[18:1];
  assign p1_add_81905_comb = p1_smul_81085_comb[18:1] + p1_smul_81530_comb;
  assign p1_concat_81907_comb = {p1_add_81531_comb, p1_smul_80667_comb[0]};
  assign p1_concat_81908_comb = {p1_add_81533_comb, p1_smul_80669_comb[0]};
  assign p1_concat_81909_comb = {p1_add_81535_comb, p1_smul_80674_comb[0]};
  assign p1_concat_81910_comb = {p1_add_81537_comb, p1_smul_80676_comb[0]};
  assign p1_concat_81911_comb = {p1_add_81539_comb, p1_smul_80677_comb[0]};
  assign p1_concat_81912_comb = {p1_add_81541_comb, p1_smul_80679_comb[0]};
  assign p1_concat_81913_comb = {p1_add_81543_comb, p1_smul_80684_comb[0]};
  assign p1_concat_81914_comb = {p1_add_81545_comb, p1_smul_80686_comb[0]};
  assign p1_concat_81923_comb = {p1_add_81563_comb, p1_smul_80689_comb[0]};
  assign p1_concat_81924_comb = {p1_add_81565_comb, p1_smul_80691_comb[0]};
  assign p1_concat_81925_comb = {p1_add_81567_comb, p1_smul_80692_comb[0]};
  assign p1_concat_81926_comb = {p1_add_81569_comb, p1_smul_80694_comb[0]};
  assign p1_concat_81927_comb = {p1_add_81571_comb, p1_smul_80699_comb[0]};
  assign p1_concat_81928_comb = {p1_add_81573_comb, p1_smul_80701_comb[0]};
  assign p1_concat_81929_comb = {p1_add_81575_comb, p1_smul_80702_comb[0]};
  assign p1_concat_81930_comb = {p1_add_81577_comb, p1_smul_80704_comb[0]};
  assign p1_add_81931_comb = p1_smul_81135_comb[18:1] + p1_smul_81580_comb;
  assign p1_add_81933_comb = p1_smul_81137_comb[18:1] + p1_smul_81582_comb;
  assign p1_add_81935_comb = p1_smul_81583_comb + p1_smul_81140_comb[18:1];
  assign p1_add_81937_comb = p1_smul_81585_comb + p1_smul_81142_comb[18:1];
  assign p1_add_81939_comb = p1_smul_81143_comb[18:1] + p1_smul_81588_comb;
  assign p1_add_81941_comb = p1_smul_81145_comb[18:1] + p1_smul_81590_comb;
  assign p1_add_81943_comb = p1_smul_81591_comb + p1_smul_81148_comb[18:1];
  assign p1_add_81945_comb = p1_smul_81593_comb + p1_smul_81150_comb[18:1];
  assign p1_add_81971_comb = p1_smul_81627_comb + p1_smul_81176_comb[18:1];
  assign p1_add_81973_comb = p1_smul_81177_comb[18:1] + p1_smul_81630_comb;
  assign p1_add_81975_comb = p1_smul_81631_comb + p1_smul_81180_comb[18:1];
  assign p1_add_81977_comb = p1_smul_81181_comb[18:1] + p1_smul_81634_comb;
  assign p1_add_81979_comb = p1_smul_81635_comb + p1_smul_81184_comb[18:1];
  assign p1_add_81981_comb = p1_smul_81185_comb[18:1] + p1_smul_81638_comb;
  assign p1_add_81983_comb = p1_smul_81639_comb + p1_smul_81188_comb[18:1];
  assign p1_add_81985_comb = p1_smul_81189_comb[18:1] + p1_smul_81642_comb;
  assign p1_concat_81987_comb = {p1_add_81643_comb, p1_smul_80779_comb[0]};
  assign p1_concat_81988_comb = {p1_add_81645_comb, p1_smul_80781_comb[0]};
  assign p1_concat_81989_comb = {p1_add_81647_comb, p1_smul_80786_comb[0]};
  assign p1_concat_81990_comb = {p1_add_81649_comb, p1_smul_80788_comb[0]};
  assign p1_concat_81991_comb = {p1_add_81651_comb, p1_smul_80789_comb[0]};
  assign p1_concat_81992_comb = {p1_add_81653_comb, p1_smul_80791_comb[0]};
  assign p1_concat_81993_comb = {p1_add_81655_comb, p1_smul_80796_comb[0]};
  assign p1_concat_81994_comb = {p1_add_81657_comb, p1_smul_80798_comb[0]};
  assign p1_concat_82003_comb = {p1_add_81675_comb, p1_smul_80801_comb[0]};
  assign p1_concat_82004_comb = {p1_add_81677_comb, p1_smul_80803_comb[0]};
  assign p1_concat_82005_comb = {p1_add_81679_comb, p1_smul_80804_comb[0]};
  assign p1_concat_82006_comb = {p1_add_81681_comb, p1_smul_80806_comb[0]};
  assign p1_concat_82007_comb = {p1_add_81683_comb, p1_smul_80811_comb[0]};
  assign p1_concat_82008_comb = {p1_add_81685_comb, p1_smul_80813_comb[0]};
  assign p1_concat_82009_comb = {p1_add_81687_comb, p1_smul_80814_comb[0]};
  assign p1_concat_82010_comb = {p1_add_81689_comb, p1_smul_80816_comb[0]};
  assign p1_add_82011_comb = p1_smul_81239_comb[18:1] + p1_smul_81692_comb;
  assign p1_add_82013_comb = p1_smul_81241_comb[18:1] + p1_smul_81694_comb;
  assign p1_add_82015_comb = p1_smul_81695_comb + p1_smul_81244_comb[18:1];
  assign p1_add_82017_comb = p1_smul_81697_comb + p1_smul_81246_comb[18:1];
  assign p1_add_82019_comb = p1_smul_81247_comb[18:1] + p1_smul_81700_comb;
  assign p1_add_82021_comb = p1_smul_81249_comb[18:1] + p1_smul_81702_comb;
  assign p1_add_82023_comb = p1_smul_81703_comb + p1_smul_81252_comb[18:1];
  assign p1_add_82025_comb = p1_smul_81705_comb + p1_smul_81254_comb[18:1];
  assign p1_add_82291_comb = {{12{p1_add_81715_comb[11]}}, p1_add_81715_comb} + {{12{p1_add_81716_comb[11]}}, p1_add_81716_comb};
  assign p1_add_82292_comb = {{12{p1_add_81717_comb[11]}}, p1_add_81717_comb} + {{12{p1_add_81718_comb[11]}}, p1_add_81718_comb};
  assign p1_add_82293_comb = {{12{p1_add_81719_comb[11]}}, p1_add_81719_comb} + {{12{p1_add_81720_comb[11]}}, p1_add_81720_comb};
  assign p1_add_82294_comb = {{12{p1_add_81721_comb[11]}}, p1_add_81721_comb} + {{12{p1_add_81722_comb[11]}}, p1_add_81722_comb};
  assign p1_add_82295_comb = {{12{p1_add_81723_comb[11]}}, p1_add_81723_comb} + {{12{p1_add_81724_comb[11]}}, p1_add_81724_comb};
  assign p1_add_82296_comb = {{12{p1_add_81725_comb[11]}}, p1_add_81725_comb} + {{12{p1_add_81726_comb[11]}}, p1_add_81726_comb};
  assign p1_add_82297_comb = {{12{p1_add_81727_comb[11]}}, p1_add_81727_comb} + {{12{p1_add_81728_comb[11]}}, p1_add_81728_comb};
  assign p1_add_82298_comb = {{12{p1_add_81729_comb[11]}}, p1_add_81729_comb} + {{12{p1_add_81730_comb[11]}}, p1_add_81730_comb};
  assign p1_add_82371_comb = {{12{p1_add_81875_comb[11]}}, p1_add_81875_comb} + {{12{p1_add_81876_comb[11]}}, p1_add_81876_comb};
  assign p1_add_82372_comb = {{12{p1_add_81877_comb[11]}}, p1_add_81877_comb} + {{12{p1_add_81878_comb[11]}}, p1_add_81878_comb};
  assign p1_add_82373_comb = {{12{p1_add_81879_comb[11]}}, p1_add_81879_comb} + {{12{p1_add_81880_comb[11]}}, p1_add_81880_comb};
  assign p1_add_82374_comb = {{12{p1_add_81881_comb[11]}}, p1_add_81881_comb} + {{12{p1_add_81882_comb[11]}}, p1_add_81882_comb};
  assign p1_add_82411_comb = {{12{p1_add_81955_comb[11]}}, p1_add_81955_comb} + {{12{p1_add_81956_comb[11]}}, p1_add_81956_comb};
  assign p1_add_82412_comb = {{12{p1_add_81957_comb[11]}}, p1_add_81957_comb} + {{12{p1_add_81958_comb[11]}}, p1_add_81958_comb};
  assign p1_add_82413_comb = {{12{p1_add_81959_comb[11]}}, p1_add_81959_comb} + {{12{p1_add_81960_comb[11]}}, p1_add_81960_comb};
  assign p1_add_82414_comb = {{12{p1_add_81961_comb[11]}}, p1_add_81961_comb} + {{12{p1_add_81962_comb[11]}}, p1_add_81962_comb};
  assign p1_sum__1118_comb = p1_sum__1324_comb + p1_sum__1325_comb;
  assign p1_sum__1111_comb = p1_sum__1310_comb + p1_sum__1311_comb;
  assign p1_sum__1104_comb = p1_sum__1296_comb + p1_sum__1297_comb;
  assign p1_sum__1097_comb = p1_sum__1282_comb + p1_sum__1283_comb;
  assign p1_sum__1124_comb = p1_sum__1336_comb + p1_sum__1337_comb;
  assign p1_sum__1091_comb = p1_sum__1270_comb + p1_sum__1271_comb;
  assign p1_sum__1129_comb = p1_sum__1346_comb + p1_sum__1347_comb;
  assign p1_sum__1086_comb = p1_sum__1260_comb + p1_sum__1261_comb;
  assign p1_add_82051_comb = {{5{p1_bit_slice_81299_comb[18]}}, p1_bit_slice_81299_comb} + {{6{p1_add_81300_comb[17]}}, p1_add_81300_comb};
  assign p1_add_82053_comb = {{6{p1_add_81301_comb[17]}}, p1_add_81301_comb} + {{5{p1_bit_slice_81302_comb[18]}}, p1_bit_slice_81302_comb};
  assign p1_add_82055_comb = {{5{p1_bit_slice_81303_comb[18]}}, p1_bit_slice_81303_comb} + {{6{p1_add_81304_comb[17]}}, p1_add_81304_comb};
  assign p1_add_82057_comb = {{6{p1_add_81305_comb[17]}}, p1_add_81305_comb} + {{5{p1_bit_slice_81306_comb[18]}}, p1_bit_slice_81306_comb};
  assign p1_add_82059_comb = {{5{p1_bit_slice_81307_comb[18]}}, p1_bit_slice_81307_comb} + {{6{p1_add_81308_comb[17]}}, p1_add_81308_comb};
  assign p1_add_82061_comb = {{6{p1_add_81309_comb[17]}}, p1_add_81309_comb} + {{5{p1_bit_slice_81310_comb[18]}}, p1_bit_slice_81310_comb};
  assign p1_add_82063_comb = {{5{p1_bit_slice_81311_comb[18]}}, p1_bit_slice_81311_comb} + {{6{p1_add_81312_comb[17]}}, p1_add_81312_comb};
  assign p1_add_82065_comb = {{6{p1_add_81313_comb[17]}}, p1_add_81313_comb} + {{5{p1_bit_slice_81314_comb[18]}}, p1_bit_slice_81314_comb};
  assign p1_concat_82067_comb = {p1_add_81747_comb, p1_smul_80876_comb[0]};
  assign p1_concat_82068_comb = {p1_add_81749_comb, p1_smul_80877_comb[0]};
  assign p1_concat_82069_comb = {p1_add_81751_comb, p1_smul_80880_comb[0]};
  assign p1_concat_82070_comb = {p1_add_81753_comb, p1_smul_80881_comb[0]};
  assign p1_concat_82071_comb = {p1_add_81755_comb, p1_smul_80884_comb[0]};
  assign p1_concat_82072_comb = {p1_add_81757_comb, p1_smul_80885_comb[0]};
  assign p1_concat_82073_comb = {p1_add_81759_comb, p1_smul_80888_comb[0]};
  assign p1_concat_82074_comb = {p1_add_81761_comb, p1_smul_80889_comb[0]};
  assign p1_concat_82075_comb = {p1_add_81763_comb, p1_smul_80892_comb[0]};
  assign p1_concat_82076_comb = {p1_add_81765_comb, p1_smul_80893_comb[0]};
  assign p1_concat_82077_comb = {p1_add_81767_comb, p1_smul_80896_comb[0]};
  assign p1_concat_82078_comb = {p1_add_81769_comb, p1_smul_80897_comb[0]};
  assign p1_concat_82079_comb = {p1_add_81771_comb, p1_smul_80900_comb[0]};
  assign p1_concat_82080_comb = {p1_add_81773_comb, p1_smul_80901_comb[0]};
  assign p1_concat_82081_comb = {p1_add_81775_comb, p1_smul_80904_comb[0]};
  assign p1_concat_82082_comb = {p1_add_81777_comb, p1_smul_80905_comb[0]};
  assign p1_sum__1756_comb = {{5{p1_concat_81779_comb[19]}}, p1_concat_81779_comb};
  assign p1_sum__1757_comb = {{5{p1_concat_81780_comb[19]}}, p1_concat_81780_comb};
  assign p1_sum__1758_comb = {{5{p1_concat_81781_comb[19]}}, p1_concat_81781_comb};
  assign p1_sum__1759_comb = {{5{p1_concat_81782_comb[19]}}, p1_concat_81782_comb};
  assign p1_sum__1732_comb = {{5{p1_concat_81783_comb[19]}}, p1_concat_81783_comb};
  assign p1_sum__1733_comb = {{5{p1_concat_81784_comb[19]}}, p1_concat_81784_comb};
  assign p1_sum__1734_comb = {{5{p1_concat_81785_comb[19]}}, p1_concat_81785_comb};
  assign p1_sum__1735_comb = {{5{p1_concat_81786_comb[19]}}, p1_concat_81786_comb};
  assign p1_sum__1704_comb = {{5{p1_concat_81787_comb[19]}}, p1_concat_81787_comb};
  assign p1_sum__1705_comb = {{5{p1_concat_81788_comb[19]}}, p1_concat_81788_comb};
  assign p1_sum__1706_comb = {{5{p1_concat_81789_comb[19]}}, p1_concat_81789_comb};
  assign p1_sum__1707_comb = {{5{p1_concat_81790_comb[19]}}, p1_concat_81790_comb};
  assign p1_sum__1676_comb = {{5{p1_concat_81791_comb[19]}}, p1_concat_81791_comb};
  assign p1_sum__1677_comb = {{5{p1_concat_81792_comb[19]}}, p1_concat_81792_comb};
  assign p1_sum__1678_comb = {{5{p1_concat_81793_comb[19]}}, p1_concat_81793_comb};
  assign p1_sum__1679_comb = {{5{p1_concat_81794_comb[19]}}, p1_concat_81794_comb};
  assign p1_sum__1712_comb = {{5{p1_concat_81811_comb[19]}}, p1_concat_81811_comb};
  assign p1_sum__1713_comb = {{5{p1_concat_81812_comb[19]}}, p1_concat_81812_comb};
  assign p1_sum__1714_comb = {{5{p1_concat_81813_comb[19]}}, p1_concat_81813_comb};
  assign p1_sum__1715_comb = {{5{p1_concat_81814_comb[19]}}, p1_concat_81814_comb};
  assign p1_sum__1684_comb = {{5{p1_concat_81815_comb[19]}}, p1_concat_81815_comb};
  assign p1_sum__1685_comb = {{5{p1_concat_81816_comb[19]}}, p1_concat_81816_comb};
  assign p1_sum__1686_comb = {{5{p1_concat_81817_comb[19]}}, p1_concat_81817_comb};
  assign p1_sum__1687_comb = {{5{p1_concat_81818_comb[19]}}, p1_concat_81818_comb};
  assign p1_sum__1656_comb = {{5{p1_concat_81819_comb[19]}}, p1_concat_81819_comb};
  assign p1_sum__1657_comb = {{5{p1_concat_81820_comb[19]}}, p1_concat_81820_comb};
  assign p1_sum__1658_comb = {{5{p1_concat_81821_comb[19]}}, p1_concat_81821_comb};
  assign p1_sum__1659_comb = {{5{p1_concat_81822_comb[19]}}, p1_concat_81822_comb};
  assign p1_sum__1632_comb = {{5{p1_concat_81823_comb[19]}}, p1_concat_81823_comb};
  assign p1_sum__1633_comb = {{5{p1_concat_81824_comb[19]}}, p1_concat_81824_comb};
  assign p1_sum__1634_comb = {{5{p1_concat_81825_comb[19]}}, p1_concat_81825_comb};
  assign p1_sum__1635_comb = {{5{p1_concat_81826_comb[19]}}, p1_concat_81826_comb};
  assign p1_concat_82131_comb = {p1_add_81827_comb, p1_smul_81003_comb[0]};
  assign p1_concat_82132_comb = {p1_add_81829_comb, p1_smul_81005_comb[0]};
  assign p1_concat_82133_comb = {p1_add_81831_comb, p1_smul_81008_comb[0]};
  assign p1_concat_82134_comb = {p1_add_81833_comb, p1_smul_81010_comb[0]};
  assign p1_concat_82135_comb = {p1_add_81835_comb, p1_smul_81011_comb[0]};
  assign p1_concat_82136_comb = {p1_add_81837_comb, p1_smul_81013_comb[0]};
  assign p1_concat_82137_comb = {p1_add_81839_comb, p1_smul_81016_comb[0]};
  assign p1_concat_82138_comb = {p1_add_81841_comb, p1_smul_81018_comb[0]};
  assign p1_concat_82139_comb = {p1_add_81843_comb, p1_smul_81019_comb[0]};
  assign p1_concat_82140_comb = {p1_add_81845_comb, p1_smul_81021_comb[0]};
  assign p1_concat_82141_comb = {p1_add_81847_comb, p1_smul_81024_comb[0]};
  assign p1_concat_82142_comb = {p1_add_81849_comb, p1_smul_81026_comb[0]};
  assign p1_concat_82143_comb = {p1_add_81851_comb, p1_smul_81027_comb[0]};
  assign p1_concat_82144_comb = {p1_add_81853_comb, p1_smul_81029_comb[0]};
  assign p1_concat_82145_comb = {p1_add_81855_comb, p1_smul_81032_comb[0]};
  assign p1_concat_82146_comb = {p1_add_81857_comb, p1_smul_81034_comb[0]};
  assign p1_add_82147_comb = {{6{p1_add_81475_comb[17]}}, p1_add_81475_comb} + {{5{p1_bit_slice_81476_comb[18]}}, p1_bit_slice_81476_comb};
  assign p1_add_82149_comb = {{5{p1_bit_slice_81477_comb[18]}}, p1_bit_slice_81477_comb} + {{6{p1_add_81478_comb[17]}}, p1_add_81478_comb};
  assign p1_add_82151_comb = {{6{p1_add_81479_comb[17]}}, p1_add_81479_comb} + {{5{p1_bit_slice_81480_comb[18]}}, p1_bit_slice_81480_comb};
  assign p1_add_82153_comb = {{5{p1_bit_slice_81481_comb[18]}}, p1_bit_slice_81481_comb} + {{6{p1_add_81482_comb[17]}}, p1_add_81482_comb};
  assign p1_add_82155_comb = {{6{p1_add_81483_comb[17]}}, p1_add_81483_comb} + {{5{p1_bit_slice_81484_comb[18]}}, p1_bit_slice_81484_comb};
  assign p1_add_82157_comb = {{5{p1_bit_slice_81485_comb[18]}}, p1_bit_slice_81485_comb} + {{6{p1_add_81486_comb[17]}}, p1_add_81486_comb};
  assign p1_add_82159_comb = {{6{p1_add_81487_comb[17]}}, p1_add_81487_comb} + {{5{p1_bit_slice_81488_comb[18]}}, p1_bit_slice_81488_comb};
  assign p1_add_82161_comb = {{5{p1_bit_slice_81489_comb[18]}}, p1_bit_slice_81489_comb} + {{6{p1_add_81490_comb[17]}}, p1_add_81490_comb};
  assign p1_add_82171_comb = {{5{p1_bit_slice_81507_comb[18]}}, p1_bit_slice_81507_comb} + {{6{p1_add_81508_comb[17]}}, p1_add_81508_comb};
  assign p1_add_82173_comb = {{6{p1_add_81509_comb[17]}}, p1_add_81509_comb} + {{5{p1_bit_slice_81510_comb[18]}}, p1_bit_slice_81510_comb};
  assign p1_add_82175_comb = {{5{p1_bit_slice_81511_comb[18]}}, p1_bit_slice_81511_comb} + {{6{p1_add_81512_comb[17]}}, p1_add_81512_comb};
  assign p1_add_82177_comb = {{6{p1_add_81513_comb[17]}}, p1_add_81513_comb} + {{5{p1_bit_slice_81514_comb[18]}}, p1_bit_slice_81514_comb};
  assign p1_concat_82179_comb = {p1_add_81891_comb, p1_smul_81072_comb[0]};
  assign p1_concat_82180_comb = {p1_add_81893_comb, p1_smul_81073_comb[0]};
  assign p1_concat_82181_comb = {p1_add_81895_comb, p1_smul_81076_comb[0]};
  assign p1_concat_82182_comb = {p1_add_81897_comb, p1_smul_81077_comb[0]};
  assign p1_concat_82183_comb = {p1_add_81899_comb, p1_smul_81080_comb[0]};
  assign p1_concat_82184_comb = {p1_add_81901_comb, p1_smul_81081_comb[0]};
  assign p1_concat_82185_comb = {p1_add_81903_comb, p1_smul_81084_comb[0]};
  assign p1_concat_82186_comb = {p1_add_81905_comb, p1_smul_81085_comb[0]};
  assign p1_sum__1776_comb = {{5{p1_concat_81907_comb[19]}}, p1_concat_81907_comb};
  assign p1_sum__1777_comb = {{5{p1_concat_81908_comb[19]}}, p1_concat_81908_comb};
  assign p1_sum__1778_comb = {{5{p1_concat_81909_comb[19]}}, p1_concat_81909_comb};
  assign p1_sum__1779_comb = {{5{p1_concat_81910_comb[19]}}, p1_concat_81910_comb};
  assign p1_sum__1648_comb = {{5{p1_concat_81911_comb[19]}}, p1_concat_81911_comb};
  assign p1_sum__1649_comb = {{5{p1_concat_81912_comb[19]}}, p1_concat_81912_comb};
  assign p1_sum__1650_comb = {{5{p1_concat_81913_comb[19]}}, p1_concat_81913_comb};
  assign p1_sum__1651_comb = {{5{p1_concat_81914_comb[19]}}, p1_concat_81914_comb};
  assign p1_sum__1740_comb = {{5{p1_concat_81923_comb[19]}}, p1_concat_81923_comb};
  assign p1_sum__1741_comb = {{5{p1_concat_81924_comb[19]}}, p1_concat_81924_comb};
  assign p1_sum__1742_comb = {{5{p1_concat_81925_comb[19]}}, p1_concat_81925_comb};
  assign p1_sum__1743_comb = {{5{p1_concat_81926_comb[19]}}, p1_concat_81926_comb};
  assign p1_sum__1612_comb = {{5{p1_concat_81927_comb[19]}}, p1_concat_81927_comb};
  assign p1_sum__1613_comb = {{5{p1_concat_81928_comb[19]}}, p1_concat_81928_comb};
  assign p1_sum__1614_comb = {{5{p1_concat_81929_comb[19]}}, p1_concat_81929_comb};
  assign p1_sum__1615_comb = {{5{p1_concat_81930_comb[19]}}, p1_concat_81930_comb};
  assign p1_concat_82211_comb = {p1_add_81931_comb, p1_smul_81135_comb[0]};
  assign p1_concat_82212_comb = {p1_add_81933_comb, p1_smul_81137_comb[0]};
  assign p1_concat_82213_comb = {p1_add_81935_comb, p1_smul_81140_comb[0]};
  assign p1_concat_82214_comb = {p1_add_81937_comb, p1_smul_81142_comb[0]};
  assign p1_concat_82215_comb = {p1_add_81939_comb, p1_smul_81143_comb[0]};
  assign p1_concat_82216_comb = {p1_add_81941_comb, p1_smul_81145_comb[0]};
  assign p1_concat_82217_comb = {p1_add_81943_comb, p1_smul_81148_comb[0]};
  assign p1_concat_82218_comb = {p1_add_81945_comb, p1_smul_81150_comb[0]};
  assign p1_add_82219_comb = {{6{p1_add_81595_comb[17]}}, p1_add_81595_comb} + {{5{p1_bit_slice_81596_comb[18]}}, p1_bit_slice_81596_comb};
  assign p1_add_82221_comb = {{5{p1_bit_slice_81597_comb[18]}}, p1_bit_slice_81597_comb} + {{6{p1_add_81598_comb[17]}}, p1_add_81598_comb};
  assign p1_add_82223_comb = {{6{p1_add_81599_comb[17]}}, p1_add_81599_comb} + {{5{p1_bit_slice_81600_comb[18]}}, p1_bit_slice_81600_comb};
  assign p1_add_82225_comb = {{5{p1_bit_slice_81601_comb[18]}}, p1_bit_slice_81601_comb} + {{6{p1_add_81602_comb[17]}}, p1_add_81602_comb};
  assign p1_add_82235_comb = {{5{p1_bit_slice_81619_comb[18]}}, p1_bit_slice_81619_comb} + {{6{p1_add_81620_comb[17]}}, p1_add_81620_comb};
  assign p1_add_82237_comb = {{6{p1_add_81621_comb[17]}}, p1_add_81621_comb} + {{5{p1_bit_slice_81622_comb[18]}}, p1_bit_slice_81622_comb};
  assign p1_add_82239_comb = {{5{p1_bit_slice_81623_comb[18]}}, p1_bit_slice_81623_comb} + {{6{p1_add_81624_comb[17]}}, p1_add_81624_comb};
  assign p1_add_82241_comb = {{6{p1_add_81625_comb[17]}}, p1_add_81625_comb} + {{5{p1_bit_slice_81626_comb[18]}}, p1_bit_slice_81626_comb};
  assign p1_concat_82243_comb = {p1_add_81971_comb, p1_smul_81176_comb[0]};
  assign p1_concat_82244_comb = {p1_add_81973_comb, p1_smul_81177_comb[0]};
  assign p1_concat_82245_comb = {p1_add_81975_comb, p1_smul_81180_comb[0]};
  assign p1_concat_82246_comb = {p1_add_81977_comb, p1_smul_81181_comb[0]};
  assign p1_concat_82247_comb = {p1_add_81979_comb, p1_smul_81184_comb[0]};
  assign p1_concat_82248_comb = {p1_add_81981_comb, p1_smul_81185_comb[0]};
  assign p1_concat_82249_comb = {p1_add_81983_comb, p1_smul_81188_comb[0]};
  assign p1_concat_82250_comb = {p1_add_81985_comb, p1_smul_81189_comb[0]};
  assign p1_sum__1792_comb = {{5{p1_concat_81987_comb[19]}}, p1_concat_81987_comb};
  assign p1_sum__1793_comb = {{5{p1_concat_81988_comb[19]}}, p1_concat_81988_comb};
  assign p1_sum__1794_comb = {{5{p1_concat_81989_comb[19]}}, p1_concat_81989_comb};
  assign p1_sum__1795_comb = {{5{p1_concat_81990_comb[19]}}, p1_concat_81990_comb};
  assign p1_sum__1624_comb = {{5{p1_concat_81991_comb[19]}}, p1_concat_81991_comb};
  assign p1_sum__1625_comb = {{5{p1_concat_81992_comb[19]}}, p1_concat_81992_comb};
  assign p1_sum__1626_comb = {{5{p1_concat_81993_comb[19]}}, p1_concat_81993_comb};
  assign p1_sum__1627_comb = {{5{p1_concat_81994_comb[19]}}, p1_concat_81994_comb};
  assign p1_sum__1764_comb = {{5{p1_concat_82003_comb[19]}}, p1_concat_82003_comb};
  assign p1_sum__1765_comb = {{5{p1_concat_82004_comb[19]}}, p1_concat_82004_comb};
  assign p1_sum__1766_comb = {{5{p1_concat_82005_comb[19]}}, p1_concat_82005_comb};
  assign p1_sum__1767_comb = {{5{p1_concat_82006_comb[19]}}, p1_concat_82006_comb};
  assign p1_sum__1596_comb = {{5{p1_concat_82007_comb[19]}}, p1_concat_82007_comb};
  assign p1_sum__1597_comb = {{5{p1_concat_82008_comb[19]}}, p1_concat_82008_comb};
  assign p1_sum__1598_comb = {{5{p1_concat_82009_comb[19]}}, p1_concat_82009_comb};
  assign p1_sum__1599_comb = {{5{p1_concat_82010_comb[19]}}, p1_concat_82010_comb};
  assign p1_concat_82275_comb = {p1_add_82011_comb, p1_smul_81239_comb[0]};
  assign p1_concat_82276_comb = {p1_add_82013_comb, p1_smul_81241_comb[0]};
  assign p1_concat_82277_comb = {p1_add_82015_comb, p1_smul_81244_comb[0]};
  assign p1_concat_82278_comb = {p1_add_82017_comb, p1_smul_81246_comb[0]};
  assign p1_concat_82279_comb = {p1_add_82019_comb, p1_smul_81247_comb[0]};
  assign p1_concat_82280_comb = {p1_add_82021_comb, p1_smul_81249_comb[0]};
  assign p1_concat_82281_comb = {p1_add_82023_comb, p1_smul_81252_comb[0]};
  assign p1_concat_82282_comb = {p1_add_82025_comb, p1_smul_81254_comb[0]};
  assign p1_add_82283_comb = {{6{p1_add_81707_comb[17]}}, p1_add_81707_comb} + {{5{p1_bit_slice_81708_comb[18]}}, p1_bit_slice_81708_comb};
  assign p1_add_82285_comb = {{5{p1_bit_slice_81709_comb[18]}}, p1_bit_slice_81709_comb} + {{6{p1_add_81710_comb[17]}}, p1_add_81710_comb};
  assign p1_add_82287_comb = {{6{p1_add_81711_comb[17]}}, p1_add_81711_comb} + {{5{p1_bit_slice_81712_comb[18]}}, p1_bit_slice_81712_comb};
  assign p1_add_82289_comb = {{5{p1_bit_slice_81713_comb[18]}}, p1_bit_slice_81713_comb} + {{6{p1_add_81714_comb[17]}}, p1_add_81714_comb};
  assign p1_add_82451_comb = p1_add_82291_comb + p1_add_82292_comb;
  assign p1_add_82453_comb = p1_add_82293_comb + p1_add_82294_comb;
  assign p1_add_82455_comb = p1_add_82295_comb + p1_add_82296_comb;
  assign p1_add_82457_comb = p1_add_82297_comb + p1_add_82298_comb;
  assign p1_add_82515_comb = p1_add_82371_comb + p1_add_82372_comb;
  assign p1_add_82517_comb = p1_add_82373_comb + p1_add_82374_comb;
  assign p1_add_82547_comb = p1_add_82411_comb + p1_add_82412_comb;
  assign p1_add_82549_comb = p1_add_82413_comb + p1_add_82414_comb;
  assign p1_add_82595_comb = p1_sum__1118_comb + 25'h000_0001;
  assign p1_add_82596_comb = p1_sum__1111_comb + 25'h000_0001;
  assign p1_add_82597_comb = p1_sum__1104_comb + 25'h000_0001;
  assign p1_add_82598_comb = p1_sum__1097_comb + 25'h000_0001;
  assign p1_add_82619_comb = p1_sum__1124_comb + 25'h000_0001;
  assign p1_add_82620_comb = p1_sum__1091_comb + 25'h000_0001;
  assign p1_add_82635_comb = p1_sum__1129_comb + 25'h000_0001;
  assign p1_add_82636_comb = p1_sum__1086_comb + 25'h000_0001;
  assign p1_sum__1348_comb = {p1_add_82051_comb, p1_add_80851_comb[0]};
  assign p1_sum__1349_comb = {p1_add_82053_comb, p1_add_80856_comb[0]};
  assign p1_sum__1340_comb = {p1_add_82055_comb, p1_add_80857_comb[0]};
  assign p1_sum__1341_comb = {p1_add_82057_comb, p1_add_80862_comb[0]};
  assign p1_sum__1330_comb = {p1_add_82059_comb, p1_add_80863_comb[0]};
  assign p1_sum__1331_comb = {p1_add_82061_comb, p1_add_80868_comb[0]};
  assign p1_sum__1318_comb = {p1_add_82063_comb, p1_add_80869_comb[0]};
  assign p1_sum__1319_comb = {p1_add_82065_comb, p1_add_80874_comb[0]};
  assign p1_sum__1334_comb = p1_sum__1756_comb + p1_sum__1757_comb;
  assign p1_sum__1335_comb = p1_sum__1758_comb + p1_sum__1759_comb;
  assign p1_sum__1322_comb = p1_sum__1732_comb + p1_sum__1733_comb;
  assign p1_sum__1323_comb = p1_sum__1734_comb + p1_sum__1735_comb;
  assign p1_sum__1308_comb = p1_sum__1704_comb + p1_sum__1705_comb;
  assign p1_sum__1309_comb = p1_sum__1706_comb + p1_sum__1707_comb;
  assign p1_sum__1294_comb = p1_sum__1676_comb + p1_sum__1677_comb;
  assign p1_sum__1295_comb = p1_sum__1678_comb + p1_sum__1679_comb;
  assign p1_sum__1312_comb = p1_sum__1712_comb + p1_sum__1713_comb;
  assign p1_sum__1313_comb = p1_sum__1714_comb + p1_sum__1715_comb;
  assign p1_sum__1298_comb = p1_sum__1684_comb + p1_sum__1685_comb;
  assign p1_sum__1299_comb = p1_sum__1686_comb + p1_sum__1687_comb;
  assign p1_sum__1284_comb = p1_sum__1656_comb + p1_sum__1657_comb;
  assign p1_sum__1285_comb = p1_sum__1658_comb + p1_sum__1659_comb;
  assign p1_sum__1272_comb = p1_sum__1632_comb + p1_sum__1633_comb;
  assign p1_sum__1273_comb = p1_sum__1634_comb + p1_sum__1635_comb;
  assign p1_sum__1288_comb = {p1_add_82147_comb, p1_add_81037_comb[0]};
  assign p1_sum__1289_comb = {p1_add_82149_comb, p1_add_81038_comb[0]};
  assign p1_sum__1276_comb = {p1_add_82151_comb, p1_add_81043_comb[0]};
  assign p1_sum__1277_comb = {p1_add_82153_comb, p1_add_81044_comb[0]};
  assign p1_sum__1266_comb = {p1_add_82155_comb, p1_add_81049_comb[0]};
  assign p1_sum__1267_comb = {p1_add_82157_comb, p1_add_81050_comb[0]};
  assign p1_sum__1258_comb = {p1_add_82159_comb, p1_add_81055_comb[0]};
  assign p1_sum__1259_comb = {p1_add_82161_comb, p1_add_81056_comb[0]};
  assign p1_sum__1354_comb = {p1_add_82171_comb, p1_add_81059_comb[0]};
  assign p1_sum__1355_comb = {p1_add_82173_comb, p1_add_81064_comb[0]};
  assign p1_sum__1304_comb = {p1_add_82175_comb, p1_add_81065_comb[0]};
  assign p1_sum__1305_comb = {p1_add_82177_comb, p1_add_81070_comb[0]};
  assign p1_sum__1344_comb = p1_sum__1776_comb + p1_sum__1777_comb;
  assign p1_sum__1345_comb = p1_sum__1778_comb + p1_sum__1779_comb;
  assign p1_sum__1280_comb = p1_sum__1648_comb + p1_sum__1649_comb;
  assign p1_sum__1281_comb = p1_sum__1650_comb + p1_sum__1651_comb;
  assign p1_sum__1326_comb = p1_sum__1740_comb + p1_sum__1741_comb;
  assign p1_sum__1327_comb = p1_sum__1742_comb + p1_sum__1743_comb;
  assign p1_sum__1262_comb = p1_sum__1612_comb + p1_sum__1613_comb;
  assign p1_sum__1263_comb = p1_sum__1614_comb + p1_sum__1615_comb;
  assign p1_sum__1302_comb = {p1_add_82219_comb, p1_add_81153_comb[0]};
  assign p1_sum__1303_comb = {p1_add_82221_comb, p1_add_81154_comb[0]};
  assign p1_sum__1252_comb = {p1_add_82223_comb, p1_add_81159_comb[0]};
  assign p1_sum__1253_comb = {p1_add_82225_comb, p1_add_81160_comb[0]};
  assign p1_sum__1358_comb = {p1_add_82235_comb, p1_add_81163_comb[0]};
  assign p1_sum__1359_comb = {p1_add_82237_comb, p1_add_81168_comb[0]};
  assign p1_sum__1290_comb = {p1_add_82239_comb, p1_add_81169_comb[0]};
  assign p1_sum__1291_comb = {p1_add_82241_comb, p1_add_81174_comb[0]};
  assign p1_sum__1352_comb = p1_sum__1792_comb + p1_sum__1793_comb;
  assign p1_sum__1353_comb = p1_sum__1794_comb + p1_sum__1795_comb;
  assign p1_sum__1268_comb = p1_sum__1624_comb + p1_sum__1625_comb;
  assign p1_sum__1269_comb = p1_sum__1626_comb + p1_sum__1627_comb;
  assign p1_sum__1338_comb = p1_sum__1764_comb + p1_sum__1765_comb;
  assign p1_sum__1339_comb = p1_sum__1766_comb + p1_sum__1767_comb;
  assign p1_sum__1254_comb = p1_sum__1596_comb + p1_sum__1597_comb;
  assign p1_sum__1255_comb = p1_sum__1598_comb + p1_sum__1599_comb;
  assign p1_sum__1316_comb = {p1_add_82283_comb, p1_add_81257_comb[0]};
  assign p1_sum__1317_comb = {p1_add_82285_comb, p1_add_81258_comb[0]};
  assign p1_sum__1248_comb = {p1_add_82287_comb, p1_add_81263_comb[0]};
  assign p1_sum__1249_comb = {p1_add_82289_comb, p1_add_81264_comb[0]};
  assign p1_umul_28108_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_82451_comb, 7'h5b);
  assign p1_umul_28110_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_82453_comb, 7'h5b);
  assign p1_umul_28112_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_82455_comb, 7'h5b);
  assign p1_umul_28114_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_82457_comb, 7'h5b);
  assign p1_umul_28106_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_82515_comb, 7'h5b);
  assign p1_umul_28116_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_82517_comb, 7'h5b);
  assign p1_umul_28104_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_82547_comb, 7'h5b);
  assign p1_umul_28118_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_82549_comb, 7'h5b);
  assign p1_bit_slice_82659_comb = p1_add_82595_comb[24:8];
  assign p1_bit_slice_82660_comb = p1_add_82596_comb[24:8];
  assign p1_bit_slice_82661_comb = p1_add_82597_comb[24:8];
  assign p1_bit_slice_82662_comb = p1_add_82598_comb[24:8];
  assign p1_bit_slice_82683_comb = p1_add_82619_comb[24:8];
  assign p1_bit_slice_82684_comb = p1_add_82620_comb[24:8];
  assign p1_bit_slice_82699_comb = p1_add_82635_comb[24:8];
  assign p1_bit_slice_82700_comb = p1_add_82636_comb[24:8];
  assign p1_sum__1130_comb = p1_sum__1348_comb + p1_sum__1349_comb;
  assign p1_sum__1126_comb = p1_sum__1340_comb + p1_sum__1341_comb;
  assign p1_sum__1121_comb = p1_sum__1330_comb + p1_sum__1331_comb;
  assign p1_sum__1115_comb = p1_sum__1318_comb + p1_sum__1319_comb;
  assign p1_add_82467_comb = {{5{p1_concat_82067_comb[18]}}, p1_concat_82067_comb} + {{5{p1_concat_82068_comb[18]}}, p1_concat_82068_comb};
  assign p1_add_82468_comb = {{5{p1_concat_82069_comb[18]}}, p1_concat_82069_comb} + {{5{p1_concat_82070_comb[18]}}, p1_concat_82070_comb};
  assign p1_add_82469_comb = {{5{p1_concat_82071_comb[18]}}, p1_concat_82071_comb} + {{5{p1_concat_82072_comb[18]}}, p1_concat_82072_comb};
  assign p1_add_82470_comb = {{5{p1_concat_82073_comb[18]}}, p1_concat_82073_comb} + {{5{p1_concat_82074_comb[18]}}, p1_concat_82074_comb};
  assign p1_add_82471_comb = {{5{p1_concat_82075_comb[18]}}, p1_concat_82075_comb} + {{5{p1_concat_82076_comb[18]}}, p1_concat_82076_comb};
  assign p1_add_82472_comb = {{5{p1_concat_82077_comb[18]}}, p1_concat_82077_comb} + {{5{p1_concat_82078_comb[18]}}, p1_concat_82078_comb};
  assign p1_add_82473_comb = {{5{p1_concat_82079_comb[18]}}, p1_concat_82079_comb} + {{5{p1_concat_82080_comb[18]}}, p1_concat_82080_comb};
  assign p1_add_82474_comb = {{5{p1_concat_82081_comb[18]}}, p1_concat_82081_comb} + {{5{p1_concat_82082_comb[18]}}, p1_concat_82082_comb};
  assign p1_sum__1123_comb = p1_sum__1334_comb + p1_sum__1335_comb;
  assign p1_sum__1117_comb = p1_sum__1322_comb + p1_sum__1323_comb;
  assign p1_sum__1110_comb = p1_sum__1308_comb + p1_sum__1309_comb;
  assign p1_sum__1103_comb = p1_sum__1294_comb + p1_sum__1295_comb;
  assign p1_sum__1112_comb = p1_sum__1312_comb + p1_sum__1313_comb;
  assign p1_sum__1105_comb = p1_sum__1298_comb + p1_sum__1299_comb;
  assign p1_sum__1098_comb = p1_sum__1284_comb + p1_sum__1285_comb;
  assign p1_sum__1092_comb = p1_sum__1272_comb + p1_sum__1273_comb;
  assign p1_add_82499_comb = {{5{p1_concat_82131_comb[18]}}, p1_concat_82131_comb} + {{5{p1_concat_82132_comb[18]}}, p1_concat_82132_comb};
  assign p1_add_82500_comb = {{5{p1_concat_82133_comb[18]}}, p1_concat_82133_comb} + {{5{p1_concat_82134_comb[18]}}, p1_concat_82134_comb};
  assign p1_add_82501_comb = {{5{p1_concat_82135_comb[18]}}, p1_concat_82135_comb} + {{5{p1_concat_82136_comb[18]}}, p1_concat_82136_comb};
  assign p1_add_82502_comb = {{5{p1_concat_82137_comb[18]}}, p1_concat_82137_comb} + {{5{p1_concat_82138_comb[18]}}, p1_concat_82138_comb};
  assign p1_add_82503_comb = {{5{p1_concat_82139_comb[18]}}, p1_concat_82139_comb} + {{5{p1_concat_82140_comb[18]}}, p1_concat_82140_comb};
  assign p1_add_82504_comb = {{5{p1_concat_82141_comb[18]}}, p1_concat_82141_comb} + {{5{p1_concat_82142_comb[18]}}, p1_concat_82142_comb};
  assign p1_add_82505_comb = {{5{p1_concat_82143_comb[18]}}, p1_concat_82143_comb} + {{5{p1_concat_82144_comb[18]}}, p1_concat_82144_comb};
  assign p1_add_82506_comb = {{5{p1_concat_82145_comb[18]}}, p1_concat_82145_comb} + {{5{p1_concat_82146_comb[18]}}, p1_concat_82146_comb};
  assign p1_sum__1100_comb = p1_sum__1288_comb + p1_sum__1289_comb;
  assign p1_sum__1094_comb = p1_sum__1276_comb + p1_sum__1277_comb;
  assign p1_sum__1089_comb = p1_sum__1266_comb + p1_sum__1267_comb;
  assign p1_sum__1085_comb = p1_sum__1258_comb + p1_sum__1259_comb;
  assign p1_sum__1133_comb = p1_sum__1354_comb + p1_sum__1355_comb;
  assign p1_sum__1108_comb = p1_sum__1304_comb + p1_sum__1305_comb;
  assign p1_add_82523_comb = {{5{p1_concat_82179_comb[18]}}, p1_concat_82179_comb} + {{5{p1_concat_82180_comb[18]}}, p1_concat_82180_comb};
  assign p1_add_82524_comb = {{5{p1_concat_82181_comb[18]}}, p1_concat_82181_comb} + {{5{p1_concat_82182_comb[18]}}, p1_concat_82182_comb};
  assign p1_add_82525_comb = {{5{p1_concat_82183_comb[18]}}, p1_concat_82183_comb} + {{5{p1_concat_82184_comb[18]}}, p1_concat_82184_comb};
  assign p1_add_82526_comb = {{5{p1_concat_82185_comb[18]}}, p1_concat_82185_comb} + {{5{p1_concat_82186_comb[18]}}, p1_concat_82186_comb};
  assign p1_sum__1128_comb = p1_sum__1344_comb + p1_sum__1345_comb;
  assign p1_sum__1096_comb = p1_sum__1280_comb + p1_sum__1281_comb;
  assign p1_sum__1119_comb = p1_sum__1326_comb + p1_sum__1327_comb;
  assign p1_sum__1087_comb = p1_sum__1262_comb + p1_sum__1263_comb;
  assign p1_add_82539_comb = {{5{p1_concat_82211_comb[18]}}, p1_concat_82211_comb} + {{5{p1_concat_82212_comb[18]}}, p1_concat_82212_comb};
  assign p1_add_82540_comb = {{5{p1_concat_82213_comb[18]}}, p1_concat_82213_comb} + {{5{p1_concat_82214_comb[18]}}, p1_concat_82214_comb};
  assign p1_add_82541_comb = {{5{p1_concat_82215_comb[18]}}, p1_concat_82215_comb} + {{5{p1_concat_82216_comb[18]}}, p1_concat_82216_comb};
  assign p1_add_82542_comb = {{5{p1_concat_82217_comb[18]}}, p1_concat_82217_comb} + {{5{p1_concat_82218_comb[18]}}, p1_concat_82218_comb};
  assign p1_sum__1107_comb = p1_sum__1302_comb + p1_sum__1303_comb;
  assign p1_sum__1082_comb = p1_sum__1252_comb + p1_sum__1253_comb;
  assign p1_sum__1135_comb = p1_sum__1358_comb + p1_sum__1359_comb;
  assign p1_sum__1101_comb = p1_sum__1290_comb + p1_sum__1291_comb;
  assign p1_add_82555_comb = {{5{p1_concat_82243_comb[18]}}, p1_concat_82243_comb} + {{5{p1_concat_82244_comb[18]}}, p1_concat_82244_comb};
  assign p1_add_82556_comb = {{5{p1_concat_82245_comb[18]}}, p1_concat_82245_comb} + {{5{p1_concat_82246_comb[18]}}, p1_concat_82246_comb};
  assign p1_add_82557_comb = {{5{p1_concat_82247_comb[18]}}, p1_concat_82247_comb} + {{5{p1_concat_82248_comb[18]}}, p1_concat_82248_comb};
  assign p1_add_82558_comb = {{5{p1_concat_82249_comb[18]}}, p1_concat_82249_comb} + {{5{p1_concat_82250_comb[18]}}, p1_concat_82250_comb};
  assign p1_sum__1132_comb = p1_sum__1352_comb + p1_sum__1353_comb;
  assign p1_sum__1090_comb = p1_sum__1268_comb + p1_sum__1269_comb;
  assign p1_sum__1125_comb = p1_sum__1338_comb + p1_sum__1339_comb;
  assign p1_sum__1083_comb = p1_sum__1254_comb + p1_sum__1255_comb;
  assign p1_add_82571_comb = {{5{p1_concat_82275_comb[18]}}, p1_concat_82275_comb} + {{5{p1_concat_82276_comb[18]}}, p1_concat_82276_comb};
  assign p1_add_82572_comb = {{5{p1_concat_82277_comb[18]}}, p1_concat_82277_comb} + {{5{p1_concat_82278_comb[18]}}, p1_concat_82278_comb};
  assign p1_add_82573_comb = {{5{p1_concat_82279_comb[18]}}, p1_concat_82279_comb} + {{5{p1_concat_82280_comb[18]}}, p1_concat_82280_comb};
  assign p1_add_82574_comb = {{5{p1_concat_82281_comb[18]}}, p1_concat_82281_comb} + {{5{p1_concat_82282_comb[18]}}, p1_concat_82282_comb};
  assign p1_sum__1114_comb = p1_sum__1316_comb + p1_sum__1317_comb;
  assign p1_sum__1080_comb = p1_sum__1248_comb + p1_sum__1249_comb;
  assign p1_bit_slice_82643_comb = p1_umul_28108_NarrowedMult__comb[23:7];
  assign p1_bit_slice_82644_comb = p1_umul_28110_NarrowedMult__comb[23:7];
  assign p1_bit_slice_82645_comb = p1_umul_28112_NarrowedMult__comb[23:7];
  assign p1_bit_slice_82646_comb = p1_umul_28114_NarrowedMult__comb[23:7];
  assign p1_bit_slice_82675_comb = p1_umul_28106_NarrowedMult__comb[23:7];
  assign p1_bit_slice_82676_comb = p1_umul_28116_NarrowedMult__comb[23:7];
  assign p1_bit_slice_82691_comb = p1_umul_28104_NarrowedMult__comb[23:7];
  assign p1_bit_slice_82692_comb = p1_umul_28118_NarrowedMult__comb[23:7];
  assign p1_add_82583_comb = p1_sum__1130_comb + 25'h000_0001;
  assign p1_add_82584_comb = p1_sum__1126_comb + 25'h000_0001;
  assign p1_add_82585_comb = p1_sum__1121_comb + 25'h000_0001;
  assign p1_add_82586_comb = p1_sum__1115_comb + 25'h000_0001;
  assign p1_add_82587_comb = p1_add_82467_comb + p1_add_82468_comb;
  assign p1_add_82588_comb = p1_add_82469_comb + p1_add_82470_comb;
  assign p1_add_82589_comb = p1_add_82471_comb + p1_add_82472_comb;
  assign p1_add_82590_comb = p1_add_82473_comb + p1_add_82474_comb;
  assign p1_add_82591_comb = p1_sum__1123_comb + 25'h000_0001;
  assign p1_add_82592_comb = p1_sum__1117_comb + 25'h000_0001;
  assign p1_add_82593_comb = p1_sum__1110_comb + 25'h000_0001;
  assign p1_add_82594_comb = p1_sum__1103_comb + 25'h000_0001;
  assign p1_add_82599_comb = p1_sum__1112_comb + 25'h000_0001;
  assign p1_add_82600_comb = p1_sum__1105_comb + 25'h000_0001;
  assign p1_add_82601_comb = p1_sum__1098_comb + 25'h000_0001;
  assign p1_add_82602_comb = p1_sum__1092_comb + 25'h000_0001;
  assign p1_add_82603_comb = p1_add_82499_comb + p1_add_82500_comb;
  assign p1_add_82604_comb = p1_add_82501_comb + p1_add_82502_comb;
  assign p1_add_82605_comb = p1_add_82503_comb + p1_add_82504_comb;
  assign p1_add_82606_comb = p1_add_82505_comb + p1_add_82506_comb;
  assign p1_add_82607_comb = p1_sum__1100_comb + 25'h000_0001;
  assign p1_add_82608_comb = p1_sum__1094_comb + 25'h000_0001;
  assign p1_add_82609_comb = p1_sum__1089_comb + 25'h000_0001;
  assign p1_add_82610_comb = p1_sum__1085_comb + 25'h000_0001;
  assign p1_add_82613_comb = p1_sum__1133_comb + 25'h000_0001;
  assign p1_add_82614_comb = p1_sum__1108_comb + 25'h000_0001;
  assign p1_add_82615_comb = p1_add_82523_comb + p1_add_82524_comb;
  assign p1_add_82616_comb = p1_add_82525_comb + p1_add_82526_comb;
  assign p1_add_82617_comb = p1_sum__1128_comb + 25'h000_0001;
  assign p1_add_82618_comb = p1_sum__1096_comb + 25'h000_0001;
  assign p1_add_82621_comb = p1_sum__1119_comb + 25'h000_0001;
  assign p1_add_82622_comb = p1_sum__1087_comb + 25'h000_0001;
  assign p1_add_82623_comb = p1_add_82539_comb + p1_add_82540_comb;
  assign p1_add_82624_comb = p1_add_82541_comb + p1_add_82542_comb;
  assign p1_add_82625_comb = p1_sum__1107_comb + 25'h000_0001;
  assign p1_add_82626_comb = p1_sum__1082_comb + 25'h000_0001;
  assign p1_add_82629_comb = p1_sum__1135_comb + 25'h000_0001;
  assign p1_add_82630_comb = p1_sum__1101_comb + 25'h000_0001;
  assign p1_add_82631_comb = p1_add_82555_comb + p1_add_82556_comb;
  assign p1_add_82632_comb = p1_add_82557_comb + p1_add_82558_comb;
  assign p1_add_82633_comb = p1_sum__1132_comb + 25'h000_0001;
  assign p1_add_82634_comb = p1_sum__1090_comb + 25'h000_0001;
  assign p1_add_82637_comb = p1_sum__1125_comb + 25'h000_0001;
  assign p1_add_82638_comb = p1_sum__1083_comb + 25'h000_0001;
  assign p1_add_82639_comb = p1_add_82571_comb + p1_add_82572_comb;
  assign p1_add_82640_comb = p1_add_82573_comb + p1_add_82574_comb;
  assign p1_add_82641_comb = p1_sum__1114_comb + 25'h000_0001;
  assign p1_add_82642_comb = p1_sum__1080_comb + 25'h000_0001;
  assign p1_add_82851_comb = {{1{p1_bit_slice_82659_comb[16]}}, p1_bit_slice_82659_comb} + 18'h0_0001;
  assign p1_add_82852_comb = {{1{p1_bit_slice_82660_comb[16]}}, p1_bit_slice_82660_comb} + 18'h0_0001;
  assign p1_add_82853_comb = {{1{p1_bit_slice_82661_comb[16]}}, p1_bit_slice_82661_comb} + 18'h0_0001;
  assign p1_add_82854_comb = {{1{p1_bit_slice_82662_comb[16]}}, p1_bit_slice_82662_comb} + 18'h0_0001;
  assign p1_add_82875_comb = {{1{p1_bit_slice_82683_comb[16]}}, p1_bit_slice_82683_comb} + 18'h0_0001;
  assign p1_add_82876_comb = {{1{p1_bit_slice_82684_comb[16]}}, p1_bit_slice_82684_comb} + 18'h0_0001;
  assign p1_add_82891_comb = {{1{p1_bit_slice_82699_comb[16]}}, p1_bit_slice_82699_comb} + 18'h0_0001;
  assign p1_add_82892_comb = {{1{p1_bit_slice_82700_comb[16]}}, p1_bit_slice_82700_comb} + 18'h0_0001;
  assign p1_bit_slice_82647_comb = p1_add_82583_comb[24:8];
  assign p1_bit_slice_82648_comb = p1_add_82584_comb[24:8];
  assign p1_bit_slice_82649_comb = p1_add_82585_comb[24:8];
  assign p1_bit_slice_82650_comb = p1_add_82586_comb[24:8];
  assign p1_bit_slice_82651_comb = p1_add_82587_comb[23:7];
  assign p1_bit_slice_82652_comb = p1_add_82588_comb[23:7];
  assign p1_bit_slice_82653_comb = p1_add_82589_comb[23:7];
  assign p1_bit_slice_82654_comb = p1_add_82590_comb[23:7];
  assign p1_bit_slice_82655_comb = p1_add_82591_comb[24:8];
  assign p1_bit_slice_82656_comb = p1_add_82592_comb[24:8];
  assign p1_bit_slice_82657_comb = p1_add_82593_comb[24:8];
  assign p1_bit_slice_82658_comb = p1_add_82594_comb[24:8];
  assign p1_bit_slice_82663_comb = p1_add_82599_comb[24:8];
  assign p1_bit_slice_82664_comb = p1_add_82600_comb[24:8];
  assign p1_bit_slice_82665_comb = p1_add_82601_comb[24:8];
  assign p1_bit_slice_82666_comb = p1_add_82602_comb[24:8];
  assign p1_bit_slice_82667_comb = p1_add_82603_comb[23:7];
  assign p1_bit_slice_82668_comb = p1_add_82604_comb[23:7];
  assign p1_bit_slice_82669_comb = p1_add_82605_comb[23:7];
  assign p1_bit_slice_82670_comb = p1_add_82606_comb[23:7];
  assign p1_bit_slice_82671_comb = p1_add_82607_comb[24:8];
  assign p1_bit_slice_82672_comb = p1_add_82608_comb[24:8];
  assign p1_bit_slice_82673_comb = p1_add_82609_comb[24:8];
  assign p1_bit_slice_82674_comb = p1_add_82610_comb[24:8];
  assign p1_bit_slice_82677_comb = p1_add_82613_comb[24:8];
  assign p1_bit_slice_82678_comb = p1_add_82614_comb[24:8];
  assign p1_bit_slice_82679_comb = p1_add_82615_comb[23:7];
  assign p1_bit_slice_82680_comb = p1_add_82616_comb[23:7];
  assign p1_bit_slice_82681_comb = p1_add_82617_comb[24:8];
  assign p1_bit_slice_82682_comb = p1_add_82618_comb[24:8];
  assign p1_bit_slice_82685_comb = p1_add_82621_comb[24:8];
  assign p1_bit_slice_82686_comb = p1_add_82622_comb[24:8];
  assign p1_bit_slice_82687_comb = p1_add_82623_comb[23:7];
  assign p1_bit_slice_82688_comb = p1_add_82624_comb[23:7];
  assign p1_bit_slice_82689_comb = p1_add_82625_comb[24:8];
  assign p1_bit_slice_82690_comb = p1_add_82626_comb[24:8];
  assign p1_bit_slice_82693_comb = p1_add_82629_comb[24:8];
  assign p1_bit_slice_82694_comb = p1_add_82630_comb[24:8];
  assign p1_bit_slice_82695_comb = p1_add_82631_comb[23:7];
  assign p1_bit_slice_82696_comb = p1_add_82632_comb[23:7];
  assign p1_bit_slice_82697_comb = p1_add_82633_comb[24:8];
  assign p1_bit_slice_82698_comb = p1_add_82634_comb[24:8];
  assign p1_bit_slice_82701_comb = p1_add_82637_comb[24:8];
  assign p1_bit_slice_82702_comb = p1_add_82638_comb[24:8];
  assign p1_bit_slice_82703_comb = p1_add_82639_comb[23:7];
  assign p1_bit_slice_82704_comb = p1_add_82640_comb[23:7];
  assign p1_bit_slice_82705_comb = p1_add_82641_comb[24:8];
  assign p1_bit_slice_82706_comb = p1_add_82642_comb[24:8];
  assign p1_add_82835_comb = {{1{p1_bit_slice_82643_comb[16]}}, p1_bit_slice_82643_comb} + 18'h0_0001;
  assign p1_add_82836_comb = {{1{p1_bit_slice_82644_comb[16]}}, p1_bit_slice_82644_comb} + 18'h0_0001;
  assign p1_add_82837_comb = {{1{p1_bit_slice_82645_comb[16]}}, p1_bit_slice_82645_comb} + 18'h0_0001;
  assign p1_add_82838_comb = {{1{p1_bit_slice_82646_comb[16]}}, p1_bit_slice_82646_comb} + 18'h0_0001;
  assign p1_add_82867_comb = {{1{p1_bit_slice_82675_comb[16]}}, p1_bit_slice_82675_comb} + 18'h0_0001;
  assign p1_add_82868_comb = {{1{p1_bit_slice_82676_comb[16]}}, p1_bit_slice_82676_comb} + 18'h0_0001;
  assign p1_add_82883_comb = {{1{p1_bit_slice_82691_comb[16]}}, p1_bit_slice_82691_comb} + 18'h0_0001;
  assign p1_add_82884_comb = {{1{p1_bit_slice_82692_comb[16]}}, p1_bit_slice_82692_comb} + 18'h0_0001;
  assign p1_bit_slice_82903_comb = p1_add_82851_comb[17:8];
  assign p1_bit_slice_82904_comb = p1_add_82852_comb[17:8];
  assign p1_bit_slice_82905_comb = p1_add_82853_comb[17:8];
  assign p1_bit_slice_82906_comb = p1_add_82854_comb[17:8];
  assign p1_bit_slice_82909_comb = p1_add_82875_comb[17:8];
  assign p1_bit_slice_82910_comb = p1_add_82876_comb[17:8];
  assign p1_bit_slice_82913_comb = p1_add_82891_comb[17:8];
  assign p1_bit_slice_82914_comb = p1_add_82892_comb[17:8];
  assign p1_bit_slice_82899_comb = p1_add_82835_comb[17:8];
  assign p1_bit_slice_82900_comb = p1_add_82836_comb[17:8];
  assign p1_bit_slice_82901_comb = p1_add_82837_comb[17:8];
  assign p1_bit_slice_82902_comb = p1_add_82838_comb[17:8];
  assign p1_bit_slice_82907_comb = p1_add_82867_comb[17:8];
  assign p1_bit_slice_82908_comb = p1_add_82868_comb[17:8];
  assign p1_bit_slice_82911_comb = p1_add_82883_comb[17:8];
  assign p1_bit_slice_82912_comb = p1_add_82884_comb[17:8];
  assign p1_add_82839_comb = {{1{p1_bit_slice_82647_comb[16]}}, p1_bit_slice_82647_comb} + 18'h0_0001;
  assign p1_add_82840_comb = {{1{p1_bit_slice_82648_comb[16]}}, p1_bit_slice_82648_comb} + 18'h0_0001;
  assign p1_add_82841_comb = {{1{p1_bit_slice_82649_comb[16]}}, p1_bit_slice_82649_comb} + 18'h0_0001;
  assign p1_add_82842_comb = {{1{p1_bit_slice_82650_comb[16]}}, p1_bit_slice_82650_comb} + 18'h0_0001;
  assign p1_add_82843_comb = {{1{p1_bit_slice_82651_comb[16]}}, p1_bit_slice_82651_comb} + 18'h0_0001;
  assign p1_add_82844_comb = {{1{p1_bit_slice_82652_comb[16]}}, p1_bit_slice_82652_comb} + 18'h0_0001;
  assign p1_add_82845_comb = {{1{p1_bit_slice_82653_comb[16]}}, p1_bit_slice_82653_comb} + 18'h0_0001;
  assign p1_add_82846_comb = {{1{p1_bit_slice_82654_comb[16]}}, p1_bit_slice_82654_comb} + 18'h0_0001;
  assign p1_add_82847_comb = {{1{p1_bit_slice_82655_comb[16]}}, p1_bit_slice_82655_comb} + 18'h0_0001;
  assign p1_add_82848_comb = {{1{p1_bit_slice_82656_comb[16]}}, p1_bit_slice_82656_comb} + 18'h0_0001;
  assign p1_add_82849_comb = {{1{p1_bit_slice_82657_comb[16]}}, p1_bit_slice_82657_comb} + 18'h0_0001;
  assign p1_add_82850_comb = {{1{p1_bit_slice_82658_comb[16]}}, p1_bit_slice_82658_comb} + 18'h0_0001;
  assign p1_add_82855_comb = {{1{p1_bit_slice_82663_comb[16]}}, p1_bit_slice_82663_comb} + 18'h0_0001;
  assign p1_add_82856_comb = {{1{p1_bit_slice_82664_comb[16]}}, p1_bit_slice_82664_comb} + 18'h0_0001;
  assign p1_add_82857_comb = {{1{p1_bit_slice_82665_comb[16]}}, p1_bit_slice_82665_comb} + 18'h0_0001;
  assign p1_add_82858_comb = {{1{p1_bit_slice_82666_comb[16]}}, p1_bit_slice_82666_comb} + 18'h0_0001;
  assign p1_add_82859_comb = {{1{p1_bit_slice_82667_comb[16]}}, p1_bit_slice_82667_comb} + 18'h0_0001;
  assign p1_add_82860_comb = {{1{p1_bit_slice_82668_comb[16]}}, p1_bit_slice_82668_comb} + 18'h0_0001;
  assign p1_add_82861_comb = {{1{p1_bit_slice_82669_comb[16]}}, p1_bit_slice_82669_comb} + 18'h0_0001;
  assign p1_add_82862_comb = {{1{p1_bit_slice_82670_comb[16]}}, p1_bit_slice_82670_comb} + 18'h0_0001;
  assign p1_add_82863_comb = {{1{p1_bit_slice_82671_comb[16]}}, p1_bit_slice_82671_comb} + 18'h0_0001;
  assign p1_add_82864_comb = {{1{p1_bit_slice_82672_comb[16]}}, p1_bit_slice_82672_comb} + 18'h0_0001;
  assign p1_add_82865_comb = {{1{p1_bit_slice_82673_comb[16]}}, p1_bit_slice_82673_comb} + 18'h0_0001;
  assign p1_add_82866_comb = {{1{p1_bit_slice_82674_comb[16]}}, p1_bit_slice_82674_comb} + 18'h0_0001;
  assign p1_add_82869_comb = {{1{p1_bit_slice_82677_comb[16]}}, p1_bit_slice_82677_comb} + 18'h0_0001;
  assign p1_add_82870_comb = {{1{p1_bit_slice_82678_comb[16]}}, p1_bit_slice_82678_comb} + 18'h0_0001;
  assign p1_add_82871_comb = {{1{p1_bit_slice_82679_comb[16]}}, p1_bit_slice_82679_comb} + 18'h0_0001;
  assign p1_add_82872_comb = {{1{p1_bit_slice_82680_comb[16]}}, p1_bit_slice_82680_comb} + 18'h0_0001;
  assign p1_add_82873_comb = {{1{p1_bit_slice_82681_comb[16]}}, p1_bit_slice_82681_comb} + 18'h0_0001;
  assign p1_add_82874_comb = {{1{p1_bit_slice_82682_comb[16]}}, p1_bit_slice_82682_comb} + 18'h0_0001;
  assign p1_add_82877_comb = {{1{p1_bit_slice_82685_comb[16]}}, p1_bit_slice_82685_comb} + 18'h0_0001;
  assign p1_add_82878_comb = {{1{p1_bit_slice_82686_comb[16]}}, p1_bit_slice_82686_comb} + 18'h0_0001;
  assign p1_add_82879_comb = {{1{p1_bit_slice_82687_comb[16]}}, p1_bit_slice_82687_comb} + 18'h0_0001;
  assign p1_add_82880_comb = {{1{p1_bit_slice_82688_comb[16]}}, p1_bit_slice_82688_comb} + 18'h0_0001;
  assign p1_add_82881_comb = {{1{p1_bit_slice_82689_comb[16]}}, p1_bit_slice_82689_comb} + 18'h0_0001;
  assign p1_add_82882_comb = {{1{p1_bit_slice_82690_comb[16]}}, p1_bit_slice_82690_comb} + 18'h0_0001;
  assign p1_add_82885_comb = {{1{p1_bit_slice_82693_comb[16]}}, p1_bit_slice_82693_comb} + 18'h0_0001;
  assign p1_add_82886_comb = {{1{p1_bit_slice_82694_comb[16]}}, p1_bit_slice_82694_comb} + 18'h0_0001;
  assign p1_add_82887_comb = {{1{p1_bit_slice_82695_comb[16]}}, p1_bit_slice_82695_comb} + 18'h0_0001;
  assign p1_add_82888_comb = {{1{p1_bit_slice_82696_comb[16]}}, p1_bit_slice_82696_comb} + 18'h0_0001;
  assign p1_add_82889_comb = {{1{p1_bit_slice_82697_comb[16]}}, p1_bit_slice_82697_comb} + 18'h0_0001;
  assign p1_add_82890_comb = {{1{p1_bit_slice_82698_comb[16]}}, p1_bit_slice_82698_comb} + 18'h0_0001;
  assign p1_add_82893_comb = {{1{p1_bit_slice_82701_comb[16]}}, p1_bit_slice_82701_comb} + 18'h0_0001;
  assign p1_add_82894_comb = {{1{p1_bit_slice_82702_comb[16]}}, p1_bit_slice_82702_comb} + 18'h0_0001;
  assign p1_add_82895_comb = {{1{p1_bit_slice_82703_comb[16]}}, p1_bit_slice_82703_comb} + 18'h0_0001;
  assign p1_add_82896_comb = {{1{p1_bit_slice_82704_comb[16]}}, p1_bit_slice_82704_comb} + 18'h0_0001;
  assign p1_add_82897_comb = {{1{p1_bit_slice_82705_comb[16]}}, p1_bit_slice_82705_comb} + 18'h0_0001;
  assign p1_add_82898_comb = {{1{p1_bit_slice_82706_comb[16]}}, p1_bit_slice_82706_comb} + 18'h0_0001;
  assign p1_sign_ext_82915_comb = {{1{p1_bit_slice_82899_comb[9]}}, p1_bit_slice_82899_comb};
  assign p1_sign_ext_82916_comb = {{1{p1_bit_slice_82900_comb[9]}}, p1_bit_slice_82900_comb};
  assign p1_sign_ext_82917_comb = {{1{p1_bit_slice_82901_comb[9]}}, p1_bit_slice_82901_comb};
  assign p1_sign_ext_82918_comb = {{1{p1_bit_slice_82902_comb[9]}}, p1_bit_slice_82902_comb};
  assign p1_sign_ext_82927_comb = {{1{p1_bit_slice_82907_comb[9]}}, p1_bit_slice_82907_comb};
  assign p1_sign_ext_82928_comb = {{1{p1_bit_slice_82908_comb[9]}}, p1_bit_slice_82908_comb};
  assign p1_sign_ext_82933_comb = {{1{p1_bit_slice_82911_comb[9]}}, p1_bit_slice_82911_comb};
  assign p1_sign_ext_82934_comb = {{1{p1_bit_slice_82912_comb[9]}}, p1_bit_slice_82912_comb};
  assign p1_bit_slice_82939_comb = p1_add_82835_comb[7:1];
  assign p1_bit_slice_82940_comb = p1_add_82836_comb[7:1];
  assign p1_bit_slice_82941_comb = p1_add_82837_comb[7:1];
  assign p1_bit_slice_82942_comb = p1_add_82838_comb[7:1];
  assign p1_add_82943_comb = {{1{p1_bit_slice_82903_comb[9]}}, p1_bit_slice_82903_comb} + 11'h001;
  assign p1_bit_slice_82944_comb = p1_add_82851_comb[7:1];
  assign p1_add_82945_comb = {{1{p1_bit_slice_82904_comb[9]}}, p1_bit_slice_82904_comb} + 11'h001;
  assign p1_bit_slice_82946_comb = p1_add_82852_comb[7:1];
  assign p1_add_82947_comb = {{1{p1_bit_slice_82905_comb[9]}}, p1_bit_slice_82905_comb} + 11'h001;
  assign p1_bit_slice_82948_comb = p1_add_82853_comb[7:1];
  assign p1_add_82949_comb = {{1{p1_bit_slice_82906_comb[9]}}, p1_bit_slice_82906_comb} + 11'h001;
  assign p1_bit_slice_82950_comb = p1_add_82854_comb[7:1];
  assign p1_bit_slice_82951_comb = p1_add_82867_comb[7:1];
  assign p1_bit_slice_82952_comb = p1_add_82868_comb[7:1];
  assign p1_add_82953_comb = {{1{p1_bit_slice_82909_comb[9]}}, p1_bit_slice_82909_comb} + 11'h001;
  assign p1_bit_slice_82954_comb = p1_add_82875_comb[7:1];
  assign p1_add_82955_comb = {{1{p1_bit_slice_82910_comb[9]}}, p1_bit_slice_82910_comb} + 11'h001;
  assign p1_bit_slice_82956_comb = p1_add_82876_comb[7:1];
  assign p1_bit_slice_82957_comb = p1_add_82883_comb[7:1];
  assign p1_bit_slice_82958_comb = p1_add_82884_comb[7:1];
  assign p1_add_82959_comb = {{1{p1_bit_slice_82913_comb[9]}}, p1_bit_slice_82913_comb} + 11'h001;
  assign p1_bit_slice_82960_comb = p1_add_82891_comb[7:1];
  assign p1_add_82961_comb = {{1{p1_bit_slice_82914_comb[9]}}, p1_bit_slice_82914_comb} + 11'h001;
  assign p1_bit_slice_82962_comb = p1_add_82892_comb[7:1];

  // Registers for pipe stage 1:
  reg [17:0] p1_add_82839;
  reg [17:0] p1_add_82840;
  reg [17:0] p1_add_82841;
  reg [17:0] p1_add_82842;
  reg [17:0] p1_add_82843;
  reg [17:0] p1_add_82844;
  reg [17:0] p1_add_82845;
  reg [17:0] p1_add_82846;
  reg [17:0] p1_add_82847;
  reg [17:0] p1_add_82848;
  reg [17:0] p1_add_82849;
  reg [17:0] p1_add_82850;
  reg [17:0] p1_add_82855;
  reg [17:0] p1_add_82856;
  reg [17:0] p1_add_82857;
  reg [17:0] p1_add_82858;
  reg [17:0] p1_add_82859;
  reg [17:0] p1_add_82860;
  reg [17:0] p1_add_82861;
  reg [17:0] p1_add_82862;
  reg [17:0] p1_add_82863;
  reg [17:0] p1_add_82864;
  reg [17:0] p1_add_82865;
  reg [17:0] p1_add_82866;
  reg [17:0] p1_add_82869;
  reg [17:0] p1_add_82870;
  reg [17:0] p1_add_82871;
  reg [17:0] p1_add_82872;
  reg [17:0] p1_add_82873;
  reg [17:0] p1_add_82874;
  reg [17:0] p1_add_82877;
  reg [17:0] p1_add_82878;
  reg [17:0] p1_add_82879;
  reg [17:0] p1_add_82880;
  reg [17:0] p1_add_82881;
  reg [17:0] p1_add_82882;
  reg [17:0] p1_add_82885;
  reg [17:0] p1_add_82886;
  reg [17:0] p1_add_82887;
  reg [17:0] p1_add_82888;
  reg [17:0] p1_add_82889;
  reg [17:0] p1_add_82890;
  reg [17:0] p1_add_82893;
  reg [17:0] p1_add_82894;
  reg [17:0] p1_add_82895;
  reg [17:0] p1_add_82896;
  reg [17:0] p1_add_82897;
  reg [17:0] p1_add_82898;
  reg [10:0] p1_sign_ext_82915;
  reg [10:0] p1_sign_ext_82916;
  reg [10:0] p1_sign_ext_82917;
  reg [10:0] p1_sign_ext_82918;
  reg [10:0] p1_sign_ext_82927;
  reg [10:0] p1_sign_ext_82928;
  reg [10:0] p1_sign_ext_82933;
  reg [10:0] p1_sign_ext_82934;
  reg [6:0] p1_bit_slice_82939;
  reg [6:0] p1_bit_slice_82940;
  reg [6:0] p1_bit_slice_82941;
  reg [6:0] p1_bit_slice_82942;
  reg [10:0] p1_add_82943;
  reg [6:0] p1_bit_slice_82944;
  reg [10:0] p1_add_82945;
  reg [6:0] p1_bit_slice_82946;
  reg [10:0] p1_add_82947;
  reg [6:0] p1_bit_slice_82948;
  reg [10:0] p1_add_82949;
  reg [6:0] p1_bit_slice_82950;
  reg [6:0] p1_bit_slice_82951;
  reg [6:0] p1_bit_slice_82952;
  reg [10:0] p1_add_82953;
  reg [6:0] p1_bit_slice_82954;
  reg [10:0] p1_add_82955;
  reg [6:0] p1_bit_slice_82956;
  reg [6:0] p1_bit_slice_82957;
  reg [6:0] p1_bit_slice_82958;
  reg [10:0] p1_add_82959;
  reg [6:0] p1_bit_slice_82960;
  reg [10:0] p1_add_82961;
  reg [6:0] p1_bit_slice_82962;
  always @ (posedge clk) begin
    p1_add_82839 <= p1_add_82839_comb;
    p1_add_82840 <= p1_add_82840_comb;
    p1_add_82841 <= p1_add_82841_comb;
    p1_add_82842 <= p1_add_82842_comb;
    p1_add_82843 <= p1_add_82843_comb;
    p1_add_82844 <= p1_add_82844_comb;
    p1_add_82845 <= p1_add_82845_comb;
    p1_add_82846 <= p1_add_82846_comb;
    p1_add_82847 <= p1_add_82847_comb;
    p1_add_82848 <= p1_add_82848_comb;
    p1_add_82849 <= p1_add_82849_comb;
    p1_add_82850 <= p1_add_82850_comb;
    p1_add_82855 <= p1_add_82855_comb;
    p1_add_82856 <= p1_add_82856_comb;
    p1_add_82857 <= p1_add_82857_comb;
    p1_add_82858 <= p1_add_82858_comb;
    p1_add_82859 <= p1_add_82859_comb;
    p1_add_82860 <= p1_add_82860_comb;
    p1_add_82861 <= p1_add_82861_comb;
    p1_add_82862 <= p1_add_82862_comb;
    p1_add_82863 <= p1_add_82863_comb;
    p1_add_82864 <= p1_add_82864_comb;
    p1_add_82865 <= p1_add_82865_comb;
    p1_add_82866 <= p1_add_82866_comb;
    p1_add_82869 <= p1_add_82869_comb;
    p1_add_82870 <= p1_add_82870_comb;
    p1_add_82871 <= p1_add_82871_comb;
    p1_add_82872 <= p1_add_82872_comb;
    p1_add_82873 <= p1_add_82873_comb;
    p1_add_82874 <= p1_add_82874_comb;
    p1_add_82877 <= p1_add_82877_comb;
    p1_add_82878 <= p1_add_82878_comb;
    p1_add_82879 <= p1_add_82879_comb;
    p1_add_82880 <= p1_add_82880_comb;
    p1_add_82881 <= p1_add_82881_comb;
    p1_add_82882 <= p1_add_82882_comb;
    p1_add_82885 <= p1_add_82885_comb;
    p1_add_82886 <= p1_add_82886_comb;
    p1_add_82887 <= p1_add_82887_comb;
    p1_add_82888 <= p1_add_82888_comb;
    p1_add_82889 <= p1_add_82889_comb;
    p1_add_82890 <= p1_add_82890_comb;
    p1_add_82893 <= p1_add_82893_comb;
    p1_add_82894 <= p1_add_82894_comb;
    p1_add_82895 <= p1_add_82895_comb;
    p1_add_82896 <= p1_add_82896_comb;
    p1_add_82897 <= p1_add_82897_comb;
    p1_add_82898 <= p1_add_82898_comb;
    p1_sign_ext_82915 <= p1_sign_ext_82915_comb;
    p1_sign_ext_82916 <= p1_sign_ext_82916_comb;
    p1_sign_ext_82917 <= p1_sign_ext_82917_comb;
    p1_sign_ext_82918 <= p1_sign_ext_82918_comb;
    p1_sign_ext_82927 <= p1_sign_ext_82927_comb;
    p1_sign_ext_82928 <= p1_sign_ext_82928_comb;
    p1_sign_ext_82933 <= p1_sign_ext_82933_comb;
    p1_sign_ext_82934 <= p1_sign_ext_82934_comb;
    p1_bit_slice_82939 <= p1_bit_slice_82939_comb;
    p1_bit_slice_82940 <= p1_bit_slice_82940_comb;
    p1_bit_slice_82941 <= p1_bit_slice_82941_comb;
    p1_bit_slice_82942 <= p1_bit_slice_82942_comb;
    p1_add_82943 <= p1_add_82943_comb;
    p1_bit_slice_82944 <= p1_bit_slice_82944_comb;
    p1_add_82945 <= p1_add_82945_comb;
    p1_bit_slice_82946 <= p1_bit_slice_82946_comb;
    p1_add_82947 <= p1_add_82947_comb;
    p1_bit_slice_82948 <= p1_bit_slice_82948_comb;
    p1_add_82949 <= p1_add_82949_comb;
    p1_bit_slice_82950 <= p1_bit_slice_82950_comb;
    p1_bit_slice_82951 <= p1_bit_slice_82951_comb;
    p1_bit_slice_82952 <= p1_bit_slice_82952_comb;
    p1_add_82953 <= p1_add_82953_comb;
    p1_bit_slice_82954 <= p1_bit_slice_82954_comb;
    p1_add_82955 <= p1_add_82955_comb;
    p1_bit_slice_82956 <= p1_bit_slice_82956_comb;
    p1_bit_slice_82957 <= p1_bit_slice_82957_comb;
    p1_bit_slice_82958 <= p1_bit_slice_82958_comb;
    p1_add_82959 <= p1_add_82959_comb;
    p1_bit_slice_82960 <= p1_bit_slice_82960_comb;
    p1_add_82961 <= p1_add_82961_comb;
    p1_bit_slice_82962 <= p1_bit_slice_82962_comb;
  end

  // ===== Pipe stage 2:
  wire [9:0] p2_bit_slice_83123_comb;
  wire [9:0] p2_bit_slice_83124_comb;
  wire [9:0] p2_bit_slice_83125_comb;
  wire [9:0] p2_bit_slice_83126_comb;
  wire [9:0] p2_bit_slice_83127_comb;
  wire [9:0] p2_bit_slice_83128_comb;
  wire [9:0] p2_bit_slice_83129_comb;
  wire [9:0] p2_bit_slice_83130_comb;
  wire [9:0] p2_bit_slice_83131_comb;
  wire [9:0] p2_bit_slice_83132_comb;
  wire [9:0] p2_bit_slice_83133_comb;
  wire [9:0] p2_bit_slice_83134_comb;
  wire [9:0] p2_bit_slice_83135_comb;
  wire [9:0] p2_bit_slice_83136_comb;
  wire [9:0] p2_bit_slice_83137_comb;
  wire [9:0] p2_bit_slice_83138_comb;
  wire [9:0] p2_bit_slice_83139_comb;
  wire [9:0] p2_bit_slice_83140_comb;
  wire [9:0] p2_bit_slice_83141_comb;
  wire [9:0] p2_bit_slice_83142_comb;
  wire [9:0] p2_bit_slice_83143_comb;
  wire [9:0] p2_bit_slice_83144_comb;
  wire [9:0] p2_bit_slice_83145_comb;
  wire [9:0] p2_bit_slice_83146_comb;
  wire [9:0] p2_bit_slice_83147_comb;
  wire [9:0] p2_bit_slice_83148_comb;
  wire [9:0] p2_bit_slice_83149_comb;
  wire [9:0] p2_bit_slice_83150_comb;
  wire [9:0] p2_bit_slice_83151_comb;
  wire [9:0] p2_bit_slice_83152_comb;
  wire [9:0] p2_bit_slice_83153_comb;
  wire [9:0] p2_bit_slice_83154_comb;
  wire [9:0] p2_bit_slice_83155_comb;
  wire [9:0] p2_bit_slice_83156_comb;
  wire [9:0] p2_bit_slice_83157_comb;
  wire [9:0] p2_bit_slice_83158_comb;
  wire [9:0] p2_bit_slice_83159_comb;
  wire [9:0] p2_bit_slice_83160_comb;
  wire [9:0] p2_bit_slice_83161_comb;
  wire [9:0] p2_bit_slice_83162_comb;
  wire [9:0] p2_bit_slice_83163_comb;
  wire [9:0] p2_bit_slice_83164_comb;
  wire [9:0] p2_bit_slice_83165_comb;
  wire [9:0] p2_bit_slice_83166_comb;
  wire [9:0] p2_bit_slice_83167_comb;
  wire [9:0] p2_bit_slice_83168_comb;
  wire [9:0] p2_bit_slice_83169_comb;
  wire [9:0] p2_bit_slice_83170_comb;
  wire [10:0] p2_add_83275_comb;
  wire [10:0] p2_add_83276_comb;
  wire [10:0] p2_add_83277_comb;
  wire [10:0] p2_add_83278_comb;
  wire [10:0] p2_add_83327_comb;
  wire [10:0] p2_add_83328_comb;
  wire [10:0] p2_add_83353_comb;
  wire [10:0] p2_add_83354_comb;
  wire [17:0] p2_concat_83427_comb;
  wire [17:0] p2_concat_83430_comb;
  wire [17:0] p2_concat_83433_comb;
  wire [17:0] p2_concat_83436_comb;
  wire [17:0] p2_concat_83499_comb;
  wire [17:0] p2_concat_83502_comb;
  wire [17:0] p2_concat_83547_comb;
  wire [17:0] p2_concat_83550_comb;
  wire [17:0] p2_concat_83379_comb;
  wire [17:0] p2_concat_83382_comb;
  wire [17:0] p2_concat_83385_comb;
  wire [17:0] p2_concat_83388_comb;
  wire [17:0] p2_concat_83475_comb;
  wire [17:0] p2_concat_83478_comb;
  wire [17:0] p2_concat_83523_comb;
  wire [17:0] p2_concat_83526_comb;
  wire [10:0] p2_add_83279_comb;
  wire [10:0] p2_add_83281_comb;
  wire [10:0] p2_add_83283_comb;
  wire [10:0] p2_add_83285_comb;
  wire [10:0] p2_add_83287_comb;
  wire [10:0] p2_add_83289_comb;
  wire [10:0] p2_add_83291_comb;
  wire [10:0] p2_add_83293_comb;
  wire [10:0] p2_add_83295_comb;
  wire [10:0] p2_add_83297_comb;
  wire [10:0] p2_add_83299_comb;
  wire [10:0] p2_add_83301_comb;
  wire [10:0] p2_add_83303_comb;
  wire [10:0] p2_add_83305_comb;
  wire [10:0] p2_add_83307_comb;
  wire [10:0] p2_add_83309_comb;
  wire [10:0] p2_add_83311_comb;
  wire [10:0] p2_add_83313_comb;
  wire [10:0] p2_add_83315_comb;
  wire [10:0] p2_add_83317_comb;
  wire [10:0] p2_add_83319_comb;
  wire [10:0] p2_add_83321_comb;
  wire [10:0] p2_add_83323_comb;
  wire [10:0] p2_add_83325_comb;
  wire [10:0] p2_add_83329_comb;
  wire [10:0] p2_add_83331_comb;
  wire [10:0] p2_add_83333_comb;
  wire [10:0] p2_add_83335_comb;
  wire [10:0] p2_add_83337_comb;
  wire [10:0] p2_add_83339_comb;
  wire [10:0] p2_add_83341_comb;
  wire [10:0] p2_add_83343_comb;
  wire [10:0] p2_add_83345_comb;
  wire [10:0] p2_add_83347_comb;
  wire [10:0] p2_add_83349_comb;
  wire [10:0] p2_add_83351_comb;
  wire [10:0] p2_add_83355_comb;
  wire [10:0] p2_add_83357_comb;
  wire [10:0] p2_add_83359_comb;
  wire [10:0] p2_add_83361_comb;
  wire [10:0] p2_add_83363_comb;
  wire [10:0] p2_add_83365_comb;
  wire [10:0] p2_add_83367_comb;
  wire [10:0] p2_add_83369_comb;
  wire [10:0] p2_add_83371_comb;
  wire [10:0] p2_add_83373_comb;
  wire [10:0] p2_add_83375_comb;
  wire [10:0] p2_add_83377_comb;
  wire [17:0] p2_concat_83391_comb;
  wire [17:0] p2_concat_83394_comb;
  wire [17:0] p2_concat_83397_comb;
  wire [17:0] p2_concat_83400_comb;
  wire [17:0] p2_concat_83403_comb;
  wire [17:0] p2_concat_83406_comb;
  wire [17:0] p2_concat_83409_comb;
  wire [17:0] p2_concat_83412_comb;
  wire [17:0] p2_concat_83415_comb;
  wire [17:0] p2_concat_83418_comb;
  wire [17:0] p2_concat_83421_comb;
  wire [17:0] p2_concat_83424_comb;
  wire [17:0] p2_concat_83439_comb;
  wire [17:0] p2_concat_83442_comb;
  wire [17:0] p2_concat_83445_comb;
  wire [17:0] p2_concat_83448_comb;
  wire [17:0] p2_concat_83451_comb;
  wire [17:0] p2_concat_83454_comb;
  wire [17:0] p2_concat_83457_comb;
  wire [17:0] p2_concat_83460_comb;
  wire [17:0] p2_concat_83463_comb;
  wire [17:0] p2_concat_83466_comb;
  wire [17:0] p2_concat_83469_comb;
  wire [17:0] p2_concat_83472_comb;
  wire [17:0] p2_concat_83481_comb;
  wire [17:0] p2_concat_83484_comb;
  wire [17:0] p2_concat_83487_comb;
  wire [17:0] p2_concat_83490_comb;
  wire [17:0] p2_concat_83493_comb;
  wire [17:0] p2_concat_83496_comb;
  wire [17:0] p2_concat_83505_comb;
  wire [17:0] p2_concat_83508_comb;
  wire [17:0] p2_concat_83511_comb;
  wire [17:0] p2_concat_83514_comb;
  wire [17:0] p2_concat_83517_comb;
  wire [17:0] p2_concat_83520_comb;
  wire [17:0] p2_concat_83529_comb;
  wire [17:0] p2_concat_83532_comb;
  wire [17:0] p2_concat_83535_comb;
  wire [17:0] p2_concat_83538_comb;
  wire [17:0] p2_concat_83541_comb;
  wire [17:0] p2_concat_83544_comb;
  wire [17:0] p2_concat_83553_comb;
  wire [17:0] p2_concat_83556_comb;
  wire [17:0] p2_concat_83559_comb;
  wire [17:0] p2_concat_83562_comb;
  wire [17:0] p2_concat_83565_comb;
  wire [17:0] p2_concat_83568_comb;
  wire [9:0] p2_clipped__44_comb;
  wire [9:0] p2_clipped__60_comb;
  wire [9:0] p2_clipped__76_comb;
  wire [9:0] p2_clipped__92_comb;
  wire [9:0] p2_clipped__28_comb;
  wire [9:0] p2_clipped__108_comb;
  wire [9:0] p2_clipped__12_comb;
  wire [9:0] p2_clipped__124_comb;
  wire [9:0] p2_clipped__40_comb;
  wire [9:0] p2_clipped__56_comb;
  wire [9:0] p2_clipped__72_comb;
  wire [9:0] p2_clipped__88_comb;
  wire [9:0] p2_clipped__24_comb;
  wire [9:0] p2_clipped__104_comb;
  wire [9:0] p2_clipped__8_comb;
  wire [9:0] p2_clipped__120_comb;
  wire [2:0] p2_bit_slice_84099_comb;
  wire [2:0] p2_bit_slice_84100_comb;
  wire [2:0] p2_bit_slice_84101_comb;
  wire [2:0] p2_bit_slice_84102_comb;
  wire [2:0] p2_bit_slice_84123_comb;
  wire [2:0] p2_bit_slice_84124_comb;
  wire [2:0] p2_bit_slice_84139_comb;
  wire [2:0] p2_bit_slice_84140_comb;
  wire [2:0] p2_bit_slice_84083_comb;
  wire [2:0] p2_bit_slice_84084_comb;
  wire [2:0] p2_bit_slice_84085_comb;
  wire [2:0] p2_bit_slice_84086_comb;
  wire [2:0] p2_bit_slice_84115_comb;
  wire [2:0] p2_bit_slice_84116_comb;
  wire [2:0] p2_bit_slice_84131_comb;
  wire [2:0] p2_bit_slice_84132_comb;
  wire [9:0] p2_clipped__41_comb;
  wire [9:0] p2_clipped__57_comb;
  wire [9:0] p2_clipped__73_comb;
  wire [9:0] p2_clipped__89_comb;
  wire [9:0] p2_clipped__42_comb;
  wire [9:0] p2_clipped__58_comb;
  wire [9:0] p2_clipped__74_comb;
  wire [9:0] p2_clipped__90_comb;
  wire [9:0] p2_clipped__43_comb;
  wire [9:0] p2_clipped__59_comb;
  wire [9:0] p2_clipped__75_comb;
  wire [9:0] p2_clipped__91_comb;
  wire [9:0] p2_clipped__45_comb;
  wire [9:0] p2_clipped__61_comb;
  wire [9:0] p2_clipped__77_comb;
  wire [9:0] p2_clipped__93_comb;
  wire [9:0] p2_clipped__46_comb;
  wire [9:0] p2_clipped__62_comb;
  wire [9:0] p2_clipped__78_comb;
  wire [9:0] p2_clipped__94_comb;
  wire [9:0] p2_clipped__47_comb;
  wire [9:0] p2_clipped__63_comb;
  wire [9:0] p2_clipped__79_comb;
  wire [9:0] p2_clipped__95_comb;
  wire [9:0] p2_clipped__25_comb;
  wire [9:0] p2_clipped__105_comb;
  wire [9:0] p2_clipped__26_comb;
  wire [9:0] p2_clipped__106_comb;
  wire [9:0] p2_clipped__27_comb;
  wire [9:0] p2_clipped__107_comb;
  wire [9:0] p2_clipped__29_comb;
  wire [9:0] p2_clipped__109_comb;
  wire [9:0] p2_clipped__30_comb;
  wire [9:0] p2_clipped__110_comb;
  wire [9:0] p2_clipped__31_comb;
  wire [9:0] p2_clipped__111_comb;
  wire [9:0] p2_clipped__9_comb;
  wire [9:0] p2_clipped__121_comb;
  wire [9:0] p2_clipped__10_comb;
  wire [9:0] p2_clipped__122_comb;
  wire [9:0] p2_clipped__11_comb;
  wire [9:0] p2_clipped__123_comb;
  wire [9:0] p2_clipped__13_comb;
  wire [9:0] p2_clipped__125_comb;
  wire [9:0] p2_clipped__14_comb;
  wire [9:0] p2_clipped__126_comb;
  wire [9:0] p2_clipped__15_comb;
  wire [9:0] p2_clipped__127_comb;
  wire [3:0] p2_add_84307_comb;
  wire [3:0] p2_add_84309_comb;
  wire [3:0] p2_add_84311_comb;
  wire [3:0] p2_add_84313_comb;
  wire [3:0] p2_add_84355_comb;
  wire [3:0] p2_add_84357_comb;
  wire [3:0] p2_add_84387_comb;
  wire [3:0] p2_add_84389_comb;
  wire [2:0] p2_bit_slice_84087_comb;
  wire [2:0] p2_bit_slice_84088_comb;
  wire [2:0] p2_bit_slice_84089_comb;
  wire [2:0] p2_bit_slice_84090_comb;
  wire [2:0] p2_bit_slice_84091_comb;
  wire [2:0] p2_bit_slice_84092_comb;
  wire [2:0] p2_bit_slice_84093_comb;
  wire [2:0] p2_bit_slice_84094_comb;
  wire [2:0] p2_bit_slice_84095_comb;
  wire [2:0] p2_bit_slice_84096_comb;
  wire [2:0] p2_bit_slice_84097_comb;
  wire [2:0] p2_bit_slice_84098_comb;
  wire [2:0] p2_bit_slice_84103_comb;
  wire [2:0] p2_bit_slice_84104_comb;
  wire [2:0] p2_bit_slice_84105_comb;
  wire [2:0] p2_bit_slice_84106_comb;
  wire [2:0] p2_bit_slice_84107_comb;
  wire [2:0] p2_bit_slice_84108_comb;
  wire [2:0] p2_bit_slice_84109_comb;
  wire [2:0] p2_bit_slice_84110_comb;
  wire [2:0] p2_bit_slice_84111_comb;
  wire [2:0] p2_bit_slice_84112_comb;
  wire [2:0] p2_bit_slice_84113_comb;
  wire [2:0] p2_bit_slice_84114_comb;
  wire [2:0] p2_bit_slice_84117_comb;
  wire [2:0] p2_bit_slice_84118_comb;
  wire [2:0] p2_bit_slice_84119_comb;
  wire [2:0] p2_bit_slice_84120_comb;
  wire [2:0] p2_bit_slice_84121_comb;
  wire [2:0] p2_bit_slice_84122_comb;
  wire [2:0] p2_bit_slice_84125_comb;
  wire [2:0] p2_bit_slice_84126_comb;
  wire [2:0] p2_bit_slice_84127_comb;
  wire [2:0] p2_bit_slice_84128_comb;
  wire [2:0] p2_bit_slice_84129_comb;
  wire [2:0] p2_bit_slice_84130_comb;
  wire [2:0] p2_bit_slice_84133_comb;
  wire [2:0] p2_bit_slice_84134_comb;
  wire [2:0] p2_bit_slice_84135_comb;
  wire [2:0] p2_bit_slice_84136_comb;
  wire [2:0] p2_bit_slice_84137_comb;
  wire [2:0] p2_bit_slice_84138_comb;
  wire [2:0] p2_bit_slice_84141_comb;
  wire [2:0] p2_bit_slice_84142_comb;
  wire [2:0] p2_bit_slice_84143_comb;
  wire [2:0] p2_bit_slice_84144_comb;
  wire [2:0] p2_bit_slice_84145_comb;
  wire [2:0] p2_bit_slice_84146_comb;
  wire [3:0] p2_add_84275_comb;
  wire [3:0] p2_add_84277_comb;
  wire [3:0] p2_add_84279_comb;
  wire [3:0] p2_add_84281_comb;
  wire [3:0] p2_add_84339_comb;
  wire [3:0] p2_add_84341_comb;
  wire [3:0] p2_add_84371_comb;
  wire [3:0] p2_add_84373_comb;
  wire [10:0] p2_concat_84419_comb;
  wire [10:0] p2_concat_84420_comb;
  wire [10:0] p2_concat_84421_comb;
  wire [10:0] p2_concat_84422_comb;
  wire [10:0] p2_concat_84443_comb;
  wire [10:0] p2_concat_84444_comb;
  wire [10:0] p2_concat_84459_comb;
  wire [10:0] p2_concat_84460_comb;
  wire [10:0] p2_concat_84403_comb;
  wire [10:0] p2_concat_84404_comb;
  wire [10:0] p2_concat_84405_comb;
  wire [10:0] p2_concat_84406_comb;
  wire [10:0] p2_concat_84435_comb;
  wire [10:0] p2_concat_84436_comb;
  wire [10:0] p2_concat_84451_comb;
  wire [10:0] p2_concat_84452_comb;
  wire [23:0] p2_sign_ext_84501_comb;
  wire [23:0] p2_sign_ext_84502_comb;
  wire [23:0] p2_sign_ext_84503_comb;
  wire [23:0] p2_sign_ext_84504_comb;
  wire [23:0] p2_sign_ext_84539_comb;
  wire [23:0] p2_sign_ext_84540_comb;
  wire [23:0] p2_sign_ext_84603_comb;
  wire [23:0] p2_sign_ext_84608_comb;
  wire [3:0] p2_add_84283_comb;
  wire [3:0] p2_add_84285_comb;
  wire [3:0] p2_add_84287_comb;
  wire [3:0] p2_add_84289_comb;
  wire [3:0] p2_add_84291_comb;
  wire [3:0] p2_add_84293_comb;
  wire [3:0] p2_add_84295_comb;
  wire [3:0] p2_add_84297_comb;
  wire [3:0] p2_add_84299_comb;
  wire [3:0] p2_add_84301_comb;
  wire [3:0] p2_add_84303_comb;
  wire [3:0] p2_add_84305_comb;
  wire [3:0] p2_add_84315_comb;
  wire [3:0] p2_add_84317_comb;
  wire [3:0] p2_add_84319_comb;
  wire [3:0] p2_add_84321_comb;
  wire [3:0] p2_add_84323_comb;
  wire [3:0] p2_add_84325_comb;
  wire [3:0] p2_add_84327_comb;
  wire [3:0] p2_add_84329_comb;
  wire [3:0] p2_add_84331_comb;
  wire [3:0] p2_add_84333_comb;
  wire [3:0] p2_add_84335_comb;
  wire [3:0] p2_add_84337_comb;
  wire [3:0] p2_add_84343_comb;
  wire [3:0] p2_add_84345_comb;
  wire [3:0] p2_add_84347_comb;
  wire [3:0] p2_add_84349_comb;
  wire [3:0] p2_add_84351_comb;
  wire [3:0] p2_add_84353_comb;
  wire [3:0] p2_add_84359_comb;
  wire [3:0] p2_add_84361_comb;
  wire [3:0] p2_add_84363_comb;
  wire [3:0] p2_add_84365_comb;
  wire [3:0] p2_add_84367_comb;
  wire [3:0] p2_add_84369_comb;
  wire [3:0] p2_add_84375_comb;
  wire [3:0] p2_add_84377_comb;
  wire [3:0] p2_add_84379_comb;
  wire [3:0] p2_add_84381_comb;
  wire [3:0] p2_add_84383_comb;
  wire [3:0] p2_add_84385_comb;
  wire [3:0] p2_add_84391_comb;
  wire [3:0] p2_add_84393_comb;
  wire [3:0] p2_add_84395_comb;
  wire [3:0] p2_add_84397_comb;
  wire [3:0] p2_add_84399_comb;
  wire [3:0] p2_add_84401_comb;
  wire [23:0] p2_sign_ext_84469_comb;
  wire [23:0] p2_sign_ext_84470_comb;
  wire [23:0] p2_sign_ext_84471_comb;
  wire [23:0] p2_sign_ext_84472_comb;
  wire [23:0] p2_sign_ext_84531_comb;
  wire [23:0] p2_sign_ext_84532_comb;
  wire [23:0] p2_sign_ext_84579_comb;
  wire [23:0] p2_sign_ext_84584_comb;
  wire [19:0] p2_smul_84707_comb;
  wire [19:0] p2_smul_84708_comb;
  wire [19:0] p2_smul_84717_comb;
  wire [19:0] p2_smul_84718_comb;
  wire [19:0] p2_smul_84859_comb;
  wire [19:0] p2_smul_84861_comb;
  wire [19:0] p2_smul_84866_comb;
  wire [19:0] p2_smul_84868_comb;
  wire [19:0] p2_smul_84941_comb;
  wire [19:0] p2_smul_84943_comb;
  wire [19:0] p2_smul_84944_comb;
  wire [19:0] p2_smul_84946_comb;
  wire [19:0] p2_smul_85063_comb;
  wire [19:0] p2_smul_85064_comb;
  wire [19:0] p2_smul_85065_comb;
  wire [19:0] p2_smul_85066_comb;
  wire [10:0] p2_concat_84407_comb;
  wire [10:0] p2_concat_84408_comb;
  wire [10:0] p2_concat_84409_comb;
  wire [10:0] p2_concat_84410_comb;
  wire [10:0] p2_concat_84411_comb;
  wire [10:0] p2_concat_84412_comb;
  wire [10:0] p2_concat_84413_comb;
  wire [10:0] p2_concat_84414_comb;
  wire [10:0] p2_concat_84415_comb;
  wire [10:0] p2_concat_84416_comb;
  wire [10:0] p2_concat_84417_comb;
  wire [10:0] p2_concat_84418_comb;
  wire [10:0] p2_concat_84423_comb;
  wire [10:0] p2_concat_84424_comb;
  wire [10:0] p2_concat_84425_comb;
  wire [10:0] p2_concat_84426_comb;
  wire [10:0] p2_concat_84427_comb;
  wire [10:0] p2_concat_84428_comb;
  wire [10:0] p2_concat_84429_comb;
  wire [10:0] p2_concat_84430_comb;
  wire [10:0] p2_concat_84431_comb;
  wire [10:0] p2_concat_84432_comb;
  wire [10:0] p2_concat_84433_comb;
  wire [10:0] p2_concat_84434_comb;
  wire [10:0] p2_concat_84437_comb;
  wire [10:0] p2_concat_84438_comb;
  wire [10:0] p2_concat_84439_comb;
  wire [10:0] p2_concat_84440_comb;
  wire [10:0] p2_concat_84441_comb;
  wire [10:0] p2_concat_84442_comb;
  wire [10:0] p2_concat_84445_comb;
  wire [10:0] p2_concat_84446_comb;
  wire [10:0] p2_concat_84447_comb;
  wire [10:0] p2_concat_84448_comb;
  wire [10:0] p2_concat_84449_comb;
  wire [10:0] p2_concat_84450_comb;
  wire [10:0] p2_concat_84453_comb;
  wire [10:0] p2_concat_84454_comb;
  wire [10:0] p2_concat_84455_comb;
  wire [10:0] p2_concat_84456_comb;
  wire [10:0] p2_concat_84457_comb;
  wire [10:0] p2_concat_84458_comb;
  wire [10:0] p2_concat_84461_comb;
  wire [10:0] p2_concat_84462_comb;
  wire [10:0] p2_concat_84463_comb;
  wire [10:0] p2_concat_84464_comb;
  wire [10:0] p2_concat_84465_comb;
  wire [10:0] p2_concat_84466_comb;
  wire [19:0] p2_smul_84659_comb;
  wire [19:0] p2_smul_84660_comb;
  wire [19:0] p2_smul_84669_comb;
  wire [19:0] p2_smul_84670_comb;
  wire [19:0] p2_smul_84819_comb;
  wire [19:0] p2_smul_84821_comb;
  wire [19:0] p2_smul_84826_comb;
  wire [19:0] p2_smul_84828_comb;
  wire [19:0] p2_smul_84901_comb;
  wire [19:0] p2_smul_84903_comb;
  wire [19:0] p2_smul_84904_comb;
  wire [19:0] p2_smul_84906_comb;
  wire [19:0] p2_smul_85015_comb;
  wire [19:0] p2_smul_85016_comb;
  wire [19:0] p2_smul_85017_comb;
  wire [19:0] p2_smul_85018_comb;
  wire [19:0] p2_add_85131_comb;
  wire [17:0] p2_smul_85132_comb;
  wire [17:0] p2_smul_85133_comb;
  wire [17:0] p2_smul_85134_comb;
  wire [17:0] p2_smul_85135_comb;
  wire [19:0] p2_add_85136_comb;
  wire [18:0] p2_smul_85188_comb;
  wire [18:0] p2_smul_85189_comb;
  wire [18:0] p2_smul_85192_comb;
  wire [18:0] p2_smul_85193_comb;
  wire [18:0] p2_smul_85252_comb;
  wire [18:0] p2_smul_85254_comb;
  wire [18:0] p2_smul_85255_comb;
  wire [18:0] p2_smul_85257_comb;
  wire [18:0] p2_smul_85379_comb;
  wire [18:0] p2_smul_85381_comb;
  wire [18:0] p2_smul_85384_comb;
  wire [18:0] p2_smul_85386_comb;
  wire [18:0] p2_smul_85443_comb;
  wire [18:0] p2_smul_85445_comb;
  wire [18:0] p2_smul_85448_comb;
  wire [18:0] p2_smul_85450_comb;
  wire [17:0] p2_smul_85499_comb;
  wire [17:0] p2_smul_85500_comb;
  wire [19:0] p2_add_85501_comb;
  wire [19:0] p2_add_85502_comb;
  wire [17:0] p2_smul_85503_comb;
  wire [17:0] p2_smul_85504_comb;
  wire [18:0] p2_smul_85747_comb;
  wire [18:0] p2_smul_85748_comb;
  wire [18:0] p2_smul_85749_comb;
  wire [18:0] p2_smul_85750_comb;
  wire [18:0] p2_smul_85751_comb;
  wire [18:0] p2_smul_85752_comb;
  wire [18:0] p2_smul_85753_comb;
  wire [18:0] p2_smul_85754_comb;
  wire [18:0] p2_smul_85779_comb;
  wire [18:0] p2_smul_85780_comb;
  wire [18:0] p2_smul_85781_comb;
  wire [18:0] p2_smul_85782_comb;
  wire [18:0] p2_smul_85783_comb;
  wire [18:0] p2_smul_85784_comb;
  wire [18:0] p2_smul_85785_comb;
  wire [18:0] p2_smul_85786_comb;
  wire [23:0] p2_sign_ext_84477_comb;
  wire [23:0] p2_sign_ext_84478_comb;
  wire [23:0] p2_sign_ext_84479_comb;
  wire [23:0] p2_sign_ext_84480_comb;
  wire [23:0] p2_sign_ext_84485_comb;
  wire [23:0] p2_sign_ext_84486_comb;
  wire [23:0] p2_sign_ext_84487_comb;
  wire [23:0] p2_sign_ext_84488_comb;
  wire [23:0] p2_sign_ext_84493_comb;
  wire [23:0] p2_sign_ext_84494_comb;
  wire [23:0] p2_sign_ext_84495_comb;
  wire [23:0] p2_sign_ext_84496_comb;
  wire [23:0] p2_sign_ext_84509_comb;
  wire [23:0] p2_sign_ext_84510_comb;
  wire [23:0] p2_sign_ext_84511_comb;
  wire [23:0] p2_sign_ext_84512_comb;
  wire [23:0] p2_sign_ext_84517_comb;
  wire [23:0] p2_sign_ext_84518_comb;
  wire [23:0] p2_sign_ext_84519_comb;
  wire [23:0] p2_sign_ext_84520_comb;
  wire [23:0] p2_sign_ext_84525_comb;
  wire [23:0] p2_sign_ext_84526_comb;
  wire [23:0] p2_sign_ext_84527_comb;
  wire [23:0] p2_sign_ext_84528_comb;
  wire [23:0] p2_sign_ext_84533_comb;
  wire [23:0] p2_sign_ext_84534_comb;
  wire [23:0] p2_sign_ext_84535_comb;
  wire [23:0] p2_sign_ext_84536_comb;
  wire [23:0] p2_sign_ext_84537_comb;
  wire [23:0] p2_sign_ext_84538_comb;
  wire [23:0] p2_sign_ext_84541_comb;
  wire [23:0] p2_sign_ext_84542_comb;
  wire [23:0] p2_sign_ext_84543_comb;
  wire [23:0] p2_sign_ext_84544_comb;
  wire [23:0] p2_sign_ext_84545_comb;
  wire [23:0] p2_sign_ext_84546_comb;
  wire [23:0] p2_sign_ext_84585_comb;
  wire [23:0] p2_sign_ext_84590_comb;
  wire [23:0] p2_sign_ext_84591_comb;
  wire [23:0] p2_sign_ext_84596_comb;
  wire [23:0] p2_sign_ext_84597_comb;
  wire [23:0] p2_sign_ext_84602_comb;
  wire [23:0] p2_sign_ext_84609_comb;
  wire [23:0] p2_sign_ext_84614_comb;
  wire [23:0] p2_sign_ext_84615_comb;
  wire [23:0] p2_sign_ext_84620_comb;
  wire [23:0] p2_sign_ext_84621_comb;
  wire [23:0] p2_sign_ext_84626_comb;
  wire [19:0] p2_add_85107_comb;
  wire [17:0] p2_smul_85108_comb;
  wire [17:0] p2_smul_85109_comb;
  wire [17:0] p2_smul_85110_comb;
  wire [17:0] p2_smul_85111_comb;
  wire [19:0] p2_add_85112_comb;
  wire [18:0] p2_smul_85156_comb;
  wire [18:0] p2_smul_85157_comb;
  wire [18:0] p2_smul_85160_comb;
  wire [18:0] p2_smul_85161_comb;
  wire [18:0] p2_smul_85220_comb;
  wire [18:0] p2_smul_85222_comb;
  wire [18:0] p2_smul_85223_comb;
  wire [18:0] p2_smul_85225_comb;
  wire [18:0] p2_smul_85347_comb;
  wire [18:0] p2_smul_85349_comb;
  wire [18:0] p2_smul_85352_comb;
  wire [18:0] p2_smul_85354_comb;
  wire [18:0] p2_smul_85411_comb;
  wire [18:0] p2_smul_85413_comb;
  wire [18:0] p2_smul_85416_comb;
  wire [18:0] p2_smul_85418_comb;
  wire [17:0] p2_smul_85475_comb;
  wire [17:0] p2_smul_85476_comb;
  wire [19:0] p2_add_85477_comb;
  wire [19:0] p2_add_85478_comb;
  wire [17:0] p2_smul_85479_comb;
  wire [17:0] p2_smul_85480_comb;
  wire [18:0] p2_bit_slice_85603_comb;
  wire [17:0] p2_add_85604_comb;
  wire [17:0] p2_add_85605_comb;
  wire [18:0] p2_bit_slice_85606_comb;
  wire [17:0] p2_smul_85651_comb;
  wire [17:0] p2_smul_85654_comb;
  wire [17:0] p2_smul_85655_comb;
  wire [17:0] p2_smul_85658_comb;
  wire [18:0] p2_add_85715_comb;
  wire [18:0] p2_add_85717_comb;
  wire [18:0] p2_add_85719_comb;
  wire [18:0] p2_add_85721_comb;
  wire [18:0] p2_smul_85755_comb;
  wire [18:0] p2_smul_85756_comb;
  wire [18:0] p2_smul_85757_comb;
  wire [18:0] p2_smul_85758_comb;
  wire [18:0] p2_smul_85759_comb;
  wire [18:0] p2_smul_85760_comb;
  wire [18:0] p2_smul_85761_comb;
  wire [18:0] p2_smul_85762_comb;
  wire [18:0] p2_smul_85763_comb;
  wire [18:0] p2_smul_85764_comb;
  wire [18:0] p2_smul_85765_comb;
  wire [18:0] p2_smul_85766_comb;
  wire [18:0] p2_smul_85767_comb;
  wire [18:0] p2_smul_85768_comb;
  wire [18:0] p2_smul_85769_comb;
  wire [18:0] p2_smul_85770_comb;
  wire [18:0] p2_smul_85771_comb;
  wire [18:0] p2_smul_85772_comb;
  wire [18:0] p2_smul_85773_comb;
  wire [18:0] p2_smul_85774_comb;
  wire [18:0] p2_smul_85775_comb;
  wire [18:0] p2_smul_85776_comb;
  wire [18:0] p2_smul_85777_comb;
  wire [18:0] p2_smul_85778_comb;
  wire [18:0] p2_smul_85787_comb;
  wire [18:0] p2_smul_85788_comb;
  wire [18:0] p2_smul_85789_comb;
  wire [18:0] p2_smul_85790_comb;
  wire [18:0] p2_smul_85791_comb;
  wire [18:0] p2_smul_85792_comb;
  wire [18:0] p2_smul_85793_comb;
  wire [18:0] p2_smul_85794_comb;
  wire [18:0] p2_smul_85795_comb;
  wire [18:0] p2_smul_85796_comb;
  wire [18:0] p2_smul_85797_comb;
  wire [18:0] p2_smul_85798_comb;
  wire [18:0] p2_smul_85799_comb;
  wire [18:0] p2_smul_85800_comb;
  wire [18:0] p2_smul_85801_comb;
  wire [18:0] p2_smul_85802_comb;
  wire [18:0] p2_smul_85803_comb;
  wire [18:0] p2_smul_85804_comb;
  wire [18:0] p2_smul_85805_comb;
  wire [18:0] p2_smul_85806_comb;
  wire [18:0] p2_smul_85807_comb;
  wire [18:0] p2_smul_85808_comb;
  wire [18:0] p2_smul_85809_comb;
  wire [18:0] p2_smul_85810_comb;
  wire [18:0] p2_add_85843_comb;
  wire [18:0] p2_add_85845_comb;
  wire [18:0] p2_add_85847_comb;
  wire [18:0] p2_add_85849_comb;
  wire [17:0] p2_smul_85908_comb;
  wire [17:0] p2_smul_85910_comb;
  wire [17:0] p2_smul_85911_comb;
  wire [17:0] p2_smul_85913_comb;
  wire [17:0] p2_add_85955_comb;
  wire [18:0] p2_bit_slice_85956_comb;
  wire [18:0] p2_bit_slice_85957_comb;
  wire [17:0] p2_add_85958_comb;
  wire [11:0] p2_add_85971_comb;
  wire [11:0] p2_add_85972_comb;
  wire [11:0] p2_add_85973_comb;
  wire [11:0] p2_add_85974_comb;
  wire [11:0] p2_add_85987_comb;
  wire [11:0] p2_add_85988_comb;
  wire [11:0] p2_add_85989_comb;
  wire [11:0] p2_add_85990_comb;
  wire [18:0] p2_add_86131_comb;
  wire [18:0] p2_add_86132_comb;
  wire [18:0] p2_add_86133_comb;
  wire [18:0] p2_add_86134_comb;
  wire [18:0] p2_add_86147_comb;
  wire [18:0] p2_add_86148_comb;
  wire [18:0] p2_add_86149_comb;
  wire [18:0] p2_add_86150_comb;
  wire [19:0] p2_smul_84671_comb;
  wire [19:0] p2_smul_84672_comb;
  wire [19:0] p2_smul_84681_comb;
  wire [19:0] p2_smul_84682_comb;
  wire [19:0] p2_smul_84683_comb;
  wire [19:0] p2_smul_84684_comb;
  wire [19:0] p2_smul_84693_comb;
  wire [19:0] p2_smul_84694_comb;
  wire [19:0] p2_smul_84695_comb;
  wire [19:0] p2_smul_84696_comb;
  wire [19:0] p2_smul_84705_comb;
  wire [19:0] p2_smul_84706_comb;
  wire [19:0] p2_smul_84719_comb;
  wire [19:0] p2_smul_84720_comb;
  wire [19:0] p2_smul_84729_comb;
  wire [19:0] p2_smul_84730_comb;
  wire [19:0] p2_smul_84731_comb;
  wire [19:0] p2_smul_84732_comb;
  wire [19:0] p2_smul_84741_comb;
  wire [19:0] p2_smul_84742_comb;
  wire [19:0] p2_smul_84743_comb;
  wire [19:0] p2_smul_84744_comb;
  wire [19:0] p2_smul_84753_comb;
  wire [19:0] p2_smul_84754_comb;
  wire [19:0] p2_smul_85027_comb;
  wire [19:0] p2_smul_85028_comb;
  wire [19:0] p2_smul_85029_comb;
  wire [19:0] p2_smul_85030_comb;
  wire [19:0] p2_smul_85039_comb;
  wire [19:0] p2_smul_85040_comb;
  wire [19:0] p2_smul_85041_comb;
  wire [19:0] p2_smul_85042_comb;
  wire [19:0] p2_smul_85051_comb;
  wire [19:0] p2_smul_85052_comb;
  wire [19:0] p2_smul_85053_comb;
  wire [19:0] p2_smul_85054_comb;
  wire [19:0] p2_smul_85075_comb;
  wire [19:0] p2_smul_85076_comb;
  wire [19:0] p2_smul_85077_comb;
  wire [19:0] p2_smul_85078_comb;
  wire [19:0] p2_smul_85087_comb;
  wire [19:0] p2_smul_85088_comb;
  wire [19:0] p2_smul_85089_comb;
  wire [19:0] p2_smul_85090_comb;
  wire [19:0] p2_smul_85099_comb;
  wire [19:0] p2_smul_85100_comb;
  wire [19:0] p2_smul_85101_comb;
  wire [19:0] p2_smul_85102_comb;
  wire [18:0] p2_bit_slice_85587_comb;
  wire [17:0] p2_add_85588_comb;
  wire [17:0] p2_add_85589_comb;
  wire [18:0] p2_bit_slice_85590_comb;
  wire [17:0] p2_smul_85619_comb;
  wire [17:0] p2_smul_85622_comb;
  wire [17:0] p2_smul_85623_comb;
  wire [17:0] p2_smul_85626_comb;
  wire [18:0] p2_add_85683_comb;
  wire [18:0] p2_add_85685_comb;
  wire [18:0] p2_add_85687_comb;
  wire [18:0] p2_add_85689_comb;
  wire [18:0] p2_add_85811_comb;
  wire [18:0] p2_add_85813_comb;
  wire [18:0] p2_add_85815_comb;
  wire [18:0] p2_add_85817_comb;
  wire [17:0] p2_smul_85876_comb;
  wire [17:0] p2_smul_85878_comb;
  wire [17:0] p2_smul_85879_comb;
  wire [17:0] p2_smul_85881_comb;
  wire [17:0] p2_add_85939_comb;
  wire [18:0] p2_bit_slice_85940_comb;
  wire [18:0] p2_bit_slice_85941_comb;
  wire [17:0] p2_add_85942_comb;
  wire [17:0] p2_add_86067_comb;
  wire [17:0] p2_add_86069_comb;
  wire [17:0] p2_add_86071_comb;
  wire [17:0] p2_add_86073_comb;
  wire [19:0] p2_concat_86115_comb;
  wire [19:0] p2_concat_86116_comb;
  wire [19:0] p2_concat_86117_comb;
  wire [19:0] p2_concat_86118_comb;
  wire [18:0] p2_add_86135_comb;
  wire [18:0] p2_add_86136_comb;
  wire [18:0] p2_add_86137_comb;
  wire [18:0] p2_add_86138_comb;
  wire [18:0] p2_add_86139_comb;
  wire [18:0] p2_add_86140_comb;
  wire [18:0] p2_add_86141_comb;
  wire [18:0] p2_add_86142_comb;
  wire [18:0] p2_add_86143_comb;
  wire [18:0] p2_add_86144_comb;
  wire [18:0] p2_add_86145_comb;
  wire [18:0] p2_add_86146_comb;
  wire [18:0] p2_add_86151_comb;
  wire [18:0] p2_add_86152_comb;
  wire [18:0] p2_add_86153_comb;
  wire [18:0] p2_add_86154_comb;
  wire [18:0] p2_add_86155_comb;
  wire [18:0] p2_add_86156_comb;
  wire [18:0] p2_add_86157_comb;
  wire [18:0] p2_add_86158_comb;
  wire [18:0] p2_add_86159_comb;
  wire [18:0] p2_add_86160_comb;
  wire [18:0] p2_add_86161_comb;
  wire [18:0] p2_add_86162_comb;
  wire [19:0] p2_concat_86179_comb;
  wire [19:0] p2_concat_86180_comb;
  wire [19:0] p2_concat_86181_comb;
  wire [19:0] p2_concat_86182_comb;
  wire [17:0] p2_add_86227_comb;
  wire [17:0] p2_add_86229_comb;
  wire [17:0] p2_add_86231_comb;
  wire [17:0] p2_add_86233_comb;
  wire [24:0] p2_sum__1568_comb;
  wire [24:0] p2_sum__1569_comb;
  wire [24:0] p2_sum__1570_comb;
  wire [24:0] p2_sum__1571_comb;
  wire [24:0] p2_sum__1456_comb;
  wire [24:0] p2_sum__1457_comb;
  wire [24:0] p2_sum__1458_comb;
  wire [24:0] p2_sum__1459_comb;
  wire [19:0] p2_smul_84829_comb;
  wire [19:0] p2_smul_84831_comb;
  wire [19:0] p2_smul_84836_comb;
  wire [19:0] p2_smul_84838_comb;
  wire [19:0] p2_smul_84839_comb;
  wire [19:0] p2_smul_84841_comb;
  wire [19:0] p2_smul_84846_comb;
  wire [19:0] p2_smul_84848_comb;
  wire [19:0] p2_smul_84849_comb;
  wire [19:0] p2_smul_84851_comb;
  wire [19:0] p2_smul_84856_comb;
  wire [19:0] p2_smul_84858_comb;
  wire [19:0] p2_smul_84869_comb;
  wire [19:0] p2_smul_84871_comb;
  wire [19:0] p2_smul_84876_comb;
  wire [19:0] p2_smul_84878_comb;
  wire [19:0] p2_smul_84879_comb;
  wire [19:0] p2_smul_84881_comb;
  wire [19:0] p2_smul_84886_comb;
  wire [19:0] p2_smul_84888_comb;
  wire [19:0] p2_smul_84889_comb;
  wire [19:0] p2_smul_84891_comb;
  wire [19:0] p2_smul_84896_comb;
  wire [19:0] p2_smul_84898_comb;
  wire [19:0] p2_smul_84911_comb;
  wire [19:0] p2_smul_84913_comb;
  wire [19:0] p2_smul_84914_comb;
  wire [19:0] p2_smul_84916_comb;
  wire [19:0] p2_smul_84921_comb;
  wire [19:0] p2_smul_84923_comb;
  wire [19:0] p2_smul_84924_comb;
  wire [19:0] p2_smul_84926_comb;
  wire [19:0] p2_smul_84931_comb;
  wire [19:0] p2_smul_84933_comb;
  wire [19:0] p2_smul_84934_comb;
  wire [19:0] p2_smul_84936_comb;
  wire [19:0] p2_smul_84951_comb;
  wire [19:0] p2_smul_84953_comb;
  wire [19:0] p2_smul_84954_comb;
  wire [19:0] p2_smul_84956_comb;
  wire [19:0] p2_smul_84961_comb;
  wire [19:0] p2_smul_84963_comb;
  wire [19:0] p2_smul_84964_comb;
  wire [19:0] p2_smul_84966_comb;
  wire [19:0] p2_smul_84971_comb;
  wire [19:0] p2_smul_84973_comb;
  wire [19:0] p2_smul_84974_comb;
  wire [19:0] p2_smul_84976_comb;
  wire [19:0] p2_add_85113_comb;
  wire [17:0] p2_smul_85114_comb;
  wire [17:0] p2_smul_85115_comb;
  wire [17:0] p2_smul_85116_comb;
  wire [17:0] p2_smul_85117_comb;
  wire [19:0] p2_add_85118_comb;
  wire [19:0] p2_add_85119_comb;
  wire [17:0] p2_smul_85120_comb;
  wire [17:0] p2_smul_85121_comb;
  wire [17:0] p2_smul_85122_comb;
  wire [17:0] p2_smul_85123_comb;
  wire [19:0] p2_add_85124_comb;
  wire [19:0] p2_add_85125_comb;
  wire [17:0] p2_smul_85126_comb;
  wire [17:0] p2_smul_85127_comb;
  wire [17:0] p2_smul_85128_comb;
  wire [17:0] p2_smul_85129_comb;
  wire [19:0] p2_add_85130_comb;
  wire [19:0] p2_add_85137_comb;
  wire [17:0] p2_smul_85138_comb;
  wire [17:0] p2_smul_85139_comb;
  wire [17:0] p2_smul_85140_comb;
  wire [17:0] p2_smul_85141_comb;
  wire [19:0] p2_add_85142_comb;
  wire [19:0] p2_add_85143_comb;
  wire [17:0] p2_smul_85144_comb;
  wire [17:0] p2_smul_85145_comb;
  wire [17:0] p2_smul_85146_comb;
  wire [17:0] p2_smul_85147_comb;
  wire [19:0] p2_add_85148_comb;
  wire [19:0] p2_add_85149_comb;
  wire [17:0] p2_smul_85150_comb;
  wire [17:0] p2_smul_85151_comb;
  wire [17:0] p2_smul_85152_comb;
  wire [17:0] p2_smul_85153_comb;
  wire [19:0] p2_add_85154_comb;
  wire [18:0] p2_smul_85164_comb;
  wire [18:0] p2_smul_85165_comb;
  wire [18:0] p2_smul_85168_comb;
  wire [18:0] p2_smul_85169_comb;
  wire [18:0] p2_smul_85172_comb;
  wire [18:0] p2_smul_85173_comb;
  wire [18:0] p2_smul_85176_comb;
  wire [18:0] p2_smul_85177_comb;
  wire [18:0] p2_smul_85180_comb;
  wire [18:0] p2_smul_85181_comb;
  wire [18:0] p2_smul_85184_comb;
  wire [18:0] p2_smul_85185_comb;
  wire [18:0] p2_smul_85196_comb;
  wire [18:0] p2_smul_85197_comb;
  wire [18:0] p2_smul_85200_comb;
  wire [18:0] p2_smul_85201_comb;
  wire [18:0] p2_smul_85204_comb;
  wire [18:0] p2_smul_85205_comb;
  wire [18:0] p2_smul_85208_comb;
  wire [18:0] p2_smul_85209_comb;
  wire [18:0] p2_smul_85212_comb;
  wire [18:0] p2_smul_85213_comb;
  wire [18:0] p2_smul_85216_comb;
  wire [18:0] p2_smul_85217_comb;
  wire [18:0] p2_smul_85419_comb;
  wire [18:0] p2_smul_85421_comb;
  wire [18:0] p2_smul_85424_comb;
  wire [18:0] p2_smul_85426_comb;
  wire [18:0] p2_smul_85427_comb;
  wire [18:0] p2_smul_85429_comb;
  wire [18:0] p2_smul_85432_comb;
  wire [18:0] p2_smul_85434_comb;
  wire [18:0] p2_smul_85435_comb;
  wire [18:0] p2_smul_85437_comb;
  wire [18:0] p2_smul_85440_comb;
  wire [18:0] p2_smul_85442_comb;
  wire [18:0] p2_smul_85451_comb;
  wire [18:0] p2_smul_85453_comb;
  wire [18:0] p2_smul_85456_comb;
  wire [18:0] p2_smul_85458_comb;
  wire [18:0] p2_smul_85459_comb;
  wire [18:0] p2_smul_85461_comb;
  wire [18:0] p2_smul_85464_comb;
  wire [18:0] p2_smul_85466_comb;
  wire [18:0] p2_smul_85467_comb;
  wire [18:0] p2_smul_85469_comb;
  wire [18:0] p2_smul_85472_comb;
  wire [18:0] p2_smul_85474_comb;
  wire [17:0] p2_smul_85481_comb;
  wire [17:0] p2_smul_85482_comb;
  wire [19:0] p2_add_85483_comb;
  wire [19:0] p2_add_85484_comb;
  wire [17:0] p2_smul_85485_comb;
  wire [17:0] p2_smul_85486_comb;
  wire [17:0] p2_smul_85487_comb;
  wire [17:0] p2_smul_85488_comb;
  wire [19:0] p2_add_85489_comb;
  wire [19:0] p2_add_85490_comb;
  wire [17:0] p2_smul_85491_comb;
  wire [17:0] p2_smul_85492_comb;
  wire [17:0] p2_smul_85493_comb;
  wire [17:0] p2_smul_85494_comb;
  wire [19:0] p2_add_85495_comb;
  wire [19:0] p2_add_85496_comb;
  wire [17:0] p2_smul_85497_comb;
  wire [17:0] p2_smul_85498_comb;
  wire [17:0] p2_smul_85505_comb;
  wire [17:0] p2_smul_85506_comb;
  wire [19:0] p2_add_85507_comb;
  wire [19:0] p2_add_85508_comb;
  wire [17:0] p2_smul_85509_comb;
  wire [17:0] p2_smul_85510_comb;
  wire [17:0] p2_smul_85511_comb;
  wire [17:0] p2_smul_85512_comb;
  wire [19:0] p2_add_85513_comb;
  wire [19:0] p2_add_85514_comb;
  wire [17:0] p2_smul_85515_comb;
  wire [17:0] p2_smul_85516_comb;
  wire [17:0] p2_smul_85517_comb;
  wire [17:0] p2_smul_85518_comb;
  wire [19:0] p2_add_85519_comb;
  wire [19:0] p2_add_85520_comb;
  wire [17:0] p2_smul_85521_comb;
  wire [17:0] p2_smul_85522_comb;
  wire [11:0] p2_add_85975_comb;
  wire [11:0] p2_add_85976_comb;
  wire [11:0] p2_add_85977_comb;
  wire [11:0] p2_add_85978_comb;
  wire [11:0] p2_add_85979_comb;
  wire [11:0] p2_add_85980_comb;
  wire [11:0] p2_add_85981_comb;
  wire [11:0] p2_add_85982_comb;
  wire [11:0] p2_add_85983_comb;
  wire [11:0] p2_add_85984_comb;
  wire [11:0] p2_add_85985_comb;
  wire [11:0] p2_add_85986_comb;
  wire [11:0] p2_add_85991_comb;
  wire [11:0] p2_add_85992_comb;
  wire [11:0] p2_add_85993_comb;
  wire [11:0] p2_add_85994_comb;
  wire [11:0] p2_add_85995_comb;
  wire [11:0] p2_add_85996_comb;
  wire [11:0] p2_add_85997_comb;
  wire [11:0] p2_add_85998_comb;
  wire [11:0] p2_add_85999_comb;
  wire [11:0] p2_add_86000_comb;
  wire [11:0] p2_add_86001_comb;
  wire [11:0] p2_add_86002_comb;
  wire [17:0] p2_add_86035_comb;
  wire [17:0] p2_add_86037_comb;
  wire [17:0] p2_add_86039_comb;
  wire [17:0] p2_add_86041_comb;
  wire [19:0] p2_concat_86099_comb;
  wire [19:0] p2_concat_86100_comb;
  wire [19:0] p2_concat_86101_comb;
  wire [19:0] p2_concat_86102_comb;
  wire [19:0] p2_concat_86163_comb;
  wire [19:0] p2_concat_86164_comb;
  wire [19:0] p2_concat_86165_comb;
  wire [19:0] p2_concat_86166_comb;
  wire [17:0] p2_add_86195_comb;
  wire [17:0] p2_add_86197_comb;
  wire [17:0] p2_add_86199_comb;
  wire [17:0] p2_add_86201_comb;
  wire [23:0] p2_add_86339_comb;
  wire [23:0] p2_add_86341_comb;
  wire [18:0] p2_concat_86371_comb;
  wire [18:0] p2_concat_86372_comb;
  wire [18:0] p2_concat_86373_comb;
  wire [18:0] p2_concat_86374_comb;
  wire [24:0] p2_sum__1460_comb;
  wire [24:0] p2_sum__1461_comb;
  wire [24:0] p2_sum__1462_comb;
  wire [24:0] p2_sum__1463_comb;
  wire [24:0] p2_sum__1540_comb;
  wire [24:0] p2_sum__1541_comb;
  wire [24:0] p2_sum__1542_comb;
  wire [24:0] p2_sum__1543_comb;
  wire [24:0] p2_sum__1512_comb;
  wire [24:0] p2_sum__1513_comb;
  wire [24:0] p2_sum__1514_comb;
  wire [24:0] p2_sum__1515_comb;
  wire [24:0] p2_sum__1484_comb;
  wire [24:0] p2_sum__1485_comb;
  wire [24:0] p2_sum__1486_comb;
  wire [24:0] p2_sum__1487_comb;
  wire [24:0] p2_sum__1428_comb;
  wire [24:0] p2_sum__1429_comb;
  wire [24:0] p2_sum__1430_comb;
  wire [24:0] p2_sum__1431_comb;
  wire [24:0] p2_sum__1400_comb;
  wire [24:0] p2_sum__1401_comb;
  wire [24:0] p2_sum__1402_comb;
  wire [24:0] p2_sum__1403_comb;
  wire [24:0] p2_sum__1372_comb;
  wire [24:0] p2_sum__1373_comb;
  wire [24:0] p2_sum__1374_comb;
  wire [24:0] p2_sum__1375_comb;
  wire [24:0] p2_sum__1452_comb;
  wire [24:0] p2_sum__1453_comb;
  wire [24:0] p2_sum__1454_comb;
  wire [24:0] p2_sum__1455_comb;
  wire [18:0] p2_concat_86451_comb;
  wire [18:0] p2_concat_86452_comb;
  wire [18:0] p2_concat_86453_comb;
  wire [18:0] p2_concat_86454_comb;
  wire [23:0] p2_add_86483_comb;
  wire [23:0] p2_add_86485_comb;
  wire [23:0] p2_add_86499_comb;
  wire [23:0] p2_add_86500_comb;
  wire [23:0] p2_add_86507_comb;
  wire [23:0] p2_add_86508_comb;
  wire [24:0] p2_sum__1240_comb;
  wire [24:0] p2_sum__1241_comb;
  wire [24:0] p2_sum__1184_comb;
  wire [24:0] p2_sum__1185_comb;
  wire [18:0] p2_smul_85228_comb;
  wire [18:0] p2_smul_85230_comb;
  wire [18:0] p2_smul_85231_comb;
  wire [18:0] p2_smul_85233_comb;
  wire [18:0] p2_smul_85236_comb;
  wire [18:0] p2_smul_85238_comb;
  wire [18:0] p2_smul_85239_comb;
  wire [18:0] p2_smul_85241_comb;
  wire [18:0] p2_smul_85244_comb;
  wire [18:0] p2_smul_85246_comb;
  wire [18:0] p2_smul_85247_comb;
  wire [18:0] p2_smul_85249_comb;
  wire [18:0] p2_smul_85260_comb;
  wire [18:0] p2_smul_85262_comb;
  wire [18:0] p2_smul_85263_comb;
  wire [18:0] p2_smul_85265_comb;
  wire [18:0] p2_smul_85268_comb;
  wire [18:0] p2_smul_85270_comb;
  wire [18:0] p2_smul_85271_comb;
  wire [18:0] p2_smul_85273_comb;
  wire [18:0] p2_smul_85276_comb;
  wire [18:0] p2_smul_85278_comb;
  wire [18:0] p2_smul_85279_comb;
  wire [18:0] p2_smul_85281_comb;
  wire [18:0] p2_smul_85355_comb;
  wire [18:0] p2_smul_85357_comb;
  wire [18:0] p2_smul_85360_comb;
  wire [18:0] p2_smul_85362_comb;
  wire [18:0] p2_smul_85363_comb;
  wire [18:0] p2_smul_85365_comb;
  wire [18:0] p2_smul_85368_comb;
  wire [18:0] p2_smul_85370_comb;
  wire [18:0] p2_smul_85371_comb;
  wire [18:0] p2_smul_85373_comb;
  wire [18:0] p2_smul_85376_comb;
  wire [18:0] p2_smul_85378_comb;
  wire [18:0] p2_smul_85387_comb;
  wire [18:0] p2_smul_85389_comb;
  wire [18:0] p2_smul_85392_comb;
  wire [18:0] p2_smul_85394_comb;
  wire [18:0] p2_smul_85395_comb;
  wire [18:0] p2_smul_85397_comb;
  wire [18:0] p2_smul_85400_comb;
  wire [18:0] p2_smul_85402_comb;
  wire [18:0] p2_smul_85403_comb;
  wire [18:0] p2_smul_85405_comb;
  wire [18:0] p2_smul_85408_comb;
  wire [18:0] p2_smul_85410_comb;
  wire [18:0] p2_bit_slice_85591_comb;
  wire [17:0] p2_add_85592_comb;
  wire [17:0] p2_add_85593_comb;
  wire [18:0] p2_bit_slice_85594_comb;
  wire [18:0] p2_bit_slice_85595_comb;
  wire [17:0] p2_add_85596_comb;
  wire [17:0] p2_add_85597_comb;
  wire [18:0] p2_bit_slice_85598_comb;
  wire [18:0] p2_bit_slice_85599_comb;
  wire [17:0] p2_add_85600_comb;
  wire [17:0] p2_add_85601_comb;
  wire [18:0] p2_bit_slice_85602_comb;
  wire [18:0] p2_bit_slice_85607_comb;
  wire [17:0] p2_add_85608_comb;
  wire [17:0] p2_add_85609_comb;
  wire [18:0] p2_bit_slice_85610_comb;
  wire [18:0] p2_bit_slice_85611_comb;
  wire [17:0] p2_add_85612_comb;
  wire [17:0] p2_add_85613_comb;
  wire [18:0] p2_bit_slice_85614_comb;
  wire [18:0] p2_bit_slice_85615_comb;
  wire [17:0] p2_add_85616_comb;
  wire [17:0] p2_add_85617_comb;
  wire [18:0] p2_bit_slice_85618_comb;
  wire [17:0] p2_smul_85627_comb;
  wire [17:0] p2_smul_85630_comb;
  wire [17:0] p2_smul_85631_comb;
  wire [17:0] p2_smul_85634_comb;
  wire [17:0] p2_smul_85635_comb;
  wire [17:0] p2_smul_85638_comb;
  wire [17:0] p2_smul_85639_comb;
  wire [17:0] p2_smul_85642_comb;
  wire [17:0] p2_smul_85643_comb;
  wire [17:0] p2_smul_85646_comb;
  wire [17:0] p2_smul_85647_comb;
  wire [17:0] p2_smul_85650_comb;
  wire [17:0] p2_smul_85659_comb;
  wire [17:0] p2_smul_85662_comb;
  wire [17:0] p2_smul_85663_comb;
  wire [17:0] p2_smul_85666_comb;
  wire [17:0] p2_smul_85667_comb;
  wire [17:0] p2_smul_85670_comb;
  wire [17:0] p2_smul_85671_comb;
  wire [17:0] p2_smul_85674_comb;
  wire [17:0] p2_smul_85675_comb;
  wire [17:0] p2_smul_85678_comb;
  wire [17:0] p2_smul_85679_comb;
  wire [17:0] p2_smul_85682_comb;
  wire [17:0] p2_smul_85884_comb;
  wire [17:0] p2_smul_85886_comb;
  wire [17:0] p2_smul_85887_comb;
  wire [17:0] p2_smul_85889_comb;
  wire [17:0] p2_smul_85892_comb;
  wire [17:0] p2_smul_85894_comb;
  wire [17:0] p2_smul_85895_comb;
  wire [17:0] p2_smul_85897_comb;
  wire [17:0] p2_smul_85900_comb;
  wire [17:0] p2_smul_85902_comb;
  wire [17:0] p2_smul_85903_comb;
  wire [17:0] p2_smul_85905_comb;
  wire [17:0] p2_smul_85916_comb;
  wire [17:0] p2_smul_85918_comb;
  wire [17:0] p2_smul_85919_comb;
  wire [17:0] p2_smul_85921_comb;
  wire [17:0] p2_smul_85924_comb;
  wire [17:0] p2_smul_85926_comb;
  wire [17:0] p2_smul_85927_comb;
  wire [17:0] p2_smul_85929_comb;
  wire [17:0] p2_smul_85932_comb;
  wire [17:0] p2_smul_85934_comb;
  wire [17:0] p2_smul_85935_comb;
  wire [17:0] p2_smul_85937_comb;
  wire [17:0] p2_add_85943_comb;
  wire [18:0] p2_bit_slice_85944_comb;
  wire [18:0] p2_bit_slice_85945_comb;
  wire [17:0] p2_add_85946_comb;
  wire [17:0] p2_add_85947_comb;
  wire [18:0] p2_bit_slice_85948_comb;
  wire [18:0] p2_bit_slice_85949_comb;
  wire [17:0] p2_add_85950_comb;
  wire [17:0] p2_add_85951_comb;
  wire [18:0] p2_bit_slice_85952_comb;
  wire [18:0] p2_bit_slice_85953_comb;
  wire [17:0] p2_add_85954_comb;
  wire [17:0] p2_add_85959_comb;
  wire [18:0] p2_bit_slice_85960_comb;
  wire [18:0] p2_bit_slice_85961_comb;
  wire [17:0] p2_add_85962_comb;
  wire [17:0] p2_add_85963_comb;
  wire [18:0] p2_bit_slice_85964_comb;
  wire [18:0] p2_bit_slice_85965_comb;
  wire [17:0] p2_add_85966_comb;
  wire [17:0] p2_add_85967_comb;
  wire [18:0] p2_bit_slice_85968_comb;
  wire [18:0] p2_bit_slice_85969_comb;
  wire [17:0] p2_add_85970_comb;
  wire [23:0] p2_add_86323_comb;
  wire [23:0] p2_add_86325_comb;
  wire [18:0] p2_concat_86355_comb;
  wire [18:0] p2_concat_86356_comb;
  wire [18:0] p2_concat_86357_comb;
  wire [18:0] p2_concat_86358_comb;
  wire [24:0] p2_sum__1572_comb;
  wire [24:0] p2_sum__1573_comb;
  wire [24:0] p2_sum__1574_comb;
  wire [24:0] p2_sum__1575_comb;
  wire [24:0] p2_sum__1564_comb;
  wire [24:0] p2_sum__1565_comb;
  wire [24:0] p2_sum__1566_comb;
  wire [24:0] p2_sum__1567_comb;
  wire [18:0] p2_concat_86435_comb;
  wire [18:0] p2_concat_86436_comb;
  wire [18:0] p2_concat_86437_comb;
  wire [18:0] p2_concat_86438_comb;
  wire [23:0] p2_add_86467_comb;
  wire [23:0] p2_add_86469_comb;
  wire [24:0] p2_sum__1190_comb;
  wire [24:0] p2_sum__1191_comb;
  wire [24:0] p2_sum__1186_comb;
  wire [24:0] p2_sum__1187_comb;
  wire [24:0] p2_sum__1226_comb;
  wire [24:0] p2_sum__1227_comb;
  wire [24:0] p2_sum__1212_comb;
  wire [24:0] p2_sum__1213_comb;
  wire [24:0] p2_sum__1198_comb;
  wire [24:0] p2_sum__1199_comb;
  wire [24:0] p2_sum__1170_comb;
  wire [24:0] p2_sum__1171_comb;
  wire [24:0] p2_sum__1156_comb;
  wire [24:0] p2_sum__1157_comb;
  wire [24:0] p2_sum__1142_comb;
  wire [24:0] p2_sum__1143_comb;
  wire [24:0] p2_sum__1182_comb;
  wire [24:0] p2_sum__1183_comb;
  wire [24:0] p2_sum__1178_comb;
  wire [24:0] p2_sum__1179_comb;
  wire [23:0] p2_add_86563_comb;
  wire [23:0] p2_add_86568_comb;
  wire [24:0] p2_sum__1076_comb;
  wire [24:0] p2_sum__1048_comb;
  wire [18:0] p2_add_85691_comb;
  wire [18:0] p2_add_85693_comb;
  wire [18:0] p2_add_85695_comb;
  wire [18:0] p2_add_85697_comb;
  wire [18:0] p2_add_85699_comb;
  wire [18:0] p2_add_85701_comb;
  wire [18:0] p2_add_85703_comb;
  wire [18:0] p2_add_85705_comb;
  wire [18:0] p2_add_85707_comb;
  wire [18:0] p2_add_85709_comb;
  wire [18:0] p2_add_85711_comb;
  wire [18:0] p2_add_85713_comb;
  wire [18:0] p2_add_85723_comb;
  wire [18:0] p2_add_85725_comb;
  wire [18:0] p2_add_85727_comb;
  wire [18:0] p2_add_85729_comb;
  wire [18:0] p2_add_85731_comb;
  wire [18:0] p2_add_85733_comb;
  wire [18:0] p2_add_85735_comb;
  wire [18:0] p2_add_85737_comb;
  wire [18:0] p2_add_85739_comb;
  wire [18:0] p2_add_85741_comb;
  wire [18:0] p2_add_85743_comb;
  wire [18:0] p2_add_85745_comb;
  wire [18:0] p2_add_85819_comb;
  wire [18:0] p2_add_85821_comb;
  wire [18:0] p2_add_85823_comb;
  wire [18:0] p2_add_85825_comb;
  wire [18:0] p2_add_85827_comb;
  wire [18:0] p2_add_85829_comb;
  wire [18:0] p2_add_85831_comb;
  wire [18:0] p2_add_85833_comb;
  wire [18:0] p2_add_85835_comb;
  wire [18:0] p2_add_85837_comb;
  wire [18:0] p2_add_85839_comb;
  wire [18:0] p2_add_85841_comb;
  wire [18:0] p2_add_85851_comb;
  wire [18:0] p2_add_85853_comb;
  wire [18:0] p2_add_85855_comb;
  wire [18:0] p2_add_85857_comb;
  wire [18:0] p2_add_85859_comb;
  wire [18:0] p2_add_85861_comb;
  wire [18:0] p2_add_85863_comb;
  wire [18:0] p2_add_85865_comb;
  wire [18:0] p2_add_85867_comb;
  wire [18:0] p2_add_85869_comb;
  wire [18:0] p2_add_85871_comb;
  wire [18:0] p2_add_85873_comb;
  wire [17:0] p2_add_86043_comb;
  wire [17:0] p2_add_86045_comb;
  wire [17:0] p2_add_86047_comb;
  wire [17:0] p2_add_86049_comb;
  wire [17:0] p2_add_86051_comb;
  wire [17:0] p2_add_86053_comb;
  wire [17:0] p2_add_86055_comb;
  wire [17:0] p2_add_86057_comb;
  wire [17:0] p2_add_86059_comb;
  wire [17:0] p2_add_86061_comb;
  wire [17:0] p2_add_86063_comb;
  wire [17:0] p2_add_86065_comb;
  wire [17:0] p2_add_86075_comb;
  wire [17:0] p2_add_86077_comb;
  wire [17:0] p2_add_86079_comb;
  wire [17:0] p2_add_86081_comb;
  wire [17:0] p2_add_86083_comb;
  wire [17:0] p2_add_86085_comb;
  wire [17:0] p2_add_86087_comb;
  wire [17:0] p2_add_86089_comb;
  wire [17:0] p2_add_86091_comb;
  wire [17:0] p2_add_86093_comb;
  wire [17:0] p2_add_86095_comb;
  wire [17:0] p2_add_86097_comb;
  wire [17:0] p2_add_86203_comb;
  wire [17:0] p2_add_86205_comb;
  wire [17:0] p2_add_86207_comb;
  wire [17:0] p2_add_86209_comb;
  wire [17:0] p2_add_86211_comb;
  wire [17:0] p2_add_86213_comb;
  wire [17:0] p2_add_86215_comb;
  wire [17:0] p2_add_86217_comb;
  wire [17:0] p2_add_86219_comb;
  wire [17:0] p2_add_86221_comb;
  wire [17:0] p2_add_86223_comb;
  wire [17:0] p2_add_86225_comb;
  wire [17:0] p2_add_86235_comb;
  wire [17:0] p2_add_86237_comb;
  wire [17:0] p2_add_86239_comb;
  wire [17:0] p2_add_86241_comb;
  wire [17:0] p2_add_86243_comb;
  wire [17:0] p2_add_86245_comb;
  wire [17:0] p2_add_86247_comb;
  wire [17:0] p2_add_86249_comb;
  wire [17:0] p2_add_86251_comb;
  wire [17:0] p2_add_86253_comb;
  wire [17:0] p2_add_86255_comb;
  wire [17:0] p2_add_86257_comb;
  wire [23:0] p2_add_86501_comb;
  wire [23:0] p2_add_86502_comb;
  wire [23:0] p2_add_86503_comb;
  wire [23:0] p2_add_86504_comb;
  wire [23:0] p2_add_86505_comb;
  wire [23:0] p2_add_86506_comb;
  wire [23:0] p2_add_86509_comb;
  wire [23:0] p2_add_86510_comb;
  wire [23:0] p2_add_86511_comb;
  wire [23:0] p2_add_86512_comb;
  wire [23:0] p2_add_86513_comb;
  wire [23:0] p2_add_86514_comb;
  wire [24:0] p2_sum__1246_comb;
  wire [24:0] p2_sum__1247_comb;
  wire [24:0] p2_sum__1242_comb;
  wire [24:0] p2_sum__1243_comb;
  wire [24:0] p2_sum__1238_comb;
  wire [24:0] p2_sum__1239_comb;
  wire [24:0] p2_sum__1234_comb;
  wire [24:0] p2_sum__1235_comb;
  wire [24:0] p2_sum__1051_comb;
  wire [23:0] p2_add_86578_comb;
  wire [23:0] p2_add_86579_comb;
  wire [24:0] p2_sum__1049_comb;
  wire [24:0] p2_sum__1069_comb;
  wire [24:0] p2_sum__1062_comb;
  wire [24:0] p2_sum__1055_comb;
  wire [24:0] p2_sum__1041_comb;
  wire [24:0] p2_sum__1034_comb;
  wire [24:0] p2_sum__1027_comb;
  wire [24:0] p2_sum__1047_comb;
  wire [23:0] p2_add_86604_comb;
  wire [23:0] p2_add_86605_comb;
  wire [24:0] p2_sum__1045_comb;
  wire [23:0] p2_umul_29016_NarrowedMult__comb;
  wire [23:0] p2_umul_29024_NarrowedMult__comb;
  wire [24:0] p2_add_86614_comb;
  wire [24:0] p2_add_86618_comb;
  wire [19:0] p2_concat_86103_comb;
  wire [19:0] p2_concat_86104_comb;
  wire [19:0] p2_concat_86105_comb;
  wire [19:0] p2_concat_86106_comb;
  wire [19:0] p2_concat_86107_comb;
  wire [19:0] p2_concat_86108_comb;
  wire [19:0] p2_concat_86109_comb;
  wire [19:0] p2_concat_86110_comb;
  wire [19:0] p2_concat_86111_comb;
  wire [19:0] p2_concat_86112_comb;
  wire [19:0] p2_concat_86113_comb;
  wire [19:0] p2_concat_86114_comb;
  wire [19:0] p2_concat_86119_comb;
  wire [19:0] p2_concat_86120_comb;
  wire [19:0] p2_concat_86121_comb;
  wire [19:0] p2_concat_86122_comb;
  wire [19:0] p2_concat_86123_comb;
  wire [19:0] p2_concat_86124_comb;
  wire [19:0] p2_concat_86125_comb;
  wire [19:0] p2_concat_86126_comb;
  wire [19:0] p2_concat_86127_comb;
  wire [19:0] p2_concat_86128_comb;
  wire [19:0] p2_concat_86129_comb;
  wire [19:0] p2_concat_86130_comb;
  wire [19:0] p2_concat_86167_comb;
  wire [19:0] p2_concat_86168_comb;
  wire [19:0] p2_concat_86169_comb;
  wire [19:0] p2_concat_86170_comb;
  wire [19:0] p2_concat_86171_comb;
  wire [19:0] p2_concat_86172_comb;
  wire [19:0] p2_concat_86173_comb;
  wire [19:0] p2_concat_86174_comb;
  wire [19:0] p2_concat_86175_comb;
  wire [19:0] p2_concat_86176_comb;
  wire [19:0] p2_concat_86177_comb;
  wire [19:0] p2_concat_86178_comb;
  wire [19:0] p2_concat_86183_comb;
  wire [19:0] p2_concat_86184_comb;
  wire [19:0] p2_concat_86185_comb;
  wire [19:0] p2_concat_86186_comb;
  wire [19:0] p2_concat_86187_comb;
  wire [19:0] p2_concat_86188_comb;
  wire [19:0] p2_concat_86189_comb;
  wire [19:0] p2_concat_86190_comb;
  wire [19:0] p2_concat_86191_comb;
  wire [19:0] p2_concat_86192_comb;
  wire [19:0] p2_concat_86193_comb;
  wire [19:0] p2_concat_86194_comb;
  wire [23:0] p2_add_86327_comb;
  wire p2_bit_slice_86328_comb;
  wire [23:0] p2_add_86329_comb;
  wire p2_bit_slice_86330_comb;
  wire [23:0] p2_add_86331_comb;
  wire p2_bit_slice_86332_comb;
  wire [23:0] p2_add_86333_comb;
  wire p2_bit_slice_86334_comb;
  wire [23:0] p2_add_86335_comb;
  wire p2_bit_slice_86336_comb;
  wire [23:0] p2_add_86337_comb;
  wire p2_bit_slice_86338_comb;
  wire [23:0] p2_add_86343_comb;
  wire p2_bit_slice_86344_comb;
  wire [23:0] p2_add_86345_comb;
  wire p2_bit_slice_86346_comb;
  wire [23:0] p2_add_86347_comb;
  wire p2_bit_slice_86348_comb;
  wire [23:0] p2_add_86349_comb;
  wire p2_bit_slice_86350_comb;
  wire [23:0] p2_add_86351_comb;
  wire p2_bit_slice_86352_comb;
  wire [23:0] p2_add_86353_comb;
  wire p2_bit_slice_86354_comb;
  wire [18:0] p2_concat_86359_comb;
  wire [18:0] p2_concat_86360_comb;
  wire [18:0] p2_concat_86361_comb;
  wire [18:0] p2_concat_86362_comb;
  wire [18:0] p2_concat_86363_comb;
  wire [18:0] p2_concat_86364_comb;
  wire [18:0] p2_concat_86365_comb;
  wire [18:0] p2_concat_86366_comb;
  wire [18:0] p2_concat_86367_comb;
  wire [18:0] p2_concat_86368_comb;
  wire [18:0] p2_concat_86369_comb;
  wire [18:0] p2_concat_86370_comb;
  wire [18:0] p2_concat_86375_comb;
  wire [18:0] p2_concat_86376_comb;
  wire [18:0] p2_concat_86377_comb;
  wire [18:0] p2_concat_86378_comb;
  wire [18:0] p2_concat_86379_comb;
  wire [18:0] p2_concat_86380_comb;
  wire [18:0] p2_concat_86381_comb;
  wire [18:0] p2_concat_86382_comb;
  wire [18:0] p2_concat_86383_comb;
  wire [18:0] p2_concat_86384_comb;
  wire [18:0] p2_concat_86385_comb;
  wire [18:0] p2_concat_86386_comb;
  wire [18:0] p2_concat_86439_comb;
  wire [18:0] p2_concat_86440_comb;
  wire [18:0] p2_concat_86441_comb;
  wire [18:0] p2_concat_86442_comb;
  wire [18:0] p2_concat_86443_comb;
  wire [18:0] p2_concat_86444_comb;
  wire [18:0] p2_concat_86445_comb;
  wire [18:0] p2_concat_86446_comb;
  wire [18:0] p2_concat_86447_comb;
  wire [18:0] p2_concat_86448_comb;
  wire [18:0] p2_concat_86449_comb;
  wire [18:0] p2_concat_86450_comb;
  wire [18:0] p2_concat_86455_comb;
  wire [18:0] p2_concat_86456_comb;
  wire [18:0] p2_concat_86457_comb;
  wire [18:0] p2_concat_86458_comb;
  wire [18:0] p2_concat_86459_comb;
  wire [18:0] p2_concat_86460_comb;
  wire [18:0] p2_concat_86461_comb;
  wire [18:0] p2_concat_86462_comb;
  wire [18:0] p2_concat_86463_comb;
  wire [18:0] p2_concat_86464_comb;
  wire [18:0] p2_concat_86465_comb;
  wire [18:0] p2_concat_86466_comb;
  wire [23:0] p2_add_86471_comb;
  wire p2_bit_slice_86472_comb;
  wire [23:0] p2_add_86473_comb;
  wire p2_bit_slice_86474_comb;
  wire [23:0] p2_add_86475_comb;
  wire p2_bit_slice_86476_comb;
  wire [23:0] p2_add_86477_comb;
  wire p2_bit_slice_86478_comb;
  wire [23:0] p2_add_86479_comb;
  wire p2_bit_slice_86480_comb;
  wire [23:0] p2_add_86481_comb;
  wire p2_bit_slice_86482_comb;
  wire [23:0] p2_add_86487_comb;
  wire p2_bit_slice_86488_comb;
  wire [23:0] p2_add_86489_comb;
  wire p2_bit_slice_86490_comb;
  wire [23:0] p2_add_86491_comb;
  wire p2_bit_slice_86492_comb;
  wire [23:0] p2_add_86493_comb;
  wire p2_bit_slice_86494_comb;
  wire [23:0] p2_add_86495_comb;
  wire p2_bit_slice_86496_comb;
  wire [23:0] p2_add_86497_comb;
  wire p2_bit_slice_86498_comb;
  wire [23:0] p2_add_86565_comb;
  wire [23:0] p2_add_86566_comb;
  wire [23:0] p2_add_86567_comb;
  wire [23:0] p2_add_86570_comb;
  wire [23:0] p2_add_86571_comb;
  wire [23:0] p2_add_86572_comb;
  wire [24:0] p2_sum__1079_comb;
  wire [23:0] p2_add_86576_comb;
  wire [23:0] p2_add_86577_comb;
  wire [24:0] p2_sum__1077_comb;
  wire [24:0] p2_sum__1075_comb;
  wire [23:0] p2_add_86602_comb;
  wire [23:0] p2_add_86603_comb;
  wire [24:0] p2_sum__1073_comb;
  wire [24:0] p2_add_86611_comb;
  wire [23:0] p2_add_86612_comb;
  wire [24:0] p2_add_86613_comb;
  wire [24:0] p2_add_86615_comb;
  wire [24:0] p2_add_86616_comb;
  wire [24:0] p2_add_86617_comb;
  wire [24:0] p2_add_86619_comb;
  wire [24:0] p2_add_86620_comb;
  wire [24:0] p2_add_86621_comb;
  wire [24:0] p2_add_86622_comb;
  wire [23:0] p2_add_86623_comb;
  wire [24:0] p2_add_86624_comb;
  wire [16:0] p2_bit_slice_86625_comb;
  wire [16:0] p2_bit_slice_86626_comb;
  wire [16:0] p2_bit_slice_86627_comb;
  wire [16:0] p2_bit_slice_86628_comb;
  assign p2_bit_slice_83123_comb = p1_add_82839[17:8];
  assign p2_bit_slice_83124_comb = p1_add_82840[17:8];
  assign p2_bit_slice_83125_comb = p1_add_82841[17:8];
  assign p2_bit_slice_83126_comb = p1_add_82842[17:8];
  assign p2_bit_slice_83127_comb = p1_add_82843[17:8];
  assign p2_bit_slice_83128_comb = p1_add_82844[17:8];
  assign p2_bit_slice_83129_comb = p1_add_82845[17:8];
  assign p2_bit_slice_83130_comb = p1_add_82846[17:8];
  assign p2_bit_slice_83131_comb = p1_add_82847[17:8];
  assign p2_bit_slice_83132_comb = p1_add_82848[17:8];
  assign p2_bit_slice_83133_comb = p1_add_82849[17:8];
  assign p2_bit_slice_83134_comb = p1_add_82850[17:8];
  assign p2_bit_slice_83135_comb = p1_add_82855[17:8];
  assign p2_bit_slice_83136_comb = p1_add_82856[17:8];
  assign p2_bit_slice_83137_comb = p1_add_82857[17:8];
  assign p2_bit_slice_83138_comb = p1_add_82858[17:8];
  assign p2_bit_slice_83139_comb = p1_add_82859[17:8];
  assign p2_bit_slice_83140_comb = p1_add_82860[17:8];
  assign p2_bit_slice_83141_comb = p1_add_82861[17:8];
  assign p2_bit_slice_83142_comb = p1_add_82862[17:8];
  assign p2_bit_slice_83143_comb = p1_add_82863[17:8];
  assign p2_bit_slice_83144_comb = p1_add_82864[17:8];
  assign p2_bit_slice_83145_comb = p1_add_82865[17:8];
  assign p2_bit_slice_83146_comb = p1_add_82866[17:8];
  assign p2_bit_slice_83147_comb = p1_add_82869[17:8];
  assign p2_bit_slice_83148_comb = p1_add_82870[17:8];
  assign p2_bit_slice_83149_comb = p1_add_82871[17:8];
  assign p2_bit_slice_83150_comb = p1_add_82872[17:8];
  assign p2_bit_slice_83151_comb = p1_add_82873[17:8];
  assign p2_bit_slice_83152_comb = p1_add_82874[17:8];
  assign p2_bit_slice_83153_comb = p1_add_82877[17:8];
  assign p2_bit_slice_83154_comb = p1_add_82878[17:8];
  assign p2_bit_slice_83155_comb = p1_add_82879[17:8];
  assign p2_bit_slice_83156_comb = p1_add_82880[17:8];
  assign p2_bit_slice_83157_comb = p1_add_82881[17:8];
  assign p2_bit_slice_83158_comb = p1_add_82882[17:8];
  assign p2_bit_slice_83159_comb = p1_add_82885[17:8];
  assign p2_bit_slice_83160_comb = p1_add_82886[17:8];
  assign p2_bit_slice_83161_comb = p1_add_82887[17:8];
  assign p2_bit_slice_83162_comb = p1_add_82888[17:8];
  assign p2_bit_slice_83163_comb = p1_add_82889[17:8];
  assign p2_bit_slice_83164_comb = p1_add_82890[17:8];
  assign p2_bit_slice_83165_comb = p1_add_82893[17:8];
  assign p2_bit_slice_83166_comb = p1_add_82894[17:8];
  assign p2_bit_slice_83167_comb = p1_add_82895[17:8];
  assign p2_bit_slice_83168_comb = p1_add_82896[17:8];
  assign p2_bit_slice_83169_comb = p1_add_82897[17:8];
  assign p2_bit_slice_83170_comb = p1_add_82898[17:8];
  assign p2_add_83275_comb = p1_sign_ext_82915 + 11'h001;
  assign p2_add_83276_comb = p1_sign_ext_82916 + 11'h001;
  assign p2_add_83277_comb = p1_sign_ext_82917 + 11'h001;
  assign p2_add_83278_comb = p1_sign_ext_82918 + 11'h001;
  assign p2_add_83327_comb = p1_sign_ext_82927 + 11'h001;
  assign p2_add_83328_comb = p1_sign_ext_82928 + 11'h001;
  assign p2_add_83353_comb = p1_sign_ext_82933 + 11'h001;
  assign p2_add_83354_comb = p1_sign_ext_82934 + 11'h001;
  assign p2_concat_83427_comb = {p1_add_82943, p1_bit_slice_82944};
  assign p2_concat_83430_comb = {p1_add_82945, p1_bit_slice_82946};
  assign p2_concat_83433_comb = {p1_add_82947, p1_bit_slice_82948};
  assign p2_concat_83436_comb = {p1_add_82949, p1_bit_slice_82950};
  assign p2_concat_83499_comb = {p1_add_82953, p1_bit_slice_82954};
  assign p2_concat_83502_comb = {p1_add_82955, p1_bit_slice_82956};
  assign p2_concat_83547_comb = {p1_add_82959, p1_bit_slice_82960};
  assign p2_concat_83550_comb = {p1_add_82961, p1_bit_slice_82962};
  assign p2_concat_83379_comb = {p2_add_83275_comb, p1_bit_slice_82939};
  assign p2_concat_83382_comb = {p2_add_83276_comb, p1_bit_slice_82940};
  assign p2_concat_83385_comb = {p2_add_83277_comb, p1_bit_slice_82941};
  assign p2_concat_83388_comb = {p2_add_83278_comb, p1_bit_slice_82942};
  assign p2_concat_83475_comb = {p2_add_83327_comb, p1_bit_slice_82951};
  assign p2_concat_83478_comb = {p2_add_83328_comb, p1_bit_slice_82952};
  assign p2_concat_83523_comb = {p2_add_83353_comb, p1_bit_slice_82957};
  assign p2_concat_83526_comb = {p2_add_83354_comb, p1_bit_slice_82958};
  assign p2_add_83279_comb = {{1{p2_bit_slice_83123_comb[9]}}, p2_bit_slice_83123_comb} + 11'h001;
  assign p2_add_83281_comb = {{1{p2_bit_slice_83124_comb[9]}}, p2_bit_slice_83124_comb} + 11'h001;
  assign p2_add_83283_comb = {{1{p2_bit_slice_83125_comb[9]}}, p2_bit_slice_83125_comb} + 11'h001;
  assign p2_add_83285_comb = {{1{p2_bit_slice_83126_comb[9]}}, p2_bit_slice_83126_comb} + 11'h001;
  assign p2_add_83287_comb = {{1{p2_bit_slice_83127_comb[9]}}, p2_bit_slice_83127_comb} + 11'h001;
  assign p2_add_83289_comb = {{1{p2_bit_slice_83128_comb[9]}}, p2_bit_slice_83128_comb} + 11'h001;
  assign p2_add_83291_comb = {{1{p2_bit_slice_83129_comb[9]}}, p2_bit_slice_83129_comb} + 11'h001;
  assign p2_add_83293_comb = {{1{p2_bit_slice_83130_comb[9]}}, p2_bit_slice_83130_comb} + 11'h001;
  assign p2_add_83295_comb = {{1{p2_bit_slice_83131_comb[9]}}, p2_bit_slice_83131_comb} + 11'h001;
  assign p2_add_83297_comb = {{1{p2_bit_slice_83132_comb[9]}}, p2_bit_slice_83132_comb} + 11'h001;
  assign p2_add_83299_comb = {{1{p2_bit_slice_83133_comb[9]}}, p2_bit_slice_83133_comb} + 11'h001;
  assign p2_add_83301_comb = {{1{p2_bit_slice_83134_comb[9]}}, p2_bit_slice_83134_comb} + 11'h001;
  assign p2_add_83303_comb = {{1{p2_bit_slice_83135_comb[9]}}, p2_bit_slice_83135_comb} + 11'h001;
  assign p2_add_83305_comb = {{1{p2_bit_slice_83136_comb[9]}}, p2_bit_slice_83136_comb} + 11'h001;
  assign p2_add_83307_comb = {{1{p2_bit_slice_83137_comb[9]}}, p2_bit_slice_83137_comb} + 11'h001;
  assign p2_add_83309_comb = {{1{p2_bit_slice_83138_comb[9]}}, p2_bit_slice_83138_comb} + 11'h001;
  assign p2_add_83311_comb = {{1{p2_bit_slice_83139_comb[9]}}, p2_bit_slice_83139_comb} + 11'h001;
  assign p2_add_83313_comb = {{1{p2_bit_slice_83140_comb[9]}}, p2_bit_slice_83140_comb} + 11'h001;
  assign p2_add_83315_comb = {{1{p2_bit_slice_83141_comb[9]}}, p2_bit_slice_83141_comb} + 11'h001;
  assign p2_add_83317_comb = {{1{p2_bit_slice_83142_comb[9]}}, p2_bit_slice_83142_comb} + 11'h001;
  assign p2_add_83319_comb = {{1{p2_bit_slice_83143_comb[9]}}, p2_bit_slice_83143_comb} + 11'h001;
  assign p2_add_83321_comb = {{1{p2_bit_slice_83144_comb[9]}}, p2_bit_slice_83144_comb} + 11'h001;
  assign p2_add_83323_comb = {{1{p2_bit_slice_83145_comb[9]}}, p2_bit_slice_83145_comb} + 11'h001;
  assign p2_add_83325_comb = {{1{p2_bit_slice_83146_comb[9]}}, p2_bit_slice_83146_comb} + 11'h001;
  assign p2_add_83329_comb = {{1{p2_bit_slice_83147_comb[9]}}, p2_bit_slice_83147_comb} + 11'h001;
  assign p2_add_83331_comb = {{1{p2_bit_slice_83148_comb[9]}}, p2_bit_slice_83148_comb} + 11'h001;
  assign p2_add_83333_comb = {{1{p2_bit_slice_83149_comb[9]}}, p2_bit_slice_83149_comb} + 11'h001;
  assign p2_add_83335_comb = {{1{p2_bit_slice_83150_comb[9]}}, p2_bit_slice_83150_comb} + 11'h001;
  assign p2_add_83337_comb = {{1{p2_bit_slice_83151_comb[9]}}, p2_bit_slice_83151_comb} + 11'h001;
  assign p2_add_83339_comb = {{1{p2_bit_slice_83152_comb[9]}}, p2_bit_slice_83152_comb} + 11'h001;
  assign p2_add_83341_comb = {{1{p2_bit_slice_83153_comb[9]}}, p2_bit_slice_83153_comb} + 11'h001;
  assign p2_add_83343_comb = {{1{p2_bit_slice_83154_comb[9]}}, p2_bit_slice_83154_comb} + 11'h001;
  assign p2_add_83345_comb = {{1{p2_bit_slice_83155_comb[9]}}, p2_bit_slice_83155_comb} + 11'h001;
  assign p2_add_83347_comb = {{1{p2_bit_slice_83156_comb[9]}}, p2_bit_slice_83156_comb} + 11'h001;
  assign p2_add_83349_comb = {{1{p2_bit_slice_83157_comb[9]}}, p2_bit_slice_83157_comb} + 11'h001;
  assign p2_add_83351_comb = {{1{p2_bit_slice_83158_comb[9]}}, p2_bit_slice_83158_comb} + 11'h001;
  assign p2_add_83355_comb = {{1{p2_bit_slice_83159_comb[9]}}, p2_bit_slice_83159_comb} + 11'h001;
  assign p2_add_83357_comb = {{1{p2_bit_slice_83160_comb[9]}}, p2_bit_slice_83160_comb} + 11'h001;
  assign p2_add_83359_comb = {{1{p2_bit_slice_83161_comb[9]}}, p2_bit_slice_83161_comb} + 11'h001;
  assign p2_add_83361_comb = {{1{p2_bit_slice_83162_comb[9]}}, p2_bit_slice_83162_comb} + 11'h001;
  assign p2_add_83363_comb = {{1{p2_bit_slice_83163_comb[9]}}, p2_bit_slice_83163_comb} + 11'h001;
  assign p2_add_83365_comb = {{1{p2_bit_slice_83164_comb[9]}}, p2_bit_slice_83164_comb} + 11'h001;
  assign p2_add_83367_comb = {{1{p2_bit_slice_83165_comb[9]}}, p2_bit_slice_83165_comb} + 11'h001;
  assign p2_add_83369_comb = {{1{p2_bit_slice_83166_comb[9]}}, p2_bit_slice_83166_comb} + 11'h001;
  assign p2_add_83371_comb = {{1{p2_bit_slice_83167_comb[9]}}, p2_bit_slice_83167_comb} + 11'h001;
  assign p2_add_83373_comb = {{1{p2_bit_slice_83168_comb[9]}}, p2_bit_slice_83168_comb} + 11'h001;
  assign p2_add_83375_comb = {{1{p2_bit_slice_83169_comb[9]}}, p2_bit_slice_83169_comb} + 11'h001;
  assign p2_add_83377_comb = {{1{p2_bit_slice_83170_comb[9]}}, p2_bit_slice_83170_comb} + 11'h001;
  assign p2_concat_83391_comb = {p2_add_83279_comb, p1_add_82839[7:1]};
  assign p2_concat_83394_comb = {p2_add_83281_comb, p1_add_82840[7:1]};
  assign p2_concat_83397_comb = {p2_add_83283_comb, p1_add_82841[7:1]};
  assign p2_concat_83400_comb = {p2_add_83285_comb, p1_add_82842[7:1]};
  assign p2_concat_83403_comb = {p2_add_83287_comb, p1_add_82843[7:1]};
  assign p2_concat_83406_comb = {p2_add_83289_comb, p1_add_82844[7:1]};
  assign p2_concat_83409_comb = {p2_add_83291_comb, p1_add_82845[7:1]};
  assign p2_concat_83412_comb = {p2_add_83293_comb, p1_add_82846[7:1]};
  assign p2_concat_83415_comb = {p2_add_83295_comb, p1_add_82847[7:1]};
  assign p2_concat_83418_comb = {p2_add_83297_comb, p1_add_82848[7:1]};
  assign p2_concat_83421_comb = {p2_add_83299_comb, p1_add_82849[7:1]};
  assign p2_concat_83424_comb = {p2_add_83301_comb, p1_add_82850[7:1]};
  assign p2_concat_83439_comb = {p2_add_83303_comb, p1_add_82855[7:1]};
  assign p2_concat_83442_comb = {p2_add_83305_comb, p1_add_82856[7:1]};
  assign p2_concat_83445_comb = {p2_add_83307_comb, p1_add_82857[7:1]};
  assign p2_concat_83448_comb = {p2_add_83309_comb, p1_add_82858[7:1]};
  assign p2_concat_83451_comb = {p2_add_83311_comb, p1_add_82859[7:1]};
  assign p2_concat_83454_comb = {p2_add_83313_comb, p1_add_82860[7:1]};
  assign p2_concat_83457_comb = {p2_add_83315_comb, p1_add_82861[7:1]};
  assign p2_concat_83460_comb = {p2_add_83317_comb, p1_add_82862[7:1]};
  assign p2_concat_83463_comb = {p2_add_83319_comb, p1_add_82863[7:1]};
  assign p2_concat_83466_comb = {p2_add_83321_comb, p1_add_82864[7:1]};
  assign p2_concat_83469_comb = {p2_add_83323_comb, p1_add_82865[7:1]};
  assign p2_concat_83472_comb = {p2_add_83325_comb, p1_add_82866[7:1]};
  assign p2_concat_83481_comb = {p2_add_83329_comb, p1_add_82869[7:1]};
  assign p2_concat_83484_comb = {p2_add_83331_comb, p1_add_82870[7:1]};
  assign p2_concat_83487_comb = {p2_add_83333_comb, p1_add_82871[7:1]};
  assign p2_concat_83490_comb = {p2_add_83335_comb, p1_add_82872[7:1]};
  assign p2_concat_83493_comb = {p2_add_83337_comb, p1_add_82873[7:1]};
  assign p2_concat_83496_comb = {p2_add_83339_comb, p1_add_82874[7:1]};
  assign p2_concat_83505_comb = {p2_add_83341_comb, p1_add_82877[7:1]};
  assign p2_concat_83508_comb = {p2_add_83343_comb, p1_add_82878[7:1]};
  assign p2_concat_83511_comb = {p2_add_83345_comb, p1_add_82879[7:1]};
  assign p2_concat_83514_comb = {p2_add_83347_comb, p1_add_82880[7:1]};
  assign p2_concat_83517_comb = {p2_add_83349_comb, p1_add_82881[7:1]};
  assign p2_concat_83520_comb = {p2_add_83351_comb, p1_add_82882[7:1]};
  assign p2_concat_83529_comb = {p2_add_83355_comb, p1_add_82885[7:1]};
  assign p2_concat_83532_comb = {p2_add_83357_comb, p1_add_82886[7:1]};
  assign p2_concat_83535_comb = {p2_add_83359_comb, p1_add_82887[7:1]};
  assign p2_concat_83538_comb = {p2_add_83361_comb, p1_add_82888[7:1]};
  assign p2_concat_83541_comb = {p2_add_83363_comb, p1_add_82889[7:1]};
  assign p2_concat_83544_comb = {p2_add_83365_comb, p1_add_82890[7:1]};
  assign p2_concat_83553_comb = {p2_add_83367_comb, p1_add_82893[7:1]};
  assign p2_concat_83556_comb = {p2_add_83369_comb, p1_add_82894[7:1]};
  assign p2_concat_83559_comb = {p2_add_83371_comb, p1_add_82895[7:1]};
  assign p2_concat_83562_comb = {p2_add_83373_comb, p1_add_82896[7:1]};
  assign p2_concat_83565_comb = {p2_add_83375_comb, p1_add_82897[7:1]};
  assign p2_concat_83568_comb = {p2_add_83377_comb, p1_add_82898[7:1]};
  assign p2_clipped__44_comb = $signed(p2_concat_83427_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83427_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p1_add_82943[2:0], p1_bit_slice_82944});
  assign p2_clipped__60_comb = $signed(p2_concat_83430_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83430_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p1_add_82945[2:0], p1_bit_slice_82946});
  assign p2_clipped__76_comb = $signed(p2_concat_83433_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83433_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p1_add_82947[2:0], p1_bit_slice_82948});
  assign p2_clipped__92_comb = $signed(p2_concat_83436_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83436_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p1_add_82949[2:0], p1_bit_slice_82950});
  assign p2_clipped__28_comb = $signed(p2_concat_83499_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83499_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p1_add_82953[2:0], p1_bit_slice_82954});
  assign p2_clipped__108_comb = $signed(p2_concat_83502_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83502_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p1_add_82955[2:0], p1_bit_slice_82956});
  assign p2_clipped__12_comb = $signed(p2_concat_83547_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83547_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p1_add_82959[2:0], p1_bit_slice_82960});
  assign p2_clipped__124_comb = $signed(p2_concat_83550_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83550_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p1_add_82961[2:0], p1_bit_slice_82962});
  assign p2_clipped__40_comb = $signed(p2_concat_83379_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83379_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83275_comb[2:0], p1_bit_slice_82939});
  assign p2_clipped__56_comb = $signed(p2_concat_83382_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83382_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83276_comb[2:0], p1_bit_slice_82940});
  assign p2_clipped__72_comb = $signed(p2_concat_83385_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83385_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83277_comb[2:0], p1_bit_slice_82941});
  assign p2_clipped__88_comb = $signed(p2_concat_83388_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83388_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83278_comb[2:0], p1_bit_slice_82942});
  assign p2_clipped__24_comb = $signed(p2_concat_83475_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83475_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83327_comb[2:0], p1_bit_slice_82951});
  assign p2_clipped__104_comb = $signed(p2_concat_83478_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83478_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83328_comb[2:0], p1_bit_slice_82952});
  assign p2_clipped__8_comb = $signed(p2_concat_83523_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83523_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83353_comb[2:0], p1_bit_slice_82957});
  assign p2_clipped__120_comb = $signed(p2_concat_83526_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83526_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83354_comb[2:0], p1_bit_slice_82958});
  assign p2_bit_slice_84099_comb = p2_clipped__44_comb[9:7];
  assign p2_bit_slice_84100_comb = p2_clipped__60_comb[9:7];
  assign p2_bit_slice_84101_comb = p2_clipped__76_comb[9:7];
  assign p2_bit_slice_84102_comb = p2_clipped__92_comb[9:7];
  assign p2_bit_slice_84123_comb = p2_clipped__28_comb[9:7];
  assign p2_bit_slice_84124_comb = p2_clipped__108_comb[9:7];
  assign p2_bit_slice_84139_comb = p2_clipped__12_comb[9:7];
  assign p2_bit_slice_84140_comb = p2_clipped__124_comb[9:7];
  assign p2_bit_slice_84083_comb = p2_clipped__40_comb[9:7];
  assign p2_bit_slice_84084_comb = p2_clipped__56_comb[9:7];
  assign p2_bit_slice_84085_comb = p2_clipped__72_comb[9:7];
  assign p2_bit_slice_84086_comb = p2_clipped__88_comb[9:7];
  assign p2_bit_slice_84115_comb = p2_clipped__24_comb[9:7];
  assign p2_bit_slice_84116_comb = p2_clipped__104_comb[9:7];
  assign p2_bit_slice_84131_comb = p2_clipped__8_comb[9:7];
  assign p2_bit_slice_84132_comb = p2_clipped__120_comb[9:7];
  assign p2_clipped__41_comb = $signed(p2_concat_83391_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83391_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83279_comb[2:0], p1_add_82839[7:1]});
  assign p2_clipped__57_comb = $signed(p2_concat_83394_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83394_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83281_comb[2:0], p1_add_82840[7:1]});
  assign p2_clipped__73_comb = $signed(p2_concat_83397_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83397_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83283_comb[2:0], p1_add_82841[7:1]});
  assign p2_clipped__89_comb = $signed(p2_concat_83400_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83400_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83285_comb[2:0], p1_add_82842[7:1]});
  assign p2_clipped__42_comb = $signed(p2_concat_83403_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83403_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83287_comb[2:0], p1_add_82843[7:1]});
  assign p2_clipped__58_comb = $signed(p2_concat_83406_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83406_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83289_comb[2:0], p1_add_82844[7:1]});
  assign p2_clipped__74_comb = $signed(p2_concat_83409_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83409_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83291_comb[2:0], p1_add_82845[7:1]});
  assign p2_clipped__90_comb = $signed(p2_concat_83412_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83412_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83293_comb[2:0], p1_add_82846[7:1]});
  assign p2_clipped__43_comb = $signed(p2_concat_83415_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83415_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83295_comb[2:0], p1_add_82847[7:1]});
  assign p2_clipped__59_comb = $signed(p2_concat_83418_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83418_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83297_comb[2:0], p1_add_82848[7:1]});
  assign p2_clipped__75_comb = $signed(p2_concat_83421_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83421_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83299_comb[2:0], p1_add_82849[7:1]});
  assign p2_clipped__91_comb = $signed(p2_concat_83424_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83424_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83301_comb[2:0], p1_add_82850[7:1]});
  assign p2_clipped__45_comb = $signed(p2_concat_83439_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83439_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83303_comb[2:0], p1_add_82855[7:1]});
  assign p2_clipped__61_comb = $signed(p2_concat_83442_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83442_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83305_comb[2:0], p1_add_82856[7:1]});
  assign p2_clipped__77_comb = $signed(p2_concat_83445_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83445_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83307_comb[2:0], p1_add_82857[7:1]});
  assign p2_clipped__93_comb = $signed(p2_concat_83448_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83448_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83309_comb[2:0], p1_add_82858[7:1]});
  assign p2_clipped__46_comb = $signed(p2_concat_83451_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83451_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83311_comb[2:0], p1_add_82859[7:1]});
  assign p2_clipped__62_comb = $signed(p2_concat_83454_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83454_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83313_comb[2:0], p1_add_82860[7:1]});
  assign p2_clipped__78_comb = $signed(p2_concat_83457_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83457_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83315_comb[2:0], p1_add_82861[7:1]});
  assign p2_clipped__94_comb = $signed(p2_concat_83460_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83460_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83317_comb[2:0], p1_add_82862[7:1]});
  assign p2_clipped__47_comb = $signed(p2_concat_83463_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83463_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83319_comb[2:0], p1_add_82863[7:1]});
  assign p2_clipped__63_comb = $signed(p2_concat_83466_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83466_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83321_comb[2:0], p1_add_82864[7:1]});
  assign p2_clipped__79_comb = $signed(p2_concat_83469_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83469_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83323_comb[2:0], p1_add_82865[7:1]});
  assign p2_clipped__95_comb = $signed(p2_concat_83472_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83472_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83325_comb[2:0], p1_add_82866[7:1]});
  assign p2_clipped__25_comb = $signed(p2_concat_83481_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83481_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83329_comb[2:0], p1_add_82869[7:1]});
  assign p2_clipped__105_comb = $signed(p2_concat_83484_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83484_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83331_comb[2:0], p1_add_82870[7:1]});
  assign p2_clipped__26_comb = $signed(p2_concat_83487_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83487_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83333_comb[2:0], p1_add_82871[7:1]});
  assign p2_clipped__106_comb = $signed(p2_concat_83490_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83490_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83335_comb[2:0], p1_add_82872[7:1]});
  assign p2_clipped__27_comb = $signed(p2_concat_83493_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83493_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83337_comb[2:0], p1_add_82873[7:1]});
  assign p2_clipped__107_comb = $signed(p2_concat_83496_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83496_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83339_comb[2:0], p1_add_82874[7:1]});
  assign p2_clipped__29_comb = $signed(p2_concat_83505_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83505_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83341_comb[2:0], p1_add_82877[7:1]});
  assign p2_clipped__109_comb = $signed(p2_concat_83508_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83508_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83343_comb[2:0], p1_add_82878[7:1]});
  assign p2_clipped__30_comb = $signed(p2_concat_83511_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83511_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83345_comb[2:0], p1_add_82879[7:1]});
  assign p2_clipped__110_comb = $signed(p2_concat_83514_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83514_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83347_comb[2:0], p1_add_82880[7:1]});
  assign p2_clipped__31_comb = $signed(p2_concat_83517_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83517_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83349_comb[2:0], p1_add_82881[7:1]});
  assign p2_clipped__111_comb = $signed(p2_concat_83520_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83520_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83351_comb[2:0], p1_add_82882[7:1]});
  assign p2_clipped__9_comb = $signed(p2_concat_83529_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83529_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83355_comb[2:0], p1_add_82885[7:1]});
  assign p2_clipped__121_comb = $signed(p2_concat_83532_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83532_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83357_comb[2:0], p1_add_82886[7:1]});
  assign p2_clipped__10_comb = $signed(p2_concat_83535_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83535_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83359_comb[2:0], p1_add_82887[7:1]});
  assign p2_clipped__122_comb = $signed(p2_concat_83538_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83538_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83361_comb[2:0], p1_add_82888[7:1]});
  assign p2_clipped__11_comb = $signed(p2_concat_83541_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83541_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83363_comb[2:0], p1_add_82889[7:1]});
  assign p2_clipped__123_comb = $signed(p2_concat_83544_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83544_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83365_comb[2:0], p1_add_82890[7:1]});
  assign p2_clipped__13_comb = $signed(p2_concat_83553_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83553_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83367_comb[2:0], p1_add_82893[7:1]});
  assign p2_clipped__125_comb = $signed(p2_concat_83556_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83556_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83369_comb[2:0], p1_add_82894[7:1]});
  assign p2_clipped__14_comb = $signed(p2_concat_83559_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83559_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83371_comb[2:0], p1_add_82895[7:1]});
  assign p2_clipped__126_comb = $signed(p2_concat_83562_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83562_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83373_comb[2:0], p1_add_82896[7:1]});
  assign p2_clipped__15_comb = $signed(p2_concat_83565_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83565_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83375_comb[2:0], p1_add_82897[7:1]});
  assign p2_clipped__127_comb = $signed(p2_concat_83568_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p2_concat_83568_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p2_add_83377_comb[2:0], p1_add_82898[7:1]});
  assign p2_add_84307_comb = {{1{p2_bit_slice_84099_comb[2]}}, p2_bit_slice_84099_comb} + 4'hf;
  assign p2_add_84309_comb = {{1{p2_bit_slice_84100_comb[2]}}, p2_bit_slice_84100_comb} + 4'hf;
  assign p2_add_84311_comb = {{1{p2_bit_slice_84101_comb[2]}}, p2_bit_slice_84101_comb} + 4'hf;
  assign p2_add_84313_comb = {{1{p2_bit_slice_84102_comb[2]}}, p2_bit_slice_84102_comb} + 4'hf;
  assign p2_add_84355_comb = {{1{p2_bit_slice_84123_comb[2]}}, p2_bit_slice_84123_comb} + 4'hf;
  assign p2_add_84357_comb = {{1{p2_bit_slice_84124_comb[2]}}, p2_bit_slice_84124_comb} + 4'hf;
  assign p2_add_84387_comb = {{1{p2_bit_slice_84139_comb[2]}}, p2_bit_slice_84139_comb} + 4'hf;
  assign p2_add_84389_comb = {{1{p2_bit_slice_84140_comb[2]}}, p2_bit_slice_84140_comb} + 4'hf;
  assign p2_bit_slice_84087_comb = p2_clipped__41_comb[9:7];
  assign p2_bit_slice_84088_comb = p2_clipped__57_comb[9:7];
  assign p2_bit_slice_84089_comb = p2_clipped__73_comb[9:7];
  assign p2_bit_slice_84090_comb = p2_clipped__89_comb[9:7];
  assign p2_bit_slice_84091_comb = p2_clipped__42_comb[9:7];
  assign p2_bit_slice_84092_comb = p2_clipped__58_comb[9:7];
  assign p2_bit_slice_84093_comb = p2_clipped__74_comb[9:7];
  assign p2_bit_slice_84094_comb = p2_clipped__90_comb[9:7];
  assign p2_bit_slice_84095_comb = p2_clipped__43_comb[9:7];
  assign p2_bit_slice_84096_comb = p2_clipped__59_comb[9:7];
  assign p2_bit_slice_84097_comb = p2_clipped__75_comb[9:7];
  assign p2_bit_slice_84098_comb = p2_clipped__91_comb[9:7];
  assign p2_bit_slice_84103_comb = p2_clipped__45_comb[9:7];
  assign p2_bit_slice_84104_comb = p2_clipped__61_comb[9:7];
  assign p2_bit_slice_84105_comb = p2_clipped__77_comb[9:7];
  assign p2_bit_slice_84106_comb = p2_clipped__93_comb[9:7];
  assign p2_bit_slice_84107_comb = p2_clipped__46_comb[9:7];
  assign p2_bit_slice_84108_comb = p2_clipped__62_comb[9:7];
  assign p2_bit_slice_84109_comb = p2_clipped__78_comb[9:7];
  assign p2_bit_slice_84110_comb = p2_clipped__94_comb[9:7];
  assign p2_bit_slice_84111_comb = p2_clipped__47_comb[9:7];
  assign p2_bit_slice_84112_comb = p2_clipped__63_comb[9:7];
  assign p2_bit_slice_84113_comb = p2_clipped__79_comb[9:7];
  assign p2_bit_slice_84114_comb = p2_clipped__95_comb[9:7];
  assign p2_bit_slice_84117_comb = p2_clipped__25_comb[9:7];
  assign p2_bit_slice_84118_comb = p2_clipped__105_comb[9:7];
  assign p2_bit_slice_84119_comb = p2_clipped__26_comb[9:7];
  assign p2_bit_slice_84120_comb = p2_clipped__106_comb[9:7];
  assign p2_bit_slice_84121_comb = p2_clipped__27_comb[9:7];
  assign p2_bit_slice_84122_comb = p2_clipped__107_comb[9:7];
  assign p2_bit_slice_84125_comb = p2_clipped__29_comb[9:7];
  assign p2_bit_slice_84126_comb = p2_clipped__109_comb[9:7];
  assign p2_bit_slice_84127_comb = p2_clipped__30_comb[9:7];
  assign p2_bit_slice_84128_comb = p2_clipped__110_comb[9:7];
  assign p2_bit_slice_84129_comb = p2_clipped__31_comb[9:7];
  assign p2_bit_slice_84130_comb = p2_clipped__111_comb[9:7];
  assign p2_bit_slice_84133_comb = p2_clipped__9_comb[9:7];
  assign p2_bit_slice_84134_comb = p2_clipped__121_comb[9:7];
  assign p2_bit_slice_84135_comb = p2_clipped__10_comb[9:7];
  assign p2_bit_slice_84136_comb = p2_clipped__122_comb[9:7];
  assign p2_bit_slice_84137_comb = p2_clipped__11_comb[9:7];
  assign p2_bit_slice_84138_comb = p2_clipped__123_comb[9:7];
  assign p2_bit_slice_84141_comb = p2_clipped__13_comb[9:7];
  assign p2_bit_slice_84142_comb = p2_clipped__125_comb[9:7];
  assign p2_bit_slice_84143_comb = p2_clipped__14_comb[9:7];
  assign p2_bit_slice_84144_comb = p2_clipped__126_comb[9:7];
  assign p2_bit_slice_84145_comb = p2_clipped__15_comb[9:7];
  assign p2_bit_slice_84146_comb = p2_clipped__127_comb[9:7];
  assign p2_add_84275_comb = {{1{p2_bit_slice_84083_comb[2]}}, p2_bit_slice_84083_comb} + 4'hf;
  assign p2_add_84277_comb = {{1{p2_bit_slice_84084_comb[2]}}, p2_bit_slice_84084_comb} + 4'hf;
  assign p2_add_84279_comb = {{1{p2_bit_slice_84085_comb[2]}}, p2_bit_slice_84085_comb} + 4'hf;
  assign p2_add_84281_comb = {{1{p2_bit_slice_84086_comb[2]}}, p2_bit_slice_84086_comb} + 4'hf;
  assign p2_add_84339_comb = {{1{p2_bit_slice_84115_comb[2]}}, p2_bit_slice_84115_comb} + 4'hf;
  assign p2_add_84341_comb = {{1{p2_bit_slice_84116_comb[2]}}, p2_bit_slice_84116_comb} + 4'hf;
  assign p2_add_84371_comb = {{1{p2_bit_slice_84131_comb[2]}}, p2_bit_slice_84131_comb} + 4'hf;
  assign p2_add_84373_comb = {{1{p2_bit_slice_84132_comb[2]}}, p2_bit_slice_84132_comb} + 4'hf;
  assign p2_concat_84419_comb = {p2_add_84307_comb, p2_clipped__44_comb[6:0]};
  assign p2_concat_84420_comb = {p2_add_84309_comb, p2_clipped__60_comb[6:0]};
  assign p2_concat_84421_comb = {p2_add_84311_comb, p2_clipped__76_comb[6:0]};
  assign p2_concat_84422_comb = {p2_add_84313_comb, p2_clipped__92_comb[6:0]};
  assign p2_concat_84443_comb = {p2_add_84355_comb, p2_clipped__28_comb[6:0]};
  assign p2_concat_84444_comb = {p2_add_84357_comb, p2_clipped__108_comb[6:0]};
  assign p2_concat_84459_comb = {p2_add_84387_comb, p2_clipped__12_comb[6:0]};
  assign p2_concat_84460_comb = {p2_add_84389_comb, p2_clipped__124_comb[6:0]};
  assign p2_concat_84403_comb = {p2_add_84275_comb, p2_clipped__40_comb[6:0]};
  assign p2_concat_84404_comb = {p2_add_84277_comb, p2_clipped__56_comb[6:0]};
  assign p2_concat_84405_comb = {p2_add_84279_comb, p2_clipped__72_comb[6:0]};
  assign p2_concat_84406_comb = {p2_add_84281_comb, p2_clipped__88_comb[6:0]};
  assign p2_concat_84435_comb = {p2_add_84339_comb, p2_clipped__24_comb[6:0]};
  assign p2_concat_84436_comb = {p2_add_84341_comb, p2_clipped__104_comb[6:0]};
  assign p2_concat_84451_comb = {p2_add_84371_comb, p2_clipped__8_comb[6:0]};
  assign p2_concat_84452_comb = {p2_add_84373_comb, p2_clipped__120_comb[6:0]};
  assign p2_sign_ext_84501_comb = {{13{p2_concat_84419_comb[10]}}, p2_concat_84419_comb};
  assign p2_sign_ext_84502_comb = {{13{p2_concat_84420_comb[10]}}, p2_concat_84420_comb};
  assign p2_sign_ext_84503_comb = {{13{p2_concat_84421_comb[10]}}, p2_concat_84421_comb};
  assign p2_sign_ext_84504_comb = {{13{p2_concat_84422_comb[10]}}, p2_concat_84422_comb};
  assign p2_sign_ext_84539_comb = {{13{p2_concat_84443_comb[10]}}, p2_concat_84443_comb};
  assign p2_sign_ext_84540_comb = {{13{p2_concat_84444_comb[10]}}, p2_concat_84444_comb};
  assign p2_sign_ext_84603_comb = {{13{p2_concat_84459_comb[10]}}, p2_concat_84459_comb};
  assign p2_sign_ext_84608_comb = {{13{p2_concat_84460_comb[10]}}, p2_concat_84460_comb};
  assign p2_add_84283_comb = {{1{p2_bit_slice_84087_comb[2]}}, p2_bit_slice_84087_comb} + 4'hf;
  assign p2_add_84285_comb = {{1{p2_bit_slice_84088_comb[2]}}, p2_bit_slice_84088_comb} + 4'hf;
  assign p2_add_84287_comb = {{1{p2_bit_slice_84089_comb[2]}}, p2_bit_slice_84089_comb} + 4'hf;
  assign p2_add_84289_comb = {{1{p2_bit_slice_84090_comb[2]}}, p2_bit_slice_84090_comb} + 4'hf;
  assign p2_add_84291_comb = {{1{p2_bit_slice_84091_comb[2]}}, p2_bit_slice_84091_comb} + 4'hf;
  assign p2_add_84293_comb = {{1{p2_bit_slice_84092_comb[2]}}, p2_bit_slice_84092_comb} + 4'hf;
  assign p2_add_84295_comb = {{1{p2_bit_slice_84093_comb[2]}}, p2_bit_slice_84093_comb} + 4'hf;
  assign p2_add_84297_comb = {{1{p2_bit_slice_84094_comb[2]}}, p2_bit_slice_84094_comb} + 4'hf;
  assign p2_add_84299_comb = {{1{p2_bit_slice_84095_comb[2]}}, p2_bit_slice_84095_comb} + 4'hf;
  assign p2_add_84301_comb = {{1{p2_bit_slice_84096_comb[2]}}, p2_bit_slice_84096_comb} + 4'hf;
  assign p2_add_84303_comb = {{1{p2_bit_slice_84097_comb[2]}}, p2_bit_slice_84097_comb} + 4'hf;
  assign p2_add_84305_comb = {{1{p2_bit_slice_84098_comb[2]}}, p2_bit_slice_84098_comb} + 4'hf;
  assign p2_add_84315_comb = {{1{p2_bit_slice_84103_comb[2]}}, p2_bit_slice_84103_comb} + 4'hf;
  assign p2_add_84317_comb = {{1{p2_bit_slice_84104_comb[2]}}, p2_bit_slice_84104_comb} + 4'hf;
  assign p2_add_84319_comb = {{1{p2_bit_slice_84105_comb[2]}}, p2_bit_slice_84105_comb} + 4'hf;
  assign p2_add_84321_comb = {{1{p2_bit_slice_84106_comb[2]}}, p2_bit_slice_84106_comb} + 4'hf;
  assign p2_add_84323_comb = {{1{p2_bit_slice_84107_comb[2]}}, p2_bit_slice_84107_comb} + 4'hf;
  assign p2_add_84325_comb = {{1{p2_bit_slice_84108_comb[2]}}, p2_bit_slice_84108_comb} + 4'hf;
  assign p2_add_84327_comb = {{1{p2_bit_slice_84109_comb[2]}}, p2_bit_slice_84109_comb} + 4'hf;
  assign p2_add_84329_comb = {{1{p2_bit_slice_84110_comb[2]}}, p2_bit_slice_84110_comb} + 4'hf;
  assign p2_add_84331_comb = {{1{p2_bit_slice_84111_comb[2]}}, p2_bit_slice_84111_comb} + 4'hf;
  assign p2_add_84333_comb = {{1{p2_bit_slice_84112_comb[2]}}, p2_bit_slice_84112_comb} + 4'hf;
  assign p2_add_84335_comb = {{1{p2_bit_slice_84113_comb[2]}}, p2_bit_slice_84113_comb} + 4'hf;
  assign p2_add_84337_comb = {{1{p2_bit_slice_84114_comb[2]}}, p2_bit_slice_84114_comb} + 4'hf;
  assign p2_add_84343_comb = {{1{p2_bit_slice_84117_comb[2]}}, p2_bit_slice_84117_comb} + 4'hf;
  assign p2_add_84345_comb = {{1{p2_bit_slice_84118_comb[2]}}, p2_bit_slice_84118_comb} + 4'hf;
  assign p2_add_84347_comb = {{1{p2_bit_slice_84119_comb[2]}}, p2_bit_slice_84119_comb} + 4'hf;
  assign p2_add_84349_comb = {{1{p2_bit_slice_84120_comb[2]}}, p2_bit_slice_84120_comb} + 4'hf;
  assign p2_add_84351_comb = {{1{p2_bit_slice_84121_comb[2]}}, p2_bit_slice_84121_comb} + 4'hf;
  assign p2_add_84353_comb = {{1{p2_bit_slice_84122_comb[2]}}, p2_bit_slice_84122_comb} + 4'hf;
  assign p2_add_84359_comb = {{1{p2_bit_slice_84125_comb[2]}}, p2_bit_slice_84125_comb} + 4'hf;
  assign p2_add_84361_comb = {{1{p2_bit_slice_84126_comb[2]}}, p2_bit_slice_84126_comb} + 4'hf;
  assign p2_add_84363_comb = {{1{p2_bit_slice_84127_comb[2]}}, p2_bit_slice_84127_comb} + 4'hf;
  assign p2_add_84365_comb = {{1{p2_bit_slice_84128_comb[2]}}, p2_bit_slice_84128_comb} + 4'hf;
  assign p2_add_84367_comb = {{1{p2_bit_slice_84129_comb[2]}}, p2_bit_slice_84129_comb} + 4'hf;
  assign p2_add_84369_comb = {{1{p2_bit_slice_84130_comb[2]}}, p2_bit_slice_84130_comb} + 4'hf;
  assign p2_add_84375_comb = {{1{p2_bit_slice_84133_comb[2]}}, p2_bit_slice_84133_comb} + 4'hf;
  assign p2_add_84377_comb = {{1{p2_bit_slice_84134_comb[2]}}, p2_bit_slice_84134_comb} + 4'hf;
  assign p2_add_84379_comb = {{1{p2_bit_slice_84135_comb[2]}}, p2_bit_slice_84135_comb} + 4'hf;
  assign p2_add_84381_comb = {{1{p2_bit_slice_84136_comb[2]}}, p2_bit_slice_84136_comb} + 4'hf;
  assign p2_add_84383_comb = {{1{p2_bit_slice_84137_comb[2]}}, p2_bit_slice_84137_comb} + 4'hf;
  assign p2_add_84385_comb = {{1{p2_bit_slice_84138_comb[2]}}, p2_bit_slice_84138_comb} + 4'hf;
  assign p2_add_84391_comb = {{1{p2_bit_slice_84141_comb[2]}}, p2_bit_slice_84141_comb} + 4'hf;
  assign p2_add_84393_comb = {{1{p2_bit_slice_84142_comb[2]}}, p2_bit_slice_84142_comb} + 4'hf;
  assign p2_add_84395_comb = {{1{p2_bit_slice_84143_comb[2]}}, p2_bit_slice_84143_comb} + 4'hf;
  assign p2_add_84397_comb = {{1{p2_bit_slice_84144_comb[2]}}, p2_bit_slice_84144_comb} + 4'hf;
  assign p2_add_84399_comb = {{1{p2_bit_slice_84145_comb[2]}}, p2_bit_slice_84145_comb} + 4'hf;
  assign p2_add_84401_comb = {{1{p2_bit_slice_84146_comb[2]}}, p2_bit_slice_84146_comb} + 4'hf;
  assign p2_sign_ext_84469_comb = {{13{p2_concat_84403_comb[10]}}, p2_concat_84403_comb};
  assign p2_sign_ext_84470_comb = {{13{p2_concat_84404_comb[10]}}, p2_concat_84404_comb};
  assign p2_sign_ext_84471_comb = {{13{p2_concat_84405_comb[10]}}, p2_concat_84405_comb};
  assign p2_sign_ext_84472_comb = {{13{p2_concat_84406_comb[10]}}, p2_concat_84406_comb};
  assign p2_sign_ext_84531_comb = {{13{p2_concat_84435_comb[10]}}, p2_concat_84435_comb};
  assign p2_sign_ext_84532_comb = {{13{p2_concat_84436_comb[10]}}, p2_concat_84436_comb};
  assign p2_sign_ext_84579_comb = {{13{p2_concat_84451_comb[10]}}, p2_concat_84451_comb};
  assign p2_sign_ext_84584_comb = {{13{p2_concat_84452_comb[10]}}, p2_concat_84452_comb};
  assign p2_smul_84707_comb = smul20b_11b_x_9b(p2_concat_84459_comb, 9'h0fb);
  assign p2_smul_84708_comb = smul20b_11b_x_9b(p2_concat_84443_comb, 9'h0d5);
  assign p2_smul_84717_comb = smul20b_11b_x_9b(p2_concat_84444_comb, 9'h12b);
  assign p2_smul_84718_comb = smul20b_11b_x_9b(p2_concat_84460_comb, 9'h105);
  assign p2_smul_84859_comb = smul20b_11b_x_9b(p2_concat_84459_comb, 9'h0d5);
  assign p2_smul_84861_comb = smul20b_11b_x_9b(p2_concat_84419_comb, 9'h105);
  assign p2_smul_84866_comb = smul20b_11b_x_9b(p2_concat_84422_comb, 9'h0fb);
  assign p2_smul_84868_comb = smul20b_11b_x_9b(p2_concat_84460_comb, 9'h12b);
  assign p2_smul_84941_comb = smul20b_11b_x_9b(p2_concat_84443_comb, 9'h105);
  assign p2_smul_84943_comb = smul20b_11b_x_9b(p2_concat_84420_comb, 9'h0d5);
  assign p2_smul_84944_comb = smul20b_11b_x_9b(p2_concat_84421_comb, 9'h0d5);
  assign p2_smul_84946_comb = smul20b_11b_x_9b(p2_concat_84444_comb, 9'h105);
  assign p2_smul_85063_comb = smul20b_11b_x_9b(p2_concat_84419_comb, 9'h0d5);
  assign p2_smul_85064_comb = smul20b_11b_x_9b(p2_concat_84420_comb, 9'h105);
  assign p2_smul_85065_comb = smul20b_11b_x_9b(p2_concat_84421_comb, 9'h105);
  assign p2_smul_85066_comb = smul20b_11b_x_9b(p2_concat_84422_comb, 9'h0d5);
  assign p2_concat_84407_comb = {p2_add_84283_comb, p2_clipped__41_comb[6:0]};
  assign p2_concat_84408_comb = {p2_add_84285_comb, p2_clipped__57_comb[6:0]};
  assign p2_concat_84409_comb = {p2_add_84287_comb, p2_clipped__73_comb[6:0]};
  assign p2_concat_84410_comb = {p2_add_84289_comb, p2_clipped__89_comb[6:0]};
  assign p2_concat_84411_comb = {p2_add_84291_comb, p2_clipped__42_comb[6:0]};
  assign p2_concat_84412_comb = {p2_add_84293_comb, p2_clipped__58_comb[6:0]};
  assign p2_concat_84413_comb = {p2_add_84295_comb, p2_clipped__74_comb[6:0]};
  assign p2_concat_84414_comb = {p2_add_84297_comb, p2_clipped__90_comb[6:0]};
  assign p2_concat_84415_comb = {p2_add_84299_comb, p2_clipped__43_comb[6:0]};
  assign p2_concat_84416_comb = {p2_add_84301_comb, p2_clipped__59_comb[6:0]};
  assign p2_concat_84417_comb = {p2_add_84303_comb, p2_clipped__75_comb[6:0]};
  assign p2_concat_84418_comb = {p2_add_84305_comb, p2_clipped__91_comb[6:0]};
  assign p2_concat_84423_comb = {p2_add_84315_comb, p2_clipped__45_comb[6:0]};
  assign p2_concat_84424_comb = {p2_add_84317_comb, p2_clipped__61_comb[6:0]};
  assign p2_concat_84425_comb = {p2_add_84319_comb, p2_clipped__77_comb[6:0]};
  assign p2_concat_84426_comb = {p2_add_84321_comb, p2_clipped__93_comb[6:0]};
  assign p2_concat_84427_comb = {p2_add_84323_comb, p2_clipped__46_comb[6:0]};
  assign p2_concat_84428_comb = {p2_add_84325_comb, p2_clipped__62_comb[6:0]};
  assign p2_concat_84429_comb = {p2_add_84327_comb, p2_clipped__78_comb[6:0]};
  assign p2_concat_84430_comb = {p2_add_84329_comb, p2_clipped__94_comb[6:0]};
  assign p2_concat_84431_comb = {p2_add_84331_comb, p2_clipped__47_comb[6:0]};
  assign p2_concat_84432_comb = {p2_add_84333_comb, p2_clipped__63_comb[6:0]};
  assign p2_concat_84433_comb = {p2_add_84335_comb, p2_clipped__79_comb[6:0]};
  assign p2_concat_84434_comb = {p2_add_84337_comb, p2_clipped__95_comb[6:0]};
  assign p2_concat_84437_comb = {p2_add_84343_comb, p2_clipped__25_comb[6:0]};
  assign p2_concat_84438_comb = {p2_add_84345_comb, p2_clipped__105_comb[6:0]};
  assign p2_concat_84439_comb = {p2_add_84347_comb, p2_clipped__26_comb[6:0]};
  assign p2_concat_84440_comb = {p2_add_84349_comb, p2_clipped__106_comb[6:0]};
  assign p2_concat_84441_comb = {p2_add_84351_comb, p2_clipped__27_comb[6:0]};
  assign p2_concat_84442_comb = {p2_add_84353_comb, p2_clipped__107_comb[6:0]};
  assign p2_concat_84445_comb = {p2_add_84359_comb, p2_clipped__29_comb[6:0]};
  assign p2_concat_84446_comb = {p2_add_84361_comb, p2_clipped__109_comb[6:0]};
  assign p2_concat_84447_comb = {p2_add_84363_comb, p2_clipped__30_comb[6:0]};
  assign p2_concat_84448_comb = {p2_add_84365_comb, p2_clipped__110_comb[6:0]};
  assign p2_concat_84449_comb = {p2_add_84367_comb, p2_clipped__31_comb[6:0]};
  assign p2_concat_84450_comb = {p2_add_84369_comb, p2_clipped__111_comb[6:0]};
  assign p2_concat_84453_comb = {p2_add_84375_comb, p2_clipped__9_comb[6:0]};
  assign p2_concat_84454_comb = {p2_add_84377_comb, p2_clipped__121_comb[6:0]};
  assign p2_concat_84455_comb = {p2_add_84379_comb, p2_clipped__10_comb[6:0]};
  assign p2_concat_84456_comb = {p2_add_84381_comb, p2_clipped__122_comb[6:0]};
  assign p2_concat_84457_comb = {p2_add_84383_comb, p2_clipped__11_comb[6:0]};
  assign p2_concat_84458_comb = {p2_add_84385_comb, p2_clipped__123_comb[6:0]};
  assign p2_concat_84461_comb = {p2_add_84391_comb, p2_clipped__13_comb[6:0]};
  assign p2_concat_84462_comb = {p2_add_84393_comb, p2_clipped__125_comb[6:0]};
  assign p2_concat_84463_comb = {p2_add_84395_comb, p2_clipped__14_comb[6:0]};
  assign p2_concat_84464_comb = {p2_add_84397_comb, p2_clipped__126_comb[6:0]};
  assign p2_concat_84465_comb = {p2_add_84399_comb, p2_clipped__15_comb[6:0]};
  assign p2_concat_84466_comb = {p2_add_84401_comb, p2_clipped__127_comb[6:0]};
  assign p2_smul_84659_comb = smul20b_11b_x_9b(p2_concat_84451_comb, 9'h0fb);
  assign p2_smul_84660_comb = smul20b_11b_x_9b(p2_concat_84435_comb, 9'h0d5);
  assign p2_smul_84669_comb = smul20b_11b_x_9b(p2_concat_84436_comb, 9'h12b);
  assign p2_smul_84670_comb = smul20b_11b_x_9b(p2_concat_84452_comb, 9'h105);
  assign p2_smul_84819_comb = smul20b_11b_x_9b(p2_concat_84451_comb, 9'h0d5);
  assign p2_smul_84821_comb = smul20b_11b_x_9b(p2_concat_84403_comb, 9'h105);
  assign p2_smul_84826_comb = smul20b_11b_x_9b(p2_concat_84406_comb, 9'h0fb);
  assign p2_smul_84828_comb = smul20b_11b_x_9b(p2_concat_84452_comb, 9'h12b);
  assign p2_smul_84901_comb = smul20b_11b_x_9b(p2_concat_84435_comb, 9'h105);
  assign p2_smul_84903_comb = smul20b_11b_x_9b(p2_concat_84404_comb, 9'h0d5);
  assign p2_smul_84904_comb = smul20b_11b_x_9b(p2_concat_84405_comb, 9'h0d5);
  assign p2_smul_84906_comb = smul20b_11b_x_9b(p2_concat_84436_comb, 9'h105);
  assign p2_smul_85015_comb = smul20b_11b_x_9b(p2_concat_84403_comb, 9'h0d5);
  assign p2_smul_85016_comb = smul20b_11b_x_9b(p2_concat_84404_comb, 9'h105);
  assign p2_smul_85017_comb = smul20b_11b_x_9b(p2_concat_84405_comb, 9'h105);
  assign p2_smul_85018_comb = smul20b_11b_x_9b(p2_concat_84406_comb, 9'h0d5);
  assign p2_add_85131_comb = p2_smul_84707_comb + p2_smul_84708_comb;
  assign p2_smul_85132_comb = smul18b_18b_x_8b(p2_sign_ext_84501_comb[17:0], 8'h47);
  assign p2_smul_85133_comb = smul18b_18b_x_6b(p2_sign_ext_84502_comb[17:0], 6'h19);
  assign p2_smul_85134_comb = smul18b_18b_x_6b(p2_sign_ext_84503_comb[17:0], 6'h27);
  assign p2_smul_85135_comb = smul18b_18b_x_8b(p2_sign_ext_84504_comb[17:0], 8'hb9);
  assign p2_add_85136_comb = p2_smul_84717_comb + p2_smul_84718_comb;
  assign p2_smul_85188_comb = smul19b_19b_x_7b(p2_sign_ext_84539_comb[18:0], 7'h31);
  assign p2_smul_85189_comb = smul19b_19b_x_7b(p2_sign_ext_84501_comb[18:0], 7'h4f);
  assign p2_smul_85192_comb = smul19b_19b_x_7b(p2_sign_ext_84504_comb[18:0], 7'h4f);
  assign p2_smul_85193_comb = smul19b_19b_x_7b(p2_sign_ext_84540_comb[18:0], 7'h31);
  assign p2_smul_85252_comb = smul19b_19b_x_6b(p2_sign_ext_84539_comb[18:0], 6'h27);
  assign p2_smul_85254_comb = smul19b_19b_x_8b(p2_sign_ext_84502_comb[18:0], 8'hb9);
  assign p2_smul_85255_comb = smul19b_19b_x_8b(p2_sign_ext_84503_comb[18:0], 8'h47);
  assign p2_smul_85257_comb = smul19b_19b_x_6b(p2_sign_ext_84540_comb[18:0], 6'h19);
  assign p2_smul_85379_comb = smul19b_19b_x_8b(p2_sign_ext_84603_comb[18:0], 8'h47);
  assign p2_smul_85381_comb = smul19b_19b_x_6b(p2_sign_ext_84501_comb[18:0], 6'h27);
  assign p2_smul_85384_comb = smul19b_19b_x_6b(p2_sign_ext_84504_comb[18:0], 6'h27);
  assign p2_smul_85386_comb = smul19b_19b_x_8b(p2_sign_ext_84608_comb[18:0], 8'h47);
  assign p2_smul_85443_comb = smul19b_19b_x_7b(p2_sign_ext_84603_comb[18:0], 7'h31);
  assign p2_smul_85445_comb = smul19b_19b_x_7b(p2_sign_ext_84501_comb[18:0], 7'h31);
  assign p2_smul_85448_comb = smul19b_19b_x_7b(p2_sign_ext_84504_comb[18:0], 7'h31);
  assign p2_smul_85450_comb = smul19b_19b_x_7b(p2_sign_ext_84608_comb[18:0], 7'h31);
  assign p2_smul_85499_comb = smul18b_18b_x_6b(p2_sign_ext_84603_comb[17:0], 6'h19);
  assign p2_smul_85500_comb = smul18b_18b_x_8b(p2_sign_ext_84539_comb[17:0], 8'hb9);
  assign p2_add_85501_comb = p2_smul_85063_comb + p2_smul_85064_comb;
  assign p2_add_85502_comb = p2_smul_85065_comb + p2_smul_85066_comb;
  assign p2_smul_85503_comb = smul18b_18b_x_8b(p2_sign_ext_84540_comb[17:0], 8'hb9);
  assign p2_smul_85504_comb = smul18b_18b_x_6b(p2_sign_ext_84608_comb[17:0], 6'h19);
  assign p2_smul_85747_comb = smul19b_11b_x_9b(p2_concat_84451_comb, 9'h0b5);
  assign p2_smul_85748_comb = smul19b_11b_x_9b(p2_concat_84435_comb, 9'h14b);
  assign p2_smul_85749_comb = smul19b_11b_x_9b(p2_concat_84403_comb, 9'h14b);
  assign p2_smul_85750_comb = smul19b_11b_x_9b(p2_concat_84404_comb, 9'h0b5);
  assign p2_smul_85751_comb = smul19b_11b_x_9b(p2_concat_84405_comb, 9'h0b5);
  assign p2_smul_85752_comb = smul19b_11b_x_9b(p2_concat_84406_comb, 9'h14b);
  assign p2_smul_85753_comb = smul19b_11b_x_9b(p2_concat_84436_comb, 9'h14b);
  assign p2_smul_85754_comb = smul19b_11b_x_9b(p2_concat_84452_comb, 9'h0b5);
  assign p2_smul_85779_comb = smul19b_11b_x_9b(p2_concat_84459_comb, 9'h0b5);
  assign p2_smul_85780_comb = smul19b_11b_x_9b(p2_concat_84443_comb, 9'h14b);
  assign p2_smul_85781_comb = smul19b_11b_x_9b(p2_concat_84419_comb, 9'h14b);
  assign p2_smul_85782_comb = smul19b_11b_x_9b(p2_concat_84420_comb, 9'h0b5);
  assign p2_smul_85783_comb = smul19b_11b_x_9b(p2_concat_84421_comb, 9'h0b5);
  assign p2_smul_85784_comb = smul19b_11b_x_9b(p2_concat_84422_comb, 9'h14b);
  assign p2_smul_85785_comb = smul19b_11b_x_9b(p2_concat_84444_comb, 9'h14b);
  assign p2_smul_85786_comb = smul19b_11b_x_9b(p2_concat_84460_comb, 9'h0b5);
  assign p2_sign_ext_84477_comb = {{13{p2_concat_84407_comb[10]}}, p2_concat_84407_comb};
  assign p2_sign_ext_84478_comb = {{13{p2_concat_84408_comb[10]}}, p2_concat_84408_comb};
  assign p2_sign_ext_84479_comb = {{13{p2_concat_84409_comb[10]}}, p2_concat_84409_comb};
  assign p2_sign_ext_84480_comb = {{13{p2_concat_84410_comb[10]}}, p2_concat_84410_comb};
  assign p2_sign_ext_84485_comb = {{13{p2_concat_84411_comb[10]}}, p2_concat_84411_comb};
  assign p2_sign_ext_84486_comb = {{13{p2_concat_84412_comb[10]}}, p2_concat_84412_comb};
  assign p2_sign_ext_84487_comb = {{13{p2_concat_84413_comb[10]}}, p2_concat_84413_comb};
  assign p2_sign_ext_84488_comb = {{13{p2_concat_84414_comb[10]}}, p2_concat_84414_comb};
  assign p2_sign_ext_84493_comb = {{13{p2_concat_84415_comb[10]}}, p2_concat_84415_comb};
  assign p2_sign_ext_84494_comb = {{13{p2_concat_84416_comb[10]}}, p2_concat_84416_comb};
  assign p2_sign_ext_84495_comb = {{13{p2_concat_84417_comb[10]}}, p2_concat_84417_comb};
  assign p2_sign_ext_84496_comb = {{13{p2_concat_84418_comb[10]}}, p2_concat_84418_comb};
  assign p2_sign_ext_84509_comb = {{13{p2_concat_84423_comb[10]}}, p2_concat_84423_comb};
  assign p2_sign_ext_84510_comb = {{13{p2_concat_84424_comb[10]}}, p2_concat_84424_comb};
  assign p2_sign_ext_84511_comb = {{13{p2_concat_84425_comb[10]}}, p2_concat_84425_comb};
  assign p2_sign_ext_84512_comb = {{13{p2_concat_84426_comb[10]}}, p2_concat_84426_comb};
  assign p2_sign_ext_84517_comb = {{13{p2_concat_84427_comb[10]}}, p2_concat_84427_comb};
  assign p2_sign_ext_84518_comb = {{13{p2_concat_84428_comb[10]}}, p2_concat_84428_comb};
  assign p2_sign_ext_84519_comb = {{13{p2_concat_84429_comb[10]}}, p2_concat_84429_comb};
  assign p2_sign_ext_84520_comb = {{13{p2_concat_84430_comb[10]}}, p2_concat_84430_comb};
  assign p2_sign_ext_84525_comb = {{13{p2_concat_84431_comb[10]}}, p2_concat_84431_comb};
  assign p2_sign_ext_84526_comb = {{13{p2_concat_84432_comb[10]}}, p2_concat_84432_comb};
  assign p2_sign_ext_84527_comb = {{13{p2_concat_84433_comb[10]}}, p2_concat_84433_comb};
  assign p2_sign_ext_84528_comb = {{13{p2_concat_84434_comb[10]}}, p2_concat_84434_comb};
  assign p2_sign_ext_84533_comb = {{13{p2_concat_84437_comb[10]}}, p2_concat_84437_comb};
  assign p2_sign_ext_84534_comb = {{13{p2_concat_84438_comb[10]}}, p2_concat_84438_comb};
  assign p2_sign_ext_84535_comb = {{13{p2_concat_84439_comb[10]}}, p2_concat_84439_comb};
  assign p2_sign_ext_84536_comb = {{13{p2_concat_84440_comb[10]}}, p2_concat_84440_comb};
  assign p2_sign_ext_84537_comb = {{13{p2_concat_84441_comb[10]}}, p2_concat_84441_comb};
  assign p2_sign_ext_84538_comb = {{13{p2_concat_84442_comb[10]}}, p2_concat_84442_comb};
  assign p2_sign_ext_84541_comb = {{13{p2_concat_84445_comb[10]}}, p2_concat_84445_comb};
  assign p2_sign_ext_84542_comb = {{13{p2_concat_84446_comb[10]}}, p2_concat_84446_comb};
  assign p2_sign_ext_84543_comb = {{13{p2_concat_84447_comb[10]}}, p2_concat_84447_comb};
  assign p2_sign_ext_84544_comb = {{13{p2_concat_84448_comb[10]}}, p2_concat_84448_comb};
  assign p2_sign_ext_84545_comb = {{13{p2_concat_84449_comb[10]}}, p2_concat_84449_comb};
  assign p2_sign_ext_84546_comb = {{13{p2_concat_84450_comb[10]}}, p2_concat_84450_comb};
  assign p2_sign_ext_84585_comb = {{13{p2_concat_84453_comb[10]}}, p2_concat_84453_comb};
  assign p2_sign_ext_84590_comb = {{13{p2_concat_84454_comb[10]}}, p2_concat_84454_comb};
  assign p2_sign_ext_84591_comb = {{13{p2_concat_84455_comb[10]}}, p2_concat_84455_comb};
  assign p2_sign_ext_84596_comb = {{13{p2_concat_84456_comb[10]}}, p2_concat_84456_comb};
  assign p2_sign_ext_84597_comb = {{13{p2_concat_84457_comb[10]}}, p2_concat_84457_comb};
  assign p2_sign_ext_84602_comb = {{13{p2_concat_84458_comb[10]}}, p2_concat_84458_comb};
  assign p2_sign_ext_84609_comb = {{13{p2_concat_84461_comb[10]}}, p2_concat_84461_comb};
  assign p2_sign_ext_84614_comb = {{13{p2_concat_84462_comb[10]}}, p2_concat_84462_comb};
  assign p2_sign_ext_84615_comb = {{13{p2_concat_84463_comb[10]}}, p2_concat_84463_comb};
  assign p2_sign_ext_84620_comb = {{13{p2_concat_84464_comb[10]}}, p2_concat_84464_comb};
  assign p2_sign_ext_84621_comb = {{13{p2_concat_84465_comb[10]}}, p2_concat_84465_comb};
  assign p2_sign_ext_84626_comb = {{13{p2_concat_84466_comb[10]}}, p2_concat_84466_comb};
  assign p2_add_85107_comb = p2_smul_84659_comb + p2_smul_84660_comb;
  assign p2_smul_85108_comb = smul18b_18b_x_8b(p2_sign_ext_84469_comb[17:0], 8'h47);
  assign p2_smul_85109_comb = smul18b_18b_x_6b(p2_sign_ext_84470_comb[17:0], 6'h19);
  assign p2_smul_85110_comb = smul18b_18b_x_6b(p2_sign_ext_84471_comb[17:0], 6'h27);
  assign p2_smul_85111_comb = smul18b_18b_x_8b(p2_sign_ext_84472_comb[17:0], 8'hb9);
  assign p2_add_85112_comb = p2_smul_84669_comb + p2_smul_84670_comb;
  assign p2_smul_85156_comb = smul19b_19b_x_7b(p2_sign_ext_84531_comb[18:0], 7'h31);
  assign p2_smul_85157_comb = smul19b_19b_x_7b(p2_sign_ext_84469_comb[18:0], 7'h4f);
  assign p2_smul_85160_comb = smul19b_19b_x_7b(p2_sign_ext_84472_comb[18:0], 7'h4f);
  assign p2_smul_85161_comb = smul19b_19b_x_7b(p2_sign_ext_84532_comb[18:0], 7'h31);
  assign p2_smul_85220_comb = smul19b_19b_x_6b(p2_sign_ext_84531_comb[18:0], 6'h27);
  assign p2_smul_85222_comb = smul19b_19b_x_8b(p2_sign_ext_84470_comb[18:0], 8'hb9);
  assign p2_smul_85223_comb = smul19b_19b_x_8b(p2_sign_ext_84471_comb[18:0], 8'h47);
  assign p2_smul_85225_comb = smul19b_19b_x_6b(p2_sign_ext_84532_comb[18:0], 6'h19);
  assign p2_smul_85347_comb = smul19b_19b_x_8b(p2_sign_ext_84579_comb[18:0], 8'h47);
  assign p2_smul_85349_comb = smul19b_19b_x_6b(p2_sign_ext_84469_comb[18:0], 6'h27);
  assign p2_smul_85352_comb = smul19b_19b_x_6b(p2_sign_ext_84472_comb[18:0], 6'h27);
  assign p2_smul_85354_comb = smul19b_19b_x_8b(p2_sign_ext_84584_comb[18:0], 8'h47);
  assign p2_smul_85411_comb = smul19b_19b_x_7b(p2_sign_ext_84579_comb[18:0], 7'h31);
  assign p2_smul_85413_comb = smul19b_19b_x_7b(p2_sign_ext_84469_comb[18:0], 7'h31);
  assign p2_smul_85416_comb = smul19b_19b_x_7b(p2_sign_ext_84472_comb[18:0], 7'h31);
  assign p2_smul_85418_comb = smul19b_19b_x_7b(p2_sign_ext_84584_comb[18:0], 7'h31);
  assign p2_smul_85475_comb = smul18b_18b_x_6b(p2_sign_ext_84579_comb[17:0], 6'h19);
  assign p2_smul_85476_comb = smul18b_18b_x_8b(p2_sign_ext_84531_comb[17:0], 8'hb9);
  assign p2_add_85477_comb = p2_smul_85015_comb + p2_smul_85016_comb;
  assign p2_add_85478_comb = p2_smul_85017_comb + p2_smul_85018_comb;
  assign p2_smul_85479_comb = smul18b_18b_x_8b(p2_sign_ext_84532_comb[17:0], 8'hb9);
  assign p2_smul_85480_comb = smul18b_18b_x_6b(p2_sign_ext_84584_comb[17:0], 6'h19);
  assign p2_bit_slice_85603_comb = p2_add_85131_comb[19:1];
  assign p2_add_85604_comb = p2_smul_85132_comb + p2_smul_85133_comb;
  assign p2_add_85605_comb = p2_smul_85134_comb + p2_smul_85135_comb;
  assign p2_bit_slice_85606_comb = p2_add_85136_comb[19:1];
  assign p2_smul_85651_comb = smul18b_18b_x_7b(p2_sign_ext_84603_comb[17:0], 7'h3b);
  assign p2_smul_85654_comb = smul18b_18b_x_7b(p2_sign_ext_84502_comb[17:0], 7'h45);
  assign p2_smul_85655_comb = smul18b_18b_x_7b(p2_sign_ext_84503_comb[17:0], 7'h45);
  assign p2_smul_85658_comb = smul18b_18b_x_7b(p2_sign_ext_84608_comb[17:0], 7'h3b);
  assign p2_add_85715_comb = p2_smul_84859_comb[19:1] + p2_smul_85252_comb;
  assign p2_add_85717_comb = p2_smul_84861_comb[19:1] + p2_smul_85254_comb;
  assign p2_add_85719_comb = p2_smul_85255_comb + p2_smul_84866_comb[19:1];
  assign p2_add_85721_comb = p2_smul_85257_comb + p2_smul_84868_comb[19:1];
  assign p2_smul_85755_comb = smul19b_11b_x_9b(p2_concat_84453_comb, 9'h0b5);
  assign p2_smul_85756_comb = smul19b_11b_x_9b(p2_concat_84437_comb, 9'h14b);
  assign p2_smul_85757_comb = smul19b_11b_x_9b(p2_concat_84407_comb, 9'h14b);
  assign p2_smul_85758_comb = smul19b_11b_x_9b(p2_concat_84408_comb, 9'h0b5);
  assign p2_smul_85759_comb = smul19b_11b_x_9b(p2_concat_84409_comb, 9'h0b5);
  assign p2_smul_85760_comb = smul19b_11b_x_9b(p2_concat_84410_comb, 9'h14b);
  assign p2_smul_85761_comb = smul19b_11b_x_9b(p2_concat_84438_comb, 9'h14b);
  assign p2_smul_85762_comb = smul19b_11b_x_9b(p2_concat_84454_comb, 9'h0b5);
  assign p2_smul_85763_comb = smul19b_11b_x_9b(p2_concat_84455_comb, 9'h0b5);
  assign p2_smul_85764_comb = smul19b_11b_x_9b(p2_concat_84439_comb, 9'h14b);
  assign p2_smul_85765_comb = smul19b_11b_x_9b(p2_concat_84411_comb, 9'h14b);
  assign p2_smul_85766_comb = smul19b_11b_x_9b(p2_concat_84412_comb, 9'h0b5);
  assign p2_smul_85767_comb = smul19b_11b_x_9b(p2_concat_84413_comb, 9'h0b5);
  assign p2_smul_85768_comb = smul19b_11b_x_9b(p2_concat_84414_comb, 9'h14b);
  assign p2_smul_85769_comb = smul19b_11b_x_9b(p2_concat_84440_comb, 9'h14b);
  assign p2_smul_85770_comb = smul19b_11b_x_9b(p2_concat_84456_comb, 9'h0b5);
  assign p2_smul_85771_comb = smul19b_11b_x_9b(p2_concat_84457_comb, 9'h0b5);
  assign p2_smul_85772_comb = smul19b_11b_x_9b(p2_concat_84441_comb, 9'h14b);
  assign p2_smul_85773_comb = smul19b_11b_x_9b(p2_concat_84415_comb, 9'h14b);
  assign p2_smul_85774_comb = smul19b_11b_x_9b(p2_concat_84416_comb, 9'h0b5);
  assign p2_smul_85775_comb = smul19b_11b_x_9b(p2_concat_84417_comb, 9'h0b5);
  assign p2_smul_85776_comb = smul19b_11b_x_9b(p2_concat_84418_comb, 9'h14b);
  assign p2_smul_85777_comb = smul19b_11b_x_9b(p2_concat_84442_comb, 9'h14b);
  assign p2_smul_85778_comb = smul19b_11b_x_9b(p2_concat_84458_comb, 9'h0b5);
  assign p2_smul_85787_comb = smul19b_11b_x_9b(p2_concat_84461_comb, 9'h0b5);
  assign p2_smul_85788_comb = smul19b_11b_x_9b(p2_concat_84445_comb, 9'h14b);
  assign p2_smul_85789_comb = smul19b_11b_x_9b(p2_concat_84423_comb, 9'h14b);
  assign p2_smul_85790_comb = smul19b_11b_x_9b(p2_concat_84424_comb, 9'h0b5);
  assign p2_smul_85791_comb = smul19b_11b_x_9b(p2_concat_84425_comb, 9'h0b5);
  assign p2_smul_85792_comb = smul19b_11b_x_9b(p2_concat_84426_comb, 9'h14b);
  assign p2_smul_85793_comb = smul19b_11b_x_9b(p2_concat_84446_comb, 9'h14b);
  assign p2_smul_85794_comb = smul19b_11b_x_9b(p2_concat_84462_comb, 9'h0b5);
  assign p2_smul_85795_comb = smul19b_11b_x_9b(p2_concat_84463_comb, 9'h0b5);
  assign p2_smul_85796_comb = smul19b_11b_x_9b(p2_concat_84447_comb, 9'h14b);
  assign p2_smul_85797_comb = smul19b_11b_x_9b(p2_concat_84427_comb, 9'h14b);
  assign p2_smul_85798_comb = smul19b_11b_x_9b(p2_concat_84428_comb, 9'h0b5);
  assign p2_smul_85799_comb = smul19b_11b_x_9b(p2_concat_84429_comb, 9'h0b5);
  assign p2_smul_85800_comb = smul19b_11b_x_9b(p2_concat_84430_comb, 9'h14b);
  assign p2_smul_85801_comb = smul19b_11b_x_9b(p2_concat_84448_comb, 9'h14b);
  assign p2_smul_85802_comb = smul19b_11b_x_9b(p2_concat_84464_comb, 9'h0b5);
  assign p2_smul_85803_comb = smul19b_11b_x_9b(p2_concat_84465_comb, 9'h0b5);
  assign p2_smul_85804_comb = smul19b_11b_x_9b(p2_concat_84449_comb, 9'h14b);
  assign p2_smul_85805_comb = smul19b_11b_x_9b(p2_concat_84431_comb, 9'h14b);
  assign p2_smul_85806_comb = smul19b_11b_x_9b(p2_concat_84432_comb, 9'h0b5);
  assign p2_smul_85807_comb = smul19b_11b_x_9b(p2_concat_84433_comb, 9'h0b5);
  assign p2_smul_85808_comb = smul19b_11b_x_9b(p2_concat_84434_comb, 9'h14b);
  assign p2_smul_85809_comb = smul19b_11b_x_9b(p2_concat_84450_comb, 9'h14b);
  assign p2_smul_85810_comb = smul19b_11b_x_9b(p2_concat_84466_comb, 9'h0b5);
  assign p2_add_85843_comb = p2_smul_85379_comb + p2_smul_84941_comb[19:1];
  assign p2_add_85845_comb = p2_smul_85381_comb + p2_smul_84943_comb[19:1];
  assign p2_add_85847_comb = p2_smul_84944_comb[19:1] + p2_smul_85384_comb;
  assign p2_add_85849_comb = p2_smul_84946_comb[19:1] + p2_smul_85386_comb;
  assign p2_smul_85908_comb = smul18b_18b_x_7b(p2_sign_ext_84539_comb[17:0], 7'h45);
  assign p2_smul_85910_comb = smul18b_18b_x_7b(p2_sign_ext_84502_comb[17:0], 7'h3b);
  assign p2_smul_85911_comb = smul18b_18b_x_7b(p2_sign_ext_84503_comb[17:0], 7'h3b);
  assign p2_smul_85913_comb = smul18b_18b_x_7b(p2_sign_ext_84540_comb[17:0], 7'h45);
  assign p2_add_85955_comb = p2_smul_85499_comb + p2_smul_85500_comb;
  assign p2_bit_slice_85956_comb = p2_add_85501_comb[19:1];
  assign p2_bit_slice_85957_comb = p2_add_85502_comb[19:1];
  assign p2_add_85958_comb = p2_smul_85503_comb + p2_smul_85504_comb;
  assign p2_add_85971_comb = p2_sign_ext_84579_comb[11:0] + p2_sign_ext_84531_comb[11:0];
  assign p2_add_85972_comb = p2_sign_ext_84469_comb[11:0] + p2_sign_ext_84470_comb[11:0];
  assign p2_add_85973_comb = p2_sign_ext_84471_comb[11:0] + p2_sign_ext_84472_comb[11:0];
  assign p2_add_85974_comb = p2_sign_ext_84532_comb[11:0] + p2_sign_ext_84584_comb[11:0];
  assign p2_add_85987_comb = p2_sign_ext_84603_comb[11:0] + p2_sign_ext_84539_comb[11:0];
  assign p2_add_85988_comb = p2_sign_ext_84501_comb[11:0] + p2_sign_ext_84502_comb[11:0];
  assign p2_add_85989_comb = p2_sign_ext_84503_comb[11:0] + p2_sign_ext_84504_comb[11:0];
  assign p2_add_85990_comb = p2_sign_ext_84540_comb[11:0] + p2_sign_ext_84608_comb[11:0];
  assign p2_add_86131_comb = p2_smul_85747_comb + p2_smul_85748_comb;
  assign p2_add_86132_comb = p2_smul_85749_comb + p2_smul_85750_comb;
  assign p2_add_86133_comb = p2_smul_85751_comb + p2_smul_85752_comb;
  assign p2_add_86134_comb = p2_smul_85753_comb + p2_smul_85754_comb;
  assign p2_add_86147_comb = p2_smul_85779_comb + p2_smul_85780_comb;
  assign p2_add_86148_comb = p2_smul_85781_comb + p2_smul_85782_comb;
  assign p2_add_86149_comb = p2_smul_85783_comb + p2_smul_85784_comb;
  assign p2_add_86150_comb = p2_smul_85785_comb + p2_smul_85786_comb;
  assign p2_smul_84671_comb = smul20b_11b_x_9b(p2_concat_84453_comb, 9'h0fb);
  assign p2_smul_84672_comb = smul20b_11b_x_9b(p2_concat_84437_comb, 9'h0d5);
  assign p2_smul_84681_comb = smul20b_11b_x_9b(p2_concat_84438_comb, 9'h12b);
  assign p2_smul_84682_comb = smul20b_11b_x_9b(p2_concat_84454_comb, 9'h105);
  assign p2_smul_84683_comb = smul20b_11b_x_9b(p2_concat_84455_comb, 9'h0fb);
  assign p2_smul_84684_comb = smul20b_11b_x_9b(p2_concat_84439_comb, 9'h0d5);
  assign p2_smul_84693_comb = smul20b_11b_x_9b(p2_concat_84440_comb, 9'h12b);
  assign p2_smul_84694_comb = smul20b_11b_x_9b(p2_concat_84456_comb, 9'h105);
  assign p2_smul_84695_comb = smul20b_11b_x_9b(p2_concat_84457_comb, 9'h0fb);
  assign p2_smul_84696_comb = smul20b_11b_x_9b(p2_concat_84441_comb, 9'h0d5);
  assign p2_smul_84705_comb = smul20b_11b_x_9b(p2_concat_84442_comb, 9'h12b);
  assign p2_smul_84706_comb = smul20b_11b_x_9b(p2_concat_84458_comb, 9'h105);
  assign p2_smul_84719_comb = smul20b_11b_x_9b(p2_concat_84461_comb, 9'h0fb);
  assign p2_smul_84720_comb = smul20b_11b_x_9b(p2_concat_84445_comb, 9'h0d5);
  assign p2_smul_84729_comb = smul20b_11b_x_9b(p2_concat_84446_comb, 9'h12b);
  assign p2_smul_84730_comb = smul20b_11b_x_9b(p2_concat_84462_comb, 9'h105);
  assign p2_smul_84731_comb = smul20b_11b_x_9b(p2_concat_84463_comb, 9'h0fb);
  assign p2_smul_84732_comb = smul20b_11b_x_9b(p2_concat_84447_comb, 9'h0d5);
  assign p2_smul_84741_comb = smul20b_11b_x_9b(p2_concat_84448_comb, 9'h12b);
  assign p2_smul_84742_comb = smul20b_11b_x_9b(p2_concat_84464_comb, 9'h105);
  assign p2_smul_84743_comb = smul20b_11b_x_9b(p2_concat_84465_comb, 9'h0fb);
  assign p2_smul_84744_comb = smul20b_11b_x_9b(p2_concat_84449_comb, 9'h0d5);
  assign p2_smul_84753_comb = smul20b_11b_x_9b(p2_concat_84450_comb, 9'h12b);
  assign p2_smul_84754_comb = smul20b_11b_x_9b(p2_concat_84466_comb, 9'h105);
  assign p2_smul_85027_comb = smul20b_11b_x_9b(p2_concat_84407_comb, 9'h0d5);
  assign p2_smul_85028_comb = smul20b_11b_x_9b(p2_concat_84408_comb, 9'h105);
  assign p2_smul_85029_comb = smul20b_11b_x_9b(p2_concat_84409_comb, 9'h105);
  assign p2_smul_85030_comb = smul20b_11b_x_9b(p2_concat_84410_comb, 9'h0d5);
  assign p2_smul_85039_comb = smul20b_11b_x_9b(p2_concat_84411_comb, 9'h0d5);
  assign p2_smul_85040_comb = smul20b_11b_x_9b(p2_concat_84412_comb, 9'h105);
  assign p2_smul_85041_comb = smul20b_11b_x_9b(p2_concat_84413_comb, 9'h105);
  assign p2_smul_85042_comb = smul20b_11b_x_9b(p2_concat_84414_comb, 9'h0d5);
  assign p2_smul_85051_comb = smul20b_11b_x_9b(p2_concat_84415_comb, 9'h0d5);
  assign p2_smul_85052_comb = smul20b_11b_x_9b(p2_concat_84416_comb, 9'h105);
  assign p2_smul_85053_comb = smul20b_11b_x_9b(p2_concat_84417_comb, 9'h105);
  assign p2_smul_85054_comb = smul20b_11b_x_9b(p2_concat_84418_comb, 9'h0d5);
  assign p2_smul_85075_comb = smul20b_11b_x_9b(p2_concat_84423_comb, 9'h0d5);
  assign p2_smul_85076_comb = smul20b_11b_x_9b(p2_concat_84424_comb, 9'h105);
  assign p2_smul_85077_comb = smul20b_11b_x_9b(p2_concat_84425_comb, 9'h105);
  assign p2_smul_85078_comb = smul20b_11b_x_9b(p2_concat_84426_comb, 9'h0d5);
  assign p2_smul_85087_comb = smul20b_11b_x_9b(p2_concat_84427_comb, 9'h0d5);
  assign p2_smul_85088_comb = smul20b_11b_x_9b(p2_concat_84428_comb, 9'h105);
  assign p2_smul_85089_comb = smul20b_11b_x_9b(p2_concat_84429_comb, 9'h105);
  assign p2_smul_85090_comb = smul20b_11b_x_9b(p2_concat_84430_comb, 9'h0d5);
  assign p2_smul_85099_comb = smul20b_11b_x_9b(p2_concat_84431_comb, 9'h0d5);
  assign p2_smul_85100_comb = smul20b_11b_x_9b(p2_concat_84432_comb, 9'h105);
  assign p2_smul_85101_comb = smul20b_11b_x_9b(p2_concat_84433_comb, 9'h105);
  assign p2_smul_85102_comb = smul20b_11b_x_9b(p2_concat_84434_comb, 9'h0d5);
  assign p2_bit_slice_85587_comb = p2_add_85107_comb[19:1];
  assign p2_add_85588_comb = p2_smul_85108_comb + p2_smul_85109_comb;
  assign p2_add_85589_comb = p2_smul_85110_comb + p2_smul_85111_comb;
  assign p2_bit_slice_85590_comb = p2_add_85112_comb[19:1];
  assign p2_smul_85619_comb = smul18b_18b_x_7b(p2_sign_ext_84579_comb[17:0], 7'h3b);
  assign p2_smul_85622_comb = smul18b_18b_x_7b(p2_sign_ext_84470_comb[17:0], 7'h45);
  assign p2_smul_85623_comb = smul18b_18b_x_7b(p2_sign_ext_84471_comb[17:0], 7'h45);
  assign p2_smul_85626_comb = smul18b_18b_x_7b(p2_sign_ext_84584_comb[17:0], 7'h3b);
  assign p2_add_85683_comb = p2_smul_84819_comb[19:1] + p2_smul_85220_comb;
  assign p2_add_85685_comb = p2_smul_84821_comb[19:1] + p2_smul_85222_comb;
  assign p2_add_85687_comb = p2_smul_85223_comb + p2_smul_84826_comb[19:1];
  assign p2_add_85689_comb = p2_smul_85225_comb + p2_smul_84828_comb[19:1];
  assign p2_add_85811_comb = p2_smul_85347_comb + p2_smul_84901_comb[19:1];
  assign p2_add_85813_comb = p2_smul_85349_comb + p2_smul_84903_comb[19:1];
  assign p2_add_85815_comb = p2_smul_84904_comb[19:1] + p2_smul_85352_comb;
  assign p2_add_85817_comb = p2_smul_84906_comb[19:1] + p2_smul_85354_comb;
  assign p2_smul_85876_comb = smul18b_18b_x_7b(p2_sign_ext_84531_comb[17:0], 7'h45);
  assign p2_smul_85878_comb = smul18b_18b_x_7b(p2_sign_ext_84470_comb[17:0], 7'h3b);
  assign p2_smul_85879_comb = smul18b_18b_x_7b(p2_sign_ext_84471_comb[17:0], 7'h3b);
  assign p2_smul_85881_comb = smul18b_18b_x_7b(p2_sign_ext_84532_comb[17:0], 7'h45);
  assign p2_add_85939_comb = p2_smul_85475_comb + p2_smul_85476_comb;
  assign p2_bit_slice_85940_comb = p2_add_85477_comb[19:1];
  assign p2_bit_slice_85941_comb = p2_add_85478_comb[19:1];
  assign p2_add_85942_comb = p2_smul_85479_comb + p2_smul_85480_comb;
  assign p2_add_86067_comb = p2_smul_85651_comb + p2_smul_85188_comb[18:1];
  assign p2_add_86069_comb = p2_smul_85189_comb[18:1] + p2_smul_85654_comb;
  assign p2_add_86071_comb = p2_smul_85655_comb + p2_smul_85192_comb[18:1];
  assign p2_add_86073_comb = p2_smul_85193_comb[18:1] + p2_smul_85658_comb;
  assign p2_concat_86115_comb = {p2_add_85715_comb, p2_smul_84859_comb[0]};
  assign p2_concat_86116_comb = {p2_add_85717_comb, p2_smul_84861_comb[0]};
  assign p2_concat_86117_comb = {p2_add_85719_comb, p2_smul_84866_comb[0]};
  assign p2_concat_86118_comb = {p2_add_85721_comb, p2_smul_84868_comb[0]};
  assign p2_add_86135_comb = p2_smul_85755_comb + p2_smul_85756_comb;
  assign p2_add_86136_comb = p2_smul_85757_comb + p2_smul_85758_comb;
  assign p2_add_86137_comb = p2_smul_85759_comb + p2_smul_85760_comb;
  assign p2_add_86138_comb = p2_smul_85761_comb + p2_smul_85762_comb;
  assign p2_add_86139_comb = p2_smul_85763_comb + p2_smul_85764_comb;
  assign p2_add_86140_comb = p2_smul_85765_comb + p2_smul_85766_comb;
  assign p2_add_86141_comb = p2_smul_85767_comb + p2_smul_85768_comb;
  assign p2_add_86142_comb = p2_smul_85769_comb + p2_smul_85770_comb;
  assign p2_add_86143_comb = p2_smul_85771_comb + p2_smul_85772_comb;
  assign p2_add_86144_comb = p2_smul_85773_comb + p2_smul_85774_comb;
  assign p2_add_86145_comb = p2_smul_85775_comb + p2_smul_85776_comb;
  assign p2_add_86146_comb = p2_smul_85777_comb + p2_smul_85778_comb;
  assign p2_add_86151_comb = p2_smul_85787_comb + p2_smul_85788_comb;
  assign p2_add_86152_comb = p2_smul_85789_comb + p2_smul_85790_comb;
  assign p2_add_86153_comb = p2_smul_85791_comb + p2_smul_85792_comb;
  assign p2_add_86154_comb = p2_smul_85793_comb + p2_smul_85794_comb;
  assign p2_add_86155_comb = p2_smul_85795_comb + p2_smul_85796_comb;
  assign p2_add_86156_comb = p2_smul_85797_comb + p2_smul_85798_comb;
  assign p2_add_86157_comb = p2_smul_85799_comb + p2_smul_85800_comb;
  assign p2_add_86158_comb = p2_smul_85801_comb + p2_smul_85802_comb;
  assign p2_add_86159_comb = p2_smul_85803_comb + p2_smul_85804_comb;
  assign p2_add_86160_comb = p2_smul_85805_comb + p2_smul_85806_comb;
  assign p2_add_86161_comb = p2_smul_85807_comb + p2_smul_85808_comb;
  assign p2_add_86162_comb = p2_smul_85809_comb + p2_smul_85810_comb;
  assign p2_concat_86179_comb = {p2_add_85843_comb, p2_smul_84941_comb[0]};
  assign p2_concat_86180_comb = {p2_add_85845_comb, p2_smul_84943_comb[0]};
  assign p2_concat_86181_comb = {p2_add_85847_comb, p2_smul_84944_comb[0]};
  assign p2_concat_86182_comb = {p2_add_85849_comb, p2_smul_84946_comb[0]};
  assign p2_add_86227_comb = p2_smul_85443_comb[18:1] + p2_smul_85908_comb;
  assign p2_add_86229_comb = p2_smul_85445_comb[18:1] + p2_smul_85910_comb;
  assign p2_add_86231_comb = p2_smul_85911_comb + p2_smul_85448_comb[18:1];
  assign p2_add_86233_comb = p2_smul_85913_comb + p2_smul_85450_comb[18:1];
  assign p2_sum__1568_comb = {{6{p2_add_86131_comb[18]}}, p2_add_86131_comb};
  assign p2_sum__1569_comb = {{6{p2_add_86132_comb[18]}}, p2_add_86132_comb};
  assign p2_sum__1570_comb = {{6{p2_add_86133_comb[18]}}, p2_add_86133_comb};
  assign p2_sum__1571_comb = {{6{p2_add_86134_comb[18]}}, p2_add_86134_comb};
  assign p2_sum__1456_comb = {{6{p2_add_86147_comb[18]}}, p2_add_86147_comb};
  assign p2_sum__1457_comb = {{6{p2_add_86148_comb[18]}}, p2_add_86148_comb};
  assign p2_sum__1458_comb = {{6{p2_add_86149_comb[18]}}, p2_add_86149_comb};
  assign p2_sum__1459_comb = {{6{p2_add_86150_comb[18]}}, p2_add_86150_comb};
  assign p2_smul_84829_comb = smul20b_11b_x_9b(p2_concat_84453_comb, 9'h0d5);
  assign p2_smul_84831_comb = smul20b_11b_x_9b(p2_concat_84407_comb, 9'h105);
  assign p2_smul_84836_comb = smul20b_11b_x_9b(p2_concat_84410_comb, 9'h0fb);
  assign p2_smul_84838_comb = smul20b_11b_x_9b(p2_concat_84454_comb, 9'h12b);
  assign p2_smul_84839_comb = smul20b_11b_x_9b(p2_concat_84455_comb, 9'h0d5);
  assign p2_smul_84841_comb = smul20b_11b_x_9b(p2_concat_84411_comb, 9'h105);
  assign p2_smul_84846_comb = smul20b_11b_x_9b(p2_concat_84414_comb, 9'h0fb);
  assign p2_smul_84848_comb = smul20b_11b_x_9b(p2_concat_84456_comb, 9'h12b);
  assign p2_smul_84849_comb = smul20b_11b_x_9b(p2_concat_84457_comb, 9'h0d5);
  assign p2_smul_84851_comb = smul20b_11b_x_9b(p2_concat_84415_comb, 9'h105);
  assign p2_smul_84856_comb = smul20b_11b_x_9b(p2_concat_84418_comb, 9'h0fb);
  assign p2_smul_84858_comb = smul20b_11b_x_9b(p2_concat_84458_comb, 9'h12b);
  assign p2_smul_84869_comb = smul20b_11b_x_9b(p2_concat_84461_comb, 9'h0d5);
  assign p2_smul_84871_comb = smul20b_11b_x_9b(p2_concat_84423_comb, 9'h105);
  assign p2_smul_84876_comb = smul20b_11b_x_9b(p2_concat_84426_comb, 9'h0fb);
  assign p2_smul_84878_comb = smul20b_11b_x_9b(p2_concat_84462_comb, 9'h12b);
  assign p2_smul_84879_comb = smul20b_11b_x_9b(p2_concat_84463_comb, 9'h0d5);
  assign p2_smul_84881_comb = smul20b_11b_x_9b(p2_concat_84427_comb, 9'h105);
  assign p2_smul_84886_comb = smul20b_11b_x_9b(p2_concat_84430_comb, 9'h0fb);
  assign p2_smul_84888_comb = smul20b_11b_x_9b(p2_concat_84464_comb, 9'h12b);
  assign p2_smul_84889_comb = smul20b_11b_x_9b(p2_concat_84465_comb, 9'h0d5);
  assign p2_smul_84891_comb = smul20b_11b_x_9b(p2_concat_84431_comb, 9'h105);
  assign p2_smul_84896_comb = smul20b_11b_x_9b(p2_concat_84434_comb, 9'h0fb);
  assign p2_smul_84898_comb = smul20b_11b_x_9b(p2_concat_84466_comb, 9'h12b);
  assign p2_smul_84911_comb = smul20b_11b_x_9b(p2_concat_84437_comb, 9'h105);
  assign p2_smul_84913_comb = smul20b_11b_x_9b(p2_concat_84408_comb, 9'h0d5);
  assign p2_smul_84914_comb = smul20b_11b_x_9b(p2_concat_84409_comb, 9'h0d5);
  assign p2_smul_84916_comb = smul20b_11b_x_9b(p2_concat_84438_comb, 9'h105);
  assign p2_smul_84921_comb = smul20b_11b_x_9b(p2_concat_84439_comb, 9'h105);
  assign p2_smul_84923_comb = smul20b_11b_x_9b(p2_concat_84412_comb, 9'h0d5);
  assign p2_smul_84924_comb = smul20b_11b_x_9b(p2_concat_84413_comb, 9'h0d5);
  assign p2_smul_84926_comb = smul20b_11b_x_9b(p2_concat_84440_comb, 9'h105);
  assign p2_smul_84931_comb = smul20b_11b_x_9b(p2_concat_84441_comb, 9'h105);
  assign p2_smul_84933_comb = smul20b_11b_x_9b(p2_concat_84416_comb, 9'h0d5);
  assign p2_smul_84934_comb = smul20b_11b_x_9b(p2_concat_84417_comb, 9'h0d5);
  assign p2_smul_84936_comb = smul20b_11b_x_9b(p2_concat_84442_comb, 9'h105);
  assign p2_smul_84951_comb = smul20b_11b_x_9b(p2_concat_84445_comb, 9'h105);
  assign p2_smul_84953_comb = smul20b_11b_x_9b(p2_concat_84424_comb, 9'h0d5);
  assign p2_smul_84954_comb = smul20b_11b_x_9b(p2_concat_84425_comb, 9'h0d5);
  assign p2_smul_84956_comb = smul20b_11b_x_9b(p2_concat_84446_comb, 9'h105);
  assign p2_smul_84961_comb = smul20b_11b_x_9b(p2_concat_84447_comb, 9'h105);
  assign p2_smul_84963_comb = smul20b_11b_x_9b(p2_concat_84428_comb, 9'h0d5);
  assign p2_smul_84964_comb = smul20b_11b_x_9b(p2_concat_84429_comb, 9'h0d5);
  assign p2_smul_84966_comb = smul20b_11b_x_9b(p2_concat_84448_comb, 9'h105);
  assign p2_smul_84971_comb = smul20b_11b_x_9b(p2_concat_84449_comb, 9'h105);
  assign p2_smul_84973_comb = smul20b_11b_x_9b(p2_concat_84432_comb, 9'h0d5);
  assign p2_smul_84974_comb = smul20b_11b_x_9b(p2_concat_84433_comb, 9'h0d5);
  assign p2_smul_84976_comb = smul20b_11b_x_9b(p2_concat_84450_comb, 9'h105);
  assign p2_add_85113_comb = p2_smul_84671_comb + p2_smul_84672_comb;
  assign p2_smul_85114_comb = smul18b_18b_x_8b(p2_sign_ext_84477_comb[17:0], 8'h47);
  assign p2_smul_85115_comb = smul18b_18b_x_6b(p2_sign_ext_84478_comb[17:0], 6'h19);
  assign p2_smul_85116_comb = smul18b_18b_x_6b(p2_sign_ext_84479_comb[17:0], 6'h27);
  assign p2_smul_85117_comb = smul18b_18b_x_8b(p2_sign_ext_84480_comb[17:0], 8'hb9);
  assign p2_add_85118_comb = p2_smul_84681_comb + p2_smul_84682_comb;
  assign p2_add_85119_comb = p2_smul_84683_comb + p2_smul_84684_comb;
  assign p2_smul_85120_comb = smul18b_18b_x_8b(p2_sign_ext_84485_comb[17:0], 8'h47);
  assign p2_smul_85121_comb = smul18b_18b_x_6b(p2_sign_ext_84486_comb[17:0], 6'h19);
  assign p2_smul_85122_comb = smul18b_18b_x_6b(p2_sign_ext_84487_comb[17:0], 6'h27);
  assign p2_smul_85123_comb = smul18b_18b_x_8b(p2_sign_ext_84488_comb[17:0], 8'hb9);
  assign p2_add_85124_comb = p2_smul_84693_comb + p2_smul_84694_comb;
  assign p2_add_85125_comb = p2_smul_84695_comb + p2_smul_84696_comb;
  assign p2_smul_85126_comb = smul18b_18b_x_8b(p2_sign_ext_84493_comb[17:0], 8'h47);
  assign p2_smul_85127_comb = smul18b_18b_x_6b(p2_sign_ext_84494_comb[17:0], 6'h19);
  assign p2_smul_85128_comb = smul18b_18b_x_6b(p2_sign_ext_84495_comb[17:0], 6'h27);
  assign p2_smul_85129_comb = smul18b_18b_x_8b(p2_sign_ext_84496_comb[17:0], 8'hb9);
  assign p2_add_85130_comb = p2_smul_84705_comb + p2_smul_84706_comb;
  assign p2_add_85137_comb = p2_smul_84719_comb + p2_smul_84720_comb;
  assign p2_smul_85138_comb = smul18b_18b_x_8b(p2_sign_ext_84509_comb[17:0], 8'h47);
  assign p2_smul_85139_comb = smul18b_18b_x_6b(p2_sign_ext_84510_comb[17:0], 6'h19);
  assign p2_smul_85140_comb = smul18b_18b_x_6b(p2_sign_ext_84511_comb[17:0], 6'h27);
  assign p2_smul_85141_comb = smul18b_18b_x_8b(p2_sign_ext_84512_comb[17:0], 8'hb9);
  assign p2_add_85142_comb = p2_smul_84729_comb + p2_smul_84730_comb;
  assign p2_add_85143_comb = p2_smul_84731_comb + p2_smul_84732_comb;
  assign p2_smul_85144_comb = smul18b_18b_x_8b(p2_sign_ext_84517_comb[17:0], 8'h47);
  assign p2_smul_85145_comb = smul18b_18b_x_6b(p2_sign_ext_84518_comb[17:0], 6'h19);
  assign p2_smul_85146_comb = smul18b_18b_x_6b(p2_sign_ext_84519_comb[17:0], 6'h27);
  assign p2_smul_85147_comb = smul18b_18b_x_8b(p2_sign_ext_84520_comb[17:0], 8'hb9);
  assign p2_add_85148_comb = p2_smul_84741_comb + p2_smul_84742_comb;
  assign p2_add_85149_comb = p2_smul_84743_comb + p2_smul_84744_comb;
  assign p2_smul_85150_comb = smul18b_18b_x_8b(p2_sign_ext_84525_comb[17:0], 8'h47);
  assign p2_smul_85151_comb = smul18b_18b_x_6b(p2_sign_ext_84526_comb[17:0], 6'h19);
  assign p2_smul_85152_comb = smul18b_18b_x_6b(p2_sign_ext_84527_comb[17:0], 6'h27);
  assign p2_smul_85153_comb = smul18b_18b_x_8b(p2_sign_ext_84528_comb[17:0], 8'hb9);
  assign p2_add_85154_comb = p2_smul_84753_comb + p2_smul_84754_comb;
  assign p2_smul_85164_comb = smul19b_19b_x_7b(p2_sign_ext_84533_comb[18:0], 7'h31);
  assign p2_smul_85165_comb = smul19b_19b_x_7b(p2_sign_ext_84477_comb[18:0], 7'h4f);
  assign p2_smul_85168_comb = smul19b_19b_x_7b(p2_sign_ext_84480_comb[18:0], 7'h4f);
  assign p2_smul_85169_comb = smul19b_19b_x_7b(p2_sign_ext_84534_comb[18:0], 7'h31);
  assign p2_smul_85172_comb = smul19b_19b_x_7b(p2_sign_ext_84535_comb[18:0], 7'h31);
  assign p2_smul_85173_comb = smul19b_19b_x_7b(p2_sign_ext_84485_comb[18:0], 7'h4f);
  assign p2_smul_85176_comb = smul19b_19b_x_7b(p2_sign_ext_84488_comb[18:0], 7'h4f);
  assign p2_smul_85177_comb = smul19b_19b_x_7b(p2_sign_ext_84536_comb[18:0], 7'h31);
  assign p2_smul_85180_comb = smul19b_19b_x_7b(p2_sign_ext_84537_comb[18:0], 7'h31);
  assign p2_smul_85181_comb = smul19b_19b_x_7b(p2_sign_ext_84493_comb[18:0], 7'h4f);
  assign p2_smul_85184_comb = smul19b_19b_x_7b(p2_sign_ext_84496_comb[18:0], 7'h4f);
  assign p2_smul_85185_comb = smul19b_19b_x_7b(p2_sign_ext_84538_comb[18:0], 7'h31);
  assign p2_smul_85196_comb = smul19b_19b_x_7b(p2_sign_ext_84541_comb[18:0], 7'h31);
  assign p2_smul_85197_comb = smul19b_19b_x_7b(p2_sign_ext_84509_comb[18:0], 7'h4f);
  assign p2_smul_85200_comb = smul19b_19b_x_7b(p2_sign_ext_84512_comb[18:0], 7'h4f);
  assign p2_smul_85201_comb = smul19b_19b_x_7b(p2_sign_ext_84542_comb[18:0], 7'h31);
  assign p2_smul_85204_comb = smul19b_19b_x_7b(p2_sign_ext_84543_comb[18:0], 7'h31);
  assign p2_smul_85205_comb = smul19b_19b_x_7b(p2_sign_ext_84517_comb[18:0], 7'h4f);
  assign p2_smul_85208_comb = smul19b_19b_x_7b(p2_sign_ext_84520_comb[18:0], 7'h4f);
  assign p2_smul_85209_comb = smul19b_19b_x_7b(p2_sign_ext_84544_comb[18:0], 7'h31);
  assign p2_smul_85212_comb = smul19b_19b_x_7b(p2_sign_ext_84545_comb[18:0], 7'h31);
  assign p2_smul_85213_comb = smul19b_19b_x_7b(p2_sign_ext_84525_comb[18:0], 7'h4f);
  assign p2_smul_85216_comb = smul19b_19b_x_7b(p2_sign_ext_84528_comb[18:0], 7'h4f);
  assign p2_smul_85217_comb = smul19b_19b_x_7b(p2_sign_ext_84546_comb[18:0], 7'h31);
  assign p2_smul_85419_comb = smul19b_19b_x_7b(p2_sign_ext_84585_comb[18:0], 7'h31);
  assign p2_smul_85421_comb = smul19b_19b_x_7b(p2_sign_ext_84477_comb[18:0], 7'h31);
  assign p2_smul_85424_comb = smul19b_19b_x_7b(p2_sign_ext_84480_comb[18:0], 7'h31);
  assign p2_smul_85426_comb = smul19b_19b_x_7b(p2_sign_ext_84590_comb[18:0], 7'h31);
  assign p2_smul_85427_comb = smul19b_19b_x_7b(p2_sign_ext_84591_comb[18:0], 7'h31);
  assign p2_smul_85429_comb = smul19b_19b_x_7b(p2_sign_ext_84485_comb[18:0], 7'h31);
  assign p2_smul_85432_comb = smul19b_19b_x_7b(p2_sign_ext_84488_comb[18:0], 7'h31);
  assign p2_smul_85434_comb = smul19b_19b_x_7b(p2_sign_ext_84596_comb[18:0], 7'h31);
  assign p2_smul_85435_comb = smul19b_19b_x_7b(p2_sign_ext_84597_comb[18:0], 7'h31);
  assign p2_smul_85437_comb = smul19b_19b_x_7b(p2_sign_ext_84493_comb[18:0], 7'h31);
  assign p2_smul_85440_comb = smul19b_19b_x_7b(p2_sign_ext_84496_comb[18:0], 7'h31);
  assign p2_smul_85442_comb = smul19b_19b_x_7b(p2_sign_ext_84602_comb[18:0], 7'h31);
  assign p2_smul_85451_comb = smul19b_19b_x_7b(p2_sign_ext_84609_comb[18:0], 7'h31);
  assign p2_smul_85453_comb = smul19b_19b_x_7b(p2_sign_ext_84509_comb[18:0], 7'h31);
  assign p2_smul_85456_comb = smul19b_19b_x_7b(p2_sign_ext_84512_comb[18:0], 7'h31);
  assign p2_smul_85458_comb = smul19b_19b_x_7b(p2_sign_ext_84614_comb[18:0], 7'h31);
  assign p2_smul_85459_comb = smul19b_19b_x_7b(p2_sign_ext_84615_comb[18:0], 7'h31);
  assign p2_smul_85461_comb = smul19b_19b_x_7b(p2_sign_ext_84517_comb[18:0], 7'h31);
  assign p2_smul_85464_comb = smul19b_19b_x_7b(p2_sign_ext_84520_comb[18:0], 7'h31);
  assign p2_smul_85466_comb = smul19b_19b_x_7b(p2_sign_ext_84620_comb[18:0], 7'h31);
  assign p2_smul_85467_comb = smul19b_19b_x_7b(p2_sign_ext_84621_comb[18:0], 7'h31);
  assign p2_smul_85469_comb = smul19b_19b_x_7b(p2_sign_ext_84525_comb[18:0], 7'h31);
  assign p2_smul_85472_comb = smul19b_19b_x_7b(p2_sign_ext_84528_comb[18:0], 7'h31);
  assign p2_smul_85474_comb = smul19b_19b_x_7b(p2_sign_ext_84626_comb[18:0], 7'h31);
  assign p2_smul_85481_comb = smul18b_18b_x_6b(p2_sign_ext_84585_comb[17:0], 6'h19);
  assign p2_smul_85482_comb = smul18b_18b_x_8b(p2_sign_ext_84533_comb[17:0], 8'hb9);
  assign p2_add_85483_comb = p2_smul_85027_comb + p2_smul_85028_comb;
  assign p2_add_85484_comb = p2_smul_85029_comb + p2_smul_85030_comb;
  assign p2_smul_85485_comb = smul18b_18b_x_8b(p2_sign_ext_84534_comb[17:0], 8'hb9);
  assign p2_smul_85486_comb = smul18b_18b_x_6b(p2_sign_ext_84590_comb[17:0], 6'h19);
  assign p2_smul_85487_comb = smul18b_18b_x_6b(p2_sign_ext_84591_comb[17:0], 6'h19);
  assign p2_smul_85488_comb = smul18b_18b_x_8b(p2_sign_ext_84535_comb[17:0], 8'hb9);
  assign p2_add_85489_comb = p2_smul_85039_comb + p2_smul_85040_comb;
  assign p2_add_85490_comb = p2_smul_85041_comb + p2_smul_85042_comb;
  assign p2_smul_85491_comb = smul18b_18b_x_8b(p2_sign_ext_84536_comb[17:0], 8'hb9);
  assign p2_smul_85492_comb = smul18b_18b_x_6b(p2_sign_ext_84596_comb[17:0], 6'h19);
  assign p2_smul_85493_comb = smul18b_18b_x_6b(p2_sign_ext_84597_comb[17:0], 6'h19);
  assign p2_smul_85494_comb = smul18b_18b_x_8b(p2_sign_ext_84537_comb[17:0], 8'hb9);
  assign p2_add_85495_comb = p2_smul_85051_comb + p2_smul_85052_comb;
  assign p2_add_85496_comb = p2_smul_85053_comb + p2_smul_85054_comb;
  assign p2_smul_85497_comb = smul18b_18b_x_8b(p2_sign_ext_84538_comb[17:0], 8'hb9);
  assign p2_smul_85498_comb = smul18b_18b_x_6b(p2_sign_ext_84602_comb[17:0], 6'h19);
  assign p2_smul_85505_comb = smul18b_18b_x_6b(p2_sign_ext_84609_comb[17:0], 6'h19);
  assign p2_smul_85506_comb = smul18b_18b_x_8b(p2_sign_ext_84541_comb[17:0], 8'hb9);
  assign p2_add_85507_comb = p2_smul_85075_comb + p2_smul_85076_comb;
  assign p2_add_85508_comb = p2_smul_85077_comb + p2_smul_85078_comb;
  assign p2_smul_85509_comb = smul18b_18b_x_8b(p2_sign_ext_84542_comb[17:0], 8'hb9);
  assign p2_smul_85510_comb = smul18b_18b_x_6b(p2_sign_ext_84614_comb[17:0], 6'h19);
  assign p2_smul_85511_comb = smul18b_18b_x_6b(p2_sign_ext_84615_comb[17:0], 6'h19);
  assign p2_smul_85512_comb = smul18b_18b_x_8b(p2_sign_ext_84543_comb[17:0], 8'hb9);
  assign p2_add_85513_comb = p2_smul_85087_comb + p2_smul_85088_comb;
  assign p2_add_85514_comb = p2_smul_85089_comb + p2_smul_85090_comb;
  assign p2_smul_85515_comb = smul18b_18b_x_8b(p2_sign_ext_84544_comb[17:0], 8'hb9);
  assign p2_smul_85516_comb = smul18b_18b_x_6b(p2_sign_ext_84620_comb[17:0], 6'h19);
  assign p2_smul_85517_comb = smul18b_18b_x_6b(p2_sign_ext_84621_comb[17:0], 6'h19);
  assign p2_smul_85518_comb = smul18b_18b_x_8b(p2_sign_ext_84545_comb[17:0], 8'hb9);
  assign p2_add_85519_comb = p2_smul_85099_comb + p2_smul_85100_comb;
  assign p2_add_85520_comb = p2_smul_85101_comb + p2_smul_85102_comb;
  assign p2_smul_85521_comb = smul18b_18b_x_8b(p2_sign_ext_84546_comb[17:0], 8'hb9);
  assign p2_smul_85522_comb = smul18b_18b_x_6b(p2_sign_ext_84626_comb[17:0], 6'h19);
  assign p2_add_85975_comb = p2_sign_ext_84585_comb[11:0] + p2_sign_ext_84533_comb[11:0];
  assign p2_add_85976_comb = p2_sign_ext_84477_comb[11:0] + p2_sign_ext_84478_comb[11:0];
  assign p2_add_85977_comb = p2_sign_ext_84479_comb[11:0] + p2_sign_ext_84480_comb[11:0];
  assign p2_add_85978_comb = p2_sign_ext_84534_comb[11:0] + p2_sign_ext_84590_comb[11:0];
  assign p2_add_85979_comb = p2_sign_ext_84591_comb[11:0] + p2_sign_ext_84535_comb[11:0];
  assign p2_add_85980_comb = p2_sign_ext_84485_comb[11:0] + p2_sign_ext_84486_comb[11:0];
  assign p2_add_85981_comb = p2_sign_ext_84487_comb[11:0] + p2_sign_ext_84488_comb[11:0];
  assign p2_add_85982_comb = p2_sign_ext_84536_comb[11:0] + p2_sign_ext_84596_comb[11:0];
  assign p2_add_85983_comb = p2_sign_ext_84597_comb[11:0] + p2_sign_ext_84537_comb[11:0];
  assign p2_add_85984_comb = p2_sign_ext_84493_comb[11:0] + p2_sign_ext_84494_comb[11:0];
  assign p2_add_85985_comb = p2_sign_ext_84495_comb[11:0] + p2_sign_ext_84496_comb[11:0];
  assign p2_add_85986_comb = p2_sign_ext_84538_comb[11:0] + p2_sign_ext_84602_comb[11:0];
  assign p2_add_85991_comb = p2_sign_ext_84609_comb[11:0] + p2_sign_ext_84541_comb[11:0];
  assign p2_add_85992_comb = p2_sign_ext_84509_comb[11:0] + p2_sign_ext_84510_comb[11:0];
  assign p2_add_85993_comb = p2_sign_ext_84511_comb[11:0] + p2_sign_ext_84512_comb[11:0];
  assign p2_add_85994_comb = p2_sign_ext_84542_comb[11:0] + p2_sign_ext_84614_comb[11:0];
  assign p2_add_85995_comb = p2_sign_ext_84615_comb[11:0] + p2_sign_ext_84543_comb[11:0];
  assign p2_add_85996_comb = p2_sign_ext_84517_comb[11:0] + p2_sign_ext_84518_comb[11:0];
  assign p2_add_85997_comb = p2_sign_ext_84519_comb[11:0] + p2_sign_ext_84520_comb[11:0];
  assign p2_add_85998_comb = p2_sign_ext_84544_comb[11:0] + p2_sign_ext_84620_comb[11:0];
  assign p2_add_85999_comb = p2_sign_ext_84621_comb[11:0] + p2_sign_ext_84545_comb[11:0];
  assign p2_add_86000_comb = p2_sign_ext_84525_comb[11:0] + p2_sign_ext_84526_comb[11:0];
  assign p2_add_86001_comb = p2_sign_ext_84527_comb[11:0] + p2_sign_ext_84528_comb[11:0];
  assign p2_add_86002_comb = p2_sign_ext_84546_comb[11:0] + p2_sign_ext_84626_comb[11:0];
  assign p2_add_86035_comb = p2_smul_85619_comb + p2_smul_85156_comb[18:1];
  assign p2_add_86037_comb = p2_smul_85157_comb[18:1] + p2_smul_85622_comb;
  assign p2_add_86039_comb = p2_smul_85623_comb + p2_smul_85160_comb[18:1];
  assign p2_add_86041_comb = p2_smul_85161_comb[18:1] + p2_smul_85626_comb;
  assign p2_concat_86099_comb = {p2_add_85683_comb, p2_smul_84819_comb[0]};
  assign p2_concat_86100_comb = {p2_add_85685_comb, p2_smul_84821_comb[0]};
  assign p2_concat_86101_comb = {p2_add_85687_comb, p2_smul_84826_comb[0]};
  assign p2_concat_86102_comb = {p2_add_85689_comb, p2_smul_84828_comb[0]};
  assign p2_concat_86163_comb = {p2_add_85811_comb, p2_smul_84901_comb[0]};
  assign p2_concat_86164_comb = {p2_add_85813_comb, p2_smul_84903_comb[0]};
  assign p2_concat_86165_comb = {p2_add_85815_comb, p2_smul_84904_comb[0]};
  assign p2_concat_86166_comb = {p2_add_85817_comb, p2_smul_84906_comb[0]};
  assign p2_add_86195_comb = p2_smul_85411_comb[18:1] + p2_smul_85876_comb;
  assign p2_add_86197_comb = p2_smul_85413_comb[18:1] + p2_smul_85878_comb;
  assign p2_add_86199_comb = p2_smul_85879_comb + p2_smul_85416_comb[18:1];
  assign p2_add_86201_comb = p2_smul_85881_comb + p2_smul_85418_comb[18:1];
  assign p2_add_86339_comb = {{5{p2_bit_slice_85603_comb[18]}}, p2_bit_slice_85603_comb} + {{6{p2_add_85604_comb[17]}}, p2_add_85604_comb};
  assign p2_add_86341_comb = {{6{p2_add_85605_comb[17]}}, p2_add_85605_comb} + {{5{p2_bit_slice_85606_comb[18]}}, p2_bit_slice_85606_comb};
  assign p2_concat_86371_comb = {p2_add_86067_comb, p2_smul_85188_comb[0]};
  assign p2_concat_86372_comb = {p2_add_86069_comb, p2_smul_85189_comb[0]};
  assign p2_concat_86373_comb = {p2_add_86071_comb, p2_smul_85192_comb[0]};
  assign p2_concat_86374_comb = {p2_add_86073_comb, p2_smul_85193_comb[0]};
  assign p2_sum__1460_comb = {{5{p2_concat_86115_comb[19]}}, p2_concat_86115_comb};
  assign p2_sum__1461_comb = {{5{p2_concat_86116_comb[19]}}, p2_concat_86116_comb};
  assign p2_sum__1462_comb = {{5{p2_concat_86117_comb[19]}}, p2_concat_86117_comb};
  assign p2_sum__1463_comb = {{5{p2_concat_86118_comb[19]}}, p2_concat_86118_comb};
  assign p2_sum__1540_comb = {{6{p2_add_86135_comb[18]}}, p2_add_86135_comb};
  assign p2_sum__1541_comb = {{6{p2_add_86136_comb[18]}}, p2_add_86136_comb};
  assign p2_sum__1542_comb = {{6{p2_add_86137_comb[18]}}, p2_add_86137_comb};
  assign p2_sum__1543_comb = {{6{p2_add_86138_comb[18]}}, p2_add_86138_comb};
  assign p2_sum__1512_comb = {{6{p2_add_86139_comb[18]}}, p2_add_86139_comb};
  assign p2_sum__1513_comb = {{6{p2_add_86140_comb[18]}}, p2_add_86140_comb};
  assign p2_sum__1514_comb = {{6{p2_add_86141_comb[18]}}, p2_add_86141_comb};
  assign p2_sum__1515_comb = {{6{p2_add_86142_comb[18]}}, p2_add_86142_comb};
  assign p2_sum__1484_comb = {{6{p2_add_86143_comb[18]}}, p2_add_86143_comb};
  assign p2_sum__1485_comb = {{6{p2_add_86144_comb[18]}}, p2_add_86144_comb};
  assign p2_sum__1486_comb = {{6{p2_add_86145_comb[18]}}, p2_add_86145_comb};
  assign p2_sum__1487_comb = {{6{p2_add_86146_comb[18]}}, p2_add_86146_comb};
  assign p2_sum__1428_comb = {{6{p2_add_86151_comb[18]}}, p2_add_86151_comb};
  assign p2_sum__1429_comb = {{6{p2_add_86152_comb[18]}}, p2_add_86152_comb};
  assign p2_sum__1430_comb = {{6{p2_add_86153_comb[18]}}, p2_add_86153_comb};
  assign p2_sum__1431_comb = {{6{p2_add_86154_comb[18]}}, p2_add_86154_comb};
  assign p2_sum__1400_comb = {{6{p2_add_86155_comb[18]}}, p2_add_86155_comb};
  assign p2_sum__1401_comb = {{6{p2_add_86156_comb[18]}}, p2_add_86156_comb};
  assign p2_sum__1402_comb = {{6{p2_add_86157_comb[18]}}, p2_add_86157_comb};
  assign p2_sum__1403_comb = {{6{p2_add_86158_comb[18]}}, p2_add_86158_comb};
  assign p2_sum__1372_comb = {{6{p2_add_86159_comb[18]}}, p2_add_86159_comb};
  assign p2_sum__1373_comb = {{6{p2_add_86160_comb[18]}}, p2_add_86160_comb};
  assign p2_sum__1374_comb = {{6{p2_add_86161_comb[18]}}, p2_add_86161_comb};
  assign p2_sum__1375_comb = {{6{p2_add_86162_comb[18]}}, p2_add_86162_comb};
  assign p2_sum__1452_comb = {{5{p2_concat_86179_comb[19]}}, p2_concat_86179_comb};
  assign p2_sum__1453_comb = {{5{p2_concat_86180_comb[19]}}, p2_concat_86180_comb};
  assign p2_sum__1454_comb = {{5{p2_concat_86181_comb[19]}}, p2_concat_86181_comb};
  assign p2_sum__1455_comb = {{5{p2_concat_86182_comb[19]}}, p2_concat_86182_comb};
  assign p2_concat_86451_comb = {p2_add_86227_comb, p2_smul_85443_comb[0]};
  assign p2_concat_86452_comb = {p2_add_86229_comb, p2_smul_85445_comb[0]};
  assign p2_concat_86453_comb = {p2_add_86231_comb, p2_smul_85448_comb[0]};
  assign p2_concat_86454_comb = {p2_add_86233_comb, p2_smul_85450_comb[0]};
  assign p2_add_86483_comb = {{6{p2_add_85955_comb[17]}}, p2_add_85955_comb} + {{5{p2_bit_slice_85956_comb[18]}}, p2_bit_slice_85956_comb};
  assign p2_add_86485_comb = {{5{p2_bit_slice_85957_comb[18]}}, p2_bit_slice_85957_comb} + {{6{p2_add_85958_comb[17]}}, p2_add_85958_comb};
  assign p2_add_86499_comb = {{12{p2_add_85971_comb[11]}}, p2_add_85971_comb} + {{12{p2_add_85972_comb[11]}}, p2_add_85972_comb};
  assign p2_add_86500_comb = {{12{p2_add_85973_comb[11]}}, p2_add_85973_comb} + {{12{p2_add_85974_comb[11]}}, p2_add_85974_comb};
  assign p2_add_86507_comb = {{12{p2_add_85987_comb[11]}}, p2_add_85987_comb} + {{12{p2_add_85988_comb[11]}}, p2_add_85988_comb};
  assign p2_add_86508_comb = {{12{p2_add_85989_comb[11]}}, p2_add_85989_comb} + {{12{p2_add_85990_comb[11]}}, p2_add_85990_comb};
  assign p2_sum__1240_comb = p2_sum__1568_comb + p2_sum__1569_comb;
  assign p2_sum__1241_comb = p2_sum__1570_comb + p2_sum__1571_comb;
  assign p2_sum__1184_comb = p2_sum__1456_comb + p2_sum__1457_comb;
  assign p2_sum__1185_comb = p2_sum__1458_comb + p2_sum__1459_comb;
  assign p2_smul_85228_comb = smul19b_19b_x_6b(p2_sign_ext_84533_comb[18:0], 6'h27);
  assign p2_smul_85230_comb = smul19b_19b_x_8b(p2_sign_ext_84478_comb[18:0], 8'hb9);
  assign p2_smul_85231_comb = smul19b_19b_x_8b(p2_sign_ext_84479_comb[18:0], 8'h47);
  assign p2_smul_85233_comb = smul19b_19b_x_6b(p2_sign_ext_84534_comb[18:0], 6'h19);
  assign p2_smul_85236_comb = smul19b_19b_x_6b(p2_sign_ext_84535_comb[18:0], 6'h27);
  assign p2_smul_85238_comb = smul19b_19b_x_8b(p2_sign_ext_84486_comb[18:0], 8'hb9);
  assign p2_smul_85239_comb = smul19b_19b_x_8b(p2_sign_ext_84487_comb[18:0], 8'h47);
  assign p2_smul_85241_comb = smul19b_19b_x_6b(p2_sign_ext_84536_comb[18:0], 6'h19);
  assign p2_smul_85244_comb = smul19b_19b_x_6b(p2_sign_ext_84537_comb[18:0], 6'h27);
  assign p2_smul_85246_comb = smul19b_19b_x_8b(p2_sign_ext_84494_comb[18:0], 8'hb9);
  assign p2_smul_85247_comb = smul19b_19b_x_8b(p2_sign_ext_84495_comb[18:0], 8'h47);
  assign p2_smul_85249_comb = smul19b_19b_x_6b(p2_sign_ext_84538_comb[18:0], 6'h19);
  assign p2_smul_85260_comb = smul19b_19b_x_6b(p2_sign_ext_84541_comb[18:0], 6'h27);
  assign p2_smul_85262_comb = smul19b_19b_x_8b(p2_sign_ext_84510_comb[18:0], 8'hb9);
  assign p2_smul_85263_comb = smul19b_19b_x_8b(p2_sign_ext_84511_comb[18:0], 8'h47);
  assign p2_smul_85265_comb = smul19b_19b_x_6b(p2_sign_ext_84542_comb[18:0], 6'h19);
  assign p2_smul_85268_comb = smul19b_19b_x_6b(p2_sign_ext_84543_comb[18:0], 6'h27);
  assign p2_smul_85270_comb = smul19b_19b_x_8b(p2_sign_ext_84518_comb[18:0], 8'hb9);
  assign p2_smul_85271_comb = smul19b_19b_x_8b(p2_sign_ext_84519_comb[18:0], 8'h47);
  assign p2_smul_85273_comb = smul19b_19b_x_6b(p2_sign_ext_84544_comb[18:0], 6'h19);
  assign p2_smul_85276_comb = smul19b_19b_x_6b(p2_sign_ext_84545_comb[18:0], 6'h27);
  assign p2_smul_85278_comb = smul19b_19b_x_8b(p2_sign_ext_84526_comb[18:0], 8'hb9);
  assign p2_smul_85279_comb = smul19b_19b_x_8b(p2_sign_ext_84527_comb[18:0], 8'h47);
  assign p2_smul_85281_comb = smul19b_19b_x_6b(p2_sign_ext_84546_comb[18:0], 6'h19);
  assign p2_smul_85355_comb = smul19b_19b_x_8b(p2_sign_ext_84585_comb[18:0], 8'h47);
  assign p2_smul_85357_comb = smul19b_19b_x_6b(p2_sign_ext_84477_comb[18:0], 6'h27);
  assign p2_smul_85360_comb = smul19b_19b_x_6b(p2_sign_ext_84480_comb[18:0], 6'h27);
  assign p2_smul_85362_comb = smul19b_19b_x_8b(p2_sign_ext_84590_comb[18:0], 8'h47);
  assign p2_smul_85363_comb = smul19b_19b_x_8b(p2_sign_ext_84591_comb[18:0], 8'h47);
  assign p2_smul_85365_comb = smul19b_19b_x_6b(p2_sign_ext_84485_comb[18:0], 6'h27);
  assign p2_smul_85368_comb = smul19b_19b_x_6b(p2_sign_ext_84488_comb[18:0], 6'h27);
  assign p2_smul_85370_comb = smul19b_19b_x_8b(p2_sign_ext_84596_comb[18:0], 8'h47);
  assign p2_smul_85371_comb = smul19b_19b_x_8b(p2_sign_ext_84597_comb[18:0], 8'h47);
  assign p2_smul_85373_comb = smul19b_19b_x_6b(p2_sign_ext_84493_comb[18:0], 6'h27);
  assign p2_smul_85376_comb = smul19b_19b_x_6b(p2_sign_ext_84496_comb[18:0], 6'h27);
  assign p2_smul_85378_comb = smul19b_19b_x_8b(p2_sign_ext_84602_comb[18:0], 8'h47);
  assign p2_smul_85387_comb = smul19b_19b_x_8b(p2_sign_ext_84609_comb[18:0], 8'h47);
  assign p2_smul_85389_comb = smul19b_19b_x_6b(p2_sign_ext_84509_comb[18:0], 6'h27);
  assign p2_smul_85392_comb = smul19b_19b_x_6b(p2_sign_ext_84512_comb[18:0], 6'h27);
  assign p2_smul_85394_comb = smul19b_19b_x_8b(p2_sign_ext_84614_comb[18:0], 8'h47);
  assign p2_smul_85395_comb = smul19b_19b_x_8b(p2_sign_ext_84615_comb[18:0], 8'h47);
  assign p2_smul_85397_comb = smul19b_19b_x_6b(p2_sign_ext_84517_comb[18:0], 6'h27);
  assign p2_smul_85400_comb = smul19b_19b_x_6b(p2_sign_ext_84520_comb[18:0], 6'h27);
  assign p2_smul_85402_comb = smul19b_19b_x_8b(p2_sign_ext_84620_comb[18:0], 8'h47);
  assign p2_smul_85403_comb = smul19b_19b_x_8b(p2_sign_ext_84621_comb[18:0], 8'h47);
  assign p2_smul_85405_comb = smul19b_19b_x_6b(p2_sign_ext_84525_comb[18:0], 6'h27);
  assign p2_smul_85408_comb = smul19b_19b_x_6b(p2_sign_ext_84528_comb[18:0], 6'h27);
  assign p2_smul_85410_comb = smul19b_19b_x_8b(p2_sign_ext_84626_comb[18:0], 8'h47);
  assign p2_bit_slice_85591_comb = p2_add_85113_comb[19:1];
  assign p2_add_85592_comb = p2_smul_85114_comb + p2_smul_85115_comb;
  assign p2_add_85593_comb = p2_smul_85116_comb + p2_smul_85117_comb;
  assign p2_bit_slice_85594_comb = p2_add_85118_comb[19:1];
  assign p2_bit_slice_85595_comb = p2_add_85119_comb[19:1];
  assign p2_add_85596_comb = p2_smul_85120_comb + p2_smul_85121_comb;
  assign p2_add_85597_comb = p2_smul_85122_comb + p2_smul_85123_comb;
  assign p2_bit_slice_85598_comb = p2_add_85124_comb[19:1];
  assign p2_bit_slice_85599_comb = p2_add_85125_comb[19:1];
  assign p2_add_85600_comb = p2_smul_85126_comb + p2_smul_85127_comb;
  assign p2_add_85601_comb = p2_smul_85128_comb + p2_smul_85129_comb;
  assign p2_bit_slice_85602_comb = p2_add_85130_comb[19:1];
  assign p2_bit_slice_85607_comb = p2_add_85137_comb[19:1];
  assign p2_add_85608_comb = p2_smul_85138_comb + p2_smul_85139_comb;
  assign p2_add_85609_comb = p2_smul_85140_comb + p2_smul_85141_comb;
  assign p2_bit_slice_85610_comb = p2_add_85142_comb[19:1];
  assign p2_bit_slice_85611_comb = p2_add_85143_comb[19:1];
  assign p2_add_85612_comb = p2_smul_85144_comb + p2_smul_85145_comb;
  assign p2_add_85613_comb = p2_smul_85146_comb + p2_smul_85147_comb;
  assign p2_bit_slice_85614_comb = p2_add_85148_comb[19:1];
  assign p2_bit_slice_85615_comb = p2_add_85149_comb[19:1];
  assign p2_add_85616_comb = p2_smul_85150_comb + p2_smul_85151_comb;
  assign p2_add_85617_comb = p2_smul_85152_comb + p2_smul_85153_comb;
  assign p2_bit_slice_85618_comb = p2_add_85154_comb[19:1];
  assign p2_smul_85627_comb = smul18b_18b_x_7b(p2_sign_ext_84585_comb[17:0], 7'h3b);
  assign p2_smul_85630_comb = smul18b_18b_x_7b(p2_sign_ext_84478_comb[17:0], 7'h45);
  assign p2_smul_85631_comb = smul18b_18b_x_7b(p2_sign_ext_84479_comb[17:0], 7'h45);
  assign p2_smul_85634_comb = smul18b_18b_x_7b(p2_sign_ext_84590_comb[17:0], 7'h3b);
  assign p2_smul_85635_comb = smul18b_18b_x_7b(p2_sign_ext_84591_comb[17:0], 7'h3b);
  assign p2_smul_85638_comb = smul18b_18b_x_7b(p2_sign_ext_84486_comb[17:0], 7'h45);
  assign p2_smul_85639_comb = smul18b_18b_x_7b(p2_sign_ext_84487_comb[17:0], 7'h45);
  assign p2_smul_85642_comb = smul18b_18b_x_7b(p2_sign_ext_84596_comb[17:0], 7'h3b);
  assign p2_smul_85643_comb = smul18b_18b_x_7b(p2_sign_ext_84597_comb[17:0], 7'h3b);
  assign p2_smul_85646_comb = smul18b_18b_x_7b(p2_sign_ext_84494_comb[17:0], 7'h45);
  assign p2_smul_85647_comb = smul18b_18b_x_7b(p2_sign_ext_84495_comb[17:0], 7'h45);
  assign p2_smul_85650_comb = smul18b_18b_x_7b(p2_sign_ext_84602_comb[17:0], 7'h3b);
  assign p2_smul_85659_comb = smul18b_18b_x_7b(p2_sign_ext_84609_comb[17:0], 7'h3b);
  assign p2_smul_85662_comb = smul18b_18b_x_7b(p2_sign_ext_84510_comb[17:0], 7'h45);
  assign p2_smul_85663_comb = smul18b_18b_x_7b(p2_sign_ext_84511_comb[17:0], 7'h45);
  assign p2_smul_85666_comb = smul18b_18b_x_7b(p2_sign_ext_84614_comb[17:0], 7'h3b);
  assign p2_smul_85667_comb = smul18b_18b_x_7b(p2_sign_ext_84615_comb[17:0], 7'h3b);
  assign p2_smul_85670_comb = smul18b_18b_x_7b(p2_sign_ext_84518_comb[17:0], 7'h45);
  assign p2_smul_85671_comb = smul18b_18b_x_7b(p2_sign_ext_84519_comb[17:0], 7'h45);
  assign p2_smul_85674_comb = smul18b_18b_x_7b(p2_sign_ext_84620_comb[17:0], 7'h3b);
  assign p2_smul_85675_comb = smul18b_18b_x_7b(p2_sign_ext_84621_comb[17:0], 7'h3b);
  assign p2_smul_85678_comb = smul18b_18b_x_7b(p2_sign_ext_84526_comb[17:0], 7'h45);
  assign p2_smul_85679_comb = smul18b_18b_x_7b(p2_sign_ext_84527_comb[17:0], 7'h45);
  assign p2_smul_85682_comb = smul18b_18b_x_7b(p2_sign_ext_84626_comb[17:0], 7'h3b);
  assign p2_smul_85884_comb = smul18b_18b_x_7b(p2_sign_ext_84533_comb[17:0], 7'h45);
  assign p2_smul_85886_comb = smul18b_18b_x_7b(p2_sign_ext_84478_comb[17:0], 7'h3b);
  assign p2_smul_85887_comb = smul18b_18b_x_7b(p2_sign_ext_84479_comb[17:0], 7'h3b);
  assign p2_smul_85889_comb = smul18b_18b_x_7b(p2_sign_ext_84534_comb[17:0], 7'h45);
  assign p2_smul_85892_comb = smul18b_18b_x_7b(p2_sign_ext_84535_comb[17:0], 7'h45);
  assign p2_smul_85894_comb = smul18b_18b_x_7b(p2_sign_ext_84486_comb[17:0], 7'h3b);
  assign p2_smul_85895_comb = smul18b_18b_x_7b(p2_sign_ext_84487_comb[17:0], 7'h3b);
  assign p2_smul_85897_comb = smul18b_18b_x_7b(p2_sign_ext_84536_comb[17:0], 7'h45);
  assign p2_smul_85900_comb = smul18b_18b_x_7b(p2_sign_ext_84537_comb[17:0], 7'h45);
  assign p2_smul_85902_comb = smul18b_18b_x_7b(p2_sign_ext_84494_comb[17:0], 7'h3b);
  assign p2_smul_85903_comb = smul18b_18b_x_7b(p2_sign_ext_84495_comb[17:0], 7'h3b);
  assign p2_smul_85905_comb = smul18b_18b_x_7b(p2_sign_ext_84538_comb[17:0], 7'h45);
  assign p2_smul_85916_comb = smul18b_18b_x_7b(p2_sign_ext_84541_comb[17:0], 7'h45);
  assign p2_smul_85918_comb = smul18b_18b_x_7b(p2_sign_ext_84510_comb[17:0], 7'h3b);
  assign p2_smul_85919_comb = smul18b_18b_x_7b(p2_sign_ext_84511_comb[17:0], 7'h3b);
  assign p2_smul_85921_comb = smul18b_18b_x_7b(p2_sign_ext_84542_comb[17:0], 7'h45);
  assign p2_smul_85924_comb = smul18b_18b_x_7b(p2_sign_ext_84543_comb[17:0], 7'h45);
  assign p2_smul_85926_comb = smul18b_18b_x_7b(p2_sign_ext_84518_comb[17:0], 7'h3b);
  assign p2_smul_85927_comb = smul18b_18b_x_7b(p2_sign_ext_84519_comb[17:0], 7'h3b);
  assign p2_smul_85929_comb = smul18b_18b_x_7b(p2_sign_ext_84544_comb[17:0], 7'h45);
  assign p2_smul_85932_comb = smul18b_18b_x_7b(p2_sign_ext_84545_comb[17:0], 7'h45);
  assign p2_smul_85934_comb = smul18b_18b_x_7b(p2_sign_ext_84526_comb[17:0], 7'h3b);
  assign p2_smul_85935_comb = smul18b_18b_x_7b(p2_sign_ext_84527_comb[17:0], 7'h3b);
  assign p2_smul_85937_comb = smul18b_18b_x_7b(p2_sign_ext_84546_comb[17:0], 7'h45);
  assign p2_add_85943_comb = p2_smul_85481_comb + p2_smul_85482_comb;
  assign p2_bit_slice_85944_comb = p2_add_85483_comb[19:1];
  assign p2_bit_slice_85945_comb = p2_add_85484_comb[19:1];
  assign p2_add_85946_comb = p2_smul_85485_comb + p2_smul_85486_comb;
  assign p2_add_85947_comb = p2_smul_85487_comb + p2_smul_85488_comb;
  assign p2_bit_slice_85948_comb = p2_add_85489_comb[19:1];
  assign p2_bit_slice_85949_comb = p2_add_85490_comb[19:1];
  assign p2_add_85950_comb = p2_smul_85491_comb + p2_smul_85492_comb;
  assign p2_add_85951_comb = p2_smul_85493_comb + p2_smul_85494_comb;
  assign p2_bit_slice_85952_comb = p2_add_85495_comb[19:1];
  assign p2_bit_slice_85953_comb = p2_add_85496_comb[19:1];
  assign p2_add_85954_comb = p2_smul_85497_comb + p2_smul_85498_comb;
  assign p2_add_85959_comb = p2_smul_85505_comb + p2_smul_85506_comb;
  assign p2_bit_slice_85960_comb = p2_add_85507_comb[19:1];
  assign p2_bit_slice_85961_comb = p2_add_85508_comb[19:1];
  assign p2_add_85962_comb = p2_smul_85509_comb + p2_smul_85510_comb;
  assign p2_add_85963_comb = p2_smul_85511_comb + p2_smul_85512_comb;
  assign p2_bit_slice_85964_comb = p2_add_85513_comb[19:1];
  assign p2_bit_slice_85965_comb = p2_add_85514_comb[19:1];
  assign p2_add_85966_comb = p2_smul_85515_comb + p2_smul_85516_comb;
  assign p2_add_85967_comb = p2_smul_85517_comb + p2_smul_85518_comb;
  assign p2_bit_slice_85968_comb = p2_add_85519_comb[19:1];
  assign p2_bit_slice_85969_comb = p2_add_85520_comb[19:1];
  assign p2_add_85970_comb = p2_smul_85521_comb + p2_smul_85522_comb;
  assign p2_add_86323_comb = {{5{p2_bit_slice_85587_comb[18]}}, p2_bit_slice_85587_comb} + {{6{p2_add_85588_comb[17]}}, p2_add_85588_comb};
  assign p2_add_86325_comb = {{6{p2_add_85589_comb[17]}}, p2_add_85589_comb} + {{5{p2_bit_slice_85590_comb[18]}}, p2_bit_slice_85590_comb};
  assign p2_concat_86355_comb = {p2_add_86035_comb, p2_smul_85156_comb[0]};
  assign p2_concat_86356_comb = {p2_add_86037_comb, p2_smul_85157_comb[0]};
  assign p2_concat_86357_comb = {p2_add_86039_comb, p2_smul_85160_comb[0]};
  assign p2_concat_86358_comb = {p2_add_86041_comb, p2_smul_85161_comb[0]};
  assign p2_sum__1572_comb = {{5{p2_concat_86099_comb[19]}}, p2_concat_86099_comb};
  assign p2_sum__1573_comb = {{5{p2_concat_86100_comb[19]}}, p2_concat_86100_comb};
  assign p2_sum__1574_comb = {{5{p2_concat_86101_comb[19]}}, p2_concat_86101_comb};
  assign p2_sum__1575_comb = {{5{p2_concat_86102_comb[19]}}, p2_concat_86102_comb};
  assign p2_sum__1564_comb = {{5{p2_concat_86163_comb[19]}}, p2_concat_86163_comb};
  assign p2_sum__1565_comb = {{5{p2_concat_86164_comb[19]}}, p2_concat_86164_comb};
  assign p2_sum__1566_comb = {{5{p2_concat_86165_comb[19]}}, p2_concat_86165_comb};
  assign p2_sum__1567_comb = {{5{p2_concat_86166_comb[19]}}, p2_concat_86166_comb};
  assign p2_concat_86435_comb = {p2_add_86195_comb, p2_smul_85411_comb[0]};
  assign p2_concat_86436_comb = {p2_add_86197_comb, p2_smul_85413_comb[0]};
  assign p2_concat_86437_comb = {p2_add_86199_comb, p2_smul_85416_comb[0]};
  assign p2_concat_86438_comb = {p2_add_86201_comb, p2_smul_85418_comb[0]};
  assign p2_add_86467_comb = {{6{p2_add_85939_comb[17]}}, p2_add_85939_comb} + {{5{p2_bit_slice_85940_comb[18]}}, p2_bit_slice_85940_comb};
  assign p2_add_86469_comb = {{5{p2_bit_slice_85941_comb[18]}}, p2_bit_slice_85941_comb} + {{6{p2_add_85942_comb[17]}}, p2_add_85942_comb};
  assign p2_sum__1190_comb = {p2_add_86339_comb, p2_add_85131_comb[0]};
  assign p2_sum__1191_comb = {p2_add_86341_comb, p2_add_85136_comb[0]};
  assign p2_sum__1186_comb = p2_sum__1460_comb + p2_sum__1461_comb;
  assign p2_sum__1187_comb = p2_sum__1462_comb + p2_sum__1463_comb;
  assign p2_sum__1226_comb = p2_sum__1540_comb + p2_sum__1541_comb;
  assign p2_sum__1227_comb = p2_sum__1542_comb + p2_sum__1543_comb;
  assign p2_sum__1212_comb = p2_sum__1512_comb + p2_sum__1513_comb;
  assign p2_sum__1213_comb = p2_sum__1514_comb + p2_sum__1515_comb;
  assign p2_sum__1198_comb = p2_sum__1484_comb + p2_sum__1485_comb;
  assign p2_sum__1199_comb = p2_sum__1486_comb + p2_sum__1487_comb;
  assign p2_sum__1170_comb = p2_sum__1428_comb + p2_sum__1429_comb;
  assign p2_sum__1171_comb = p2_sum__1430_comb + p2_sum__1431_comb;
  assign p2_sum__1156_comb = p2_sum__1400_comb + p2_sum__1401_comb;
  assign p2_sum__1157_comb = p2_sum__1402_comb + p2_sum__1403_comb;
  assign p2_sum__1142_comb = p2_sum__1372_comb + p2_sum__1373_comb;
  assign p2_sum__1143_comb = p2_sum__1374_comb + p2_sum__1375_comb;
  assign p2_sum__1182_comb = p2_sum__1452_comb + p2_sum__1453_comb;
  assign p2_sum__1183_comb = p2_sum__1454_comb + p2_sum__1455_comb;
  assign p2_sum__1178_comb = {p2_add_86483_comb, p2_add_85501_comb[0]};
  assign p2_sum__1179_comb = {p2_add_86485_comb, p2_add_85502_comb[0]};
  assign p2_add_86563_comb = p2_add_86499_comb + p2_add_86500_comb;
  assign p2_add_86568_comb = p2_add_86507_comb + p2_add_86508_comb;
  assign p2_sum__1076_comb = p2_sum__1240_comb + p2_sum__1241_comb;
  assign p2_sum__1048_comb = p2_sum__1184_comb + p2_sum__1185_comb;
  assign p2_add_85691_comb = p2_smul_84829_comb[19:1] + p2_smul_85228_comb;
  assign p2_add_85693_comb = p2_smul_84831_comb[19:1] + p2_smul_85230_comb;
  assign p2_add_85695_comb = p2_smul_85231_comb + p2_smul_84836_comb[19:1];
  assign p2_add_85697_comb = p2_smul_85233_comb + p2_smul_84838_comb[19:1];
  assign p2_add_85699_comb = p2_smul_84839_comb[19:1] + p2_smul_85236_comb;
  assign p2_add_85701_comb = p2_smul_84841_comb[19:1] + p2_smul_85238_comb;
  assign p2_add_85703_comb = p2_smul_85239_comb + p2_smul_84846_comb[19:1];
  assign p2_add_85705_comb = p2_smul_85241_comb + p2_smul_84848_comb[19:1];
  assign p2_add_85707_comb = p2_smul_84849_comb[19:1] + p2_smul_85244_comb;
  assign p2_add_85709_comb = p2_smul_84851_comb[19:1] + p2_smul_85246_comb;
  assign p2_add_85711_comb = p2_smul_85247_comb + p2_smul_84856_comb[19:1];
  assign p2_add_85713_comb = p2_smul_85249_comb + p2_smul_84858_comb[19:1];
  assign p2_add_85723_comb = p2_smul_84869_comb[19:1] + p2_smul_85260_comb;
  assign p2_add_85725_comb = p2_smul_84871_comb[19:1] + p2_smul_85262_comb;
  assign p2_add_85727_comb = p2_smul_85263_comb + p2_smul_84876_comb[19:1];
  assign p2_add_85729_comb = p2_smul_85265_comb + p2_smul_84878_comb[19:1];
  assign p2_add_85731_comb = p2_smul_84879_comb[19:1] + p2_smul_85268_comb;
  assign p2_add_85733_comb = p2_smul_84881_comb[19:1] + p2_smul_85270_comb;
  assign p2_add_85735_comb = p2_smul_85271_comb + p2_smul_84886_comb[19:1];
  assign p2_add_85737_comb = p2_smul_85273_comb + p2_smul_84888_comb[19:1];
  assign p2_add_85739_comb = p2_smul_84889_comb[19:1] + p2_smul_85276_comb;
  assign p2_add_85741_comb = p2_smul_84891_comb[19:1] + p2_smul_85278_comb;
  assign p2_add_85743_comb = p2_smul_85279_comb + p2_smul_84896_comb[19:1];
  assign p2_add_85745_comb = p2_smul_85281_comb + p2_smul_84898_comb[19:1];
  assign p2_add_85819_comb = p2_smul_85355_comb + p2_smul_84911_comb[19:1];
  assign p2_add_85821_comb = p2_smul_85357_comb + p2_smul_84913_comb[19:1];
  assign p2_add_85823_comb = p2_smul_84914_comb[19:1] + p2_smul_85360_comb;
  assign p2_add_85825_comb = p2_smul_84916_comb[19:1] + p2_smul_85362_comb;
  assign p2_add_85827_comb = p2_smul_85363_comb + p2_smul_84921_comb[19:1];
  assign p2_add_85829_comb = p2_smul_85365_comb + p2_smul_84923_comb[19:1];
  assign p2_add_85831_comb = p2_smul_84924_comb[19:1] + p2_smul_85368_comb;
  assign p2_add_85833_comb = p2_smul_84926_comb[19:1] + p2_smul_85370_comb;
  assign p2_add_85835_comb = p2_smul_85371_comb + p2_smul_84931_comb[19:1];
  assign p2_add_85837_comb = p2_smul_85373_comb + p2_smul_84933_comb[19:1];
  assign p2_add_85839_comb = p2_smul_84934_comb[19:1] + p2_smul_85376_comb;
  assign p2_add_85841_comb = p2_smul_84936_comb[19:1] + p2_smul_85378_comb;
  assign p2_add_85851_comb = p2_smul_85387_comb + p2_smul_84951_comb[19:1];
  assign p2_add_85853_comb = p2_smul_85389_comb + p2_smul_84953_comb[19:1];
  assign p2_add_85855_comb = p2_smul_84954_comb[19:1] + p2_smul_85392_comb;
  assign p2_add_85857_comb = p2_smul_84956_comb[19:1] + p2_smul_85394_comb;
  assign p2_add_85859_comb = p2_smul_85395_comb + p2_smul_84961_comb[19:1];
  assign p2_add_85861_comb = p2_smul_85397_comb + p2_smul_84963_comb[19:1];
  assign p2_add_85863_comb = p2_smul_84964_comb[19:1] + p2_smul_85400_comb;
  assign p2_add_85865_comb = p2_smul_84966_comb[19:1] + p2_smul_85402_comb;
  assign p2_add_85867_comb = p2_smul_85403_comb + p2_smul_84971_comb[19:1];
  assign p2_add_85869_comb = p2_smul_85405_comb + p2_smul_84973_comb[19:1];
  assign p2_add_85871_comb = p2_smul_84974_comb[19:1] + p2_smul_85408_comb;
  assign p2_add_85873_comb = p2_smul_84976_comb[19:1] + p2_smul_85410_comb;
  assign p2_add_86043_comb = p2_smul_85627_comb + p2_smul_85164_comb[18:1];
  assign p2_add_86045_comb = p2_smul_85165_comb[18:1] + p2_smul_85630_comb;
  assign p2_add_86047_comb = p2_smul_85631_comb + p2_smul_85168_comb[18:1];
  assign p2_add_86049_comb = p2_smul_85169_comb[18:1] + p2_smul_85634_comb;
  assign p2_add_86051_comb = p2_smul_85635_comb + p2_smul_85172_comb[18:1];
  assign p2_add_86053_comb = p2_smul_85173_comb[18:1] + p2_smul_85638_comb;
  assign p2_add_86055_comb = p2_smul_85639_comb + p2_smul_85176_comb[18:1];
  assign p2_add_86057_comb = p2_smul_85177_comb[18:1] + p2_smul_85642_comb;
  assign p2_add_86059_comb = p2_smul_85643_comb + p2_smul_85180_comb[18:1];
  assign p2_add_86061_comb = p2_smul_85181_comb[18:1] + p2_smul_85646_comb;
  assign p2_add_86063_comb = p2_smul_85647_comb + p2_smul_85184_comb[18:1];
  assign p2_add_86065_comb = p2_smul_85185_comb[18:1] + p2_smul_85650_comb;
  assign p2_add_86075_comb = p2_smul_85659_comb + p2_smul_85196_comb[18:1];
  assign p2_add_86077_comb = p2_smul_85197_comb[18:1] + p2_smul_85662_comb;
  assign p2_add_86079_comb = p2_smul_85663_comb + p2_smul_85200_comb[18:1];
  assign p2_add_86081_comb = p2_smul_85201_comb[18:1] + p2_smul_85666_comb;
  assign p2_add_86083_comb = p2_smul_85667_comb + p2_smul_85204_comb[18:1];
  assign p2_add_86085_comb = p2_smul_85205_comb[18:1] + p2_smul_85670_comb;
  assign p2_add_86087_comb = p2_smul_85671_comb + p2_smul_85208_comb[18:1];
  assign p2_add_86089_comb = p2_smul_85209_comb[18:1] + p2_smul_85674_comb;
  assign p2_add_86091_comb = p2_smul_85675_comb + p2_smul_85212_comb[18:1];
  assign p2_add_86093_comb = p2_smul_85213_comb[18:1] + p2_smul_85678_comb;
  assign p2_add_86095_comb = p2_smul_85679_comb + p2_smul_85216_comb[18:1];
  assign p2_add_86097_comb = p2_smul_85217_comb[18:1] + p2_smul_85682_comb;
  assign p2_add_86203_comb = p2_smul_85419_comb[18:1] + p2_smul_85884_comb;
  assign p2_add_86205_comb = p2_smul_85421_comb[18:1] + p2_smul_85886_comb;
  assign p2_add_86207_comb = p2_smul_85887_comb + p2_smul_85424_comb[18:1];
  assign p2_add_86209_comb = p2_smul_85889_comb + p2_smul_85426_comb[18:1];
  assign p2_add_86211_comb = p2_smul_85427_comb[18:1] + p2_smul_85892_comb;
  assign p2_add_86213_comb = p2_smul_85429_comb[18:1] + p2_smul_85894_comb;
  assign p2_add_86215_comb = p2_smul_85895_comb + p2_smul_85432_comb[18:1];
  assign p2_add_86217_comb = p2_smul_85897_comb + p2_smul_85434_comb[18:1];
  assign p2_add_86219_comb = p2_smul_85435_comb[18:1] + p2_smul_85900_comb;
  assign p2_add_86221_comb = p2_smul_85437_comb[18:1] + p2_smul_85902_comb;
  assign p2_add_86223_comb = p2_smul_85903_comb + p2_smul_85440_comb[18:1];
  assign p2_add_86225_comb = p2_smul_85905_comb + p2_smul_85442_comb[18:1];
  assign p2_add_86235_comb = p2_smul_85451_comb[18:1] + p2_smul_85916_comb;
  assign p2_add_86237_comb = p2_smul_85453_comb[18:1] + p2_smul_85918_comb;
  assign p2_add_86239_comb = p2_smul_85919_comb + p2_smul_85456_comb[18:1];
  assign p2_add_86241_comb = p2_smul_85921_comb + p2_smul_85458_comb[18:1];
  assign p2_add_86243_comb = p2_smul_85459_comb[18:1] + p2_smul_85924_comb;
  assign p2_add_86245_comb = p2_smul_85461_comb[18:1] + p2_smul_85926_comb;
  assign p2_add_86247_comb = p2_smul_85927_comb + p2_smul_85464_comb[18:1];
  assign p2_add_86249_comb = p2_smul_85929_comb + p2_smul_85466_comb[18:1];
  assign p2_add_86251_comb = p2_smul_85467_comb[18:1] + p2_smul_85932_comb;
  assign p2_add_86253_comb = p2_smul_85469_comb[18:1] + p2_smul_85934_comb;
  assign p2_add_86255_comb = p2_smul_85935_comb + p2_smul_85472_comb[18:1];
  assign p2_add_86257_comb = p2_smul_85937_comb + p2_smul_85474_comb[18:1];
  assign p2_add_86501_comb = {{12{p2_add_85975_comb[11]}}, p2_add_85975_comb} + {{12{p2_add_85976_comb[11]}}, p2_add_85976_comb};
  assign p2_add_86502_comb = {{12{p2_add_85977_comb[11]}}, p2_add_85977_comb} + {{12{p2_add_85978_comb[11]}}, p2_add_85978_comb};
  assign p2_add_86503_comb = {{12{p2_add_85979_comb[11]}}, p2_add_85979_comb} + {{12{p2_add_85980_comb[11]}}, p2_add_85980_comb};
  assign p2_add_86504_comb = {{12{p2_add_85981_comb[11]}}, p2_add_85981_comb} + {{12{p2_add_85982_comb[11]}}, p2_add_85982_comb};
  assign p2_add_86505_comb = {{12{p2_add_85983_comb[11]}}, p2_add_85983_comb} + {{12{p2_add_85984_comb[11]}}, p2_add_85984_comb};
  assign p2_add_86506_comb = {{12{p2_add_85985_comb[11]}}, p2_add_85985_comb} + {{12{p2_add_85986_comb[11]}}, p2_add_85986_comb};
  assign p2_add_86509_comb = {{12{p2_add_85991_comb[11]}}, p2_add_85991_comb} + {{12{p2_add_85992_comb[11]}}, p2_add_85992_comb};
  assign p2_add_86510_comb = {{12{p2_add_85993_comb[11]}}, p2_add_85993_comb} + {{12{p2_add_85994_comb[11]}}, p2_add_85994_comb};
  assign p2_add_86511_comb = {{12{p2_add_85995_comb[11]}}, p2_add_85995_comb} + {{12{p2_add_85996_comb[11]}}, p2_add_85996_comb};
  assign p2_add_86512_comb = {{12{p2_add_85997_comb[11]}}, p2_add_85997_comb} + {{12{p2_add_85998_comb[11]}}, p2_add_85998_comb};
  assign p2_add_86513_comb = {{12{p2_add_85999_comb[11]}}, p2_add_85999_comb} + {{12{p2_add_86000_comb[11]}}, p2_add_86000_comb};
  assign p2_add_86514_comb = {{12{p2_add_86001_comb[11]}}, p2_add_86001_comb} + {{12{p2_add_86002_comb[11]}}, p2_add_86002_comb};
  assign p2_sum__1246_comb = {p2_add_86323_comb, p2_add_85107_comb[0]};
  assign p2_sum__1247_comb = {p2_add_86325_comb, p2_add_85112_comb[0]};
  assign p2_sum__1242_comb = p2_sum__1572_comb + p2_sum__1573_comb;
  assign p2_sum__1243_comb = p2_sum__1574_comb + p2_sum__1575_comb;
  assign p2_sum__1238_comb = p2_sum__1564_comb + p2_sum__1565_comb;
  assign p2_sum__1239_comb = p2_sum__1566_comb + p2_sum__1567_comb;
  assign p2_sum__1234_comb = {p2_add_86467_comb, p2_add_85477_comb[0]};
  assign p2_sum__1235_comb = {p2_add_86469_comb, p2_add_85478_comb[0]};
  assign p2_sum__1051_comb = p2_sum__1190_comb + p2_sum__1191_comb;
  assign p2_add_86578_comb = {{5{p2_concat_86371_comb[18]}}, p2_concat_86371_comb} + {{5{p2_concat_86372_comb[18]}}, p2_concat_86372_comb};
  assign p2_add_86579_comb = {{5{p2_concat_86373_comb[18]}}, p2_concat_86373_comb} + {{5{p2_concat_86374_comb[18]}}, p2_concat_86374_comb};
  assign p2_sum__1049_comb = p2_sum__1186_comb + p2_sum__1187_comb;
  assign p2_sum__1069_comb = p2_sum__1226_comb + p2_sum__1227_comb;
  assign p2_sum__1062_comb = p2_sum__1212_comb + p2_sum__1213_comb;
  assign p2_sum__1055_comb = p2_sum__1198_comb + p2_sum__1199_comb;
  assign p2_sum__1041_comb = p2_sum__1170_comb + p2_sum__1171_comb;
  assign p2_sum__1034_comb = p2_sum__1156_comb + p2_sum__1157_comb;
  assign p2_sum__1027_comb = p2_sum__1142_comb + p2_sum__1143_comb;
  assign p2_sum__1047_comb = p2_sum__1182_comb + p2_sum__1183_comb;
  assign p2_add_86604_comb = {{5{p2_concat_86451_comb[18]}}, p2_concat_86451_comb} + {{5{p2_concat_86452_comb[18]}}, p2_concat_86452_comb};
  assign p2_add_86605_comb = {{5{p2_concat_86453_comb[18]}}, p2_concat_86453_comb} + {{5{p2_concat_86454_comb[18]}}, p2_concat_86454_comb};
  assign p2_sum__1045_comb = p2_sum__1178_comb + p2_sum__1179_comb;
  assign p2_umul_29016_NarrowedMult__comb = umul24b_24b_x_7b(p2_add_86563_comb, 7'h5b);
  assign p2_umul_29024_NarrowedMult__comb = umul24b_24b_x_7b(p2_add_86568_comb, 7'h5b);
  assign p2_add_86614_comb = p2_sum__1076_comb + 25'h000_0001;
  assign p2_add_86618_comb = p2_sum__1048_comb + 25'h000_0001;
  assign p2_concat_86103_comb = {p2_add_85691_comb, p2_smul_84829_comb[0]};
  assign p2_concat_86104_comb = {p2_add_85693_comb, p2_smul_84831_comb[0]};
  assign p2_concat_86105_comb = {p2_add_85695_comb, p2_smul_84836_comb[0]};
  assign p2_concat_86106_comb = {p2_add_85697_comb, p2_smul_84838_comb[0]};
  assign p2_concat_86107_comb = {p2_add_85699_comb, p2_smul_84839_comb[0]};
  assign p2_concat_86108_comb = {p2_add_85701_comb, p2_smul_84841_comb[0]};
  assign p2_concat_86109_comb = {p2_add_85703_comb, p2_smul_84846_comb[0]};
  assign p2_concat_86110_comb = {p2_add_85705_comb, p2_smul_84848_comb[0]};
  assign p2_concat_86111_comb = {p2_add_85707_comb, p2_smul_84849_comb[0]};
  assign p2_concat_86112_comb = {p2_add_85709_comb, p2_smul_84851_comb[0]};
  assign p2_concat_86113_comb = {p2_add_85711_comb, p2_smul_84856_comb[0]};
  assign p2_concat_86114_comb = {p2_add_85713_comb, p2_smul_84858_comb[0]};
  assign p2_concat_86119_comb = {p2_add_85723_comb, p2_smul_84869_comb[0]};
  assign p2_concat_86120_comb = {p2_add_85725_comb, p2_smul_84871_comb[0]};
  assign p2_concat_86121_comb = {p2_add_85727_comb, p2_smul_84876_comb[0]};
  assign p2_concat_86122_comb = {p2_add_85729_comb, p2_smul_84878_comb[0]};
  assign p2_concat_86123_comb = {p2_add_85731_comb, p2_smul_84879_comb[0]};
  assign p2_concat_86124_comb = {p2_add_85733_comb, p2_smul_84881_comb[0]};
  assign p2_concat_86125_comb = {p2_add_85735_comb, p2_smul_84886_comb[0]};
  assign p2_concat_86126_comb = {p2_add_85737_comb, p2_smul_84888_comb[0]};
  assign p2_concat_86127_comb = {p2_add_85739_comb, p2_smul_84889_comb[0]};
  assign p2_concat_86128_comb = {p2_add_85741_comb, p2_smul_84891_comb[0]};
  assign p2_concat_86129_comb = {p2_add_85743_comb, p2_smul_84896_comb[0]};
  assign p2_concat_86130_comb = {p2_add_85745_comb, p2_smul_84898_comb[0]};
  assign p2_concat_86167_comb = {p2_add_85819_comb, p2_smul_84911_comb[0]};
  assign p2_concat_86168_comb = {p2_add_85821_comb, p2_smul_84913_comb[0]};
  assign p2_concat_86169_comb = {p2_add_85823_comb, p2_smul_84914_comb[0]};
  assign p2_concat_86170_comb = {p2_add_85825_comb, p2_smul_84916_comb[0]};
  assign p2_concat_86171_comb = {p2_add_85827_comb, p2_smul_84921_comb[0]};
  assign p2_concat_86172_comb = {p2_add_85829_comb, p2_smul_84923_comb[0]};
  assign p2_concat_86173_comb = {p2_add_85831_comb, p2_smul_84924_comb[0]};
  assign p2_concat_86174_comb = {p2_add_85833_comb, p2_smul_84926_comb[0]};
  assign p2_concat_86175_comb = {p2_add_85835_comb, p2_smul_84931_comb[0]};
  assign p2_concat_86176_comb = {p2_add_85837_comb, p2_smul_84933_comb[0]};
  assign p2_concat_86177_comb = {p2_add_85839_comb, p2_smul_84934_comb[0]};
  assign p2_concat_86178_comb = {p2_add_85841_comb, p2_smul_84936_comb[0]};
  assign p2_concat_86183_comb = {p2_add_85851_comb, p2_smul_84951_comb[0]};
  assign p2_concat_86184_comb = {p2_add_85853_comb, p2_smul_84953_comb[0]};
  assign p2_concat_86185_comb = {p2_add_85855_comb, p2_smul_84954_comb[0]};
  assign p2_concat_86186_comb = {p2_add_85857_comb, p2_smul_84956_comb[0]};
  assign p2_concat_86187_comb = {p2_add_85859_comb, p2_smul_84961_comb[0]};
  assign p2_concat_86188_comb = {p2_add_85861_comb, p2_smul_84963_comb[0]};
  assign p2_concat_86189_comb = {p2_add_85863_comb, p2_smul_84964_comb[0]};
  assign p2_concat_86190_comb = {p2_add_85865_comb, p2_smul_84966_comb[0]};
  assign p2_concat_86191_comb = {p2_add_85867_comb, p2_smul_84971_comb[0]};
  assign p2_concat_86192_comb = {p2_add_85869_comb, p2_smul_84973_comb[0]};
  assign p2_concat_86193_comb = {p2_add_85871_comb, p2_smul_84974_comb[0]};
  assign p2_concat_86194_comb = {p2_add_85873_comb, p2_smul_84976_comb[0]};
  assign p2_add_86327_comb = {{5{p2_bit_slice_85591_comb[18]}}, p2_bit_slice_85591_comb} + {{6{p2_add_85592_comb[17]}}, p2_add_85592_comb};
  assign p2_bit_slice_86328_comb = p2_add_85113_comb[0];
  assign p2_add_86329_comb = {{6{p2_add_85593_comb[17]}}, p2_add_85593_comb} + {{5{p2_bit_slice_85594_comb[18]}}, p2_bit_slice_85594_comb};
  assign p2_bit_slice_86330_comb = p2_add_85118_comb[0];
  assign p2_add_86331_comb = {{5{p2_bit_slice_85595_comb[18]}}, p2_bit_slice_85595_comb} + {{6{p2_add_85596_comb[17]}}, p2_add_85596_comb};
  assign p2_bit_slice_86332_comb = p2_add_85119_comb[0];
  assign p2_add_86333_comb = {{6{p2_add_85597_comb[17]}}, p2_add_85597_comb} + {{5{p2_bit_slice_85598_comb[18]}}, p2_bit_slice_85598_comb};
  assign p2_bit_slice_86334_comb = p2_add_85124_comb[0];
  assign p2_add_86335_comb = {{5{p2_bit_slice_85599_comb[18]}}, p2_bit_slice_85599_comb} + {{6{p2_add_85600_comb[17]}}, p2_add_85600_comb};
  assign p2_bit_slice_86336_comb = p2_add_85125_comb[0];
  assign p2_add_86337_comb = {{6{p2_add_85601_comb[17]}}, p2_add_85601_comb} + {{5{p2_bit_slice_85602_comb[18]}}, p2_bit_slice_85602_comb};
  assign p2_bit_slice_86338_comb = p2_add_85130_comb[0];
  assign p2_add_86343_comb = {{5{p2_bit_slice_85607_comb[18]}}, p2_bit_slice_85607_comb} + {{6{p2_add_85608_comb[17]}}, p2_add_85608_comb};
  assign p2_bit_slice_86344_comb = p2_add_85137_comb[0];
  assign p2_add_86345_comb = {{6{p2_add_85609_comb[17]}}, p2_add_85609_comb} + {{5{p2_bit_slice_85610_comb[18]}}, p2_bit_slice_85610_comb};
  assign p2_bit_slice_86346_comb = p2_add_85142_comb[0];
  assign p2_add_86347_comb = {{5{p2_bit_slice_85611_comb[18]}}, p2_bit_slice_85611_comb} + {{6{p2_add_85612_comb[17]}}, p2_add_85612_comb};
  assign p2_bit_slice_86348_comb = p2_add_85143_comb[0];
  assign p2_add_86349_comb = {{6{p2_add_85613_comb[17]}}, p2_add_85613_comb} + {{5{p2_bit_slice_85614_comb[18]}}, p2_bit_slice_85614_comb};
  assign p2_bit_slice_86350_comb = p2_add_85148_comb[0];
  assign p2_add_86351_comb = {{5{p2_bit_slice_85615_comb[18]}}, p2_bit_slice_85615_comb} + {{6{p2_add_85616_comb[17]}}, p2_add_85616_comb};
  assign p2_bit_slice_86352_comb = p2_add_85149_comb[0];
  assign p2_add_86353_comb = {{6{p2_add_85617_comb[17]}}, p2_add_85617_comb} + {{5{p2_bit_slice_85618_comb[18]}}, p2_bit_slice_85618_comb};
  assign p2_bit_slice_86354_comb = p2_add_85154_comb[0];
  assign p2_concat_86359_comb = {p2_add_86043_comb, p2_smul_85164_comb[0]};
  assign p2_concat_86360_comb = {p2_add_86045_comb, p2_smul_85165_comb[0]};
  assign p2_concat_86361_comb = {p2_add_86047_comb, p2_smul_85168_comb[0]};
  assign p2_concat_86362_comb = {p2_add_86049_comb, p2_smul_85169_comb[0]};
  assign p2_concat_86363_comb = {p2_add_86051_comb, p2_smul_85172_comb[0]};
  assign p2_concat_86364_comb = {p2_add_86053_comb, p2_smul_85173_comb[0]};
  assign p2_concat_86365_comb = {p2_add_86055_comb, p2_smul_85176_comb[0]};
  assign p2_concat_86366_comb = {p2_add_86057_comb, p2_smul_85177_comb[0]};
  assign p2_concat_86367_comb = {p2_add_86059_comb, p2_smul_85180_comb[0]};
  assign p2_concat_86368_comb = {p2_add_86061_comb, p2_smul_85181_comb[0]};
  assign p2_concat_86369_comb = {p2_add_86063_comb, p2_smul_85184_comb[0]};
  assign p2_concat_86370_comb = {p2_add_86065_comb, p2_smul_85185_comb[0]};
  assign p2_concat_86375_comb = {p2_add_86075_comb, p2_smul_85196_comb[0]};
  assign p2_concat_86376_comb = {p2_add_86077_comb, p2_smul_85197_comb[0]};
  assign p2_concat_86377_comb = {p2_add_86079_comb, p2_smul_85200_comb[0]};
  assign p2_concat_86378_comb = {p2_add_86081_comb, p2_smul_85201_comb[0]};
  assign p2_concat_86379_comb = {p2_add_86083_comb, p2_smul_85204_comb[0]};
  assign p2_concat_86380_comb = {p2_add_86085_comb, p2_smul_85205_comb[0]};
  assign p2_concat_86381_comb = {p2_add_86087_comb, p2_smul_85208_comb[0]};
  assign p2_concat_86382_comb = {p2_add_86089_comb, p2_smul_85209_comb[0]};
  assign p2_concat_86383_comb = {p2_add_86091_comb, p2_smul_85212_comb[0]};
  assign p2_concat_86384_comb = {p2_add_86093_comb, p2_smul_85213_comb[0]};
  assign p2_concat_86385_comb = {p2_add_86095_comb, p2_smul_85216_comb[0]};
  assign p2_concat_86386_comb = {p2_add_86097_comb, p2_smul_85217_comb[0]};
  assign p2_concat_86439_comb = {p2_add_86203_comb, p2_smul_85419_comb[0]};
  assign p2_concat_86440_comb = {p2_add_86205_comb, p2_smul_85421_comb[0]};
  assign p2_concat_86441_comb = {p2_add_86207_comb, p2_smul_85424_comb[0]};
  assign p2_concat_86442_comb = {p2_add_86209_comb, p2_smul_85426_comb[0]};
  assign p2_concat_86443_comb = {p2_add_86211_comb, p2_smul_85427_comb[0]};
  assign p2_concat_86444_comb = {p2_add_86213_comb, p2_smul_85429_comb[0]};
  assign p2_concat_86445_comb = {p2_add_86215_comb, p2_smul_85432_comb[0]};
  assign p2_concat_86446_comb = {p2_add_86217_comb, p2_smul_85434_comb[0]};
  assign p2_concat_86447_comb = {p2_add_86219_comb, p2_smul_85435_comb[0]};
  assign p2_concat_86448_comb = {p2_add_86221_comb, p2_smul_85437_comb[0]};
  assign p2_concat_86449_comb = {p2_add_86223_comb, p2_smul_85440_comb[0]};
  assign p2_concat_86450_comb = {p2_add_86225_comb, p2_smul_85442_comb[0]};
  assign p2_concat_86455_comb = {p2_add_86235_comb, p2_smul_85451_comb[0]};
  assign p2_concat_86456_comb = {p2_add_86237_comb, p2_smul_85453_comb[0]};
  assign p2_concat_86457_comb = {p2_add_86239_comb, p2_smul_85456_comb[0]};
  assign p2_concat_86458_comb = {p2_add_86241_comb, p2_smul_85458_comb[0]};
  assign p2_concat_86459_comb = {p2_add_86243_comb, p2_smul_85459_comb[0]};
  assign p2_concat_86460_comb = {p2_add_86245_comb, p2_smul_85461_comb[0]};
  assign p2_concat_86461_comb = {p2_add_86247_comb, p2_smul_85464_comb[0]};
  assign p2_concat_86462_comb = {p2_add_86249_comb, p2_smul_85466_comb[0]};
  assign p2_concat_86463_comb = {p2_add_86251_comb, p2_smul_85467_comb[0]};
  assign p2_concat_86464_comb = {p2_add_86253_comb, p2_smul_85469_comb[0]};
  assign p2_concat_86465_comb = {p2_add_86255_comb, p2_smul_85472_comb[0]};
  assign p2_concat_86466_comb = {p2_add_86257_comb, p2_smul_85474_comb[0]};
  assign p2_add_86471_comb = {{6{p2_add_85943_comb[17]}}, p2_add_85943_comb} + {{5{p2_bit_slice_85944_comb[18]}}, p2_bit_slice_85944_comb};
  assign p2_bit_slice_86472_comb = p2_add_85483_comb[0];
  assign p2_add_86473_comb = {{5{p2_bit_slice_85945_comb[18]}}, p2_bit_slice_85945_comb} + {{6{p2_add_85946_comb[17]}}, p2_add_85946_comb};
  assign p2_bit_slice_86474_comb = p2_add_85484_comb[0];
  assign p2_add_86475_comb = {{6{p2_add_85947_comb[17]}}, p2_add_85947_comb} + {{5{p2_bit_slice_85948_comb[18]}}, p2_bit_slice_85948_comb};
  assign p2_bit_slice_86476_comb = p2_add_85489_comb[0];
  assign p2_add_86477_comb = {{5{p2_bit_slice_85949_comb[18]}}, p2_bit_slice_85949_comb} + {{6{p2_add_85950_comb[17]}}, p2_add_85950_comb};
  assign p2_bit_slice_86478_comb = p2_add_85490_comb[0];
  assign p2_add_86479_comb = {{6{p2_add_85951_comb[17]}}, p2_add_85951_comb} + {{5{p2_bit_slice_85952_comb[18]}}, p2_bit_slice_85952_comb};
  assign p2_bit_slice_86480_comb = p2_add_85495_comb[0];
  assign p2_add_86481_comb = {{5{p2_bit_slice_85953_comb[18]}}, p2_bit_slice_85953_comb} + {{6{p2_add_85954_comb[17]}}, p2_add_85954_comb};
  assign p2_bit_slice_86482_comb = p2_add_85496_comb[0];
  assign p2_add_86487_comb = {{6{p2_add_85959_comb[17]}}, p2_add_85959_comb} + {{5{p2_bit_slice_85960_comb[18]}}, p2_bit_slice_85960_comb};
  assign p2_bit_slice_86488_comb = p2_add_85507_comb[0];
  assign p2_add_86489_comb = {{5{p2_bit_slice_85961_comb[18]}}, p2_bit_slice_85961_comb} + {{6{p2_add_85962_comb[17]}}, p2_add_85962_comb};
  assign p2_bit_slice_86490_comb = p2_add_85508_comb[0];
  assign p2_add_86491_comb = {{6{p2_add_85963_comb[17]}}, p2_add_85963_comb} + {{5{p2_bit_slice_85964_comb[18]}}, p2_bit_slice_85964_comb};
  assign p2_bit_slice_86492_comb = p2_add_85513_comb[0];
  assign p2_add_86493_comb = {{5{p2_bit_slice_85965_comb[18]}}, p2_bit_slice_85965_comb} + {{6{p2_add_85966_comb[17]}}, p2_add_85966_comb};
  assign p2_bit_slice_86494_comb = p2_add_85514_comb[0];
  assign p2_add_86495_comb = {{6{p2_add_85967_comb[17]}}, p2_add_85967_comb} + {{5{p2_bit_slice_85968_comb[18]}}, p2_bit_slice_85968_comb};
  assign p2_bit_slice_86496_comb = p2_add_85519_comb[0];
  assign p2_add_86497_comb = {{5{p2_bit_slice_85969_comb[18]}}, p2_bit_slice_85969_comb} + {{6{p2_add_85970_comb[17]}}, p2_add_85970_comb};
  assign p2_bit_slice_86498_comb = p2_add_85520_comb[0];
  assign p2_add_86565_comb = p2_add_86501_comb + p2_add_86502_comb;
  assign p2_add_86566_comb = p2_add_86503_comb + p2_add_86504_comb;
  assign p2_add_86567_comb = p2_add_86505_comb + p2_add_86506_comb;
  assign p2_add_86570_comb = p2_add_86509_comb + p2_add_86510_comb;
  assign p2_add_86571_comb = p2_add_86511_comb + p2_add_86512_comb;
  assign p2_add_86572_comb = p2_add_86513_comb + p2_add_86514_comb;
  assign p2_sum__1079_comb = p2_sum__1246_comb + p2_sum__1247_comb;
  assign p2_add_86576_comb = {{5{p2_concat_86355_comb[18]}}, p2_concat_86355_comb} + {{5{p2_concat_86356_comb[18]}}, p2_concat_86356_comb};
  assign p2_add_86577_comb = {{5{p2_concat_86357_comb[18]}}, p2_concat_86357_comb} + {{5{p2_concat_86358_comb[18]}}, p2_concat_86358_comb};
  assign p2_sum__1077_comb = p2_sum__1242_comb + p2_sum__1243_comb;
  assign p2_sum__1075_comb = p2_sum__1238_comb + p2_sum__1239_comb;
  assign p2_add_86602_comb = {{5{p2_concat_86435_comb[18]}}, p2_concat_86435_comb} + {{5{p2_concat_86436_comb[18]}}, p2_concat_86436_comb};
  assign p2_add_86603_comb = {{5{p2_concat_86437_comb[18]}}, p2_concat_86437_comb} + {{5{p2_concat_86438_comb[18]}}, p2_concat_86438_comb};
  assign p2_sum__1073_comb = p2_sum__1234_comb + p2_sum__1235_comb;
  assign p2_add_86611_comb = p2_sum__1051_comb + 25'h000_0001;
  assign p2_add_86612_comb = p2_add_86578_comb + p2_add_86579_comb;
  assign p2_add_86613_comb = p2_sum__1049_comb + 25'h000_0001;
  assign p2_add_86615_comb = p2_sum__1069_comb + 25'h000_0001;
  assign p2_add_86616_comb = p2_sum__1062_comb + 25'h000_0001;
  assign p2_add_86617_comb = p2_sum__1055_comb + 25'h000_0001;
  assign p2_add_86619_comb = p2_sum__1041_comb + 25'h000_0001;
  assign p2_add_86620_comb = p2_sum__1034_comb + 25'h000_0001;
  assign p2_add_86621_comb = p2_sum__1027_comb + 25'h000_0001;
  assign p2_add_86622_comb = p2_sum__1047_comb + 25'h000_0001;
  assign p2_add_86623_comb = p2_add_86604_comb + p2_add_86605_comb;
  assign p2_add_86624_comb = p2_sum__1045_comb + 25'h000_0001;
  assign p2_bit_slice_86625_comb = p2_umul_29016_NarrowedMult__comb[23:7];
  assign p2_bit_slice_86626_comb = p2_umul_29024_NarrowedMult__comb[23:7];
  assign p2_bit_slice_86627_comb = p2_add_86614_comb[24:8];
  assign p2_bit_slice_86628_comb = p2_add_86618_comb[24:8];

  // Registers for pipe stage 2:
  reg [19:0] p2_concat_86103;
  reg [19:0] p2_concat_86104;
  reg [19:0] p2_concat_86105;
  reg [19:0] p2_concat_86106;
  reg [19:0] p2_concat_86107;
  reg [19:0] p2_concat_86108;
  reg [19:0] p2_concat_86109;
  reg [19:0] p2_concat_86110;
  reg [19:0] p2_concat_86111;
  reg [19:0] p2_concat_86112;
  reg [19:0] p2_concat_86113;
  reg [19:0] p2_concat_86114;
  reg [19:0] p2_concat_86119;
  reg [19:0] p2_concat_86120;
  reg [19:0] p2_concat_86121;
  reg [19:0] p2_concat_86122;
  reg [19:0] p2_concat_86123;
  reg [19:0] p2_concat_86124;
  reg [19:0] p2_concat_86125;
  reg [19:0] p2_concat_86126;
  reg [19:0] p2_concat_86127;
  reg [19:0] p2_concat_86128;
  reg [19:0] p2_concat_86129;
  reg [19:0] p2_concat_86130;
  reg [19:0] p2_concat_86167;
  reg [19:0] p2_concat_86168;
  reg [19:0] p2_concat_86169;
  reg [19:0] p2_concat_86170;
  reg [19:0] p2_concat_86171;
  reg [19:0] p2_concat_86172;
  reg [19:0] p2_concat_86173;
  reg [19:0] p2_concat_86174;
  reg [19:0] p2_concat_86175;
  reg [19:0] p2_concat_86176;
  reg [19:0] p2_concat_86177;
  reg [19:0] p2_concat_86178;
  reg [19:0] p2_concat_86183;
  reg [19:0] p2_concat_86184;
  reg [19:0] p2_concat_86185;
  reg [19:0] p2_concat_86186;
  reg [19:0] p2_concat_86187;
  reg [19:0] p2_concat_86188;
  reg [19:0] p2_concat_86189;
  reg [19:0] p2_concat_86190;
  reg [19:0] p2_concat_86191;
  reg [19:0] p2_concat_86192;
  reg [19:0] p2_concat_86193;
  reg [19:0] p2_concat_86194;
  reg [23:0] p2_add_86327;
  reg p2_bit_slice_86328;
  reg [23:0] p2_add_86329;
  reg p2_bit_slice_86330;
  reg [23:0] p2_add_86331;
  reg p2_bit_slice_86332;
  reg [23:0] p2_add_86333;
  reg p2_bit_slice_86334;
  reg [23:0] p2_add_86335;
  reg p2_bit_slice_86336;
  reg [23:0] p2_add_86337;
  reg p2_bit_slice_86338;
  reg [23:0] p2_add_86343;
  reg p2_bit_slice_86344;
  reg [23:0] p2_add_86345;
  reg p2_bit_slice_86346;
  reg [23:0] p2_add_86347;
  reg p2_bit_slice_86348;
  reg [23:0] p2_add_86349;
  reg p2_bit_slice_86350;
  reg [23:0] p2_add_86351;
  reg p2_bit_slice_86352;
  reg [23:0] p2_add_86353;
  reg p2_bit_slice_86354;
  reg [18:0] p2_concat_86359;
  reg [18:0] p2_concat_86360;
  reg [18:0] p2_concat_86361;
  reg [18:0] p2_concat_86362;
  reg [18:0] p2_concat_86363;
  reg [18:0] p2_concat_86364;
  reg [18:0] p2_concat_86365;
  reg [18:0] p2_concat_86366;
  reg [18:0] p2_concat_86367;
  reg [18:0] p2_concat_86368;
  reg [18:0] p2_concat_86369;
  reg [18:0] p2_concat_86370;
  reg [18:0] p2_concat_86375;
  reg [18:0] p2_concat_86376;
  reg [18:0] p2_concat_86377;
  reg [18:0] p2_concat_86378;
  reg [18:0] p2_concat_86379;
  reg [18:0] p2_concat_86380;
  reg [18:0] p2_concat_86381;
  reg [18:0] p2_concat_86382;
  reg [18:0] p2_concat_86383;
  reg [18:0] p2_concat_86384;
  reg [18:0] p2_concat_86385;
  reg [18:0] p2_concat_86386;
  reg [18:0] p2_concat_86439;
  reg [18:0] p2_concat_86440;
  reg [18:0] p2_concat_86441;
  reg [18:0] p2_concat_86442;
  reg [18:0] p2_concat_86443;
  reg [18:0] p2_concat_86444;
  reg [18:0] p2_concat_86445;
  reg [18:0] p2_concat_86446;
  reg [18:0] p2_concat_86447;
  reg [18:0] p2_concat_86448;
  reg [18:0] p2_concat_86449;
  reg [18:0] p2_concat_86450;
  reg [18:0] p2_concat_86455;
  reg [18:0] p2_concat_86456;
  reg [18:0] p2_concat_86457;
  reg [18:0] p2_concat_86458;
  reg [18:0] p2_concat_86459;
  reg [18:0] p2_concat_86460;
  reg [18:0] p2_concat_86461;
  reg [18:0] p2_concat_86462;
  reg [18:0] p2_concat_86463;
  reg [18:0] p2_concat_86464;
  reg [18:0] p2_concat_86465;
  reg [18:0] p2_concat_86466;
  reg [23:0] p2_add_86471;
  reg p2_bit_slice_86472;
  reg [23:0] p2_add_86473;
  reg p2_bit_slice_86474;
  reg [23:0] p2_add_86475;
  reg p2_bit_slice_86476;
  reg [23:0] p2_add_86477;
  reg p2_bit_slice_86478;
  reg [23:0] p2_add_86479;
  reg p2_bit_slice_86480;
  reg [23:0] p2_add_86481;
  reg p2_bit_slice_86482;
  reg [23:0] p2_add_86487;
  reg p2_bit_slice_86488;
  reg [23:0] p2_add_86489;
  reg p2_bit_slice_86490;
  reg [23:0] p2_add_86491;
  reg p2_bit_slice_86492;
  reg [23:0] p2_add_86493;
  reg p2_bit_slice_86494;
  reg [23:0] p2_add_86495;
  reg p2_bit_slice_86496;
  reg [23:0] p2_add_86497;
  reg p2_bit_slice_86498;
  reg [23:0] p2_add_86565;
  reg [23:0] p2_add_86566;
  reg [23:0] p2_add_86567;
  reg [23:0] p2_add_86570;
  reg [23:0] p2_add_86571;
  reg [23:0] p2_add_86572;
  reg [24:0] p2_sum__1079;
  reg [23:0] p2_add_86576;
  reg [23:0] p2_add_86577;
  reg [24:0] p2_sum__1077;
  reg [24:0] p2_sum__1075;
  reg [23:0] p2_add_86602;
  reg [23:0] p2_add_86603;
  reg [24:0] p2_sum__1073;
  reg [24:0] p2_add_86611;
  reg [23:0] p2_add_86612;
  reg [24:0] p2_add_86613;
  reg [24:0] p2_add_86615;
  reg [24:0] p2_add_86616;
  reg [24:0] p2_add_86617;
  reg [24:0] p2_add_86619;
  reg [24:0] p2_add_86620;
  reg [24:0] p2_add_86621;
  reg [24:0] p2_add_86622;
  reg [23:0] p2_add_86623;
  reg [24:0] p2_add_86624;
  reg [16:0] p2_bit_slice_86625;
  reg [16:0] p2_bit_slice_86626;
  reg [16:0] p2_bit_slice_86627;
  reg [16:0] p2_bit_slice_86628;
  always @ (posedge clk) begin
    p2_concat_86103 <= p2_concat_86103_comb;
    p2_concat_86104 <= p2_concat_86104_comb;
    p2_concat_86105 <= p2_concat_86105_comb;
    p2_concat_86106 <= p2_concat_86106_comb;
    p2_concat_86107 <= p2_concat_86107_comb;
    p2_concat_86108 <= p2_concat_86108_comb;
    p2_concat_86109 <= p2_concat_86109_comb;
    p2_concat_86110 <= p2_concat_86110_comb;
    p2_concat_86111 <= p2_concat_86111_comb;
    p2_concat_86112 <= p2_concat_86112_comb;
    p2_concat_86113 <= p2_concat_86113_comb;
    p2_concat_86114 <= p2_concat_86114_comb;
    p2_concat_86119 <= p2_concat_86119_comb;
    p2_concat_86120 <= p2_concat_86120_comb;
    p2_concat_86121 <= p2_concat_86121_comb;
    p2_concat_86122 <= p2_concat_86122_comb;
    p2_concat_86123 <= p2_concat_86123_comb;
    p2_concat_86124 <= p2_concat_86124_comb;
    p2_concat_86125 <= p2_concat_86125_comb;
    p2_concat_86126 <= p2_concat_86126_comb;
    p2_concat_86127 <= p2_concat_86127_comb;
    p2_concat_86128 <= p2_concat_86128_comb;
    p2_concat_86129 <= p2_concat_86129_comb;
    p2_concat_86130 <= p2_concat_86130_comb;
    p2_concat_86167 <= p2_concat_86167_comb;
    p2_concat_86168 <= p2_concat_86168_comb;
    p2_concat_86169 <= p2_concat_86169_comb;
    p2_concat_86170 <= p2_concat_86170_comb;
    p2_concat_86171 <= p2_concat_86171_comb;
    p2_concat_86172 <= p2_concat_86172_comb;
    p2_concat_86173 <= p2_concat_86173_comb;
    p2_concat_86174 <= p2_concat_86174_comb;
    p2_concat_86175 <= p2_concat_86175_comb;
    p2_concat_86176 <= p2_concat_86176_comb;
    p2_concat_86177 <= p2_concat_86177_comb;
    p2_concat_86178 <= p2_concat_86178_comb;
    p2_concat_86183 <= p2_concat_86183_comb;
    p2_concat_86184 <= p2_concat_86184_comb;
    p2_concat_86185 <= p2_concat_86185_comb;
    p2_concat_86186 <= p2_concat_86186_comb;
    p2_concat_86187 <= p2_concat_86187_comb;
    p2_concat_86188 <= p2_concat_86188_comb;
    p2_concat_86189 <= p2_concat_86189_comb;
    p2_concat_86190 <= p2_concat_86190_comb;
    p2_concat_86191 <= p2_concat_86191_comb;
    p2_concat_86192 <= p2_concat_86192_comb;
    p2_concat_86193 <= p2_concat_86193_comb;
    p2_concat_86194 <= p2_concat_86194_comb;
    p2_add_86327 <= p2_add_86327_comb;
    p2_bit_slice_86328 <= p2_bit_slice_86328_comb;
    p2_add_86329 <= p2_add_86329_comb;
    p2_bit_slice_86330 <= p2_bit_slice_86330_comb;
    p2_add_86331 <= p2_add_86331_comb;
    p2_bit_slice_86332 <= p2_bit_slice_86332_comb;
    p2_add_86333 <= p2_add_86333_comb;
    p2_bit_slice_86334 <= p2_bit_slice_86334_comb;
    p2_add_86335 <= p2_add_86335_comb;
    p2_bit_slice_86336 <= p2_bit_slice_86336_comb;
    p2_add_86337 <= p2_add_86337_comb;
    p2_bit_slice_86338 <= p2_bit_slice_86338_comb;
    p2_add_86343 <= p2_add_86343_comb;
    p2_bit_slice_86344 <= p2_bit_slice_86344_comb;
    p2_add_86345 <= p2_add_86345_comb;
    p2_bit_slice_86346 <= p2_bit_slice_86346_comb;
    p2_add_86347 <= p2_add_86347_comb;
    p2_bit_slice_86348 <= p2_bit_slice_86348_comb;
    p2_add_86349 <= p2_add_86349_comb;
    p2_bit_slice_86350 <= p2_bit_slice_86350_comb;
    p2_add_86351 <= p2_add_86351_comb;
    p2_bit_slice_86352 <= p2_bit_slice_86352_comb;
    p2_add_86353 <= p2_add_86353_comb;
    p2_bit_slice_86354 <= p2_bit_slice_86354_comb;
    p2_concat_86359 <= p2_concat_86359_comb;
    p2_concat_86360 <= p2_concat_86360_comb;
    p2_concat_86361 <= p2_concat_86361_comb;
    p2_concat_86362 <= p2_concat_86362_comb;
    p2_concat_86363 <= p2_concat_86363_comb;
    p2_concat_86364 <= p2_concat_86364_comb;
    p2_concat_86365 <= p2_concat_86365_comb;
    p2_concat_86366 <= p2_concat_86366_comb;
    p2_concat_86367 <= p2_concat_86367_comb;
    p2_concat_86368 <= p2_concat_86368_comb;
    p2_concat_86369 <= p2_concat_86369_comb;
    p2_concat_86370 <= p2_concat_86370_comb;
    p2_concat_86375 <= p2_concat_86375_comb;
    p2_concat_86376 <= p2_concat_86376_comb;
    p2_concat_86377 <= p2_concat_86377_comb;
    p2_concat_86378 <= p2_concat_86378_comb;
    p2_concat_86379 <= p2_concat_86379_comb;
    p2_concat_86380 <= p2_concat_86380_comb;
    p2_concat_86381 <= p2_concat_86381_comb;
    p2_concat_86382 <= p2_concat_86382_comb;
    p2_concat_86383 <= p2_concat_86383_comb;
    p2_concat_86384 <= p2_concat_86384_comb;
    p2_concat_86385 <= p2_concat_86385_comb;
    p2_concat_86386 <= p2_concat_86386_comb;
    p2_concat_86439 <= p2_concat_86439_comb;
    p2_concat_86440 <= p2_concat_86440_comb;
    p2_concat_86441 <= p2_concat_86441_comb;
    p2_concat_86442 <= p2_concat_86442_comb;
    p2_concat_86443 <= p2_concat_86443_comb;
    p2_concat_86444 <= p2_concat_86444_comb;
    p2_concat_86445 <= p2_concat_86445_comb;
    p2_concat_86446 <= p2_concat_86446_comb;
    p2_concat_86447 <= p2_concat_86447_comb;
    p2_concat_86448 <= p2_concat_86448_comb;
    p2_concat_86449 <= p2_concat_86449_comb;
    p2_concat_86450 <= p2_concat_86450_comb;
    p2_concat_86455 <= p2_concat_86455_comb;
    p2_concat_86456 <= p2_concat_86456_comb;
    p2_concat_86457 <= p2_concat_86457_comb;
    p2_concat_86458 <= p2_concat_86458_comb;
    p2_concat_86459 <= p2_concat_86459_comb;
    p2_concat_86460 <= p2_concat_86460_comb;
    p2_concat_86461 <= p2_concat_86461_comb;
    p2_concat_86462 <= p2_concat_86462_comb;
    p2_concat_86463 <= p2_concat_86463_comb;
    p2_concat_86464 <= p2_concat_86464_comb;
    p2_concat_86465 <= p2_concat_86465_comb;
    p2_concat_86466 <= p2_concat_86466_comb;
    p2_add_86471 <= p2_add_86471_comb;
    p2_bit_slice_86472 <= p2_bit_slice_86472_comb;
    p2_add_86473 <= p2_add_86473_comb;
    p2_bit_slice_86474 <= p2_bit_slice_86474_comb;
    p2_add_86475 <= p2_add_86475_comb;
    p2_bit_slice_86476 <= p2_bit_slice_86476_comb;
    p2_add_86477 <= p2_add_86477_comb;
    p2_bit_slice_86478 <= p2_bit_slice_86478_comb;
    p2_add_86479 <= p2_add_86479_comb;
    p2_bit_slice_86480 <= p2_bit_slice_86480_comb;
    p2_add_86481 <= p2_add_86481_comb;
    p2_bit_slice_86482 <= p2_bit_slice_86482_comb;
    p2_add_86487 <= p2_add_86487_comb;
    p2_bit_slice_86488 <= p2_bit_slice_86488_comb;
    p2_add_86489 <= p2_add_86489_comb;
    p2_bit_slice_86490 <= p2_bit_slice_86490_comb;
    p2_add_86491 <= p2_add_86491_comb;
    p2_bit_slice_86492 <= p2_bit_slice_86492_comb;
    p2_add_86493 <= p2_add_86493_comb;
    p2_bit_slice_86494 <= p2_bit_slice_86494_comb;
    p2_add_86495 <= p2_add_86495_comb;
    p2_bit_slice_86496 <= p2_bit_slice_86496_comb;
    p2_add_86497 <= p2_add_86497_comb;
    p2_bit_slice_86498 <= p2_bit_slice_86498_comb;
    p2_add_86565 <= p2_add_86565_comb;
    p2_add_86566 <= p2_add_86566_comb;
    p2_add_86567 <= p2_add_86567_comb;
    p2_add_86570 <= p2_add_86570_comb;
    p2_add_86571 <= p2_add_86571_comb;
    p2_add_86572 <= p2_add_86572_comb;
    p2_sum__1079 <= p2_sum__1079_comb;
    p2_add_86576 <= p2_add_86576_comb;
    p2_add_86577 <= p2_add_86577_comb;
    p2_sum__1077 <= p2_sum__1077_comb;
    p2_sum__1075 <= p2_sum__1075_comb;
    p2_add_86602 <= p2_add_86602_comb;
    p2_add_86603 <= p2_add_86603_comb;
    p2_sum__1073 <= p2_sum__1073_comb;
    p2_add_86611 <= p2_add_86611_comb;
    p2_add_86612 <= p2_add_86612_comb;
    p2_add_86613 <= p2_add_86613_comb;
    p2_add_86615 <= p2_add_86615_comb;
    p2_add_86616 <= p2_add_86616_comb;
    p2_add_86617 <= p2_add_86617_comb;
    p2_add_86619 <= p2_add_86619_comb;
    p2_add_86620 <= p2_add_86620_comb;
    p2_add_86621 <= p2_add_86621_comb;
    p2_add_86622 <= p2_add_86622_comb;
    p2_add_86623 <= p2_add_86623_comb;
    p2_add_86624 <= p2_add_86624_comb;
    p2_bit_slice_86625 <= p2_bit_slice_86625_comb;
    p2_bit_slice_86626 <= p2_bit_slice_86626_comb;
    p2_bit_slice_86627 <= p2_bit_slice_86627_comb;
    p2_bit_slice_86628 <= p2_bit_slice_86628_comb;
  end

  // ===== Pipe stage 3:
  wire [24:0] p3_sum__1544_comb;
  wire [24:0] p3_sum__1545_comb;
  wire [24:0] p3_sum__1546_comb;
  wire [24:0] p3_sum__1547_comb;
  wire [24:0] p3_sum__1516_comb;
  wire [24:0] p3_sum__1517_comb;
  wire [24:0] p3_sum__1518_comb;
  wire [24:0] p3_sum__1519_comb;
  wire [24:0] p3_sum__1488_comb;
  wire [24:0] p3_sum__1489_comb;
  wire [24:0] p3_sum__1490_comb;
  wire [24:0] p3_sum__1491_comb;
  wire [24:0] p3_sum__1432_comb;
  wire [24:0] p3_sum__1433_comb;
  wire [24:0] p3_sum__1434_comb;
  wire [24:0] p3_sum__1435_comb;
  wire [24:0] p3_sum__1404_comb;
  wire [24:0] p3_sum__1405_comb;
  wire [24:0] p3_sum__1406_comb;
  wire [24:0] p3_sum__1407_comb;
  wire [24:0] p3_sum__1376_comb;
  wire [24:0] p3_sum__1377_comb;
  wire [24:0] p3_sum__1378_comb;
  wire [24:0] p3_sum__1379_comb;
  wire [24:0] p3_sum__1536_comb;
  wire [24:0] p3_sum__1537_comb;
  wire [24:0] p3_sum__1538_comb;
  wire [24:0] p3_sum__1539_comb;
  wire [24:0] p3_sum__1508_comb;
  wire [24:0] p3_sum__1509_comb;
  wire [24:0] p3_sum__1510_comb;
  wire [24:0] p3_sum__1511_comb;
  wire [24:0] p3_sum__1480_comb;
  wire [24:0] p3_sum__1481_comb;
  wire [24:0] p3_sum__1482_comb;
  wire [24:0] p3_sum__1483_comb;
  wire [24:0] p3_sum__1424_comb;
  wire [24:0] p3_sum__1425_comb;
  wire [24:0] p3_sum__1426_comb;
  wire [24:0] p3_sum__1427_comb;
  wire [24:0] p3_sum__1396_comb;
  wire [24:0] p3_sum__1397_comb;
  wire [24:0] p3_sum__1398_comb;
  wire [24:0] p3_sum__1399_comb;
  wire [24:0] p3_sum__1368_comb;
  wire [24:0] p3_sum__1369_comb;
  wire [24:0] p3_sum__1370_comb;
  wire [24:0] p3_sum__1371_comb;
  wire [24:0] p3_sum__1232_comb;
  wire [24:0] p3_sum__1233_comb;
  wire [24:0] p3_sum__1218_comb;
  wire [24:0] p3_sum__1219_comb;
  wire [24:0] p3_sum__1204_comb;
  wire [24:0] p3_sum__1205_comb;
  wire [24:0] p3_sum__1176_comb;
  wire [24:0] p3_sum__1177_comb;
  wire [24:0] p3_sum__1162_comb;
  wire [24:0] p3_sum__1163_comb;
  wire [24:0] p3_sum__1148_comb;
  wire [24:0] p3_sum__1149_comb;
  wire [24:0] p3_sum__1228_comb;
  wire [24:0] p3_sum__1229_comb;
  wire [24:0] p3_sum__1214_comb;
  wire [24:0] p3_sum__1215_comb;
  wire [24:0] p3_sum__1200_comb;
  wire [24:0] p3_sum__1201_comb;
  wire [24:0] p3_sum__1172_comb;
  wire [24:0] p3_sum__1173_comb;
  wire [24:0] p3_sum__1158_comb;
  wire [24:0] p3_sum__1159_comb;
  wire [24:0] p3_sum__1144_comb;
  wire [24:0] p3_sum__1145_comb;
  wire [24:0] p3_sum__1224_comb;
  wire [24:0] p3_sum__1225_comb;
  wire [24:0] p3_sum__1210_comb;
  wire [24:0] p3_sum__1211_comb;
  wire [24:0] p3_sum__1196_comb;
  wire [24:0] p3_sum__1197_comb;
  wire [24:0] p3_sum__1168_comb;
  wire [24:0] p3_sum__1169_comb;
  wire [24:0] p3_sum__1154_comb;
  wire [24:0] p3_sum__1155_comb;
  wire [24:0] p3_sum__1140_comb;
  wire [24:0] p3_sum__1141_comb;
  wire [24:0] p3_sum__1220_comb;
  wire [24:0] p3_sum__1221_comb;
  wire [24:0] p3_sum__1206_comb;
  wire [24:0] p3_sum__1207_comb;
  wire [24:0] p3_sum__1192_comb;
  wire [24:0] p3_sum__1193_comb;
  wire [24:0] p3_sum__1164_comb;
  wire [24:0] p3_sum__1165_comb;
  wire [24:0] p3_sum__1150_comb;
  wire [24:0] p3_sum__1151_comb;
  wire [24:0] p3_sum__1136_comb;
  wire [24:0] p3_sum__1137_comb;
  wire [24:0] p3_sum__1072_comb;
  wire [24:0] p3_sum__1065_comb;
  wire [24:0] p3_sum__1058_comb;
  wire [24:0] p3_sum__1044_comb;
  wire [24:0] p3_sum__1037_comb;
  wire [24:0] p3_sum__1030_comb;
  wire [23:0] p3_add_87140_comb;
  wire [23:0] p3_add_87141_comb;
  wire [23:0] p3_add_87142_comb;
  wire [23:0] p3_add_87143_comb;
  wire [23:0] p3_add_87144_comb;
  wire [23:0] p3_add_87145_comb;
  wire [23:0] p3_add_87146_comb;
  wire [23:0] p3_add_87147_comb;
  wire [23:0] p3_add_87148_comb;
  wire [23:0] p3_add_87149_comb;
  wire [23:0] p3_add_87150_comb;
  wire [23:0] p3_add_87151_comb;
  wire [24:0] p3_sum__1070_comb;
  wire [24:0] p3_sum__1063_comb;
  wire [24:0] p3_sum__1056_comb;
  wire [24:0] p3_sum__1042_comb;
  wire [24:0] p3_sum__1035_comb;
  wire [24:0] p3_sum__1028_comb;
  wire [24:0] p3_sum__1068_comb;
  wire [24:0] p3_sum__1061_comb;
  wire [24:0] p3_sum__1054_comb;
  wire [24:0] p3_sum__1040_comb;
  wire [24:0] p3_sum__1033_comb;
  wire [24:0] p3_sum__1026_comb;
  wire [23:0] p3_add_87178_comb;
  wire [23:0] p3_add_87179_comb;
  wire [23:0] p3_add_87180_comb;
  wire [23:0] p3_add_87181_comb;
  wire [23:0] p3_add_87182_comb;
  wire [23:0] p3_add_87183_comb;
  wire [23:0] p3_add_87184_comb;
  wire [23:0] p3_add_87185_comb;
  wire [23:0] p3_add_87186_comb;
  wire [23:0] p3_add_87187_comb;
  wire [23:0] p3_add_87188_comb;
  wire [23:0] p3_add_87189_comb;
  wire [24:0] p3_sum__1066_comb;
  wire [24:0] p3_sum__1059_comb;
  wire [24:0] p3_sum__1052_comb;
  wire [24:0] p3_sum__1038_comb;
  wire [24:0] p3_sum__1031_comb;
  wire [24:0] p3_sum__1024_comb;
  wire [23:0] p3_umul_29018_NarrowedMult__comb;
  wire [23:0] p3_umul_29020_NarrowedMult__comb;
  wire [23:0] p3_umul_29022_NarrowedMult__comb;
  wire [23:0] p3_umul_29026_NarrowedMult__comb;
  wire [23:0] p3_umul_29028_NarrowedMult__comb;
  wire [23:0] p3_umul_29030_NarrowedMult__comb;
  wire [24:0] p3_add_87209_comb;
  wire [24:0] p3_add_87210_comb;
  wire [24:0] p3_add_87211_comb;
  wire [24:0] p3_add_87212_comb;
  wire [24:0] p3_add_87213_comb;
  wire [24:0] p3_add_87214_comb;
  wire [24:0] p3_add_87215_comb;
  wire [23:0] p3_add_87216_comb;
  wire [23:0] p3_add_87217_comb;
  wire [23:0] p3_add_87218_comb;
  wire [23:0] p3_add_87219_comb;
  wire [23:0] p3_add_87220_comb;
  wire [23:0] p3_add_87221_comb;
  wire [23:0] p3_add_87222_comb;
  wire [24:0] p3_add_87223_comb;
  wire [24:0] p3_add_87224_comb;
  wire [24:0] p3_add_87225_comb;
  wire [24:0] p3_add_87226_comb;
  wire [24:0] p3_add_87227_comb;
  wire [24:0] p3_add_87228_comb;
  wire [24:0] p3_add_87229_comb;
  wire [24:0] p3_add_87230_comb;
  wire [24:0] p3_add_87231_comb;
  wire [24:0] p3_add_87232_comb;
  wire [24:0] p3_add_87233_comb;
  wire [24:0] p3_add_87234_comb;
  wire [24:0] p3_add_87235_comb;
  wire [24:0] p3_add_87236_comb;
  wire [23:0] p3_add_87237_comb;
  wire [23:0] p3_add_87238_comb;
  wire [23:0] p3_add_87239_comb;
  wire [23:0] p3_add_87240_comb;
  wire [23:0] p3_add_87241_comb;
  wire [23:0] p3_add_87242_comb;
  wire [23:0] p3_add_87243_comb;
  wire [24:0] p3_add_87244_comb;
  wire [24:0] p3_add_87245_comb;
  wire [24:0] p3_add_87246_comb;
  wire [24:0] p3_add_87247_comb;
  wire [24:0] p3_add_87248_comb;
  wire [24:0] p3_add_87249_comb;
  wire [24:0] p3_add_87250_comb;
  wire [16:0] p3_bit_slice_87251_comb;
  wire [16:0] p3_bit_slice_87252_comb;
  wire [16:0] p3_bit_slice_87253_comb;
  wire [16:0] p3_bit_slice_87254_comb;
  wire [16:0] p3_bit_slice_87255_comb;
  wire [16:0] p3_bit_slice_87256_comb;
  wire [16:0] p3_bit_slice_87257_comb;
  wire [16:0] p3_bit_slice_87258_comb;
  wire [16:0] p3_bit_slice_87259_comb;
  wire [16:0] p3_bit_slice_87260_comb;
  wire [16:0] p3_bit_slice_87261_comb;
  wire [16:0] p3_bit_slice_87262_comb;
  wire [16:0] p3_bit_slice_87263_comb;
  wire [16:0] p3_bit_slice_87264_comb;
  wire [16:0] p3_bit_slice_87265_comb;
  wire [16:0] p3_bit_slice_87266_comb;
  wire [16:0] p3_bit_slice_87267_comb;
  wire [16:0] p3_bit_slice_87268_comb;
  wire [16:0] p3_bit_slice_87269_comb;
  wire [16:0] p3_bit_slice_87270_comb;
  wire [16:0] p3_bit_slice_87271_comb;
  wire [16:0] p3_bit_slice_87272_comb;
  wire [16:0] p3_bit_slice_87273_comb;
  wire [16:0] p3_bit_slice_87274_comb;
  wire [16:0] p3_bit_slice_87275_comb;
  wire [16:0] p3_bit_slice_87276_comb;
  wire [16:0] p3_bit_slice_87277_comb;
  wire [16:0] p3_bit_slice_87278_comb;
  wire [16:0] p3_bit_slice_87279_comb;
  wire [16:0] p3_bit_slice_87280_comb;
  wire [16:0] p3_bit_slice_87281_comb;
  wire [16:0] p3_bit_slice_87282_comb;
  wire [16:0] p3_bit_slice_87283_comb;
  wire [16:0] p3_bit_slice_87284_comb;
  wire [16:0] p3_bit_slice_87285_comb;
  wire [16:0] p3_bit_slice_87286_comb;
  wire [16:0] p3_bit_slice_87287_comb;
  wire [16:0] p3_bit_slice_87288_comb;
  wire [16:0] p3_bit_slice_87289_comb;
  wire [16:0] p3_bit_slice_87290_comb;
  wire [16:0] p3_bit_slice_87291_comb;
  wire [16:0] p3_bit_slice_87292_comb;
  wire [16:0] p3_bit_slice_87293_comb;
  wire [16:0] p3_bit_slice_87294_comb;
  wire [16:0] p3_bit_slice_87295_comb;
  wire [16:0] p3_bit_slice_87296_comb;
  wire [16:0] p3_bit_slice_87297_comb;
  wire [16:0] p3_bit_slice_87298_comb;
  wire [16:0] p3_bit_slice_87299_comb;
  wire [16:0] p3_bit_slice_87300_comb;
  wire [16:0] p3_bit_slice_87301_comb;
  wire [16:0] p3_bit_slice_87302_comb;
  wire [16:0] p3_bit_slice_87303_comb;
  wire [16:0] p3_bit_slice_87304_comb;
  wire [16:0] p3_bit_slice_87305_comb;
  wire [16:0] p3_bit_slice_87306_comb;
  wire [16:0] p3_bit_slice_87307_comb;
  wire [16:0] p3_bit_slice_87308_comb;
  wire [16:0] p3_bit_slice_87309_comb;
  wire [16:0] p3_bit_slice_87310_comb;
  wire [17:0] p3_add_87439_comb;
  wire [17:0] p3_add_87440_comb;
  wire [17:0] p3_add_87441_comb;
  wire [17:0] p3_add_87442_comb;
  wire [17:0] p3_add_87443_comb;
  wire [17:0] p3_add_87444_comb;
  wire [17:0] p3_add_87445_comb;
  wire [17:0] p3_add_87446_comb;
  wire [17:0] p3_add_87447_comb;
  wire [17:0] p3_add_87448_comb;
  wire [17:0] p3_add_87449_comb;
  wire [17:0] p3_add_87450_comb;
  wire [17:0] p3_add_87451_comb;
  wire [17:0] p3_add_87452_comb;
  wire [17:0] p3_add_87453_comb;
  wire [17:0] p3_add_87454_comb;
  wire [17:0] p3_add_87455_comb;
  wire [17:0] p3_add_87456_comb;
  wire [17:0] p3_add_87457_comb;
  wire [17:0] p3_add_87458_comb;
  wire [17:0] p3_add_87459_comb;
  wire [17:0] p3_add_87460_comb;
  wire [17:0] p3_add_87461_comb;
  wire [17:0] p3_add_87462_comb;
  wire [17:0] p3_add_87463_comb;
  wire [17:0] p3_add_87464_comb;
  wire [17:0] p3_add_87465_comb;
  wire [17:0] p3_add_87466_comb;
  wire [17:0] p3_add_87467_comb;
  wire [17:0] p3_add_87468_comb;
  wire [17:0] p3_add_87469_comb;
  wire [17:0] p3_add_87470_comb;
  wire [17:0] p3_add_87471_comb;
  wire [17:0] p3_add_87472_comb;
  wire [17:0] p3_add_87473_comb;
  wire [17:0] p3_add_87474_comb;
  wire [17:0] p3_add_87475_comb;
  wire [17:0] p3_add_87476_comb;
  wire [17:0] p3_add_87477_comb;
  wire [17:0] p3_add_87478_comb;
  wire [17:0] p3_add_87479_comb;
  wire [17:0] p3_add_87480_comb;
  wire [17:0] p3_add_87481_comb;
  wire [17:0] p3_add_87482_comb;
  wire [17:0] p3_add_87483_comb;
  wire [17:0] p3_add_87484_comb;
  wire [17:0] p3_add_87485_comb;
  wire [17:0] p3_add_87486_comb;
  wire [17:0] p3_add_87487_comb;
  wire [17:0] p3_add_87488_comb;
  wire [17:0] p3_add_87489_comb;
  wire [17:0] p3_add_87490_comb;
  wire [17:0] p3_add_87491_comb;
  wire [17:0] p3_add_87492_comb;
  wire [17:0] p3_add_87493_comb;
  wire [17:0] p3_add_87494_comb;
  wire [17:0] p3_add_87495_comb;
  wire [17:0] p3_add_87496_comb;
  wire [17:0] p3_add_87497_comb;
  wire [17:0] p3_add_87498_comb;
  wire [17:0] p3_add_87499_comb;
  wire [17:0] p3_add_87500_comb;
  wire [17:0] p3_add_87501_comb;
  wire [17:0] p3_add_87502_comb;
  wire [9:0] p3_bit_slice_87503_comb;
  wire [9:0] p3_bit_slice_87504_comb;
  wire [9:0] p3_bit_slice_87505_comb;
  wire [9:0] p3_bit_slice_87506_comb;
  wire [9:0] p3_bit_slice_87507_comb;
  wire [9:0] p3_bit_slice_87508_comb;
  wire [9:0] p3_bit_slice_87509_comb;
  wire [9:0] p3_bit_slice_87510_comb;
  wire [9:0] p3_bit_slice_87511_comb;
  wire [9:0] p3_bit_slice_87512_comb;
  wire [9:0] p3_bit_slice_87513_comb;
  wire [9:0] p3_bit_slice_87514_comb;
  wire [9:0] p3_bit_slice_87515_comb;
  wire [9:0] p3_bit_slice_87516_comb;
  wire [9:0] p3_bit_slice_87517_comb;
  wire [9:0] p3_bit_slice_87518_comb;
  wire [9:0] p3_bit_slice_87519_comb;
  wire [9:0] p3_bit_slice_87520_comb;
  wire [9:0] p3_bit_slice_87521_comb;
  wire [9:0] p3_bit_slice_87522_comb;
  wire [9:0] p3_bit_slice_87523_comb;
  wire [9:0] p3_bit_slice_87524_comb;
  wire [9:0] p3_bit_slice_87525_comb;
  wire [9:0] p3_bit_slice_87526_comb;
  wire [9:0] p3_bit_slice_87527_comb;
  wire [9:0] p3_bit_slice_87528_comb;
  wire [9:0] p3_bit_slice_87529_comb;
  wire [9:0] p3_bit_slice_87530_comb;
  wire [9:0] p3_bit_slice_87531_comb;
  wire [9:0] p3_bit_slice_87532_comb;
  wire [9:0] p3_bit_slice_87533_comb;
  wire [9:0] p3_bit_slice_87534_comb;
  wire [9:0] p3_bit_slice_87535_comb;
  wire [9:0] p3_bit_slice_87536_comb;
  wire [9:0] p3_bit_slice_87537_comb;
  wire [9:0] p3_bit_slice_87538_comb;
  wire [9:0] p3_bit_slice_87539_comb;
  wire [9:0] p3_bit_slice_87540_comb;
  wire [9:0] p3_bit_slice_87541_comb;
  wire [9:0] p3_bit_slice_87542_comb;
  wire [9:0] p3_bit_slice_87543_comb;
  wire [9:0] p3_bit_slice_87544_comb;
  wire [9:0] p3_bit_slice_87545_comb;
  wire [9:0] p3_bit_slice_87546_comb;
  wire [9:0] p3_bit_slice_87547_comb;
  wire [9:0] p3_bit_slice_87548_comb;
  wire [9:0] p3_bit_slice_87549_comb;
  wire [9:0] p3_bit_slice_87550_comb;
  wire [9:0] p3_bit_slice_87551_comb;
  wire [9:0] p3_bit_slice_87552_comb;
  wire [9:0] p3_bit_slice_87553_comb;
  wire [9:0] p3_bit_slice_87554_comb;
  wire [9:0] p3_bit_slice_87555_comb;
  wire [9:0] p3_bit_slice_87556_comb;
  wire [9:0] p3_bit_slice_87557_comb;
  wire [9:0] p3_bit_slice_87558_comb;
  wire [9:0] p3_bit_slice_87559_comb;
  wire [9:0] p3_bit_slice_87560_comb;
  wire [9:0] p3_bit_slice_87561_comb;
  wire [9:0] p3_bit_slice_87562_comb;
  wire [9:0] p3_bit_slice_87563_comb;
  wire [9:0] p3_bit_slice_87564_comb;
  wire [9:0] p3_bit_slice_87565_comb;
  wire [9:0] p3_bit_slice_87566_comb;
  wire [10:0] p3_add_87695_comb;
  wire [10:0] p3_add_87697_comb;
  wire [10:0] p3_add_87699_comb;
  wire [10:0] p3_add_87701_comb;
  wire [10:0] p3_add_87703_comb;
  wire [10:0] p3_add_87705_comb;
  wire [10:0] p3_add_87707_comb;
  wire [10:0] p3_add_87709_comb;
  wire [10:0] p3_add_87711_comb;
  wire [10:0] p3_add_87713_comb;
  wire [10:0] p3_add_87715_comb;
  wire [10:0] p3_add_87717_comb;
  wire [10:0] p3_add_87719_comb;
  wire [10:0] p3_add_87721_comb;
  wire [10:0] p3_add_87723_comb;
  wire [10:0] p3_add_87725_comb;
  wire [10:0] p3_add_87727_comb;
  wire [10:0] p3_add_87729_comb;
  wire [10:0] p3_add_87731_comb;
  wire [10:0] p3_add_87733_comb;
  wire [10:0] p3_add_87735_comb;
  wire [10:0] p3_add_87737_comb;
  wire [10:0] p3_add_87739_comb;
  wire [10:0] p3_add_87741_comb;
  wire [10:0] p3_add_87743_comb;
  wire [10:0] p3_add_87745_comb;
  wire [10:0] p3_add_87747_comb;
  wire [10:0] p3_add_87749_comb;
  wire [10:0] p3_add_87751_comb;
  wire [10:0] p3_add_87753_comb;
  wire [10:0] p3_add_87755_comb;
  wire [10:0] p3_add_87757_comb;
  wire [10:0] p3_add_87759_comb;
  wire [10:0] p3_add_87761_comb;
  wire [10:0] p3_add_87763_comb;
  wire [10:0] p3_add_87765_comb;
  wire [10:0] p3_add_87767_comb;
  wire [10:0] p3_add_87769_comb;
  wire [10:0] p3_add_87771_comb;
  wire [10:0] p3_add_87773_comb;
  wire [10:0] p3_add_87775_comb;
  wire [10:0] p3_add_87777_comb;
  wire [10:0] p3_add_87779_comb;
  wire [10:0] p3_add_87781_comb;
  wire [10:0] p3_add_87783_comb;
  wire [10:0] p3_add_87785_comb;
  wire [10:0] p3_add_87787_comb;
  wire [10:0] p3_add_87789_comb;
  wire [10:0] p3_add_87791_comb;
  wire [10:0] p3_add_87793_comb;
  wire [10:0] p3_add_87795_comb;
  wire [10:0] p3_add_87797_comb;
  wire [10:0] p3_add_87799_comb;
  wire [10:0] p3_add_87801_comb;
  wire [10:0] p3_add_87803_comb;
  wire [10:0] p3_add_87805_comb;
  wire [10:0] p3_add_87807_comb;
  wire [10:0] p3_add_87809_comb;
  wire [10:0] p3_add_87811_comb;
  wire [10:0] p3_add_87813_comb;
  wire [10:0] p3_add_87815_comb;
  wire [10:0] p3_add_87817_comb;
  wire [10:0] p3_add_87819_comb;
  wire [10:0] p3_add_87821_comb;
  wire [17:0] p3_concat_87823_comb;
  wire [17:0] p3_concat_87826_comb;
  wire [17:0] p3_concat_87829_comb;
  wire [17:0] p3_concat_87832_comb;
  wire [17:0] p3_concat_87835_comb;
  wire [17:0] p3_concat_87838_comb;
  wire [17:0] p3_concat_87841_comb;
  wire [17:0] p3_concat_87844_comb;
  wire [17:0] p3_concat_87847_comb;
  wire [17:0] p3_concat_87850_comb;
  wire [17:0] p3_concat_87853_comb;
  wire [17:0] p3_concat_87856_comb;
  wire [17:0] p3_concat_87859_comb;
  wire [17:0] p3_concat_87862_comb;
  wire [17:0] p3_concat_87865_comb;
  wire [17:0] p3_concat_87868_comb;
  wire [17:0] p3_concat_87871_comb;
  wire [17:0] p3_concat_87874_comb;
  wire [17:0] p3_concat_87877_comb;
  wire [17:0] p3_concat_87880_comb;
  wire [17:0] p3_concat_87883_comb;
  wire [17:0] p3_concat_87886_comb;
  wire [17:0] p3_concat_87889_comb;
  wire [17:0] p3_concat_87892_comb;
  wire [17:0] p3_concat_87895_comb;
  wire [17:0] p3_concat_87898_comb;
  wire [17:0] p3_concat_87901_comb;
  wire [17:0] p3_concat_87904_comb;
  wire [17:0] p3_concat_87907_comb;
  wire [17:0] p3_concat_87910_comb;
  wire [17:0] p3_concat_87913_comb;
  wire [17:0] p3_concat_87916_comb;
  wire [17:0] p3_concat_87919_comb;
  wire [17:0] p3_concat_87922_comb;
  wire [17:0] p3_concat_87925_comb;
  wire [17:0] p3_concat_87928_comb;
  wire [17:0] p3_concat_87931_comb;
  wire [17:0] p3_concat_87934_comb;
  wire [17:0] p3_concat_87937_comb;
  wire [17:0] p3_concat_87940_comb;
  wire [17:0] p3_concat_87943_comb;
  wire [17:0] p3_concat_87946_comb;
  wire [17:0] p3_concat_87949_comb;
  wire [17:0] p3_concat_87952_comb;
  wire [17:0] p3_concat_87955_comb;
  wire [17:0] p3_concat_87958_comb;
  wire [17:0] p3_concat_87961_comb;
  wire [17:0] p3_concat_87964_comb;
  wire [17:0] p3_concat_87967_comb;
  wire [17:0] p3_concat_87970_comb;
  wire [17:0] p3_concat_87973_comb;
  wire [17:0] p3_concat_87976_comb;
  wire [17:0] p3_concat_87979_comb;
  wire [17:0] p3_concat_87982_comb;
  wire [17:0] p3_concat_87985_comb;
  wire [17:0] p3_concat_87988_comb;
  wire [17:0] p3_concat_87991_comb;
  wire [17:0] p3_concat_87994_comb;
  wire [17:0] p3_concat_87997_comb;
  wire [17:0] p3_concat_88000_comb;
  wire [17:0] p3_concat_88003_comb;
  wire [17:0] p3_concat_88006_comb;
  wire [17:0] p3_concat_88009_comb;
  wire [17:0] p3_concat_88012_comb;
  wire [9:0] p3_clipped__136_comb;
  wire [9:0] p3_clipped__152_comb;
  wire [9:0] p3_clipped__168_comb;
  wire [9:0] p3_clipped__184_comb;
  wire [9:0] p3_clipped__200_comb;
  wire [9:0] p3_clipped__216_comb;
  wire [9:0] p3_clipped__232_comb;
  wire [9:0] p3_clipped__248_comb;
  wire [9:0] p3_clipped__137_comb;
  wire [9:0] p3_clipped__153_comb;
  wire [9:0] p3_clipped__169_comb;
  wire [9:0] p3_clipped__185_comb;
  wire [9:0] p3_clipped__201_comb;
  wire [9:0] p3_clipped__217_comb;
  wire [9:0] p3_clipped__233_comb;
  wire [9:0] p3_clipped__249_comb;
  wire [9:0] p3_clipped__138_comb;
  wire [9:0] p3_clipped__154_comb;
  wire [9:0] p3_clipped__170_comb;
  wire [9:0] p3_clipped__186_comb;
  wire [9:0] p3_clipped__202_comb;
  wire [9:0] p3_clipped__218_comb;
  wire [9:0] p3_clipped__234_comb;
  wire [9:0] p3_clipped__250_comb;
  wire [9:0] p3_clipped__139_comb;
  wire [9:0] p3_clipped__155_comb;
  wire [9:0] p3_clipped__171_comb;
  wire [9:0] p3_clipped__187_comb;
  wire [9:0] p3_clipped__203_comb;
  wire [9:0] p3_clipped__219_comb;
  wire [9:0] p3_clipped__235_comb;
  wire [9:0] p3_clipped__251_comb;
  wire [9:0] p3_clipped__140_comb;
  wire [9:0] p3_clipped__156_comb;
  wire [9:0] p3_clipped__172_comb;
  wire [9:0] p3_clipped__188_comb;
  wire [9:0] p3_clipped__204_comb;
  wire [9:0] p3_clipped__220_comb;
  wire [9:0] p3_clipped__236_comb;
  wire [9:0] p3_clipped__252_comb;
  wire [9:0] p3_clipped__141_comb;
  wire [9:0] p3_clipped__157_comb;
  wire [9:0] p3_clipped__173_comb;
  wire [9:0] p3_clipped__189_comb;
  wire [9:0] p3_clipped__205_comb;
  wire [9:0] p3_clipped__221_comb;
  wire [9:0] p3_clipped__237_comb;
  wire [9:0] p3_clipped__253_comb;
  wire [9:0] p3_clipped__142_comb;
  wire [9:0] p3_clipped__158_comb;
  wire [9:0] p3_clipped__174_comb;
  wire [9:0] p3_clipped__190_comb;
  wire [9:0] p3_clipped__206_comb;
  wire [9:0] p3_clipped__222_comb;
  wire [9:0] p3_clipped__238_comb;
  wire [9:0] p3_clipped__254_comb;
  wire [9:0] p3_clipped__143_comb;
  wire [9:0] p3_clipped__159_comb;
  wire [9:0] p3_clipped__175_comb;
  wire [9:0] p3_clipped__191_comb;
  wire [9:0] p3_clipped__207_comb;
  wire [9:0] p3_clipped__223_comb;
  wire [9:0] p3_clipped__239_comb;
  wire [9:0] p3_clipped__255_comb;
  wire [9:0] p3_array_88527_comb[0:7];
  wire [9:0] p3_array_88528_comb[0:7];
  wire [9:0] p3_array_88529_comb[0:7];
  wire [9:0] p3_array_88530_comb[0:7];
  wire [9:0] p3_array_88531_comb[0:7];
  wire [9:0] p3_array_88532_comb[0:7];
  wire [9:0] p3_array_88533_comb[0:7];
  wire [9:0] p3_array_88534_comb[0:7];
  wire [9:0] p3_col_transformed_comb[0:7][0:7];
  assign p3_sum__1544_comb = {{5{p2_concat_86103[19]}}, p2_concat_86103};
  assign p3_sum__1545_comb = {{5{p2_concat_86104[19]}}, p2_concat_86104};
  assign p3_sum__1546_comb = {{5{p2_concat_86105[19]}}, p2_concat_86105};
  assign p3_sum__1547_comb = {{5{p2_concat_86106[19]}}, p2_concat_86106};
  assign p3_sum__1516_comb = {{5{p2_concat_86107[19]}}, p2_concat_86107};
  assign p3_sum__1517_comb = {{5{p2_concat_86108[19]}}, p2_concat_86108};
  assign p3_sum__1518_comb = {{5{p2_concat_86109[19]}}, p2_concat_86109};
  assign p3_sum__1519_comb = {{5{p2_concat_86110[19]}}, p2_concat_86110};
  assign p3_sum__1488_comb = {{5{p2_concat_86111[19]}}, p2_concat_86111};
  assign p3_sum__1489_comb = {{5{p2_concat_86112[19]}}, p2_concat_86112};
  assign p3_sum__1490_comb = {{5{p2_concat_86113[19]}}, p2_concat_86113};
  assign p3_sum__1491_comb = {{5{p2_concat_86114[19]}}, p2_concat_86114};
  assign p3_sum__1432_comb = {{5{p2_concat_86119[19]}}, p2_concat_86119};
  assign p3_sum__1433_comb = {{5{p2_concat_86120[19]}}, p2_concat_86120};
  assign p3_sum__1434_comb = {{5{p2_concat_86121[19]}}, p2_concat_86121};
  assign p3_sum__1435_comb = {{5{p2_concat_86122[19]}}, p2_concat_86122};
  assign p3_sum__1404_comb = {{5{p2_concat_86123[19]}}, p2_concat_86123};
  assign p3_sum__1405_comb = {{5{p2_concat_86124[19]}}, p2_concat_86124};
  assign p3_sum__1406_comb = {{5{p2_concat_86125[19]}}, p2_concat_86125};
  assign p3_sum__1407_comb = {{5{p2_concat_86126[19]}}, p2_concat_86126};
  assign p3_sum__1376_comb = {{5{p2_concat_86127[19]}}, p2_concat_86127};
  assign p3_sum__1377_comb = {{5{p2_concat_86128[19]}}, p2_concat_86128};
  assign p3_sum__1378_comb = {{5{p2_concat_86129[19]}}, p2_concat_86129};
  assign p3_sum__1379_comb = {{5{p2_concat_86130[19]}}, p2_concat_86130};
  assign p3_sum__1536_comb = {{5{p2_concat_86167[19]}}, p2_concat_86167};
  assign p3_sum__1537_comb = {{5{p2_concat_86168[19]}}, p2_concat_86168};
  assign p3_sum__1538_comb = {{5{p2_concat_86169[19]}}, p2_concat_86169};
  assign p3_sum__1539_comb = {{5{p2_concat_86170[19]}}, p2_concat_86170};
  assign p3_sum__1508_comb = {{5{p2_concat_86171[19]}}, p2_concat_86171};
  assign p3_sum__1509_comb = {{5{p2_concat_86172[19]}}, p2_concat_86172};
  assign p3_sum__1510_comb = {{5{p2_concat_86173[19]}}, p2_concat_86173};
  assign p3_sum__1511_comb = {{5{p2_concat_86174[19]}}, p2_concat_86174};
  assign p3_sum__1480_comb = {{5{p2_concat_86175[19]}}, p2_concat_86175};
  assign p3_sum__1481_comb = {{5{p2_concat_86176[19]}}, p2_concat_86176};
  assign p3_sum__1482_comb = {{5{p2_concat_86177[19]}}, p2_concat_86177};
  assign p3_sum__1483_comb = {{5{p2_concat_86178[19]}}, p2_concat_86178};
  assign p3_sum__1424_comb = {{5{p2_concat_86183[19]}}, p2_concat_86183};
  assign p3_sum__1425_comb = {{5{p2_concat_86184[19]}}, p2_concat_86184};
  assign p3_sum__1426_comb = {{5{p2_concat_86185[19]}}, p2_concat_86185};
  assign p3_sum__1427_comb = {{5{p2_concat_86186[19]}}, p2_concat_86186};
  assign p3_sum__1396_comb = {{5{p2_concat_86187[19]}}, p2_concat_86187};
  assign p3_sum__1397_comb = {{5{p2_concat_86188[19]}}, p2_concat_86188};
  assign p3_sum__1398_comb = {{5{p2_concat_86189[19]}}, p2_concat_86189};
  assign p3_sum__1399_comb = {{5{p2_concat_86190[19]}}, p2_concat_86190};
  assign p3_sum__1368_comb = {{5{p2_concat_86191[19]}}, p2_concat_86191};
  assign p3_sum__1369_comb = {{5{p2_concat_86192[19]}}, p2_concat_86192};
  assign p3_sum__1370_comb = {{5{p2_concat_86193[19]}}, p2_concat_86193};
  assign p3_sum__1371_comb = {{5{p2_concat_86194[19]}}, p2_concat_86194};
  assign p3_sum__1232_comb = {p2_add_86327, p2_bit_slice_86328};
  assign p3_sum__1233_comb = {p2_add_86329, p2_bit_slice_86330};
  assign p3_sum__1218_comb = {p2_add_86331, p2_bit_slice_86332};
  assign p3_sum__1219_comb = {p2_add_86333, p2_bit_slice_86334};
  assign p3_sum__1204_comb = {p2_add_86335, p2_bit_slice_86336};
  assign p3_sum__1205_comb = {p2_add_86337, p2_bit_slice_86338};
  assign p3_sum__1176_comb = {p2_add_86343, p2_bit_slice_86344};
  assign p3_sum__1177_comb = {p2_add_86345, p2_bit_slice_86346};
  assign p3_sum__1162_comb = {p2_add_86347, p2_bit_slice_86348};
  assign p3_sum__1163_comb = {p2_add_86349, p2_bit_slice_86350};
  assign p3_sum__1148_comb = {p2_add_86351, p2_bit_slice_86352};
  assign p3_sum__1149_comb = {p2_add_86353, p2_bit_slice_86354};
  assign p3_sum__1228_comb = p3_sum__1544_comb + p3_sum__1545_comb;
  assign p3_sum__1229_comb = p3_sum__1546_comb + p3_sum__1547_comb;
  assign p3_sum__1214_comb = p3_sum__1516_comb + p3_sum__1517_comb;
  assign p3_sum__1215_comb = p3_sum__1518_comb + p3_sum__1519_comb;
  assign p3_sum__1200_comb = p3_sum__1488_comb + p3_sum__1489_comb;
  assign p3_sum__1201_comb = p3_sum__1490_comb + p3_sum__1491_comb;
  assign p3_sum__1172_comb = p3_sum__1432_comb + p3_sum__1433_comb;
  assign p3_sum__1173_comb = p3_sum__1434_comb + p3_sum__1435_comb;
  assign p3_sum__1158_comb = p3_sum__1404_comb + p3_sum__1405_comb;
  assign p3_sum__1159_comb = p3_sum__1406_comb + p3_sum__1407_comb;
  assign p3_sum__1144_comb = p3_sum__1376_comb + p3_sum__1377_comb;
  assign p3_sum__1145_comb = p3_sum__1378_comb + p3_sum__1379_comb;
  assign p3_sum__1224_comb = p3_sum__1536_comb + p3_sum__1537_comb;
  assign p3_sum__1225_comb = p3_sum__1538_comb + p3_sum__1539_comb;
  assign p3_sum__1210_comb = p3_sum__1508_comb + p3_sum__1509_comb;
  assign p3_sum__1211_comb = p3_sum__1510_comb + p3_sum__1511_comb;
  assign p3_sum__1196_comb = p3_sum__1480_comb + p3_sum__1481_comb;
  assign p3_sum__1197_comb = p3_sum__1482_comb + p3_sum__1483_comb;
  assign p3_sum__1168_comb = p3_sum__1424_comb + p3_sum__1425_comb;
  assign p3_sum__1169_comb = p3_sum__1426_comb + p3_sum__1427_comb;
  assign p3_sum__1154_comb = p3_sum__1396_comb + p3_sum__1397_comb;
  assign p3_sum__1155_comb = p3_sum__1398_comb + p3_sum__1399_comb;
  assign p3_sum__1140_comb = p3_sum__1368_comb + p3_sum__1369_comb;
  assign p3_sum__1141_comb = p3_sum__1370_comb + p3_sum__1371_comb;
  assign p3_sum__1220_comb = {p2_add_86471, p2_bit_slice_86472};
  assign p3_sum__1221_comb = {p2_add_86473, p2_bit_slice_86474};
  assign p3_sum__1206_comb = {p2_add_86475, p2_bit_slice_86476};
  assign p3_sum__1207_comb = {p2_add_86477, p2_bit_slice_86478};
  assign p3_sum__1192_comb = {p2_add_86479, p2_bit_slice_86480};
  assign p3_sum__1193_comb = {p2_add_86481, p2_bit_slice_86482};
  assign p3_sum__1164_comb = {p2_add_86487, p2_bit_slice_86488};
  assign p3_sum__1165_comb = {p2_add_86489, p2_bit_slice_86490};
  assign p3_sum__1150_comb = {p2_add_86491, p2_bit_slice_86492};
  assign p3_sum__1151_comb = {p2_add_86493, p2_bit_slice_86494};
  assign p3_sum__1136_comb = {p2_add_86495, p2_bit_slice_86496};
  assign p3_sum__1137_comb = {p2_add_86497, p2_bit_slice_86498};
  assign p3_sum__1072_comb = p3_sum__1232_comb + p3_sum__1233_comb;
  assign p3_sum__1065_comb = p3_sum__1218_comb + p3_sum__1219_comb;
  assign p3_sum__1058_comb = p3_sum__1204_comb + p3_sum__1205_comb;
  assign p3_sum__1044_comb = p3_sum__1176_comb + p3_sum__1177_comb;
  assign p3_sum__1037_comb = p3_sum__1162_comb + p3_sum__1163_comb;
  assign p3_sum__1030_comb = p3_sum__1148_comb + p3_sum__1149_comb;
  assign p3_add_87140_comb = {{5{p2_concat_86359[18]}}, p2_concat_86359} + {{5{p2_concat_86360[18]}}, p2_concat_86360};
  assign p3_add_87141_comb = {{5{p2_concat_86361[18]}}, p2_concat_86361} + {{5{p2_concat_86362[18]}}, p2_concat_86362};
  assign p3_add_87142_comb = {{5{p2_concat_86363[18]}}, p2_concat_86363} + {{5{p2_concat_86364[18]}}, p2_concat_86364};
  assign p3_add_87143_comb = {{5{p2_concat_86365[18]}}, p2_concat_86365} + {{5{p2_concat_86366[18]}}, p2_concat_86366};
  assign p3_add_87144_comb = {{5{p2_concat_86367[18]}}, p2_concat_86367} + {{5{p2_concat_86368[18]}}, p2_concat_86368};
  assign p3_add_87145_comb = {{5{p2_concat_86369[18]}}, p2_concat_86369} + {{5{p2_concat_86370[18]}}, p2_concat_86370};
  assign p3_add_87146_comb = {{5{p2_concat_86375[18]}}, p2_concat_86375} + {{5{p2_concat_86376[18]}}, p2_concat_86376};
  assign p3_add_87147_comb = {{5{p2_concat_86377[18]}}, p2_concat_86377} + {{5{p2_concat_86378[18]}}, p2_concat_86378};
  assign p3_add_87148_comb = {{5{p2_concat_86379[18]}}, p2_concat_86379} + {{5{p2_concat_86380[18]}}, p2_concat_86380};
  assign p3_add_87149_comb = {{5{p2_concat_86381[18]}}, p2_concat_86381} + {{5{p2_concat_86382[18]}}, p2_concat_86382};
  assign p3_add_87150_comb = {{5{p2_concat_86383[18]}}, p2_concat_86383} + {{5{p2_concat_86384[18]}}, p2_concat_86384};
  assign p3_add_87151_comb = {{5{p2_concat_86385[18]}}, p2_concat_86385} + {{5{p2_concat_86386[18]}}, p2_concat_86386};
  assign p3_sum__1070_comb = p3_sum__1228_comb + p3_sum__1229_comb;
  assign p3_sum__1063_comb = p3_sum__1214_comb + p3_sum__1215_comb;
  assign p3_sum__1056_comb = p3_sum__1200_comb + p3_sum__1201_comb;
  assign p3_sum__1042_comb = p3_sum__1172_comb + p3_sum__1173_comb;
  assign p3_sum__1035_comb = p3_sum__1158_comb + p3_sum__1159_comb;
  assign p3_sum__1028_comb = p3_sum__1144_comb + p3_sum__1145_comb;
  assign p3_sum__1068_comb = p3_sum__1224_comb + p3_sum__1225_comb;
  assign p3_sum__1061_comb = p3_sum__1210_comb + p3_sum__1211_comb;
  assign p3_sum__1054_comb = p3_sum__1196_comb + p3_sum__1197_comb;
  assign p3_sum__1040_comb = p3_sum__1168_comb + p3_sum__1169_comb;
  assign p3_sum__1033_comb = p3_sum__1154_comb + p3_sum__1155_comb;
  assign p3_sum__1026_comb = p3_sum__1140_comb + p3_sum__1141_comb;
  assign p3_add_87178_comb = {{5{p2_concat_86439[18]}}, p2_concat_86439} + {{5{p2_concat_86440[18]}}, p2_concat_86440};
  assign p3_add_87179_comb = {{5{p2_concat_86441[18]}}, p2_concat_86441} + {{5{p2_concat_86442[18]}}, p2_concat_86442};
  assign p3_add_87180_comb = {{5{p2_concat_86443[18]}}, p2_concat_86443} + {{5{p2_concat_86444[18]}}, p2_concat_86444};
  assign p3_add_87181_comb = {{5{p2_concat_86445[18]}}, p2_concat_86445} + {{5{p2_concat_86446[18]}}, p2_concat_86446};
  assign p3_add_87182_comb = {{5{p2_concat_86447[18]}}, p2_concat_86447} + {{5{p2_concat_86448[18]}}, p2_concat_86448};
  assign p3_add_87183_comb = {{5{p2_concat_86449[18]}}, p2_concat_86449} + {{5{p2_concat_86450[18]}}, p2_concat_86450};
  assign p3_add_87184_comb = {{5{p2_concat_86455[18]}}, p2_concat_86455} + {{5{p2_concat_86456[18]}}, p2_concat_86456};
  assign p3_add_87185_comb = {{5{p2_concat_86457[18]}}, p2_concat_86457} + {{5{p2_concat_86458[18]}}, p2_concat_86458};
  assign p3_add_87186_comb = {{5{p2_concat_86459[18]}}, p2_concat_86459} + {{5{p2_concat_86460[18]}}, p2_concat_86460};
  assign p3_add_87187_comb = {{5{p2_concat_86461[18]}}, p2_concat_86461} + {{5{p2_concat_86462[18]}}, p2_concat_86462};
  assign p3_add_87188_comb = {{5{p2_concat_86463[18]}}, p2_concat_86463} + {{5{p2_concat_86464[18]}}, p2_concat_86464};
  assign p3_add_87189_comb = {{5{p2_concat_86465[18]}}, p2_concat_86465} + {{5{p2_concat_86466[18]}}, p2_concat_86466};
  assign p3_sum__1066_comb = p3_sum__1220_comb + p3_sum__1221_comb;
  assign p3_sum__1059_comb = p3_sum__1206_comb + p3_sum__1207_comb;
  assign p3_sum__1052_comb = p3_sum__1192_comb + p3_sum__1193_comb;
  assign p3_sum__1038_comb = p3_sum__1164_comb + p3_sum__1165_comb;
  assign p3_sum__1031_comb = p3_sum__1150_comb + p3_sum__1151_comb;
  assign p3_sum__1024_comb = p3_sum__1136_comb + p3_sum__1137_comb;
  assign p3_umul_29018_NarrowedMult__comb = umul24b_24b_x_7b(p2_add_86565, 7'h5b);
  assign p3_umul_29020_NarrowedMult__comb = umul24b_24b_x_7b(p2_add_86566, 7'h5b);
  assign p3_umul_29022_NarrowedMult__comb = umul24b_24b_x_7b(p2_add_86567, 7'h5b);
  assign p3_umul_29026_NarrowedMult__comb = umul24b_24b_x_7b(p2_add_86570, 7'h5b);
  assign p3_umul_29028_NarrowedMult__comb = umul24b_24b_x_7b(p2_add_86571, 7'h5b);
  assign p3_umul_29030_NarrowedMult__comb = umul24b_24b_x_7b(p2_add_86572, 7'h5b);
  assign p3_add_87209_comb = p2_sum__1079 + 25'h000_0001;
  assign p3_add_87210_comb = p3_sum__1072_comb + 25'h000_0001;
  assign p3_add_87211_comb = p3_sum__1065_comb + 25'h000_0001;
  assign p3_add_87212_comb = p3_sum__1058_comb + 25'h000_0001;
  assign p3_add_87213_comb = p3_sum__1044_comb + 25'h000_0001;
  assign p3_add_87214_comb = p3_sum__1037_comb + 25'h000_0001;
  assign p3_add_87215_comb = p3_sum__1030_comb + 25'h000_0001;
  assign p3_add_87216_comb = p2_add_86576 + p2_add_86577;
  assign p3_add_87217_comb = p3_add_87140_comb + p3_add_87141_comb;
  assign p3_add_87218_comb = p3_add_87142_comb + p3_add_87143_comb;
  assign p3_add_87219_comb = p3_add_87144_comb + p3_add_87145_comb;
  assign p3_add_87220_comb = p3_add_87146_comb + p3_add_87147_comb;
  assign p3_add_87221_comb = p3_add_87148_comb + p3_add_87149_comb;
  assign p3_add_87222_comb = p3_add_87150_comb + p3_add_87151_comb;
  assign p3_add_87223_comb = p2_sum__1077 + 25'h000_0001;
  assign p3_add_87224_comb = p3_sum__1070_comb + 25'h000_0001;
  assign p3_add_87225_comb = p3_sum__1063_comb + 25'h000_0001;
  assign p3_add_87226_comb = p3_sum__1056_comb + 25'h000_0001;
  assign p3_add_87227_comb = p3_sum__1042_comb + 25'h000_0001;
  assign p3_add_87228_comb = p3_sum__1035_comb + 25'h000_0001;
  assign p3_add_87229_comb = p3_sum__1028_comb + 25'h000_0001;
  assign p3_add_87230_comb = p2_sum__1075 + 25'h000_0001;
  assign p3_add_87231_comb = p3_sum__1068_comb + 25'h000_0001;
  assign p3_add_87232_comb = p3_sum__1061_comb + 25'h000_0001;
  assign p3_add_87233_comb = p3_sum__1054_comb + 25'h000_0001;
  assign p3_add_87234_comb = p3_sum__1040_comb + 25'h000_0001;
  assign p3_add_87235_comb = p3_sum__1033_comb + 25'h000_0001;
  assign p3_add_87236_comb = p3_sum__1026_comb + 25'h000_0001;
  assign p3_add_87237_comb = p2_add_86602 + p2_add_86603;
  assign p3_add_87238_comb = p3_add_87178_comb + p3_add_87179_comb;
  assign p3_add_87239_comb = p3_add_87180_comb + p3_add_87181_comb;
  assign p3_add_87240_comb = p3_add_87182_comb + p3_add_87183_comb;
  assign p3_add_87241_comb = p3_add_87184_comb + p3_add_87185_comb;
  assign p3_add_87242_comb = p3_add_87186_comb + p3_add_87187_comb;
  assign p3_add_87243_comb = p3_add_87188_comb + p3_add_87189_comb;
  assign p3_add_87244_comb = p2_sum__1073 + 25'h000_0001;
  assign p3_add_87245_comb = p3_sum__1066_comb + 25'h000_0001;
  assign p3_add_87246_comb = p3_sum__1059_comb + 25'h000_0001;
  assign p3_add_87247_comb = p3_sum__1052_comb + 25'h000_0001;
  assign p3_add_87248_comb = p3_sum__1038_comb + 25'h000_0001;
  assign p3_add_87249_comb = p3_sum__1031_comb + 25'h000_0001;
  assign p3_add_87250_comb = p3_sum__1024_comb + 25'h000_0001;
  assign p3_bit_slice_87251_comb = p3_umul_29018_NarrowedMult__comb[23:7];
  assign p3_bit_slice_87252_comb = p3_umul_29020_NarrowedMult__comb[23:7];
  assign p3_bit_slice_87253_comb = p3_umul_29022_NarrowedMult__comb[23:7];
  assign p3_bit_slice_87254_comb = p3_umul_29026_NarrowedMult__comb[23:7];
  assign p3_bit_slice_87255_comb = p3_umul_29028_NarrowedMult__comb[23:7];
  assign p3_bit_slice_87256_comb = p3_umul_29030_NarrowedMult__comb[23:7];
  assign p3_bit_slice_87257_comb = p3_add_87209_comb[24:8];
  assign p3_bit_slice_87258_comb = p3_add_87210_comb[24:8];
  assign p3_bit_slice_87259_comb = p3_add_87211_comb[24:8];
  assign p3_bit_slice_87260_comb = p3_add_87212_comb[24:8];
  assign p3_bit_slice_87261_comb = p2_add_86611[24:8];
  assign p3_bit_slice_87262_comb = p3_add_87213_comb[24:8];
  assign p3_bit_slice_87263_comb = p3_add_87214_comb[24:8];
  assign p3_bit_slice_87264_comb = p3_add_87215_comb[24:8];
  assign p3_bit_slice_87265_comb = p3_add_87216_comb[23:7];
  assign p3_bit_slice_87266_comb = p3_add_87217_comb[23:7];
  assign p3_bit_slice_87267_comb = p3_add_87218_comb[23:7];
  assign p3_bit_slice_87268_comb = p3_add_87219_comb[23:7];
  assign p3_bit_slice_87269_comb = p2_add_86612[23:7];
  assign p3_bit_slice_87270_comb = p3_add_87220_comb[23:7];
  assign p3_bit_slice_87271_comb = p3_add_87221_comb[23:7];
  assign p3_bit_slice_87272_comb = p3_add_87222_comb[23:7];
  assign p3_bit_slice_87273_comb = p3_add_87223_comb[24:8];
  assign p3_bit_slice_87274_comb = p3_add_87224_comb[24:8];
  assign p3_bit_slice_87275_comb = p3_add_87225_comb[24:8];
  assign p3_bit_slice_87276_comb = p3_add_87226_comb[24:8];
  assign p3_bit_slice_87277_comb = p2_add_86613[24:8];
  assign p3_bit_slice_87278_comb = p3_add_87227_comb[24:8];
  assign p3_bit_slice_87279_comb = p3_add_87228_comb[24:8];
  assign p3_bit_slice_87280_comb = p3_add_87229_comb[24:8];
  assign p3_bit_slice_87281_comb = p2_add_86615[24:8];
  assign p3_bit_slice_87282_comb = p2_add_86616[24:8];
  assign p3_bit_slice_87283_comb = p2_add_86617[24:8];
  assign p3_bit_slice_87284_comb = p2_add_86619[24:8];
  assign p3_bit_slice_87285_comb = p2_add_86620[24:8];
  assign p3_bit_slice_87286_comb = p2_add_86621[24:8];
  assign p3_bit_slice_87287_comb = p3_add_87230_comb[24:8];
  assign p3_bit_slice_87288_comb = p3_add_87231_comb[24:8];
  assign p3_bit_slice_87289_comb = p3_add_87232_comb[24:8];
  assign p3_bit_slice_87290_comb = p3_add_87233_comb[24:8];
  assign p3_bit_slice_87291_comb = p2_add_86622[24:8];
  assign p3_bit_slice_87292_comb = p3_add_87234_comb[24:8];
  assign p3_bit_slice_87293_comb = p3_add_87235_comb[24:8];
  assign p3_bit_slice_87294_comb = p3_add_87236_comb[24:8];
  assign p3_bit_slice_87295_comb = p3_add_87237_comb[23:7];
  assign p3_bit_slice_87296_comb = p3_add_87238_comb[23:7];
  assign p3_bit_slice_87297_comb = p3_add_87239_comb[23:7];
  assign p3_bit_slice_87298_comb = p3_add_87240_comb[23:7];
  assign p3_bit_slice_87299_comb = p2_add_86623[23:7];
  assign p3_bit_slice_87300_comb = p3_add_87241_comb[23:7];
  assign p3_bit_slice_87301_comb = p3_add_87242_comb[23:7];
  assign p3_bit_slice_87302_comb = p3_add_87243_comb[23:7];
  assign p3_bit_slice_87303_comb = p3_add_87244_comb[24:8];
  assign p3_bit_slice_87304_comb = p3_add_87245_comb[24:8];
  assign p3_bit_slice_87305_comb = p3_add_87246_comb[24:8];
  assign p3_bit_slice_87306_comb = p3_add_87247_comb[24:8];
  assign p3_bit_slice_87307_comb = p2_add_86624[24:8];
  assign p3_bit_slice_87308_comb = p3_add_87248_comb[24:8];
  assign p3_bit_slice_87309_comb = p3_add_87249_comb[24:8];
  assign p3_bit_slice_87310_comb = p3_add_87250_comb[24:8];
  assign p3_add_87439_comb = {{1{p2_bit_slice_86625[16]}}, p2_bit_slice_86625} + 18'h0_0001;
  assign p3_add_87440_comb = {{1{p3_bit_slice_87251_comb[16]}}, p3_bit_slice_87251_comb} + 18'h0_0001;
  assign p3_add_87441_comb = {{1{p3_bit_slice_87252_comb[16]}}, p3_bit_slice_87252_comb} + 18'h0_0001;
  assign p3_add_87442_comb = {{1{p3_bit_slice_87253_comb[16]}}, p3_bit_slice_87253_comb} + 18'h0_0001;
  assign p3_add_87443_comb = {{1{p2_bit_slice_86626[16]}}, p2_bit_slice_86626} + 18'h0_0001;
  assign p3_add_87444_comb = {{1{p3_bit_slice_87254_comb[16]}}, p3_bit_slice_87254_comb} + 18'h0_0001;
  assign p3_add_87445_comb = {{1{p3_bit_slice_87255_comb[16]}}, p3_bit_slice_87255_comb} + 18'h0_0001;
  assign p3_add_87446_comb = {{1{p3_bit_slice_87256_comb[16]}}, p3_bit_slice_87256_comb} + 18'h0_0001;
  assign p3_add_87447_comb = {{1{p3_bit_slice_87257_comb[16]}}, p3_bit_slice_87257_comb} + 18'h0_0001;
  assign p3_add_87448_comb = {{1{p3_bit_slice_87258_comb[16]}}, p3_bit_slice_87258_comb} + 18'h0_0001;
  assign p3_add_87449_comb = {{1{p3_bit_slice_87259_comb[16]}}, p3_bit_slice_87259_comb} + 18'h0_0001;
  assign p3_add_87450_comb = {{1{p3_bit_slice_87260_comb[16]}}, p3_bit_slice_87260_comb} + 18'h0_0001;
  assign p3_add_87451_comb = {{1{p3_bit_slice_87261_comb[16]}}, p3_bit_slice_87261_comb} + 18'h0_0001;
  assign p3_add_87452_comb = {{1{p3_bit_slice_87262_comb[16]}}, p3_bit_slice_87262_comb} + 18'h0_0001;
  assign p3_add_87453_comb = {{1{p3_bit_slice_87263_comb[16]}}, p3_bit_slice_87263_comb} + 18'h0_0001;
  assign p3_add_87454_comb = {{1{p3_bit_slice_87264_comb[16]}}, p3_bit_slice_87264_comb} + 18'h0_0001;
  assign p3_add_87455_comb = {{1{p3_bit_slice_87265_comb[16]}}, p3_bit_slice_87265_comb} + 18'h0_0001;
  assign p3_add_87456_comb = {{1{p3_bit_slice_87266_comb[16]}}, p3_bit_slice_87266_comb} + 18'h0_0001;
  assign p3_add_87457_comb = {{1{p3_bit_slice_87267_comb[16]}}, p3_bit_slice_87267_comb} + 18'h0_0001;
  assign p3_add_87458_comb = {{1{p3_bit_slice_87268_comb[16]}}, p3_bit_slice_87268_comb} + 18'h0_0001;
  assign p3_add_87459_comb = {{1{p3_bit_slice_87269_comb[16]}}, p3_bit_slice_87269_comb} + 18'h0_0001;
  assign p3_add_87460_comb = {{1{p3_bit_slice_87270_comb[16]}}, p3_bit_slice_87270_comb} + 18'h0_0001;
  assign p3_add_87461_comb = {{1{p3_bit_slice_87271_comb[16]}}, p3_bit_slice_87271_comb} + 18'h0_0001;
  assign p3_add_87462_comb = {{1{p3_bit_slice_87272_comb[16]}}, p3_bit_slice_87272_comb} + 18'h0_0001;
  assign p3_add_87463_comb = {{1{p3_bit_slice_87273_comb[16]}}, p3_bit_slice_87273_comb} + 18'h0_0001;
  assign p3_add_87464_comb = {{1{p3_bit_slice_87274_comb[16]}}, p3_bit_slice_87274_comb} + 18'h0_0001;
  assign p3_add_87465_comb = {{1{p3_bit_slice_87275_comb[16]}}, p3_bit_slice_87275_comb} + 18'h0_0001;
  assign p3_add_87466_comb = {{1{p3_bit_slice_87276_comb[16]}}, p3_bit_slice_87276_comb} + 18'h0_0001;
  assign p3_add_87467_comb = {{1{p3_bit_slice_87277_comb[16]}}, p3_bit_slice_87277_comb} + 18'h0_0001;
  assign p3_add_87468_comb = {{1{p3_bit_slice_87278_comb[16]}}, p3_bit_slice_87278_comb} + 18'h0_0001;
  assign p3_add_87469_comb = {{1{p3_bit_slice_87279_comb[16]}}, p3_bit_slice_87279_comb} + 18'h0_0001;
  assign p3_add_87470_comb = {{1{p3_bit_slice_87280_comb[16]}}, p3_bit_slice_87280_comb} + 18'h0_0001;
  assign p3_add_87471_comb = {{1{p2_bit_slice_86627[16]}}, p2_bit_slice_86627} + 18'h0_0001;
  assign p3_add_87472_comb = {{1{p3_bit_slice_87281_comb[16]}}, p3_bit_slice_87281_comb} + 18'h0_0001;
  assign p3_add_87473_comb = {{1{p3_bit_slice_87282_comb[16]}}, p3_bit_slice_87282_comb} + 18'h0_0001;
  assign p3_add_87474_comb = {{1{p3_bit_slice_87283_comb[16]}}, p3_bit_slice_87283_comb} + 18'h0_0001;
  assign p3_add_87475_comb = {{1{p2_bit_slice_86628[16]}}, p2_bit_slice_86628} + 18'h0_0001;
  assign p3_add_87476_comb = {{1{p3_bit_slice_87284_comb[16]}}, p3_bit_slice_87284_comb} + 18'h0_0001;
  assign p3_add_87477_comb = {{1{p3_bit_slice_87285_comb[16]}}, p3_bit_slice_87285_comb} + 18'h0_0001;
  assign p3_add_87478_comb = {{1{p3_bit_slice_87286_comb[16]}}, p3_bit_slice_87286_comb} + 18'h0_0001;
  assign p3_add_87479_comb = {{1{p3_bit_slice_87287_comb[16]}}, p3_bit_slice_87287_comb} + 18'h0_0001;
  assign p3_add_87480_comb = {{1{p3_bit_slice_87288_comb[16]}}, p3_bit_slice_87288_comb} + 18'h0_0001;
  assign p3_add_87481_comb = {{1{p3_bit_slice_87289_comb[16]}}, p3_bit_slice_87289_comb} + 18'h0_0001;
  assign p3_add_87482_comb = {{1{p3_bit_slice_87290_comb[16]}}, p3_bit_slice_87290_comb} + 18'h0_0001;
  assign p3_add_87483_comb = {{1{p3_bit_slice_87291_comb[16]}}, p3_bit_slice_87291_comb} + 18'h0_0001;
  assign p3_add_87484_comb = {{1{p3_bit_slice_87292_comb[16]}}, p3_bit_slice_87292_comb} + 18'h0_0001;
  assign p3_add_87485_comb = {{1{p3_bit_slice_87293_comb[16]}}, p3_bit_slice_87293_comb} + 18'h0_0001;
  assign p3_add_87486_comb = {{1{p3_bit_slice_87294_comb[16]}}, p3_bit_slice_87294_comb} + 18'h0_0001;
  assign p3_add_87487_comb = {{1{p3_bit_slice_87295_comb[16]}}, p3_bit_slice_87295_comb} + 18'h0_0001;
  assign p3_add_87488_comb = {{1{p3_bit_slice_87296_comb[16]}}, p3_bit_slice_87296_comb} + 18'h0_0001;
  assign p3_add_87489_comb = {{1{p3_bit_slice_87297_comb[16]}}, p3_bit_slice_87297_comb} + 18'h0_0001;
  assign p3_add_87490_comb = {{1{p3_bit_slice_87298_comb[16]}}, p3_bit_slice_87298_comb} + 18'h0_0001;
  assign p3_add_87491_comb = {{1{p3_bit_slice_87299_comb[16]}}, p3_bit_slice_87299_comb} + 18'h0_0001;
  assign p3_add_87492_comb = {{1{p3_bit_slice_87300_comb[16]}}, p3_bit_slice_87300_comb} + 18'h0_0001;
  assign p3_add_87493_comb = {{1{p3_bit_slice_87301_comb[16]}}, p3_bit_slice_87301_comb} + 18'h0_0001;
  assign p3_add_87494_comb = {{1{p3_bit_slice_87302_comb[16]}}, p3_bit_slice_87302_comb} + 18'h0_0001;
  assign p3_add_87495_comb = {{1{p3_bit_slice_87303_comb[16]}}, p3_bit_slice_87303_comb} + 18'h0_0001;
  assign p3_add_87496_comb = {{1{p3_bit_slice_87304_comb[16]}}, p3_bit_slice_87304_comb} + 18'h0_0001;
  assign p3_add_87497_comb = {{1{p3_bit_slice_87305_comb[16]}}, p3_bit_slice_87305_comb} + 18'h0_0001;
  assign p3_add_87498_comb = {{1{p3_bit_slice_87306_comb[16]}}, p3_bit_slice_87306_comb} + 18'h0_0001;
  assign p3_add_87499_comb = {{1{p3_bit_slice_87307_comb[16]}}, p3_bit_slice_87307_comb} + 18'h0_0001;
  assign p3_add_87500_comb = {{1{p3_bit_slice_87308_comb[16]}}, p3_bit_slice_87308_comb} + 18'h0_0001;
  assign p3_add_87501_comb = {{1{p3_bit_slice_87309_comb[16]}}, p3_bit_slice_87309_comb} + 18'h0_0001;
  assign p3_add_87502_comb = {{1{p3_bit_slice_87310_comb[16]}}, p3_bit_slice_87310_comb} + 18'h0_0001;
  assign p3_bit_slice_87503_comb = p3_add_87439_comb[17:8];
  assign p3_bit_slice_87504_comb = p3_add_87440_comb[17:8];
  assign p3_bit_slice_87505_comb = p3_add_87441_comb[17:8];
  assign p3_bit_slice_87506_comb = p3_add_87442_comb[17:8];
  assign p3_bit_slice_87507_comb = p3_add_87443_comb[17:8];
  assign p3_bit_slice_87508_comb = p3_add_87444_comb[17:8];
  assign p3_bit_slice_87509_comb = p3_add_87445_comb[17:8];
  assign p3_bit_slice_87510_comb = p3_add_87446_comb[17:8];
  assign p3_bit_slice_87511_comb = p3_add_87447_comb[17:8];
  assign p3_bit_slice_87512_comb = p3_add_87448_comb[17:8];
  assign p3_bit_slice_87513_comb = p3_add_87449_comb[17:8];
  assign p3_bit_slice_87514_comb = p3_add_87450_comb[17:8];
  assign p3_bit_slice_87515_comb = p3_add_87451_comb[17:8];
  assign p3_bit_slice_87516_comb = p3_add_87452_comb[17:8];
  assign p3_bit_slice_87517_comb = p3_add_87453_comb[17:8];
  assign p3_bit_slice_87518_comb = p3_add_87454_comb[17:8];
  assign p3_bit_slice_87519_comb = p3_add_87455_comb[17:8];
  assign p3_bit_slice_87520_comb = p3_add_87456_comb[17:8];
  assign p3_bit_slice_87521_comb = p3_add_87457_comb[17:8];
  assign p3_bit_slice_87522_comb = p3_add_87458_comb[17:8];
  assign p3_bit_slice_87523_comb = p3_add_87459_comb[17:8];
  assign p3_bit_slice_87524_comb = p3_add_87460_comb[17:8];
  assign p3_bit_slice_87525_comb = p3_add_87461_comb[17:8];
  assign p3_bit_slice_87526_comb = p3_add_87462_comb[17:8];
  assign p3_bit_slice_87527_comb = p3_add_87463_comb[17:8];
  assign p3_bit_slice_87528_comb = p3_add_87464_comb[17:8];
  assign p3_bit_slice_87529_comb = p3_add_87465_comb[17:8];
  assign p3_bit_slice_87530_comb = p3_add_87466_comb[17:8];
  assign p3_bit_slice_87531_comb = p3_add_87467_comb[17:8];
  assign p3_bit_slice_87532_comb = p3_add_87468_comb[17:8];
  assign p3_bit_slice_87533_comb = p3_add_87469_comb[17:8];
  assign p3_bit_slice_87534_comb = p3_add_87470_comb[17:8];
  assign p3_bit_slice_87535_comb = p3_add_87471_comb[17:8];
  assign p3_bit_slice_87536_comb = p3_add_87472_comb[17:8];
  assign p3_bit_slice_87537_comb = p3_add_87473_comb[17:8];
  assign p3_bit_slice_87538_comb = p3_add_87474_comb[17:8];
  assign p3_bit_slice_87539_comb = p3_add_87475_comb[17:8];
  assign p3_bit_slice_87540_comb = p3_add_87476_comb[17:8];
  assign p3_bit_slice_87541_comb = p3_add_87477_comb[17:8];
  assign p3_bit_slice_87542_comb = p3_add_87478_comb[17:8];
  assign p3_bit_slice_87543_comb = p3_add_87479_comb[17:8];
  assign p3_bit_slice_87544_comb = p3_add_87480_comb[17:8];
  assign p3_bit_slice_87545_comb = p3_add_87481_comb[17:8];
  assign p3_bit_slice_87546_comb = p3_add_87482_comb[17:8];
  assign p3_bit_slice_87547_comb = p3_add_87483_comb[17:8];
  assign p3_bit_slice_87548_comb = p3_add_87484_comb[17:8];
  assign p3_bit_slice_87549_comb = p3_add_87485_comb[17:8];
  assign p3_bit_slice_87550_comb = p3_add_87486_comb[17:8];
  assign p3_bit_slice_87551_comb = p3_add_87487_comb[17:8];
  assign p3_bit_slice_87552_comb = p3_add_87488_comb[17:8];
  assign p3_bit_slice_87553_comb = p3_add_87489_comb[17:8];
  assign p3_bit_slice_87554_comb = p3_add_87490_comb[17:8];
  assign p3_bit_slice_87555_comb = p3_add_87491_comb[17:8];
  assign p3_bit_slice_87556_comb = p3_add_87492_comb[17:8];
  assign p3_bit_slice_87557_comb = p3_add_87493_comb[17:8];
  assign p3_bit_slice_87558_comb = p3_add_87494_comb[17:8];
  assign p3_bit_slice_87559_comb = p3_add_87495_comb[17:8];
  assign p3_bit_slice_87560_comb = p3_add_87496_comb[17:8];
  assign p3_bit_slice_87561_comb = p3_add_87497_comb[17:8];
  assign p3_bit_slice_87562_comb = p3_add_87498_comb[17:8];
  assign p3_bit_slice_87563_comb = p3_add_87499_comb[17:8];
  assign p3_bit_slice_87564_comb = p3_add_87500_comb[17:8];
  assign p3_bit_slice_87565_comb = p3_add_87501_comb[17:8];
  assign p3_bit_slice_87566_comb = p3_add_87502_comb[17:8];
  assign p3_add_87695_comb = {{1{p3_bit_slice_87503_comb[9]}}, p3_bit_slice_87503_comb} + 11'h001;
  assign p3_add_87697_comb = {{1{p3_bit_slice_87504_comb[9]}}, p3_bit_slice_87504_comb} + 11'h001;
  assign p3_add_87699_comb = {{1{p3_bit_slice_87505_comb[9]}}, p3_bit_slice_87505_comb} + 11'h001;
  assign p3_add_87701_comb = {{1{p3_bit_slice_87506_comb[9]}}, p3_bit_slice_87506_comb} + 11'h001;
  assign p3_add_87703_comb = {{1{p3_bit_slice_87507_comb[9]}}, p3_bit_slice_87507_comb} + 11'h001;
  assign p3_add_87705_comb = {{1{p3_bit_slice_87508_comb[9]}}, p3_bit_slice_87508_comb} + 11'h001;
  assign p3_add_87707_comb = {{1{p3_bit_slice_87509_comb[9]}}, p3_bit_slice_87509_comb} + 11'h001;
  assign p3_add_87709_comb = {{1{p3_bit_slice_87510_comb[9]}}, p3_bit_slice_87510_comb} + 11'h001;
  assign p3_add_87711_comb = {{1{p3_bit_slice_87511_comb[9]}}, p3_bit_slice_87511_comb} + 11'h001;
  assign p3_add_87713_comb = {{1{p3_bit_slice_87512_comb[9]}}, p3_bit_slice_87512_comb} + 11'h001;
  assign p3_add_87715_comb = {{1{p3_bit_slice_87513_comb[9]}}, p3_bit_slice_87513_comb} + 11'h001;
  assign p3_add_87717_comb = {{1{p3_bit_slice_87514_comb[9]}}, p3_bit_slice_87514_comb} + 11'h001;
  assign p3_add_87719_comb = {{1{p3_bit_slice_87515_comb[9]}}, p3_bit_slice_87515_comb} + 11'h001;
  assign p3_add_87721_comb = {{1{p3_bit_slice_87516_comb[9]}}, p3_bit_slice_87516_comb} + 11'h001;
  assign p3_add_87723_comb = {{1{p3_bit_slice_87517_comb[9]}}, p3_bit_slice_87517_comb} + 11'h001;
  assign p3_add_87725_comb = {{1{p3_bit_slice_87518_comb[9]}}, p3_bit_slice_87518_comb} + 11'h001;
  assign p3_add_87727_comb = {{1{p3_bit_slice_87519_comb[9]}}, p3_bit_slice_87519_comb} + 11'h001;
  assign p3_add_87729_comb = {{1{p3_bit_slice_87520_comb[9]}}, p3_bit_slice_87520_comb} + 11'h001;
  assign p3_add_87731_comb = {{1{p3_bit_slice_87521_comb[9]}}, p3_bit_slice_87521_comb} + 11'h001;
  assign p3_add_87733_comb = {{1{p3_bit_slice_87522_comb[9]}}, p3_bit_slice_87522_comb} + 11'h001;
  assign p3_add_87735_comb = {{1{p3_bit_slice_87523_comb[9]}}, p3_bit_slice_87523_comb} + 11'h001;
  assign p3_add_87737_comb = {{1{p3_bit_slice_87524_comb[9]}}, p3_bit_slice_87524_comb} + 11'h001;
  assign p3_add_87739_comb = {{1{p3_bit_slice_87525_comb[9]}}, p3_bit_slice_87525_comb} + 11'h001;
  assign p3_add_87741_comb = {{1{p3_bit_slice_87526_comb[9]}}, p3_bit_slice_87526_comb} + 11'h001;
  assign p3_add_87743_comb = {{1{p3_bit_slice_87527_comb[9]}}, p3_bit_slice_87527_comb} + 11'h001;
  assign p3_add_87745_comb = {{1{p3_bit_slice_87528_comb[9]}}, p3_bit_slice_87528_comb} + 11'h001;
  assign p3_add_87747_comb = {{1{p3_bit_slice_87529_comb[9]}}, p3_bit_slice_87529_comb} + 11'h001;
  assign p3_add_87749_comb = {{1{p3_bit_slice_87530_comb[9]}}, p3_bit_slice_87530_comb} + 11'h001;
  assign p3_add_87751_comb = {{1{p3_bit_slice_87531_comb[9]}}, p3_bit_slice_87531_comb} + 11'h001;
  assign p3_add_87753_comb = {{1{p3_bit_slice_87532_comb[9]}}, p3_bit_slice_87532_comb} + 11'h001;
  assign p3_add_87755_comb = {{1{p3_bit_slice_87533_comb[9]}}, p3_bit_slice_87533_comb} + 11'h001;
  assign p3_add_87757_comb = {{1{p3_bit_slice_87534_comb[9]}}, p3_bit_slice_87534_comb} + 11'h001;
  assign p3_add_87759_comb = {{1{p3_bit_slice_87535_comb[9]}}, p3_bit_slice_87535_comb} + 11'h001;
  assign p3_add_87761_comb = {{1{p3_bit_slice_87536_comb[9]}}, p3_bit_slice_87536_comb} + 11'h001;
  assign p3_add_87763_comb = {{1{p3_bit_slice_87537_comb[9]}}, p3_bit_slice_87537_comb} + 11'h001;
  assign p3_add_87765_comb = {{1{p3_bit_slice_87538_comb[9]}}, p3_bit_slice_87538_comb} + 11'h001;
  assign p3_add_87767_comb = {{1{p3_bit_slice_87539_comb[9]}}, p3_bit_slice_87539_comb} + 11'h001;
  assign p3_add_87769_comb = {{1{p3_bit_slice_87540_comb[9]}}, p3_bit_slice_87540_comb} + 11'h001;
  assign p3_add_87771_comb = {{1{p3_bit_slice_87541_comb[9]}}, p3_bit_slice_87541_comb} + 11'h001;
  assign p3_add_87773_comb = {{1{p3_bit_slice_87542_comb[9]}}, p3_bit_slice_87542_comb} + 11'h001;
  assign p3_add_87775_comb = {{1{p3_bit_slice_87543_comb[9]}}, p3_bit_slice_87543_comb} + 11'h001;
  assign p3_add_87777_comb = {{1{p3_bit_slice_87544_comb[9]}}, p3_bit_slice_87544_comb} + 11'h001;
  assign p3_add_87779_comb = {{1{p3_bit_slice_87545_comb[9]}}, p3_bit_slice_87545_comb} + 11'h001;
  assign p3_add_87781_comb = {{1{p3_bit_slice_87546_comb[9]}}, p3_bit_slice_87546_comb} + 11'h001;
  assign p3_add_87783_comb = {{1{p3_bit_slice_87547_comb[9]}}, p3_bit_slice_87547_comb} + 11'h001;
  assign p3_add_87785_comb = {{1{p3_bit_slice_87548_comb[9]}}, p3_bit_slice_87548_comb} + 11'h001;
  assign p3_add_87787_comb = {{1{p3_bit_slice_87549_comb[9]}}, p3_bit_slice_87549_comb} + 11'h001;
  assign p3_add_87789_comb = {{1{p3_bit_slice_87550_comb[9]}}, p3_bit_slice_87550_comb} + 11'h001;
  assign p3_add_87791_comb = {{1{p3_bit_slice_87551_comb[9]}}, p3_bit_slice_87551_comb} + 11'h001;
  assign p3_add_87793_comb = {{1{p3_bit_slice_87552_comb[9]}}, p3_bit_slice_87552_comb} + 11'h001;
  assign p3_add_87795_comb = {{1{p3_bit_slice_87553_comb[9]}}, p3_bit_slice_87553_comb} + 11'h001;
  assign p3_add_87797_comb = {{1{p3_bit_slice_87554_comb[9]}}, p3_bit_slice_87554_comb} + 11'h001;
  assign p3_add_87799_comb = {{1{p3_bit_slice_87555_comb[9]}}, p3_bit_slice_87555_comb} + 11'h001;
  assign p3_add_87801_comb = {{1{p3_bit_slice_87556_comb[9]}}, p3_bit_slice_87556_comb} + 11'h001;
  assign p3_add_87803_comb = {{1{p3_bit_slice_87557_comb[9]}}, p3_bit_slice_87557_comb} + 11'h001;
  assign p3_add_87805_comb = {{1{p3_bit_slice_87558_comb[9]}}, p3_bit_slice_87558_comb} + 11'h001;
  assign p3_add_87807_comb = {{1{p3_bit_slice_87559_comb[9]}}, p3_bit_slice_87559_comb} + 11'h001;
  assign p3_add_87809_comb = {{1{p3_bit_slice_87560_comb[9]}}, p3_bit_slice_87560_comb} + 11'h001;
  assign p3_add_87811_comb = {{1{p3_bit_slice_87561_comb[9]}}, p3_bit_slice_87561_comb} + 11'h001;
  assign p3_add_87813_comb = {{1{p3_bit_slice_87562_comb[9]}}, p3_bit_slice_87562_comb} + 11'h001;
  assign p3_add_87815_comb = {{1{p3_bit_slice_87563_comb[9]}}, p3_bit_slice_87563_comb} + 11'h001;
  assign p3_add_87817_comb = {{1{p3_bit_slice_87564_comb[9]}}, p3_bit_slice_87564_comb} + 11'h001;
  assign p3_add_87819_comb = {{1{p3_bit_slice_87565_comb[9]}}, p3_bit_slice_87565_comb} + 11'h001;
  assign p3_add_87821_comb = {{1{p3_bit_slice_87566_comb[9]}}, p3_bit_slice_87566_comb} + 11'h001;
  assign p3_concat_87823_comb = {p3_add_87695_comb, p3_add_87439_comb[7:1]};
  assign p3_concat_87826_comb = {p3_add_87697_comb, p3_add_87440_comb[7:1]};
  assign p3_concat_87829_comb = {p3_add_87699_comb, p3_add_87441_comb[7:1]};
  assign p3_concat_87832_comb = {p3_add_87701_comb, p3_add_87442_comb[7:1]};
  assign p3_concat_87835_comb = {p3_add_87703_comb, p3_add_87443_comb[7:1]};
  assign p3_concat_87838_comb = {p3_add_87705_comb, p3_add_87444_comb[7:1]};
  assign p3_concat_87841_comb = {p3_add_87707_comb, p3_add_87445_comb[7:1]};
  assign p3_concat_87844_comb = {p3_add_87709_comb, p3_add_87446_comb[7:1]};
  assign p3_concat_87847_comb = {p3_add_87711_comb, p3_add_87447_comb[7:1]};
  assign p3_concat_87850_comb = {p3_add_87713_comb, p3_add_87448_comb[7:1]};
  assign p3_concat_87853_comb = {p3_add_87715_comb, p3_add_87449_comb[7:1]};
  assign p3_concat_87856_comb = {p3_add_87717_comb, p3_add_87450_comb[7:1]};
  assign p3_concat_87859_comb = {p3_add_87719_comb, p3_add_87451_comb[7:1]};
  assign p3_concat_87862_comb = {p3_add_87721_comb, p3_add_87452_comb[7:1]};
  assign p3_concat_87865_comb = {p3_add_87723_comb, p3_add_87453_comb[7:1]};
  assign p3_concat_87868_comb = {p3_add_87725_comb, p3_add_87454_comb[7:1]};
  assign p3_concat_87871_comb = {p3_add_87727_comb, p3_add_87455_comb[7:1]};
  assign p3_concat_87874_comb = {p3_add_87729_comb, p3_add_87456_comb[7:1]};
  assign p3_concat_87877_comb = {p3_add_87731_comb, p3_add_87457_comb[7:1]};
  assign p3_concat_87880_comb = {p3_add_87733_comb, p3_add_87458_comb[7:1]};
  assign p3_concat_87883_comb = {p3_add_87735_comb, p3_add_87459_comb[7:1]};
  assign p3_concat_87886_comb = {p3_add_87737_comb, p3_add_87460_comb[7:1]};
  assign p3_concat_87889_comb = {p3_add_87739_comb, p3_add_87461_comb[7:1]};
  assign p3_concat_87892_comb = {p3_add_87741_comb, p3_add_87462_comb[7:1]};
  assign p3_concat_87895_comb = {p3_add_87743_comb, p3_add_87463_comb[7:1]};
  assign p3_concat_87898_comb = {p3_add_87745_comb, p3_add_87464_comb[7:1]};
  assign p3_concat_87901_comb = {p3_add_87747_comb, p3_add_87465_comb[7:1]};
  assign p3_concat_87904_comb = {p3_add_87749_comb, p3_add_87466_comb[7:1]};
  assign p3_concat_87907_comb = {p3_add_87751_comb, p3_add_87467_comb[7:1]};
  assign p3_concat_87910_comb = {p3_add_87753_comb, p3_add_87468_comb[7:1]};
  assign p3_concat_87913_comb = {p3_add_87755_comb, p3_add_87469_comb[7:1]};
  assign p3_concat_87916_comb = {p3_add_87757_comb, p3_add_87470_comb[7:1]};
  assign p3_concat_87919_comb = {p3_add_87759_comb, p3_add_87471_comb[7:1]};
  assign p3_concat_87922_comb = {p3_add_87761_comb, p3_add_87472_comb[7:1]};
  assign p3_concat_87925_comb = {p3_add_87763_comb, p3_add_87473_comb[7:1]};
  assign p3_concat_87928_comb = {p3_add_87765_comb, p3_add_87474_comb[7:1]};
  assign p3_concat_87931_comb = {p3_add_87767_comb, p3_add_87475_comb[7:1]};
  assign p3_concat_87934_comb = {p3_add_87769_comb, p3_add_87476_comb[7:1]};
  assign p3_concat_87937_comb = {p3_add_87771_comb, p3_add_87477_comb[7:1]};
  assign p3_concat_87940_comb = {p3_add_87773_comb, p3_add_87478_comb[7:1]};
  assign p3_concat_87943_comb = {p3_add_87775_comb, p3_add_87479_comb[7:1]};
  assign p3_concat_87946_comb = {p3_add_87777_comb, p3_add_87480_comb[7:1]};
  assign p3_concat_87949_comb = {p3_add_87779_comb, p3_add_87481_comb[7:1]};
  assign p3_concat_87952_comb = {p3_add_87781_comb, p3_add_87482_comb[7:1]};
  assign p3_concat_87955_comb = {p3_add_87783_comb, p3_add_87483_comb[7:1]};
  assign p3_concat_87958_comb = {p3_add_87785_comb, p3_add_87484_comb[7:1]};
  assign p3_concat_87961_comb = {p3_add_87787_comb, p3_add_87485_comb[7:1]};
  assign p3_concat_87964_comb = {p3_add_87789_comb, p3_add_87486_comb[7:1]};
  assign p3_concat_87967_comb = {p3_add_87791_comb, p3_add_87487_comb[7:1]};
  assign p3_concat_87970_comb = {p3_add_87793_comb, p3_add_87488_comb[7:1]};
  assign p3_concat_87973_comb = {p3_add_87795_comb, p3_add_87489_comb[7:1]};
  assign p3_concat_87976_comb = {p3_add_87797_comb, p3_add_87490_comb[7:1]};
  assign p3_concat_87979_comb = {p3_add_87799_comb, p3_add_87491_comb[7:1]};
  assign p3_concat_87982_comb = {p3_add_87801_comb, p3_add_87492_comb[7:1]};
  assign p3_concat_87985_comb = {p3_add_87803_comb, p3_add_87493_comb[7:1]};
  assign p3_concat_87988_comb = {p3_add_87805_comb, p3_add_87494_comb[7:1]};
  assign p3_concat_87991_comb = {p3_add_87807_comb, p3_add_87495_comb[7:1]};
  assign p3_concat_87994_comb = {p3_add_87809_comb, p3_add_87496_comb[7:1]};
  assign p3_concat_87997_comb = {p3_add_87811_comb, p3_add_87497_comb[7:1]};
  assign p3_concat_88000_comb = {p3_add_87813_comb, p3_add_87498_comb[7:1]};
  assign p3_concat_88003_comb = {p3_add_87815_comb, p3_add_87499_comb[7:1]};
  assign p3_concat_88006_comb = {p3_add_87817_comb, p3_add_87500_comb[7:1]};
  assign p3_concat_88009_comb = {p3_add_87819_comb, p3_add_87501_comb[7:1]};
  assign p3_concat_88012_comb = {p3_add_87821_comb, p3_add_87502_comb[7:1]};
  assign p3_clipped__136_comb = $signed(p3_concat_87823_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87823_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87695_comb[2:0], p3_add_87439_comb[7:1]});
  assign p3_clipped__152_comb = $signed(p3_concat_87826_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87826_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87697_comb[2:0], p3_add_87440_comb[7:1]});
  assign p3_clipped__168_comb = $signed(p3_concat_87829_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87829_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87699_comb[2:0], p3_add_87441_comb[7:1]});
  assign p3_clipped__184_comb = $signed(p3_concat_87832_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87832_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87701_comb[2:0], p3_add_87442_comb[7:1]});
  assign p3_clipped__200_comb = $signed(p3_concat_87835_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87835_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87703_comb[2:0], p3_add_87443_comb[7:1]});
  assign p3_clipped__216_comb = $signed(p3_concat_87838_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87838_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87705_comb[2:0], p3_add_87444_comb[7:1]});
  assign p3_clipped__232_comb = $signed(p3_concat_87841_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87841_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87707_comb[2:0], p3_add_87445_comb[7:1]});
  assign p3_clipped__248_comb = $signed(p3_concat_87844_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87844_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87709_comb[2:0], p3_add_87446_comb[7:1]});
  assign p3_clipped__137_comb = $signed(p3_concat_87847_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87847_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87711_comb[2:0], p3_add_87447_comb[7:1]});
  assign p3_clipped__153_comb = $signed(p3_concat_87850_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87850_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87713_comb[2:0], p3_add_87448_comb[7:1]});
  assign p3_clipped__169_comb = $signed(p3_concat_87853_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87853_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87715_comb[2:0], p3_add_87449_comb[7:1]});
  assign p3_clipped__185_comb = $signed(p3_concat_87856_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87856_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87717_comb[2:0], p3_add_87450_comb[7:1]});
  assign p3_clipped__201_comb = $signed(p3_concat_87859_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87859_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87719_comb[2:0], p3_add_87451_comb[7:1]});
  assign p3_clipped__217_comb = $signed(p3_concat_87862_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87862_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87721_comb[2:0], p3_add_87452_comb[7:1]});
  assign p3_clipped__233_comb = $signed(p3_concat_87865_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87865_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87723_comb[2:0], p3_add_87453_comb[7:1]});
  assign p3_clipped__249_comb = $signed(p3_concat_87868_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87868_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87725_comb[2:0], p3_add_87454_comb[7:1]});
  assign p3_clipped__138_comb = $signed(p3_concat_87871_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87871_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87727_comb[2:0], p3_add_87455_comb[7:1]});
  assign p3_clipped__154_comb = $signed(p3_concat_87874_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87874_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87729_comb[2:0], p3_add_87456_comb[7:1]});
  assign p3_clipped__170_comb = $signed(p3_concat_87877_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87877_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87731_comb[2:0], p3_add_87457_comb[7:1]});
  assign p3_clipped__186_comb = $signed(p3_concat_87880_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87880_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87733_comb[2:0], p3_add_87458_comb[7:1]});
  assign p3_clipped__202_comb = $signed(p3_concat_87883_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87883_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87735_comb[2:0], p3_add_87459_comb[7:1]});
  assign p3_clipped__218_comb = $signed(p3_concat_87886_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87886_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87737_comb[2:0], p3_add_87460_comb[7:1]});
  assign p3_clipped__234_comb = $signed(p3_concat_87889_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87889_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87739_comb[2:0], p3_add_87461_comb[7:1]});
  assign p3_clipped__250_comb = $signed(p3_concat_87892_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87892_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87741_comb[2:0], p3_add_87462_comb[7:1]});
  assign p3_clipped__139_comb = $signed(p3_concat_87895_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87895_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87743_comb[2:0], p3_add_87463_comb[7:1]});
  assign p3_clipped__155_comb = $signed(p3_concat_87898_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87898_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87745_comb[2:0], p3_add_87464_comb[7:1]});
  assign p3_clipped__171_comb = $signed(p3_concat_87901_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87901_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87747_comb[2:0], p3_add_87465_comb[7:1]});
  assign p3_clipped__187_comb = $signed(p3_concat_87904_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87904_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87749_comb[2:0], p3_add_87466_comb[7:1]});
  assign p3_clipped__203_comb = $signed(p3_concat_87907_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87907_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87751_comb[2:0], p3_add_87467_comb[7:1]});
  assign p3_clipped__219_comb = $signed(p3_concat_87910_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87910_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87753_comb[2:0], p3_add_87468_comb[7:1]});
  assign p3_clipped__235_comb = $signed(p3_concat_87913_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87913_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87755_comb[2:0], p3_add_87469_comb[7:1]});
  assign p3_clipped__251_comb = $signed(p3_concat_87916_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87916_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87757_comb[2:0], p3_add_87470_comb[7:1]});
  assign p3_clipped__140_comb = $signed(p3_concat_87919_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87919_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87759_comb[2:0], p3_add_87471_comb[7:1]});
  assign p3_clipped__156_comb = $signed(p3_concat_87922_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87922_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87761_comb[2:0], p3_add_87472_comb[7:1]});
  assign p3_clipped__172_comb = $signed(p3_concat_87925_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87925_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87763_comb[2:0], p3_add_87473_comb[7:1]});
  assign p3_clipped__188_comb = $signed(p3_concat_87928_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87928_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87765_comb[2:0], p3_add_87474_comb[7:1]});
  assign p3_clipped__204_comb = $signed(p3_concat_87931_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87931_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87767_comb[2:0], p3_add_87475_comb[7:1]});
  assign p3_clipped__220_comb = $signed(p3_concat_87934_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87934_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87769_comb[2:0], p3_add_87476_comb[7:1]});
  assign p3_clipped__236_comb = $signed(p3_concat_87937_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87937_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87771_comb[2:0], p3_add_87477_comb[7:1]});
  assign p3_clipped__252_comb = $signed(p3_concat_87940_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87940_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87773_comb[2:0], p3_add_87478_comb[7:1]});
  assign p3_clipped__141_comb = $signed(p3_concat_87943_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87943_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87775_comb[2:0], p3_add_87479_comb[7:1]});
  assign p3_clipped__157_comb = $signed(p3_concat_87946_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87946_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87777_comb[2:0], p3_add_87480_comb[7:1]});
  assign p3_clipped__173_comb = $signed(p3_concat_87949_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87949_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87779_comb[2:0], p3_add_87481_comb[7:1]});
  assign p3_clipped__189_comb = $signed(p3_concat_87952_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87952_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87781_comb[2:0], p3_add_87482_comb[7:1]});
  assign p3_clipped__205_comb = $signed(p3_concat_87955_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87955_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87783_comb[2:0], p3_add_87483_comb[7:1]});
  assign p3_clipped__221_comb = $signed(p3_concat_87958_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87958_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87785_comb[2:0], p3_add_87484_comb[7:1]});
  assign p3_clipped__237_comb = $signed(p3_concat_87961_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87961_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87787_comb[2:0], p3_add_87485_comb[7:1]});
  assign p3_clipped__253_comb = $signed(p3_concat_87964_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87964_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87789_comb[2:0], p3_add_87486_comb[7:1]});
  assign p3_clipped__142_comb = $signed(p3_concat_87967_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87967_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87791_comb[2:0], p3_add_87487_comb[7:1]});
  assign p3_clipped__158_comb = $signed(p3_concat_87970_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87970_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87793_comb[2:0], p3_add_87488_comb[7:1]});
  assign p3_clipped__174_comb = $signed(p3_concat_87973_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87973_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87795_comb[2:0], p3_add_87489_comb[7:1]});
  assign p3_clipped__190_comb = $signed(p3_concat_87976_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87976_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87797_comb[2:0], p3_add_87490_comb[7:1]});
  assign p3_clipped__206_comb = $signed(p3_concat_87979_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87979_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87799_comb[2:0], p3_add_87491_comb[7:1]});
  assign p3_clipped__222_comb = $signed(p3_concat_87982_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87982_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87801_comb[2:0], p3_add_87492_comb[7:1]});
  assign p3_clipped__238_comb = $signed(p3_concat_87985_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87985_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87803_comb[2:0], p3_add_87493_comb[7:1]});
  assign p3_clipped__254_comb = $signed(p3_concat_87988_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87988_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87805_comb[2:0], p3_add_87494_comb[7:1]});
  assign p3_clipped__143_comb = $signed(p3_concat_87991_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87991_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87807_comb[2:0], p3_add_87495_comb[7:1]});
  assign p3_clipped__159_comb = $signed(p3_concat_87994_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87994_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87809_comb[2:0], p3_add_87496_comb[7:1]});
  assign p3_clipped__175_comb = $signed(p3_concat_87997_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_87997_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87811_comb[2:0], p3_add_87497_comb[7:1]});
  assign p3_clipped__191_comb = $signed(p3_concat_88000_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_88000_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87813_comb[2:0], p3_add_87498_comb[7:1]});
  assign p3_clipped__207_comb = $signed(p3_concat_88003_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_88003_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87815_comb[2:0], p3_add_87499_comb[7:1]});
  assign p3_clipped__223_comb = $signed(p3_concat_88006_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_88006_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87817_comb[2:0], p3_add_87500_comb[7:1]});
  assign p3_clipped__239_comb = $signed(p3_concat_88009_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_88009_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87819_comb[2:0], p3_add_87501_comb[7:1]});
  assign p3_clipped__255_comb = $signed(p3_concat_88012_comb) < $signed(18'h3_fe01) ? 10'h201 : ($signed(p3_concat_88012_comb) > $signed(18'h0_01ff) ? 10'h1ff : {p3_add_87821_comb[2:0], p3_add_87502_comb[7:1]});
  assign p3_array_88527_comb[0] = p3_clipped__136_comb;
  assign p3_array_88527_comb[1] = p3_clipped__152_comb;
  assign p3_array_88527_comb[2] = p3_clipped__168_comb;
  assign p3_array_88527_comb[3] = p3_clipped__184_comb;
  assign p3_array_88527_comb[4] = p3_clipped__200_comb;
  assign p3_array_88527_comb[5] = p3_clipped__216_comb;
  assign p3_array_88527_comb[6] = p3_clipped__232_comb;
  assign p3_array_88527_comb[7] = p3_clipped__248_comb;
  assign p3_array_88528_comb[0] = p3_clipped__137_comb;
  assign p3_array_88528_comb[1] = p3_clipped__153_comb;
  assign p3_array_88528_comb[2] = p3_clipped__169_comb;
  assign p3_array_88528_comb[3] = p3_clipped__185_comb;
  assign p3_array_88528_comb[4] = p3_clipped__201_comb;
  assign p3_array_88528_comb[5] = p3_clipped__217_comb;
  assign p3_array_88528_comb[6] = p3_clipped__233_comb;
  assign p3_array_88528_comb[7] = p3_clipped__249_comb;
  assign p3_array_88529_comb[0] = p3_clipped__138_comb;
  assign p3_array_88529_comb[1] = p3_clipped__154_comb;
  assign p3_array_88529_comb[2] = p3_clipped__170_comb;
  assign p3_array_88529_comb[3] = p3_clipped__186_comb;
  assign p3_array_88529_comb[4] = p3_clipped__202_comb;
  assign p3_array_88529_comb[5] = p3_clipped__218_comb;
  assign p3_array_88529_comb[6] = p3_clipped__234_comb;
  assign p3_array_88529_comb[7] = p3_clipped__250_comb;
  assign p3_array_88530_comb[0] = p3_clipped__139_comb;
  assign p3_array_88530_comb[1] = p3_clipped__155_comb;
  assign p3_array_88530_comb[2] = p3_clipped__171_comb;
  assign p3_array_88530_comb[3] = p3_clipped__187_comb;
  assign p3_array_88530_comb[4] = p3_clipped__203_comb;
  assign p3_array_88530_comb[5] = p3_clipped__219_comb;
  assign p3_array_88530_comb[6] = p3_clipped__235_comb;
  assign p3_array_88530_comb[7] = p3_clipped__251_comb;
  assign p3_array_88531_comb[0] = p3_clipped__140_comb;
  assign p3_array_88531_comb[1] = p3_clipped__156_comb;
  assign p3_array_88531_comb[2] = p3_clipped__172_comb;
  assign p3_array_88531_comb[3] = p3_clipped__188_comb;
  assign p3_array_88531_comb[4] = p3_clipped__204_comb;
  assign p3_array_88531_comb[5] = p3_clipped__220_comb;
  assign p3_array_88531_comb[6] = p3_clipped__236_comb;
  assign p3_array_88531_comb[7] = p3_clipped__252_comb;
  assign p3_array_88532_comb[0] = p3_clipped__141_comb;
  assign p3_array_88532_comb[1] = p3_clipped__157_comb;
  assign p3_array_88532_comb[2] = p3_clipped__173_comb;
  assign p3_array_88532_comb[3] = p3_clipped__189_comb;
  assign p3_array_88532_comb[4] = p3_clipped__205_comb;
  assign p3_array_88532_comb[5] = p3_clipped__221_comb;
  assign p3_array_88532_comb[6] = p3_clipped__237_comb;
  assign p3_array_88532_comb[7] = p3_clipped__253_comb;
  assign p3_array_88533_comb[0] = p3_clipped__142_comb;
  assign p3_array_88533_comb[1] = p3_clipped__158_comb;
  assign p3_array_88533_comb[2] = p3_clipped__174_comb;
  assign p3_array_88533_comb[3] = p3_clipped__190_comb;
  assign p3_array_88533_comb[4] = p3_clipped__206_comb;
  assign p3_array_88533_comb[5] = p3_clipped__222_comb;
  assign p3_array_88533_comb[6] = p3_clipped__238_comb;
  assign p3_array_88533_comb[7] = p3_clipped__254_comb;
  assign p3_array_88534_comb[0] = p3_clipped__143_comb;
  assign p3_array_88534_comb[1] = p3_clipped__159_comb;
  assign p3_array_88534_comb[2] = p3_clipped__175_comb;
  assign p3_array_88534_comb[3] = p3_clipped__191_comb;
  assign p3_array_88534_comb[4] = p3_clipped__207_comb;
  assign p3_array_88534_comb[5] = p3_clipped__223_comb;
  assign p3_array_88534_comb[6] = p3_clipped__239_comb;
  assign p3_array_88534_comb[7] = p3_clipped__255_comb;
  assign p3_col_transformed_comb[0][0] = p3_array_88527_comb[0];
  assign p3_col_transformed_comb[0][1] = p3_array_88527_comb[1];
  assign p3_col_transformed_comb[0][2] = p3_array_88527_comb[2];
  assign p3_col_transformed_comb[0][3] = p3_array_88527_comb[3];
  assign p3_col_transformed_comb[0][4] = p3_array_88527_comb[4];
  assign p3_col_transformed_comb[0][5] = p3_array_88527_comb[5];
  assign p3_col_transformed_comb[0][6] = p3_array_88527_comb[6];
  assign p3_col_transformed_comb[0][7] = p3_array_88527_comb[7];
  assign p3_col_transformed_comb[1][0] = p3_array_88528_comb[0];
  assign p3_col_transformed_comb[1][1] = p3_array_88528_comb[1];
  assign p3_col_transformed_comb[1][2] = p3_array_88528_comb[2];
  assign p3_col_transformed_comb[1][3] = p3_array_88528_comb[3];
  assign p3_col_transformed_comb[1][4] = p3_array_88528_comb[4];
  assign p3_col_transformed_comb[1][5] = p3_array_88528_comb[5];
  assign p3_col_transformed_comb[1][6] = p3_array_88528_comb[6];
  assign p3_col_transformed_comb[1][7] = p3_array_88528_comb[7];
  assign p3_col_transformed_comb[2][0] = p3_array_88529_comb[0];
  assign p3_col_transformed_comb[2][1] = p3_array_88529_comb[1];
  assign p3_col_transformed_comb[2][2] = p3_array_88529_comb[2];
  assign p3_col_transformed_comb[2][3] = p3_array_88529_comb[3];
  assign p3_col_transformed_comb[2][4] = p3_array_88529_comb[4];
  assign p3_col_transformed_comb[2][5] = p3_array_88529_comb[5];
  assign p3_col_transformed_comb[2][6] = p3_array_88529_comb[6];
  assign p3_col_transformed_comb[2][7] = p3_array_88529_comb[7];
  assign p3_col_transformed_comb[3][0] = p3_array_88530_comb[0];
  assign p3_col_transformed_comb[3][1] = p3_array_88530_comb[1];
  assign p3_col_transformed_comb[3][2] = p3_array_88530_comb[2];
  assign p3_col_transformed_comb[3][3] = p3_array_88530_comb[3];
  assign p3_col_transformed_comb[3][4] = p3_array_88530_comb[4];
  assign p3_col_transformed_comb[3][5] = p3_array_88530_comb[5];
  assign p3_col_transformed_comb[3][6] = p3_array_88530_comb[6];
  assign p3_col_transformed_comb[3][7] = p3_array_88530_comb[7];
  assign p3_col_transformed_comb[4][0] = p3_array_88531_comb[0];
  assign p3_col_transformed_comb[4][1] = p3_array_88531_comb[1];
  assign p3_col_transformed_comb[4][2] = p3_array_88531_comb[2];
  assign p3_col_transformed_comb[4][3] = p3_array_88531_comb[3];
  assign p3_col_transformed_comb[4][4] = p3_array_88531_comb[4];
  assign p3_col_transformed_comb[4][5] = p3_array_88531_comb[5];
  assign p3_col_transformed_comb[4][6] = p3_array_88531_comb[6];
  assign p3_col_transformed_comb[4][7] = p3_array_88531_comb[7];
  assign p3_col_transformed_comb[5][0] = p3_array_88532_comb[0];
  assign p3_col_transformed_comb[5][1] = p3_array_88532_comb[1];
  assign p3_col_transformed_comb[5][2] = p3_array_88532_comb[2];
  assign p3_col_transformed_comb[5][3] = p3_array_88532_comb[3];
  assign p3_col_transformed_comb[5][4] = p3_array_88532_comb[4];
  assign p3_col_transformed_comb[5][5] = p3_array_88532_comb[5];
  assign p3_col_transformed_comb[5][6] = p3_array_88532_comb[6];
  assign p3_col_transformed_comb[5][7] = p3_array_88532_comb[7];
  assign p3_col_transformed_comb[6][0] = p3_array_88533_comb[0];
  assign p3_col_transformed_comb[6][1] = p3_array_88533_comb[1];
  assign p3_col_transformed_comb[6][2] = p3_array_88533_comb[2];
  assign p3_col_transformed_comb[6][3] = p3_array_88533_comb[3];
  assign p3_col_transformed_comb[6][4] = p3_array_88533_comb[4];
  assign p3_col_transformed_comb[6][5] = p3_array_88533_comb[5];
  assign p3_col_transformed_comb[6][6] = p3_array_88533_comb[6];
  assign p3_col_transformed_comb[6][7] = p3_array_88533_comb[7];
  assign p3_col_transformed_comb[7][0] = p3_array_88534_comb[0];
  assign p3_col_transformed_comb[7][1] = p3_array_88534_comb[1];
  assign p3_col_transformed_comb[7][2] = p3_array_88534_comb[2];
  assign p3_col_transformed_comb[7][3] = p3_array_88534_comb[3];
  assign p3_col_transformed_comb[7][4] = p3_array_88534_comb[4];
  assign p3_col_transformed_comb[7][5] = p3_array_88534_comb[5];
  assign p3_col_transformed_comb[7][6] = p3_array_88534_comb[6];
  assign p3_col_transformed_comb[7][7] = p3_array_88534_comb[7];

  // Registers for pipe stage 3:
  reg [9:0] p3_col_transformed[0:7][0:7];
  always @ (posedge clk) begin
    p3_col_transformed[0][0] <= p3_col_transformed_comb[0][0];
    p3_col_transformed[0][1] <= p3_col_transformed_comb[0][1];
    p3_col_transformed[0][2] <= p3_col_transformed_comb[0][2];
    p3_col_transformed[0][3] <= p3_col_transformed_comb[0][3];
    p3_col_transformed[0][4] <= p3_col_transformed_comb[0][4];
    p3_col_transformed[0][5] <= p3_col_transformed_comb[0][5];
    p3_col_transformed[0][6] <= p3_col_transformed_comb[0][6];
    p3_col_transformed[0][7] <= p3_col_transformed_comb[0][7];
    p3_col_transformed[1][0] <= p3_col_transformed_comb[1][0];
    p3_col_transformed[1][1] <= p3_col_transformed_comb[1][1];
    p3_col_transformed[1][2] <= p3_col_transformed_comb[1][2];
    p3_col_transformed[1][3] <= p3_col_transformed_comb[1][3];
    p3_col_transformed[1][4] <= p3_col_transformed_comb[1][4];
    p3_col_transformed[1][5] <= p3_col_transformed_comb[1][5];
    p3_col_transformed[1][6] <= p3_col_transformed_comb[1][6];
    p3_col_transformed[1][7] <= p3_col_transformed_comb[1][7];
    p3_col_transformed[2][0] <= p3_col_transformed_comb[2][0];
    p3_col_transformed[2][1] <= p3_col_transformed_comb[2][1];
    p3_col_transformed[2][2] <= p3_col_transformed_comb[2][2];
    p3_col_transformed[2][3] <= p3_col_transformed_comb[2][3];
    p3_col_transformed[2][4] <= p3_col_transformed_comb[2][4];
    p3_col_transformed[2][5] <= p3_col_transformed_comb[2][5];
    p3_col_transformed[2][6] <= p3_col_transformed_comb[2][6];
    p3_col_transformed[2][7] <= p3_col_transformed_comb[2][7];
    p3_col_transformed[3][0] <= p3_col_transformed_comb[3][0];
    p3_col_transformed[3][1] <= p3_col_transformed_comb[3][1];
    p3_col_transformed[3][2] <= p3_col_transformed_comb[3][2];
    p3_col_transformed[3][3] <= p3_col_transformed_comb[3][3];
    p3_col_transformed[3][4] <= p3_col_transformed_comb[3][4];
    p3_col_transformed[3][5] <= p3_col_transformed_comb[3][5];
    p3_col_transformed[3][6] <= p3_col_transformed_comb[3][6];
    p3_col_transformed[3][7] <= p3_col_transformed_comb[3][7];
    p3_col_transformed[4][0] <= p3_col_transformed_comb[4][0];
    p3_col_transformed[4][1] <= p3_col_transformed_comb[4][1];
    p3_col_transformed[4][2] <= p3_col_transformed_comb[4][2];
    p3_col_transformed[4][3] <= p3_col_transformed_comb[4][3];
    p3_col_transformed[4][4] <= p3_col_transformed_comb[4][4];
    p3_col_transformed[4][5] <= p3_col_transformed_comb[4][5];
    p3_col_transformed[4][6] <= p3_col_transformed_comb[4][6];
    p3_col_transformed[4][7] <= p3_col_transformed_comb[4][7];
    p3_col_transformed[5][0] <= p3_col_transformed_comb[5][0];
    p3_col_transformed[5][1] <= p3_col_transformed_comb[5][1];
    p3_col_transformed[5][2] <= p3_col_transformed_comb[5][2];
    p3_col_transformed[5][3] <= p3_col_transformed_comb[5][3];
    p3_col_transformed[5][4] <= p3_col_transformed_comb[5][4];
    p3_col_transformed[5][5] <= p3_col_transformed_comb[5][5];
    p3_col_transformed[5][6] <= p3_col_transformed_comb[5][6];
    p3_col_transformed[5][7] <= p3_col_transformed_comb[5][7];
    p3_col_transformed[6][0] <= p3_col_transformed_comb[6][0];
    p3_col_transformed[6][1] <= p3_col_transformed_comb[6][1];
    p3_col_transformed[6][2] <= p3_col_transformed_comb[6][2];
    p3_col_transformed[6][3] <= p3_col_transformed_comb[6][3];
    p3_col_transformed[6][4] <= p3_col_transformed_comb[6][4];
    p3_col_transformed[6][5] <= p3_col_transformed_comb[6][5];
    p3_col_transformed[6][6] <= p3_col_transformed_comb[6][6];
    p3_col_transformed[6][7] <= p3_col_transformed_comb[6][7];
    p3_col_transformed[7][0] <= p3_col_transformed_comb[7][0];
    p3_col_transformed[7][1] <= p3_col_transformed_comb[7][1];
    p3_col_transformed[7][2] <= p3_col_transformed_comb[7][2];
    p3_col_transformed[7][3] <= p3_col_transformed_comb[7][3];
    p3_col_transformed[7][4] <= p3_col_transformed_comb[7][4];
    p3_col_transformed[7][5] <= p3_col_transformed_comb[7][5];
    p3_col_transformed[7][6] <= p3_col_transformed_comb[7][6];
    p3_col_transformed[7][7] <= p3_col_transformed_comb[7][7];
  end
  assign out = {{p3_col_transformed[7][7], p3_col_transformed[7][6], p3_col_transformed[7][5], p3_col_transformed[7][4], p3_col_transformed[7][3], p3_col_transformed[7][2], p3_col_transformed[7][1], p3_col_transformed[7][0]}, {p3_col_transformed[6][7], p3_col_transformed[6][6], p3_col_transformed[6][5], p3_col_transformed[6][4], p3_col_transformed[6][3], p3_col_transformed[6][2], p3_col_transformed[6][1], p3_col_transformed[6][0]}, {p3_col_transformed[5][7], p3_col_transformed[5][6], p3_col_transformed[5][5], p3_col_transformed[5][4], p3_col_transformed[5][3], p3_col_transformed[5][2], p3_col_transformed[5][1], p3_col_transformed[5][0]}, {p3_col_transformed[4][7], p3_col_transformed[4][6], p3_col_transformed[4][5], p3_col_transformed[4][4], p3_col_transformed[4][3], p3_col_transformed[4][2], p3_col_transformed[4][1], p3_col_transformed[4][0]}, {p3_col_transformed[3][7], p3_col_transformed[3][6], p3_col_transformed[3][5], p3_col_transformed[3][4], p3_col_transformed[3][3], p3_col_transformed[3][2], p3_col_transformed[3][1], p3_col_transformed[3][0]}, {p3_col_transformed[2][7], p3_col_transformed[2][6], p3_col_transformed[2][5], p3_col_transformed[2][4], p3_col_transformed[2][3], p3_col_transformed[2][2], p3_col_transformed[2][1], p3_col_transformed[2][0]}, {p3_col_transformed[1][7], p3_col_transformed[1][6], p3_col_transformed[1][5], p3_col_transformed[1][4], p3_col_transformed[1][3], p3_col_transformed[1][2], p3_col_transformed[1][1], p3_col_transformed[1][0]}, {p3_col_transformed[0][7], p3_col_transformed[0][6], p3_col_transformed[0][5], p3_col_transformed[0][4], p3_col_transformed[0][3], p3_col_transformed[0][2], p3_col_transformed[0][1], p3_col_transformed[0][0]}};
endmodule
