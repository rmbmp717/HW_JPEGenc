module Huffman_ACenc(
  input wire clk,
  input wire [511:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [35:0] out
);
  wire [4:0] literal_9083[0:251];
  assign literal_9083[0] = 5'h02;
  assign literal_9083[1] = 5'h02;
  assign literal_9083[2] = 5'h03;
  assign literal_9083[3] = 5'h04;
  assign literal_9083[4] = 5'h05;
  assign literal_9083[5] = 5'h07;
  assign literal_9083[6] = 5'h08;
  assign literal_9083[7] = 5'h0e;
  assign literal_9083[8] = 5'h10;
  assign literal_9083[9] = 5'h10;
  assign literal_9083[10] = 5'h10;
  assign literal_9083[11] = 5'h00;
  assign literal_9083[12] = 5'h00;
  assign literal_9083[13] = 5'h00;
  assign literal_9083[14] = 5'h00;
  assign literal_9083[15] = 5'h00;
  assign literal_9083[16] = 5'h00;
  assign literal_9083[17] = 5'h03;
  assign literal_9083[18] = 5'h06;
  assign literal_9083[19] = 5'h07;
  assign literal_9083[20] = 5'h09;
  assign literal_9083[21] = 5'h0b;
  assign literal_9083[22] = 5'h0d;
  assign literal_9083[23] = 5'h10;
  assign literal_9083[24] = 5'h10;
  assign literal_9083[25] = 5'h10;
  assign literal_9083[26] = 5'h10;
  assign literal_9083[27] = 5'h00;
  assign literal_9083[28] = 5'h00;
  assign literal_9083[29] = 5'h00;
  assign literal_9083[30] = 5'h00;
  assign literal_9083[31] = 5'h00;
  assign literal_9083[32] = 5'h00;
  assign literal_9083[33] = 5'h05;
  assign literal_9083[34] = 5'h07;
  assign literal_9083[35] = 5'h0a;
  assign literal_9083[36] = 5'h0c;
  assign literal_9083[37] = 5'h0d;
  assign literal_9083[38] = 5'h10;
  assign literal_9083[39] = 5'h10;
  assign literal_9083[40] = 5'h10;
  assign literal_9083[41] = 5'h10;
  assign literal_9083[42] = 5'h10;
  assign literal_9083[43] = 5'h00;
  assign literal_9083[44] = 5'h00;
  assign literal_9083[45] = 5'h00;
  assign literal_9083[46] = 5'h00;
  assign literal_9083[47] = 5'h00;
  assign literal_9083[48] = 5'h00;
  assign literal_9083[49] = 5'h06;
  assign literal_9083[50] = 5'h08;
  assign literal_9083[51] = 5'h0b;
  assign literal_9083[52] = 5'h0c;
  assign literal_9083[53] = 5'h0f;
  assign literal_9083[54] = 5'h10;
  assign literal_9083[55] = 5'h10;
  assign literal_9083[56] = 5'h10;
  assign literal_9083[57] = 5'h10;
  assign literal_9083[58] = 5'h10;
  assign literal_9083[59] = 5'h00;
  assign literal_9083[60] = 5'h00;
  assign literal_9083[61] = 5'h00;
  assign literal_9083[62] = 5'h00;
  assign literal_9083[63] = 5'h00;
  assign literal_9083[64] = 5'h00;
  assign literal_9083[65] = 5'h06;
  assign literal_9083[66] = 5'h0a;
  assign literal_9083[67] = 5'h0c;
  assign literal_9083[68] = 5'h0f;
  assign literal_9083[69] = 5'h10;
  assign literal_9083[70] = 5'h10;
  assign literal_9083[71] = 5'h10;
  assign literal_9083[72] = 5'h10;
  assign literal_9083[73] = 5'h10;
  assign literal_9083[74] = 5'h10;
  assign literal_9083[75] = 5'h00;
  assign literal_9083[76] = 5'h00;
  assign literal_9083[77] = 5'h00;
  assign literal_9083[78] = 5'h00;
  assign literal_9083[79] = 5'h00;
  assign literal_9083[80] = 5'h00;
  assign literal_9083[81] = 5'h07;
  assign literal_9083[82] = 5'h0b;
  assign literal_9083[83] = 5'h0d;
  assign literal_9083[84] = 5'h10;
  assign literal_9083[85] = 5'h10;
  assign literal_9083[86] = 5'h10;
  assign literal_9083[87] = 5'h10;
  assign literal_9083[88] = 5'h10;
  assign literal_9083[89] = 5'h10;
  assign literal_9083[90] = 5'h10;
  assign literal_9083[91] = 5'h00;
  assign literal_9083[92] = 5'h00;
  assign literal_9083[93] = 5'h00;
  assign literal_9083[94] = 5'h00;
  assign literal_9083[95] = 5'h00;
  assign literal_9083[96] = 5'h00;
  assign literal_9083[97] = 5'h07;
  assign literal_9083[98] = 5'h0b;
  assign literal_9083[99] = 5'h0d;
  assign literal_9083[100] = 5'h10;
  assign literal_9083[101] = 5'h10;
  assign literal_9083[102] = 5'h10;
  assign literal_9083[103] = 5'h10;
  assign literal_9083[104] = 5'h10;
  assign literal_9083[105] = 5'h10;
  assign literal_9083[106] = 5'h10;
  assign literal_9083[107] = 5'h00;
  assign literal_9083[108] = 5'h00;
  assign literal_9083[109] = 5'h00;
  assign literal_9083[110] = 5'h00;
  assign literal_9083[111] = 5'h00;
  assign literal_9083[112] = 5'h00;
  assign literal_9083[113] = 5'h08;
  assign literal_9083[114] = 5'h0b;
  assign literal_9083[115] = 5'h0e;
  assign literal_9083[116] = 5'h10;
  assign literal_9083[117] = 5'h10;
  assign literal_9083[118] = 5'h10;
  assign literal_9083[119] = 5'h10;
  assign literal_9083[120] = 5'h10;
  assign literal_9083[121] = 5'h10;
  assign literal_9083[122] = 5'h10;
  assign literal_9083[123] = 5'h00;
  assign literal_9083[124] = 5'h00;
  assign literal_9083[125] = 5'h00;
  assign literal_9083[126] = 5'h00;
  assign literal_9083[127] = 5'h00;
  assign literal_9083[128] = 5'h00;
  assign literal_9083[129] = 5'h08;
  assign literal_9083[130] = 5'h0c;
  assign literal_9083[131] = 5'h10;
  assign literal_9083[132] = 5'h10;
  assign literal_9083[133] = 5'h10;
  assign literal_9083[134] = 5'h10;
  assign literal_9083[135] = 5'h10;
  assign literal_9083[136] = 5'h10;
  assign literal_9083[137] = 5'h10;
  assign literal_9083[138] = 5'h10;
  assign literal_9083[139] = 5'h00;
  assign literal_9083[140] = 5'h00;
  assign literal_9083[141] = 5'h00;
  assign literal_9083[142] = 5'h00;
  assign literal_9083[143] = 5'h00;
  assign literal_9083[144] = 5'h00;
  assign literal_9083[145] = 5'h08;
  assign literal_9083[146] = 5'h0d;
  assign literal_9083[147] = 5'h10;
  assign literal_9083[148] = 5'h10;
  assign literal_9083[149] = 5'h10;
  assign literal_9083[150] = 5'h10;
  assign literal_9083[151] = 5'h10;
  assign literal_9083[152] = 5'h10;
  assign literal_9083[153] = 5'h10;
  assign literal_9083[154] = 5'h10;
  assign literal_9083[155] = 5'h00;
  assign literal_9083[156] = 5'h00;
  assign literal_9083[157] = 5'h00;
  assign literal_9083[158] = 5'h00;
  assign literal_9083[159] = 5'h00;
  assign literal_9083[160] = 5'h00;
  assign literal_9083[161] = 5'h09;
  assign literal_9083[162] = 5'h0d;
  assign literal_9083[163] = 5'h10;
  assign literal_9083[164] = 5'h10;
  assign literal_9083[165] = 5'h10;
  assign literal_9083[166] = 5'h10;
  assign literal_9083[167] = 5'h10;
  assign literal_9083[168] = 5'h10;
  assign literal_9083[169] = 5'h10;
  assign literal_9083[170] = 5'h10;
  assign literal_9083[171] = 5'h00;
  assign literal_9083[172] = 5'h00;
  assign literal_9083[173] = 5'h00;
  assign literal_9083[174] = 5'h00;
  assign literal_9083[175] = 5'h00;
  assign literal_9083[176] = 5'h00;
  assign literal_9083[177] = 5'h09;
  assign literal_9083[178] = 5'h0d;
  assign literal_9083[179] = 5'h10;
  assign literal_9083[180] = 5'h10;
  assign literal_9083[181] = 5'h10;
  assign literal_9083[182] = 5'h10;
  assign literal_9083[183] = 5'h10;
  assign literal_9083[184] = 5'h10;
  assign literal_9083[185] = 5'h10;
  assign literal_9083[186] = 5'h10;
  assign literal_9083[187] = 5'h00;
  assign literal_9083[188] = 5'h00;
  assign literal_9083[189] = 5'h00;
  assign literal_9083[190] = 5'h00;
  assign literal_9083[191] = 5'h00;
  assign literal_9083[192] = 5'h00;
  assign literal_9083[193] = 5'h0a;
  assign literal_9083[194] = 5'h0d;
  assign literal_9083[195] = 5'h10;
  assign literal_9083[196] = 5'h10;
  assign literal_9083[197] = 5'h10;
  assign literal_9083[198] = 5'h10;
  assign literal_9083[199] = 5'h10;
  assign literal_9083[200] = 5'h10;
  assign literal_9083[201] = 5'h10;
  assign literal_9083[202] = 5'h10;
  assign literal_9083[203] = 5'h00;
  assign literal_9083[204] = 5'h00;
  assign literal_9083[205] = 5'h00;
  assign literal_9083[206] = 5'h00;
  assign literal_9083[207] = 5'h00;
  assign literal_9083[208] = 5'h00;
  assign literal_9083[209] = 5'h0a;
  assign literal_9083[210] = 5'h0e;
  assign literal_9083[211] = 5'h10;
  assign literal_9083[212] = 5'h10;
  assign literal_9083[213] = 5'h10;
  assign literal_9083[214] = 5'h10;
  assign literal_9083[215] = 5'h10;
  assign literal_9083[216] = 5'h10;
  assign literal_9083[217] = 5'h10;
  assign literal_9083[218] = 5'h10;
  assign literal_9083[219] = 5'h00;
  assign literal_9083[220] = 5'h00;
  assign literal_9083[221] = 5'h00;
  assign literal_9083[222] = 5'h00;
  assign literal_9083[223] = 5'h00;
  assign literal_9083[224] = 5'h00;
  assign literal_9083[225] = 5'h0a;
  assign literal_9083[226] = 5'h0f;
  assign literal_9083[227] = 5'h10;
  assign literal_9083[228] = 5'h10;
  assign literal_9083[229] = 5'h10;
  assign literal_9083[230] = 5'h10;
  assign literal_9083[231] = 5'h10;
  assign literal_9083[232] = 5'h10;
  assign literal_9083[233] = 5'h10;
  assign literal_9083[234] = 5'h10;
  assign literal_9083[235] = 5'h00;
  assign literal_9083[236] = 5'h00;
  assign literal_9083[237] = 5'h00;
  assign literal_9083[238] = 5'h00;
  assign literal_9083[239] = 5'h00;
  assign literal_9083[240] = 5'h09;
  assign literal_9083[241] = 5'h0b;
  assign literal_9083[242] = 5'h10;
  assign literal_9083[243] = 5'h10;
  assign literal_9083[244] = 5'h10;
  assign literal_9083[245] = 5'h10;
  assign literal_9083[246] = 5'h10;
  assign literal_9083[247] = 5'h10;
  assign literal_9083[248] = 5'h10;
  assign literal_9083[249] = 5'h10;
  assign literal_9083[250] = 5'h10;
  assign literal_9083[251] = 5'h00;
  wire [4:0] literal_9085[0:251];
  assign literal_9085[0] = 5'h04;
  assign literal_9085[1] = 5'h02;
  assign literal_9085[2] = 5'h02;
  assign literal_9085[3] = 5'h03;
  assign literal_9085[4] = 5'h04;
  assign literal_9085[5] = 5'h05;
  assign literal_9085[6] = 5'h07;
  assign literal_9085[7] = 5'h09;
  assign literal_9085[8] = 5'h00;
  assign literal_9085[9] = 5'h00;
  assign literal_9085[10] = 5'h00;
  assign literal_9085[11] = 5'h00;
  assign literal_9085[12] = 5'h00;
  assign literal_9085[13] = 5'h00;
  assign literal_9085[14] = 5'h00;
  assign literal_9085[15] = 5'h00;
  assign literal_9085[16] = 5'h00;
  assign literal_9085[17] = 5'h04;
  assign literal_9085[18] = 5'h05;
  assign literal_9085[19] = 5'h07;
  assign literal_9085[20] = 5'h09;
  assign literal_9085[21] = 5'h0a;
  assign literal_9085[22] = 5'h0b;
  assign literal_9085[23] = 5'h10;
  assign literal_9085[24] = 5'h00;
  assign literal_9085[25] = 5'h00;
  assign literal_9085[26] = 5'h00;
  assign literal_9085[27] = 5'h00;
  assign literal_9085[28] = 5'h00;
  assign literal_9085[29] = 5'h00;
  assign literal_9085[30] = 5'h00;
  assign literal_9085[31] = 5'h00;
  assign literal_9085[32] = 5'h00;
  assign literal_9085[33] = 5'h05;
  assign literal_9085[34] = 5'h08;
  assign literal_9085[35] = 5'h0a;
  assign literal_9085[36] = 5'h0c;
  assign literal_9085[37] = 5'h00;
  assign literal_9085[38] = 5'h00;
  assign literal_9085[39] = 5'h00;
  assign literal_9085[40] = 5'h00;
  assign literal_9085[41] = 5'h00;
  assign literal_9085[42] = 5'h00;
  assign literal_9085[43] = 5'h00;
  assign literal_9085[44] = 5'h00;
  assign literal_9085[45] = 5'h00;
  assign literal_9085[46] = 5'h00;
  assign literal_9085[47] = 5'h00;
  assign literal_9085[48] = 5'h00;
  assign literal_9085[49] = 5'h06;
  assign literal_9085[50] = 5'h09;
  assign literal_9085[51] = 5'h00;
  assign literal_9085[52] = 5'h0c;
  assign literal_9085[53] = 5'h10;
  assign literal_9085[54] = 5'h10;
  assign literal_9085[55] = 5'h10;
  assign literal_9085[56] = 5'h10;
  assign literal_9085[57] = 5'h10;
  assign literal_9085[58] = 5'h00;
  assign literal_9085[59] = 5'h00;
  assign literal_9085[60] = 5'h00;
  assign literal_9085[61] = 5'h00;
  assign literal_9085[62] = 5'h00;
  assign literal_9085[63] = 5'h00;
  assign literal_9085[64] = 5'h00;
  assign literal_9085[65] = 5'h06;
  assign literal_9085[66] = 5'h0a;
  assign literal_9085[67] = 5'h0e;
  assign literal_9085[68] = 5'h10;
  assign literal_9085[69] = 5'h10;
  assign literal_9085[70] = 5'h10;
  assign literal_9085[71] = 5'h10;
  assign literal_9085[72] = 5'h10;
  assign literal_9085[73] = 5'h10;
  assign literal_9085[74] = 5'h00;
  assign literal_9085[75] = 5'h00;
  assign literal_9085[76] = 5'h00;
  assign literal_9085[77] = 5'h00;
  assign literal_9085[78] = 5'h00;
  assign literal_9085[79] = 5'h00;
  assign literal_9085[80] = 5'h00;
  assign literal_9085[81] = 5'h07;
  assign literal_9085[82] = 5'h0a;
  assign literal_9085[83] = 5'h0e;
  assign literal_9085[84] = 5'h10;
  assign literal_9085[85] = 5'h10;
  assign literal_9085[86] = 5'h10;
  assign literal_9085[87] = 5'h10;
  assign literal_9085[88] = 5'h10;
  assign literal_9085[89] = 5'h10;
  assign literal_9085[90] = 5'h00;
  assign literal_9085[91] = 5'h00;
  assign literal_9085[92] = 5'h00;
  assign literal_9085[93] = 5'h00;
  assign literal_9085[94] = 5'h00;
  assign literal_9085[95] = 5'h00;
  assign literal_9085[96] = 5'h00;
  assign literal_9085[97] = 5'h07;
  assign literal_9085[98] = 5'h0c;
  assign literal_9085[99] = 5'h0f;
  assign literal_9085[100] = 5'h10;
  assign literal_9085[101] = 5'h10;
  assign literal_9085[102] = 5'h10;
  assign literal_9085[103] = 5'h10;
  assign literal_9085[104] = 5'h10;
  assign literal_9085[105] = 5'h10;
  assign literal_9085[106] = 5'h10;
  assign literal_9085[107] = 5'h10;
  assign literal_9085[108] = 5'h00;
  assign literal_9085[109] = 5'h00;
  assign literal_9085[110] = 5'h00;
  assign literal_9085[111] = 5'h00;
  assign literal_9085[112] = 5'h00;
  assign literal_9085[113] = 5'h08;
  assign literal_9085[114] = 5'h0c;
  assign literal_9085[115] = 5'h10;
  assign literal_9085[116] = 5'h10;
  assign literal_9085[117] = 5'h10;
  assign literal_9085[118] = 5'h10;
  assign literal_9085[119] = 5'h10;
  assign literal_9085[120] = 5'h10;
  assign literal_9085[121] = 5'h10;
  assign literal_9085[122] = 5'h10;
  assign literal_9085[123] = 5'h00;
  assign literal_9085[124] = 5'h00;
  assign literal_9085[125] = 5'h00;
  assign literal_9085[126] = 5'h00;
  assign literal_9085[127] = 5'h00;
  assign literal_9085[128] = 5'h00;
  assign literal_9085[129] = 5'h09;
  assign literal_9085[130] = 5'h0d;
  assign literal_9085[131] = 5'h10;
  assign literal_9085[132] = 5'h10;
  assign literal_9085[133] = 5'h00;
  assign literal_9085[134] = 5'h10;
  assign literal_9085[135] = 5'h10;
  assign literal_9085[136] = 5'h10;
  assign literal_9085[137] = 5'h10;
  assign literal_9085[138] = 5'h00;
  assign literal_9085[139] = 5'h00;
  assign literal_9085[140] = 5'h00;
  assign literal_9085[141] = 5'h00;
  assign literal_9085[142] = 5'h00;
  assign literal_9085[143] = 5'h00;
  assign literal_9085[144] = 5'h00;
  assign literal_9085[145] = 5'h09;
  assign literal_9085[146] = 5'h0f;
  assign literal_9085[147] = 5'h10;
  assign literal_9085[148] = 5'h10;
  assign literal_9085[149] = 5'h10;
  assign literal_9085[150] = 5'h10;
  assign literal_9085[151] = 5'h10;
  assign literal_9085[152] = 5'h10;
  assign literal_9085[153] = 5'h10;
  assign literal_9085[154] = 5'h10;
  assign literal_9085[155] = 5'h00;
  assign literal_9085[156] = 5'h00;
  assign literal_9085[157] = 5'h00;
  assign literal_9085[158] = 5'h00;
  assign literal_9085[159] = 5'h00;
  assign literal_9085[160] = 5'h00;
  assign literal_9085[161] = 5'h09;
  assign literal_9085[162] = 5'h0f;
  assign literal_9085[163] = 5'h10;
  assign literal_9085[164] = 5'h10;
  assign literal_9085[165] = 5'h10;
  assign literal_9085[166] = 5'h10;
  assign literal_9085[167] = 5'h10;
  assign literal_9085[168] = 5'h10;
  assign literal_9085[169] = 5'h10;
  assign literal_9085[170] = 5'h00;
  assign literal_9085[171] = 5'h00;
  assign literal_9085[172] = 5'h00;
  assign literal_9085[173] = 5'h00;
  assign literal_9085[174] = 5'h00;
  assign literal_9085[175] = 5'h00;
  assign literal_9085[176] = 5'h00;
  assign literal_9085[177] = 5'h0a;
  assign literal_9085[178] = 5'h0f;
  assign literal_9085[179] = 5'h10;
  assign literal_9085[180] = 5'h10;
  assign literal_9085[181] = 5'h10;
  assign literal_9085[182] = 5'h10;
  assign literal_9085[183] = 5'h10;
  assign literal_9085[184] = 5'h10;
  assign literal_9085[185] = 5'h10;
  assign literal_9085[186] = 5'h00;
  assign literal_9085[187] = 5'h00;
  assign literal_9085[188] = 5'h00;
  assign literal_9085[189] = 5'h00;
  assign literal_9085[190] = 5'h00;
  assign literal_9085[191] = 5'h00;
  assign literal_9085[192] = 5'h00;
  assign literal_9085[193] = 5'h0a;
  assign literal_9085[194] = 5'h10;
  assign literal_9085[195] = 5'h10;
  assign literal_9085[196] = 5'h10;
  assign literal_9085[197] = 5'h10;
  assign literal_9085[198] = 5'h10;
  assign literal_9085[199] = 5'h10;
  assign literal_9085[200] = 5'h10;
  assign literal_9085[201] = 5'h10;
  assign literal_9085[202] = 5'h00;
  assign literal_9085[203] = 5'h00;
  assign literal_9085[204] = 5'h00;
  assign literal_9085[205] = 5'h00;
  assign literal_9085[206] = 5'h00;
  assign literal_9085[207] = 5'h00;
  assign literal_9085[208] = 5'h00;
  assign literal_9085[209] = 5'h0a;
  assign literal_9085[210] = 5'h10;
  assign literal_9085[211] = 5'h10;
  assign literal_9085[212] = 5'h10;
  assign literal_9085[213] = 5'h10;
  assign literal_9085[214] = 5'h10;
  assign literal_9085[215] = 5'h10;
  assign literal_9085[216] = 5'h10;
  assign literal_9085[217] = 5'h10;
  assign literal_9085[218] = 5'h00;
  assign literal_9085[219] = 5'h00;
  assign literal_9085[220] = 5'h00;
  assign literal_9085[221] = 5'h00;
  assign literal_9085[222] = 5'h00;
  assign literal_9085[223] = 5'h00;
  assign literal_9085[224] = 5'h00;
  assign literal_9085[225] = 5'h0b;
  assign literal_9085[226] = 5'h10;
  assign literal_9085[227] = 5'h10;
  assign literal_9085[228] = 5'h10;
  assign literal_9085[229] = 5'h10;
  assign literal_9085[230] = 5'h10;
  assign literal_9085[231] = 5'h10;
  assign literal_9085[232] = 5'h10;
  assign literal_9085[233] = 5'h10;
  assign literal_9085[234] = 5'h00;
  assign literal_9085[235] = 5'h00;
  assign literal_9085[236] = 5'h00;
  assign literal_9085[237] = 5'h00;
  assign literal_9085[238] = 5'h00;
  assign literal_9085[239] = 5'h00;
  assign literal_9085[240] = 5'h0c;
  assign literal_9085[241] = 5'h0d;
  assign literal_9085[242] = 5'h10;
  assign literal_9085[243] = 5'h10;
  assign literal_9085[244] = 5'h10;
  assign literal_9085[245] = 5'h10;
  assign literal_9085[246] = 5'h10;
  assign literal_9085[247] = 5'h10;
  assign literal_9085[248] = 5'h10;
  assign literal_9085[249] = 5'h10;
  assign literal_9085[250] = 5'h10;
  assign literal_9085[251] = 5'h00;
  wire [15:0] literal_9086[0:251];
  assign literal_9086[0] = 16'h0001;
  assign literal_9086[1] = 16'h0000;
  assign literal_9086[2] = 16'h0004;
  assign literal_9086[3] = 16'h000c;
  assign literal_9086[4] = 16'h001a;
  assign literal_9086[5] = 16'h0076;
  assign literal_9086[6] = 16'h00f6;
  assign literal_9086[7] = 16'h3fe0;
  assign literal_9086[8] = 16'hff96;
  assign literal_9086[9] = 16'hff97;
  assign literal_9086[10] = 16'hff98;
  assign literal_9086[11] = 16'h0000;
  assign literal_9086[12] = 16'h0000;
  assign literal_9086[13] = 16'h0000;
  assign literal_9086[14] = 16'h0000;
  assign literal_9086[15] = 16'h0000;
  assign literal_9086[16] = 16'h0000;
  assign literal_9086[17] = 16'h0005;
  assign literal_9086[18] = 16'h0038;
  assign literal_9086[19] = 16'h0078;
  assign literal_9086[20] = 16'h01f9;
  assign literal_9086[21] = 16'h07f2;
  assign literal_9086[22] = 16'h1fe8;
  assign literal_9086[23] = 16'hff93;
  assign literal_9086[24] = 16'hff99;
  assign literal_9086[25] = 16'hff9a;
  assign literal_9086[26] = 16'hff9e;
  assign literal_9086[27] = 16'h0000;
  assign literal_9086[28] = 16'h0000;
  assign literal_9086[29] = 16'h0000;
  assign literal_9086[30] = 16'h0000;
  assign literal_9086[31] = 16'h0000;
  assign literal_9086[32] = 16'h0000;
  assign literal_9086[33] = 16'h001b;
  assign literal_9086[34] = 16'h007a;
  assign literal_9086[35] = 16'h03f7;
  assign literal_9086[36] = 16'h0ff0;
  assign literal_9086[37] = 16'h1feb;
  assign literal_9086[38] = 16'hff9b;
  assign literal_9086[39] = 16'hff9f;
  assign literal_9086[40] = 16'hffa8;
  assign literal_9086[41] = 16'hffa9;
  assign literal_9086[42] = 16'hfff1;
  assign literal_9086[43] = 16'h0000;
  assign literal_9086[44] = 16'h0000;
  assign literal_9086[45] = 16'h0000;
  assign literal_9086[46] = 16'h0000;
  assign literal_9086[47] = 16'h0000;
  assign literal_9086[48] = 16'h0000;
  assign literal_9086[49] = 16'h0039;
  assign literal_9086[50] = 16'h00fa;
  assign literal_9086[51] = 16'h07f7;
  assign literal_9086[52] = 16'h0ff1;
  assign literal_9086[53] = 16'h7fc6;
  assign literal_9086[54] = 16'hff9c;
  assign literal_9086[55] = 16'hffa3;
  assign literal_9086[56] = 16'hffd7;
  assign literal_9086[57] = 16'hffe4;
  assign literal_9086[58] = 16'hfff2;
  assign literal_9086[59] = 16'h0000;
  assign literal_9086[60] = 16'h0000;
  assign literal_9086[61] = 16'h0000;
  assign literal_9086[62] = 16'h0000;
  assign literal_9086[63] = 16'h0000;
  assign literal_9086[64] = 16'h0000;
  assign literal_9086[65] = 16'h003a;
  assign literal_9086[66] = 16'h03f8;
  assign literal_9086[67] = 16'h0ff2;
  assign literal_9086[68] = 16'h7fc8;
  assign literal_9086[69] = 16'hff9d;
  assign literal_9086[70] = 16'hffbf;
  assign literal_9086[71] = 16'hffcb;
  assign literal_9086[72] = 16'hffd8;
  assign literal_9086[73] = 16'hffe5;
  assign literal_9086[74] = 16'hfff3;
  assign literal_9086[75] = 16'h0000;
  assign literal_9086[76] = 16'h0000;
  assign literal_9086[77] = 16'h0000;
  assign literal_9086[78] = 16'h0000;
  assign literal_9086[79] = 16'h0000;
  assign literal_9086[80] = 16'h0000;
  assign literal_9086[81] = 16'h0077;
  assign literal_9086[82] = 16'h07f3;
  assign literal_9086[83] = 16'h1fea;
  assign literal_9086[84] = 16'hff94;
  assign literal_9086[85] = 16'hffa2;
  assign literal_9086[86] = 16'hffc0;
  assign literal_9086[87] = 16'hffcc;
  assign literal_9086[88] = 16'hffd9;
  assign literal_9086[89] = 16'hffe6;
  assign literal_9086[90] = 16'hfff4;
  assign literal_9086[91] = 16'h0000;
  assign literal_9086[92] = 16'h0000;
  assign literal_9086[93] = 16'h0000;
  assign literal_9086[94] = 16'h0000;
  assign literal_9086[95] = 16'h0000;
  assign literal_9086[96] = 16'h0000;
  assign literal_9086[97] = 16'h0079;
  assign literal_9086[98] = 16'h07f4;
  assign literal_9086[99] = 16'h1fed;
  assign literal_9086[100] = 16'hffa0;
  assign literal_9086[101] = 16'hffb5;
  assign literal_9086[102] = 16'hffc1;
  assign literal_9086[103] = 16'hffcd;
  assign literal_9086[104] = 16'hffda;
  assign literal_9086[105] = 16'hffe7;
  assign literal_9086[106] = 16'hfff5;
  assign literal_9086[107] = 16'h0000;
  assign literal_9086[108] = 16'h0000;
  assign literal_9086[109] = 16'h0000;
  assign literal_9086[110] = 16'h0000;
  assign literal_9086[111] = 16'h0000;
  assign literal_9086[112] = 16'h0000;
  assign literal_9086[113] = 16'h00f7;
  assign literal_9086[114] = 16'h07f5;
  assign literal_9086[115] = 16'h3fe1;
  assign literal_9086[116] = 16'hffa1;
  assign literal_9086[117] = 16'hffb6;
  assign literal_9086[118] = 16'hffc2;
  assign literal_9086[119] = 16'hffce;
  assign literal_9086[120] = 16'hffdb;
  assign literal_9086[121] = 16'hffe8;
  assign literal_9086[122] = 16'hfff6;
  assign literal_9086[123] = 16'h0000;
  assign literal_9086[124] = 16'h0000;
  assign literal_9086[125] = 16'h0000;
  assign literal_9086[126] = 16'h0000;
  assign literal_9086[127] = 16'h0000;
  assign literal_9086[128] = 16'h0000;
  assign literal_9086[129] = 16'h00f8;
  assign literal_9086[130] = 16'h0ff3;
  assign literal_9086[131] = 16'hff92;
  assign literal_9086[132] = 16'hffad;
  assign literal_9086[133] = 16'hffb7;
  assign literal_9086[134] = 16'hffc3;
  assign literal_9086[135] = 16'hffcf;
  assign literal_9086[136] = 16'hffdc;
  assign literal_9086[137] = 16'hffe9;
  assign literal_9086[138] = 16'hfff7;
  assign literal_9086[139] = 16'h0000;
  assign literal_9086[140] = 16'h0000;
  assign literal_9086[141] = 16'h0000;
  assign literal_9086[142] = 16'h0000;
  assign literal_9086[143] = 16'h0000;
  assign literal_9086[144] = 16'h0000;
  assign literal_9086[145] = 16'h00f9;
  assign literal_9086[146] = 16'h1fe9;
  assign literal_9086[147] = 16'hff95;
  assign literal_9086[148] = 16'hffae;
  assign literal_9086[149] = 16'hffb8;
  assign literal_9086[150] = 16'hffc4;
  assign literal_9086[151] = 16'hffd0;
  assign literal_9086[152] = 16'hffdd;
  assign literal_9086[153] = 16'hffea;
  assign literal_9086[154] = 16'hfff8;
  assign literal_9086[155] = 16'h0000;
  assign literal_9086[156] = 16'h0000;
  assign literal_9086[157] = 16'h0000;
  assign literal_9086[158] = 16'h0000;
  assign literal_9086[159] = 16'h0000;
  assign literal_9086[160] = 16'h0000;
  assign literal_9086[161] = 16'h01f6;
  assign literal_9086[162] = 16'h1fec;
  assign literal_9086[163] = 16'hffa5;
  assign literal_9086[164] = 16'hffaf;
  assign literal_9086[165] = 16'hffb9;
  assign literal_9086[166] = 16'hffc5;
  assign literal_9086[167] = 16'hffd1;
  assign literal_9086[168] = 16'hffde;
  assign literal_9086[169] = 16'hffeb;
  assign literal_9086[170] = 16'hfff9;
  assign literal_9086[171] = 16'h0000;
  assign literal_9086[172] = 16'h0000;
  assign literal_9086[173] = 16'h0000;
  assign literal_9086[174] = 16'h0000;
  assign literal_9086[175] = 16'h0000;
  assign literal_9086[176] = 16'h0000;
  assign literal_9086[177] = 16'h01f7;
  assign literal_9086[178] = 16'h1fee;
  assign literal_9086[179] = 16'hffa6;
  assign literal_9086[180] = 16'hffb0;
  assign literal_9086[181] = 16'hffba;
  assign literal_9086[182] = 16'hffc6;
  assign literal_9086[183] = 16'hffd2;
  assign literal_9086[184] = 16'hffdf;
  assign literal_9086[185] = 16'hffec;
  assign literal_9086[186] = 16'hfffa;
  assign literal_9086[187] = 16'h0000;
  assign literal_9086[188] = 16'h0000;
  assign literal_9086[189] = 16'h0000;
  assign literal_9086[190] = 16'h0000;
  assign literal_9086[191] = 16'h0000;
  assign literal_9086[192] = 16'h0000;
  assign literal_9086[193] = 16'h03f4;
  assign literal_9086[194] = 16'h1fef;
  assign literal_9086[195] = 16'hffa7;
  assign literal_9086[196] = 16'hffb1;
  assign literal_9086[197] = 16'hffbb;
  assign literal_9086[198] = 16'hffc7;
  assign literal_9086[199] = 16'hffd3;
  assign literal_9086[200] = 16'hffe0;
  assign literal_9086[201] = 16'hffed;
  assign literal_9086[202] = 16'hfffb;
  assign literal_9086[203] = 16'h0000;
  assign literal_9086[204] = 16'h0000;
  assign literal_9086[205] = 16'h0000;
  assign literal_9086[206] = 16'h0000;
  assign literal_9086[207] = 16'h0000;
  assign literal_9086[208] = 16'h0000;
  assign literal_9086[209] = 16'h03f5;
  assign literal_9086[210] = 16'h3fe2;
  assign literal_9086[211] = 16'hffaa;
  assign literal_9086[212] = 16'hffb2;
  assign literal_9086[213] = 16'hffbc;
  assign literal_9086[214] = 16'hffc8;
  assign literal_9086[215] = 16'hffd4;
  assign literal_9086[216] = 16'hffe1;
  assign literal_9086[217] = 16'hffee;
  assign literal_9086[218] = 16'hfffc;
  assign literal_9086[219] = 16'h0000;
  assign literal_9086[220] = 16'h0000;
  assign literal_9086[221] = 16'h0000;
  assign literal_9086[222] = 16'h0000;
  assign literal_9086[223] = 16'h0000;
  assign literal_9086[224] = 16'h0000;
  assign literal_9086[225] = 16'h03f6;
  assign literal_9086[226] = 16'h7fc7;
  assign literal_9086[227] = 16'hffab;
  assign literal_9086[228] = 16'hffb3;
  assign literal_9086[229] = 16'hffbd;
  assign literal_9086[230] = 16'hffc9;
  assign literal_9086[231] = 16'hffd5;
  assign literal_9086[232] = 16'hffe2;
  assign literal_9086[233] = 16'hffef;
  assign literal_9086[234] = 16'hfffd;
  assign literal_9086[235] = 16'h0000;
  assign literal_9086[236] = 16'h0000;
  assign literal_9086[237] = 16'h0000;
  assign literal_9086[238] = 16'h0000;
  assign literal_9086[239] = 16'h0000;
  assign literal_9086[240] = 16'h01f8;
  assign literal_9086[241] = 16'h07f6;
  assign literal_9086[242] = 16'hffa4;
  assign literal_9086[243] = 16'hffac;
  assign literal_9086[244] = 16'hffb4;
  assign literal_9086[245] = 16'hffbe;
  assign literal_9086[246] = 16'hffca;
  assign literal_9086[247] = 16'hffd6;
  assign literal_9086[248] = 16'hffe3;
  assign literal_9086[249] = 16'hfff0;
  assign literal_9086[250] = 16'hfffe;
  assign literal_9086[251] = 16'h0000;
  wire [15:0] literal_9087[0:251];
  assign literal_9087[0] = 16'h000c;
  assign literal_9087[1] = 16'h0000;
  assign literal_9087[2] = 16'h0001;
  assign literal_9087[3] = 16'h0004;
  assign literal_9087[4] = 16'h000b;
  assign literal_9087[5] = 16'h001a;
  assign literal_9087[6] = 16'h0079;
  assign literal_9087[7] = 16'h01f9;
  assign literal_9087[8] = 16'h0000;
  assign literal_9087[9] = 16'h0000;
  assign literal_9087[10] = 16'h0000;
  assign literal_9087[11] = 16'h0000;
  assign literal_9087[12] = 16'h0000;
  assign literal_9087[13] = 16'h0000;
  assign literal_9087[14] = 16'h0000;
  assign literal_9087[15] = 16'h0000;
  assign literal_9087[16] = 16'h0000;
  assign literal_9087[17] = 16'h000a;
  assign literal_9087[18] = 16'h001c;
  assign literal_9087[19] = 16'h007a;
  assign literal_9087[20] = 16'h01f5;
  assign literal_9087[21] = 16'h03f4;
  assign literal_9087[22] = 16'h07f8;
  assign literal_9087[23] = 16'hff95;
  assign literal_9087[24] = 16'h0000;
  assign literal_9087[25] = 16'h0000;
  assign literal_9087[26] = 16'h0000;
  assign literal_9087[27] = 16'h0000;
  assign literal_9087[28] = 16'h0000;
  assign literal_9087[29] = 16'h0000;
  assign literal_9087[30] = 16'h0000;
  assign literal_9087[31] = 16'h0000;
  assign literal_9087[32] = 16'h0000;
  assign literal_9087[33] = 16'h001b;
  assign literal_9087[34] = 16'h00f8;
  assign literal_9087[35] = 16'h03f7;
  assign literal_9087[36] = 16'h0ff4;
  assign literal_9087[37] = 16'h0000;
  assign literal_9087[38] = 16'h0000;
  assign literal_9087[39] = 16'h0000;
  assign literal_9087[40] = 16'h0000;
  assign literal_9087[41] = 16'h0000;
  assign literal_9087[42] = 16'h0000;
  assign literal_9087[43] = 16'h0000;
  assign literal_9087[44] = 16'h0000;
  assign literal_9087[45] = 16'h0000;
  assign literal_9087[46] = 16'h0000;
  assign literal_9087[47] = 16'h0000;
  assign literal_9087[48] = 16'h0000;
  assign literal_9087[49] = 16'h003a;
  assign literal_9087[50] = 16'h01f6;
  assign literal_9087[51] = 16'h0000;
  assign literal_9087[52] = 16'h0ff5;
  assign literal_9087[53] = 16'hff8e;
  assign literal_9087[54] = 16'hff96;
  assign literal_9087[55] = 16'hffc9;
  assign literal_9087[56] = 16'hffd6;
  assign literal_9087[57] = 16'hffe4;
  assign literal_9087[58] = 16'h0000;
  assign literal_9087[59] = 16'h0000;
  assign literal_9087[60] = 16'h0000;
  assign literal_9087[61] = 16'h0000;
  assign literal_9087[62] = 16'h0000;
  assign literal_9087[63] = 16'h0000;
  assign literal_9087[64] = 16'h0000;
  assign literal_9087[65] = 16'h003b;
  assign literal_9087[66] = 16'h03f6;
  assign literal_9087[67] = 16'hff5d;
  assign literal_9087[68] = 16'hff8f;
  assign literal_9087[69] = 16'hffa5;
  assign literal_9087[70] = 16'hffa6;
  assign literal_9087[71] = 16'hffca;
  assign literal_9087[72] = 16'hffd7;
  assign literal_9087[73] = 16'hfff3;
  assign literal_9087[74] = 16'h0000;
  assign literal_9087[75] = 16'h0000;
  assign literal_9087[76] = 16'h0000;
  assign literal_9087[77] = 16'h0000;
  assign literal_9087[78] = 16'h0000;
  assign literal_9087[79] = 16'h0000;
  assign literal_9087[80] = 16'h0000;
  assign literal_9087[81] = 16'h0078;
  assign literal_9087[82] = 16'h03f9;
  assign literal_9087[83] = 16'hff5f;
  assign literal_9087[84] = 16'hff96;
  assign literal_9087[85] = 16'hffab;
  assign literal_9087[86] = 16'hffa9;
  assign literal_9087[87] = 16'hffcb;
  assign literal_9087[88] = 16'hffd7;
  assign literal_9087[89] = 16'hffe6;
  assign literal_9087[90] = 16'h0000;
  assign literal_9087[91] = 16'h0000;
  assign literal_9087[92] = 16'h0000;
  assign literal_9087[93] = 16'h0000;
  assign literal_9087[94] = 16'h0000;
  assign literal_9087[95] = 16'h0000;
  assign literal_9087[96] = 16'h0000;
  assign literal_9087[97] = 16'h007b;
  assign literal_9087[98] = 16'h0ff2;
  assign literal_9087[99] = 16'hff85;
  assign literal_9087[100] = 16'hff97;
  assign literal_9087[101] = 16'hffb5;
  assign literal_9087[102] = 16'hffbf;
  assign literal_9087[103] = 16'hffcc;
  assign literal_9087[104] = 16'hffd9;
  assign literal_9087[105] = 16'hffe7;
  assign literal_9087[106] = 16'hfff5;
  assign literal_9087[107] = 16'hfff5;
  assign literal_9087[108] = 16'h0000;
  assign literal_9087[109] = 16'h0000;
  assign literal_9087[110] = 16'h0000;
  assign literal_9087[111] = 16'h0000;
  assign literal_9087[112] = 16'h0000;
  assign literal_9087[113] = 16'h00f9;
  assign literal_9087[114] = 16'h0ff5;
  assign literal_9087[115] = 16'hff8c;
  assign literal_9087[116] = 16'hff98;
  assign literal_9087[117] = 16'hffb6;
  assign literal_9087[118] = 16'hffc0;
  assign literal_9087[119] = 16'hffcd;
  assign literal_9087[120] = 16'hffda;
  assign literal_9087[121] = 16'hffe8;
  assign literal_9087[122] = 16'hfff6;
  assign literal_9087[123] = 16'h0000;
  assign literal_9087[124] = 16'h0000;
  assign literal_9087[125] = 16'h0000;
  assign literal_9087[126] = 16'h0000;
  assign literal_9087[127] = 16'h0000;
  assign literal_9087[128] = 16'h0000;
  assign literal_9087[129] = 16'h01f4;
  assign literal_9087[130] = 16'h3fd4;
  assign literal_9087[131] = 16'hff9e;
  assign literal_9087[132] = 16'hffa3;
  assign literal_9087[133] = 16'h0000;
  assign literal_9087[134] = 16'hffc1;
  assign literal_9087[135] = 16'hffce;
  assign literal_9087[136] = 16'hffdb;
  assign literal_9087[137] = 16'hffe9;
  assign literal_9087[138] = 16'h0000;
  assign literal_9087[139] = 16'h0000;
  assign literal_9087[140] = 16'h0000;
  assign literal_9087[141] = 16'h0000;
  assign literal_9087[142] = 16'h0000;
  assign literal_9087[143] = 16'h0000;
  assign literal_9087[144] = 16'h0000;
  assign literal_9087[145] = 16'h01f7;
  assign literal_9087[146] = 16'h7fc0;
  assign literal_9087[147] = 16'hff91;
  assign literal_9087[148] = 16'hffa4;
  assign literal_9087[149] = 16'hffb8;
  assign literal_9087[150] = 16'hffc2;
  assign literal_9087[151] = 16'hffcf;
  assign literal_9087[152] = 16'hffdc;
  assign literal_9087[153] = 16'hffea;
  assign literal_9087[154] = 16'hfff8;
  assign literal_9087[155] = 16'h0000;
  assign literal_9087[156] = 16'h0000;
  assign literal_9087[157] = 16'h0000;
  assign literal_9087[158] = 16'h0000;
  assign literal_9087[159] = 16'h0000;
  assign literal_9087[160] = 16'h0000;
  assign literal_9087[161] = 16'h01f8;
  assign literal_9087[162] = 16'h7fc1;
  assign literal_9087[163] = 16'hff92;
  assign literal_9087[164] = 16'hffa7;
  assign literal_9087[165] = 16'hffb9;
  assign literal_9087[166] = 16'hffc3;
  assign literal_9087[167] = 16'hffd0;
  assign literal_9087[168] = 16'hffdd;
  assign literal_9087[169] = 16'hffeb;
  assign literal_9087[170] = 16'h0000;
  assign literal_9087[171] = 16'h0000;
  assign literal_9087[172] = 16'h0000;
  assign literal_9087[173] = 16'h0000;
  assign literal_9087[174] = 16'h0000;
  assign literal_9087[175] = 16'h0000;
  assign literal_9087[176] = 16'h0000;
  assign literal_9087[177] = 16'h03f5;
  assign literal_9087[178] = 16'hff84;
  assign literal_9087[179] = 16'hff93;
  assign literal_9087[180] = 16'hffa8;
  assign literal_9087[181] = 16'hffba;
  assign literal_9087[182] = 16'hffc4;
  assign literal_9087[183] = 16'hffd1;
  assign literal_9087[184] = 16'hffde;
  assign literal_9087[185] = 16'hffeb;
  assign literal_9087[186] = 16'h0000;
  assign literal_9087[187] = 16'h0000;
  assign literal_9087[188] = 16'h0000;
  assign literal_9087[189] = 16'h0000;
  assign literal_9087[190] = 16'h0000;
  assign literal_9087[191] = 16'h0000;
  assign literal_9087[192] = 16'h0000;
  assign literal_9087[193] = 16'h03f8;
  assign literal_9087[194] = 16'hff8d;
  assign literal_9087[195] = 16'hff99;
  assign literal_9087[196] = 16'hffb1;
  assign literal_9087[197] = 16'hffbb;
  assign literal_9087[198] = 16'hffc5;
  assign literal_9087[199] = 16'hffd2;
  assign literal_9087[200] = 16'hffdf;
  assign literal_9087[201] = 16'hffed;
  assign literal_9087[202] = 16'h0000;
  assign literal_9087[203] = 16'h0000;
  assign literal_9087[204] = 16'h0000;
  assign literal_9087[205] = 16'h0000;
  assign literal_9087[206] = 16'h0000;
  assign literal_9087[207] = 16'h0000;
  assign literal_9087[208] = 16'h0000;
  assign literal_9087[209] = 16'h03fa;
  assign literal_9087[210] = 16'hff9a;
  assign literal_9087[211] = 16'hffaa;
  assign literal_9087[212] = 16'hffb2;
  assign literal_9087[213] = 16'hffbc;
  assign literal_9087[214] = 16'hffc6;
  assign literal_9087[215] = 16'hffd3;
  assign literal_9087[216] = 16'hffe0;
  assign literal_9087[217] = 16'hffee;
  assign literal_9087[218] = 16'h0000;
  assign literal_9087[219] = 16'h0000;
  assign literal_9087[220] = 16'h0000;
  assign literal_9087[221] = 16'h0000;
  assign literal_9087[222] = 16'h0000;
  assign literal_9087[223] = 16'h0000;
  assign literal_9087[224] = 16'h0000;
  assign literal_9087[225] = 16'h07f6;
  assign literal_9087[226] = 16'hff9b;
  assign literal_9087[227] = 16'hffaf;
  assign literal_9087[228] = 16'hffb3;
  assign literal_9087[229] = 16'hffbd;
  assign literal_9087[230] = 16'hffc7;
  assign literal_9087[231] = 16'hffd4;
  assign literal_9087[232] = 16'hffe1;
  assign literal_9087[233] = 16'hffef;
  assign literal_9087[234] = 16'h0000;
  assign literal_9087[235] = 16'h0000;
  assign literal_9087[236] = 16'h0000;
  assign literal_9087[237] = 16'h0000;
  assign literal_9087[238] = 16'h0000;
  assign literal_9087[239] = 16'h0000;
  assign literal_9087[240] = 16'h0ff3;
  assign literal_9087[241] = 16'h3fd5;
  assign literal_9087[242] = 16'hffae;
  assign literal_9087[243] = 16'hffb0;
  assign literal_9087[244] = 16'hffb4;
  assign literal_9087[245] = 16'hffbe;
  assign literal_9087[246] = 16'hffc8;
  assign literal_9087[247] = 16'hffd5;
  assign literal_9087[248] = 16'hffe2;
  assign literal_9087[249] = 16'hfff0;
  assign literal_9087[250] = 16'hfffe;
  assign literal_9087[251] = 16'h0000;
  wire [7:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[7:0];
  assign matrix_unflattened[0][1] = matrix[15:8];
  assign matrix_unflattened[0][2] = matrix[23:16];
  assign matrix_unflattened[0][3] = matrix[31:24];
  assign matrix_unflattened[0][4] = matrix[39:32];
  assign matrix_unflattened[0][5] = matrix[47:40];
  assign matrix_unflattened[0][6] = matrix[55:48];
  assign matrix_unflattened[0][7] = matrix[63:56];
  assign matrix_unflattened[1][0] = matrix[71:64];
  assign matrix_unflattened[1][1] = matrix[79:72];
  assign matrix_unflattened[1][2] = matrix[87:80];
  assign matrix_unflattened[1][3] = matrix[95:88];
  assign matrix_unflattened[1][4] = matrix[103:96];
  assign matrix_unflattened[1][5] = matrix[111:104];
  assign matrix_unflattened[1][6] = matrix[119:112];
  assign matrix_unflattened[1][7] = matrix[127:120];
  assign matrix_unflattened[2][0] = matrix[135:128];
  assign matrix_unflattened[2][1] = matrix[143:136];
  assign matrix_unflattened[2][2] = matrix[151:144];
  assign matrix_unflattened[2][3] = matrix[159:152];
  assign matrix_unflattened[2][4] = matrix[167:160];
  assign matrix_unflattened[2][5] = matrix[175:168];
  assign matrix_unflattened[2][6] = matrix[183:176];
  assign matrix_unflattened[2][7] = matrix[191:184];
  assign matrix_unflattened[3][0] = matrix[199:192];
  assign matrix_unflattened[3][1] = matrix[207:200];
  assign matrix_unflattened[3][2] = matrix[215:208];
  assign matrix_unflattened[3][3] = matrix[223:216];
  assign matrix_unflattened[3][4] = matrix[231:224];
  assign matrix_unflattened[3][5] = matrix[239:232];
  assign matrix_unflattened[3][6] = matrix[247:240];
  assign matrix_unflattened[3][7] = matrix[255:248];
  assign matrix_unflattened[4][0] = matrix[263:256];
  assign matrix_unflattened[4][1] = matrix[271:264];
  assign matrix_unflattened[4][2] = matrix[279:272];
  assign matrix_unflattened[4][3] = matrix[287:280];
  assign matrix_unflattened[4][4] = matrix[295:288];
  assign matrix_unflattened[4][5] = matrix[303:296];
  assign matrix_unflattened[4][6] = matrix[311:304];
  assign matrix_unflattened[4][7] = matrix[319:312];
  assign matrix_unflattened[5][0] = matrix[327:320];
  assign matrix_unflattened[5][1] = matrix[335:328];
  assign matrix_unflattened[5][2] = matrix[343:336];
  assign matrix_unflattened[5][3] = matrix[351:344];
  assign matrix_unflattened[5][4] = matrix[359:352];
  assign matrix_unflattened[5][5] = matrix[367:360];
  assign matrix_unflattened[5][6] = matrix[375:368];
  assign matrix_unflattened[5][7] = matrix[383:376];
  assign matrix_unflattened[6][0] = matrix[391:384];
  assign matrix_unflattened[6][1] = matrix[399:392];
  assign matrix_unflattened[6][2] = matrix[407:400];
  assign matrix_unflattened[6][3] = matrix[415:408];
  assign matrix_unflattened[6][4] = matrix[423:416];
  assign matrix_unflattened[6][5] = matrix[431:424];
  assign matrix_unflattened[6][6] = matrix[439:432];
  assign matrix_unflattened[6][7] = matrix[447:440];
  assign matrix_unflattened[7][0] = matrix[455:448];
  assign matrix_unflattened[7][1] = matrix[463:456];
  assign matrix_unflattened[7][2] = matrix[471:464];
  assign matrix_unflattened[7][3] = matrix[479:472];
  assign matrix_unflattened[7][4] = matrix[487:480];
  assign matrix_unflattened[7][5] = matrix[495:488];
  assign matrix_unflattened[7][6] = matrix[503:496];
  assign matrix_unflattened[7][7] = matrix[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_row0_comb[0:7];
  wire [7:0] p1_row1_comb[0:7];
  wire [7:0] p1_array_concat_8212_comb[0:15];
  wire [7:0] p1_row2_comb[0:7];
  wire [7:0] p1_array_concat_8215_comb[0:23];
  wire [7:0] p1_row3_comb[0:7];
  wire [2:0] p1_idx_u8__4_squeezed_comb;
  wire [7:0] p1_array_concat_8218_comb[0:31];
  wire [7:0] p1_row4_comb[0:7];
  wire [2:0] p1_idx_u8__5_squeezed_comb;
  wire [7:0] p1_array_concat_8221_comb[0:39];
  wire [7:0] p1_row5_comb[0:7];
  wire [2:0] p1_idx_u8__6_squeezed_comb;
  wire [7:0] p1_idx_u8__13_comb;
  wire [7:0] p1_array_concat_8227_comb[0:47];
  wire [7:0] p1_row6_comb[0:7];
  wire [2:0] p1_idx_u8__7_squeezed_comb;
  wire [6:0] p1_add_8230_comb;
  wire [7:0] p1_actual_index__13_comb;
  wire [7:0] p1_array_concat_8234_comb[0:55];
  wire [7:0] p1_row7_comb[0:7];
  wire [5:0] p1_add_8239_comb;
  wire [7:0] p1_flat_comb[0:63];
  wire [7:0] p1_actual_index__14_comb;
  wire [7:0] p1_idx_u8__1_comb;
  wire [7:0] p1_idx_u8__3_comb;
  wire [7:0] p1_idx_u8__5_comb;
  wire [7:0] p1_idx_u8__7_comb;
  wire [7:0] p1_idx_u8__9_comb;
  wire [7:0] p1_idx_u8__11_comb;
  wire [7:0] p1_actual_index__12_comb;
  wire [7:0] p1_actual_index__1_comb;
  wire [6:0] p1_add_8350_comb;
  wire [7:0] p1_actual_index__3_comb;
  wire [5:0] p1_add_8333_comb;
  wire [7:0] p1_actual_index__5_comb;
  wire [6:0] p1_add_8316_comb;
  wire [7:0] p1_actual_index__7_comb;
  wire [7:0] p1_actual_index__9_comb;
  wire [6:0] p1_add_8263_comb;
  wire [7:0] p1_actual_index__11_comb;
  wire [7:0] p1_idx_u8__15_comb;
  wire [7:0] p1_idx_u8__17_comb;
  wire [7:0] p1_idx_u8__19_comb;
  wire [7:0] p1_idx_u8__21_comb;
  wire [7:0] p1_idx_u8__23_comb;
  wire [7:0] p1_idx_u8__25_comb;
  wire [7:0] p1_idx_u8__27_comb;
  wire [7:0] p1_idx_u8__29_comb;
  wire [7:0] p1_idx_u8__31_comb;
  wire [7:0] p1_idx_u8__33_comb;
  wire [7:0] p1_idx_u8__35_comb;
  wire [7:0] p1_idx_u8__37_comb;
  wire [7:0] p1_idx_u8__39_comb;
  wire [7:0] p1_idx_u8__41_comb;
  wire [7:0] p1_idx_u8__43_comb;
  wire [7:0] p1_idx_u8__45_comb;
  wire [7:0] p1_idx_u8__47_comb;
  wire [7:0] p1_idx_u8__49_comb;
  wire [7:0] p1_idx_u8__51_comb;
  wire [7:0] p1_idx_u8__53_comb;
  wire [7:0] p1_idx_u8__55_comb;
  wire [7:0] p1_idx_u8__57_comb;
  wire [7:0] p1_idx_u8__59_comb;
  wire [7:0] p1_idx_u8__61_comb;
  wire [7:0] p1_and_8258_comb;
  wire [4:0] p1_add_8282_comb;
  wire [7:0] p1_actual_index__15_comb;
  wire [3:0] p1_add_8453_comb;
  wire [7:0] p1_actual_index__17_comb;
  wire [6:0] p1_add_8455_comb;
  wire [7:0] p1_actual_index__19_comb;
  wire [5:0] p1_add_8457_comb;
  wire [7:0] p1_actual_index__21_comb;
  wire [6:0] p1_add_8459_comb;
  wire [7:0] p1_actual_index__23_comb;
  wire [4:0] p1_add_8461_comb;
  wire [7:0] p1_actual_index__25_comb;
  wire [6:0] p1_add_8463_comb;
  wire [7:0] p1_actual_index__27_comb;
  wire [5:0] p1_add_8465_comb;
  wire [7:0] p1_actual_index__29_comb;
  wire [6:0] p1_add_8467_comb;
  wire [7:0] p1_actual_index__31_comb;
  wire [2:0] p1_add_8469_comb;
  wire [7:0] p1_actual_index__33_comb;
  wire [6:0] p1_add_8471_comb;
  wire [7:0] p1_actual_index__35_comb;
  wire [5:0] p1_add_8473_comb;
  wire [7:0] p1_actual_index__37_comb;
  wire [6:0] p1_add_8475_comb;
  wire [7:0] p1_actual_index__39_comb;
  wire [4:0] p1_add_8477_comb;
  wire [7:0] p1_actual_index__41_comb;
  wire [6:0] p1_add_8479_comb;
  wire [7:0] p1_actual_index__43_comb;
  wire [5:0] p1_add_8481_comb;
  wire [7:0] p1_actual_index__45_comb;
  wire [6:0] p1_add_8483_comb;
  wire [7:0] p1_actual_index__47_comb;
  wire [3:0] p1_add_8485_comb;
  wire [7:0] p1_actual_index__49_comb;
  wire [6:0] p1_add_8487_comb;
  wire [7:0] p1_actual_index__51_comb;
  wire [5:0] p1_add_8489_comb;
  wire [7:0] p1_actual_index__53_comb;
  wire [6:0] p1_add_8491_comb;
  wire [7:0] p1_actual_index__55_comb;
  wire [4:0] p1_add_8493_comb;
  wire [7:0] p1_actual_index__57_comb;
  wire [6:0] p1_add_8495_comb;
  wire [7:0] p1_actual_index__59_comb;
  wire [5:0] p1_add_8497_comb;
  wire [7:0] p1_actual_index__61_comb;
  wire [6:0] p1_add_8499_comb;
  wire [7:0] p1_and_8266_comb;
  wire p1_eq_8269_comb;
  wire [7:0] p1_and_8270_comb;
  wire [7:0] p1_actual_index__2_comb;
  wire [7:0] p1_actual_index__4_comb;
  wire [7:0] p1_actual_index__6_comb;
  wire [7:0] p1_actual_index__10_comb;
  wire p1_ne_8278_comb;
  wire [1:0] p1_idx_u8__1_squeezed_comb;
  wire p1_eq_8281_comb;
  wire [7:0] p1_actual_index__8_comb;
  wire [7:0] p1_actual_index__16_comb;
  wire [7:0] p1_actual_index__18_comb;
  wire [7:0] p1_actual_index__20_comb;
  wire [7:0] p1_actual_index__22_comb;
  wire [7:0] p1_actual_index__24_comb;
  wire [7:0] p1_actual_index__26_comb;
  wire [7:0] p1_actual_index__28_comb;
  wire [7:0] p1_actual_index__30_comb;
  wire [7:0] p1_actual_index__32_comb;
  wire [7:0] p1_actual_index__34_comb;
  wire [7:0] p1_actual_index__36_comb;
  wire [7:0] p1_actual_index__38_comb;
  wire [7:0] p1_actual_index__40_comb;
  wire [7:0] p1_actual_index__42_comb;
  wire [7:0] p1_actual_index__44_comb;
  wire [7:0] p1_actual_index__46_comb;
  wire [7:0] p1_actual_index__48_comb;
  wire [7:0] p1_actual_index__50_comb;
  wire [7:0] p1_actual_index__52_comb;
  wire [7:0] p1_actual_index__54_comb;
  wire [7:0] p1_actual_index__56_comb;
  wire [7:0] p1_actual_index__58_comb;
  wire [7:0] p1_actual_index__60_comb;
  wire [7:0] p1_actual_index__62_comb;
  wire [7:0] p1_and_8394_comb;
  wire [7:0] p1_and_8396_comb;
  wire [7:0] p1_and_8391_comb;
  wire [7:0] p1_and_8384_comb;
  wire [7:0] p1_and_8377_comb;
  wire [7:0] p1_and_8366_comb;
  wire [7:0] p1_and_8357_comb;
  wire [7:0] p1_and_8347_comb;
  wire [7:0] p1_and_8319_comb;
  wire [7:0] p1_and_8308_comb;
  wire [7:0] p1_and_8298_comb;
  wire p1_ne_8399_comb;
  wire p1_ne_8400_comb;
  wire p1_ne_8398_comb;
  wire p1_ne_8393_comb;
  wire p1_ne_8386_comb;
  wire p1_ne_8379_comb;
  wire p1_ne_8368_comb;
  wire p1_ne_8359_comb;
  wire [7:0] p1_and_8323_comb;
  wire p1_ne_8330_comb;
  wire p1_ne_8321_comb;
  wire p1_ne_8310_comb;
  wire p1_not_8401_comb;
  wire p1_eq_8331_comb;
  wire [2:0] p1_sel_8322_comb;
  wire p1_and_8921_comb;
  wire [7:0] p1_value_comb;
  assign p1_row0_comb[0] = p0_matrix[3'h0][0];
  assign p1_row0_comb[1] = p0_matrix[3'h0][1];
  assign p1_row0_comb[2] = p0_matrix[3'h0][2];
  assign p1_row0_comb[3] = p0_matrix[3'h0][3];
  assign p1_row0_comb[4] = p0_matrix[3'h0][4];
  assign p1_row0_comb[5] = p0_matrix[3'h0][5];
  assign p1_row0_comb[6] = p0_matrix[3'h0][6];
  assign p1_row0_comb[7] = p0_matrix[3'h0][7];
  assign p1_row1_comb[0] = p0_matrix[3'h1][0];
  assign p1_row1_comb[1] = p0_matrix[3'h1][1];
  assign p1_row1_comb[2] = p0_matrix[3'h1][2];
  assign p1_row1_comb[3] = p0_matrix[3'h1][3];
  assign p1_row1_comb[4] = p0_matrix[3'h1][4];
  assign p1_row1_comb[5] = p0_matrix[3'h1][5];
  assign p1_row1_comb[6] = p0_matrix[3'h1][6];
  assign p1_row1_comb[7] = p0_matrix[3'h1][7];
  assign p1_array_concat_8212_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_8212_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_8212_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_8212_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_8212_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_8212_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_8212_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_8212_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_8212_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_8212_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_8212_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_8212_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_8212_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_8212_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_8212_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_8212_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_8215_comb[0] = p1_array_concat_8212_comb[0];
  assign p1_array_concat_8215_comb[1] = p1_array_concat_8212_comb[1];
  assign p1_array_concat_8215_comb[2] = p1_array_concat_8212_comb[2];
  assign p1_array_concat_8215_comb[3] = p1_array_concat_8212_comb[3];
  assign p1_array_concat_8215_comb[4] = p1_array_concat_8212_comb[4];
  assign p1_array_concat_8215_comb[5] = p1_array_concat_8212_comb[5];
  assign p1_array_concat_8215_comb[6] = p1_array_concat_8212_comb[6];
  assign p1_array_concat_8215_comb[7] = p1_array_concat_8212_comb[7];
  assign p1_array_concat_8215_comb[8] = p1_array_concat_8212_comb[8];
  assign p1_array_concat_8215_comb[9] = p1_array_concat_8212_comb[9];
  assign p1_array_concat_8215_comb[10] = p1_array_concat_8212_comb[10];
  assign p1_array_concat_8215_comb[11] = p1_array_concat_8212_comb[11];
  assign p1_array_concat_8215_comb[12] = p1_array_concat_8212_comb[12];
  assign p1_array_concat_8215_comb[13] = p1_array_concat_8212_comb[13];
  assign p1_array_concat_8215_comb[14] = p1_array_concat_8212_comb[14];
  assign p1_array_concat_8215_comb[15] = p1_array_concat_8212_comb[15];
  assign p1_array_concat_8215_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_8215_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_8215_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_8215_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_8215_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_8215_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_8215_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_8215_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_idx_u8__4_squeezed_comb = 3'h4;
  assign p1_array_concat_8218_comb[0] = p1_array_concat_8215_comb[0];
  assign p1_array_concat_8218_comb[1] = p1_array_concat_8215_comb[1];
  assign p1_array_concat_8218_comb[2] = p1_array_concat_8215_comb[2];
  assign p1_array_concat_8218_comb[3] = p1_array_concat_8215_comb[3];
  assign p1_array_concat_8218_comb[4] = p1_array_concat_8215_comb[4];
  assign p1_array_concat_8218_comb[5] = p1_array_concat_8215_comb[5];
  assign p1_array_concat_8218_comb[6] = p1_array_concat_8215_comb[6];
  assign p1_array_concat_8218_comb[7] = p1_array_concat_8215_comb[7];
  assign p1_array_concat_8218_comb[8] = p1_array_concat_8215_comb[8];
  assign p1_array_concat_8218_comb[9] = p1_array_concat_8215_comb[9];
  assign p1_array_concat_8218_comb[10] = p1_array_concat_8215_comb[10];
  assign p1_array_concat_8218_comb[11] = p1_array_concat_8215_comb[11];
  assign p1_array_concat_8218_comb[12] = p1_array_concat_8215_comb[12];
  assign p1_array_concat_8218_comb[13] = p1_array_concat_8215_comb[13];
  assign p1_array_concat_8218_comb[14] = p1_array_concat_8215_comb[14];
  assign p1_array_concat_8218_comb[15] = p1_array_concat_8215_comb[15];
  assign p1_array_concat_8218_comb[16] = p1_array_concat_8215_comb[16];
  assign p1_array_concat_8218_comb[17] = p1_array_concat_8215_comb[17];
  assign p1_array_concat_8218_comb[18] = p1_array_concat_8215_comb[18];
  assign p1_array_concat_8218_comb[19] = p1_array_concat_8215_comb[19];
  assign p1_array_concat_8218_comb[20] = p1_array_concat_8215_comb[20];
  assign p1_array_concat_8218_comb[21] = p1_array_concat_8215_comb[21];
  assign p1_array_concat_8218_comb[22] = p1_array_concat_8215_comb[22];
  assign p1_array_concat_8218_comb[23] = p1_array_concat_8215_comb[23];
  assign p1_array_concat_8218_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_8218_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_8218_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_8218_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_8218_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_8218_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_8218_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_8218_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[p1_idx_u8__4_squeezed_comb][0];
  assign p1_row4_comb[1] = p0_matrix[p1_idx_u8__4_squeezed_comb][1];
  assign p1_row4_comb[2] = p0_matrix[p1_idx_u8__4_squeezed_comb][2];
  assign p1_row4_comb[3] = p0_matrix[p1_idx_u8__4_squeezed_comb][3];
  assign p1_row4_comb[4] = p0_matrix[p1_idx_u8__4_squeezed_comb][4];
  assign p1_row4_comb[5] = p0_matrix[p1_idx_u8__4_squeezed_comb][5];
  assign p1_row4_comb[6] = p0_matrix[p1_idx_u8__4_squeezed_comb][6];
  assign p1_row4_comb[7] = p0_matrix[p1_idx_u8__4_squeezed_comb][7];
  assign p1_idx_u8__5_squeezed_comb = 3'h5;
  assign p1_array_concat_8221_comb[0] = p1_array_concat_8218_comb[0];
  assign p1_array_concat_8221_comb[1] = p1_array_concat_8218_comb[1];
  assign p1_array_concat_8221_comb[2] = p1_array_concat_8218_comb[2];
  assign p1_array_concat_8221_comb[3] = p1_array_concat_8218_comb[3];
  assign p1_array_concat_8221_comb[4] = p1_array_concat_8218_comb[4];
  assign p1_array_concat_8221_comb[5] = p1_array_concat_8218_comb[5];
  assign p1_array_concat_8221_comb[6] = p1_array_concat_8218_comb[6];
  assign p1_array_concat_8221_comb[7] = p1_array_concat_8218_comb[7];
  assign p1_array_concat_8221_comb[8] = p1_array_concat_8218_comb[8];
  assign p1_array_concat_8221_comb[9] = p1_array_concat_8218_comb[9];
  assign p1_array_concat_8221_comb[10] = p1_array_concat_8218_comb[10];
  assign p1_array_concat_8221_comb[11] = p1_array_concat_8218_comb[11];
  assign p1_array_concat_8221_comb[12] = p1_array_concat_8218_comb[12];
  assign p1_array_concat_8221_comb[13] = p1_array_concat_8218_comb[13];
  assign p1_array_concat_8221_comb[14] = p1_array_concat_8218_comb[14];
  assign p1_array_concat_8221_comb[15] = p1_array_concat_8218_comb[15];
  assign p1_array_concat_8221_comb[16] = p1_array_concat_8218_comb[16];
  assign p1_array_concat_8221_comb[17] = p1_array_concat_8218_comb[17];
  assign p1_array_concat_8221_comb[18] = p1_array_concat_8218_comb[18];
  assign p1_array_concat_8221_comb[19] = p1_array_concat_8218_comb[19];
  assign p1_array_concat_8221_comb[20] = p1_array_concat_8218_comb[20];
  assign p1_array_concat_8221_comb[21] = p1_array_concat_8218_comb[21];
  assign p1_array_concat_8221_comb[22] = p1_array_concat_8218_comb[22];
  assign p1_array_concat_8221_comb[23] = p1_array_concat_8218_comb[23];
  assign p1_array_concat_8221_comb[24] = p1_array_concat_8218_comb[24];
  assign p1_array_concat_8221_comb[25] = p1_array_concat_8218_comb[25];
  assign p1_array_concat_8221_comb[26] = p1_array_concat_8218_comb[26];
  assign p1_array_concat_8221_comb[27] = p1_array_concat_8218_comb[27];
  assign p1_array_concat_8221_comb[28] = p1_array_concat_8218_comb[28];
  assign p1_array_concat_8221_comb[29] = p1_array_concat_8218_comb[29];
  assign p1_array_concat_8221_comb[30] = p1_array_concat_8218_comb[30];
  assign p1_array_concat_8221_comb[31] = p1_array_concat_8218_comb[31];
  assign p1_array_concat_8221_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_8221_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_8221_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_8221_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_8221_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_8221_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_8221_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_8221_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[p1_idx_u8__5_squeezed_comb][0];
  assign p1_row5_comb[1] = p0_matrix[p1_idx_u8__5_squeezed_comb][1];
  assign p1_row5_comb[2] = p0_matrix[p1_idx_u8__5_squeezed_comb][2];
  assign p1_row5_comb[3] = p0_matrix[p1_idx_u8__5_squeezed_comb][3];
  assign p1_row5_comb[4] = p0_matrix[p1_idx_u8__5_squeezed_comb][4];
  assign p1_row5_comb[5] = p0_matrix[p1_idx_u8__5_squeezed_comb][5];
  assign p1_row5_comb[6] = p0_matrix[p1_idx_u8__5_squeezed_comb][6];
  assign p1_row5_comb[7] = p0_matrix[p1_idx_u8__5_squeezed_comb][7];
  assign p1_idx_u8__6_squeezed_comb = 3'h6;
  assign p1_idx_u8__13_comb = 8'h0d;
  assign p1_array_concat_8227_comb[0] = p1_array_concat_8221_comb[0];
  assign p1_array_concat_8227_comb[1] = p1_array_concat_8221_comb[1];
  assign p1_array_concat_8227_comb[2] = p1_array_concat_8221_comb[2];
  assign p1_array_concat_8227_comb[3] = p1_array_concat_8221_comb[3];
  assign p1_array_concat_8227_comb[4] = p1_array_concat_8221_comb[4];
  assign p1_array_concat_8227_comb[5] = p1_array_concat_8221_comb[5];
  assign p1_array_concat_8227_comb[6] = p1_array_concat_8221_comb[6];
  assign p1_array_concat_8227_comb[7] = p1_array_concat_8221_comb[7];
  assign p1_array_concat_8227_comb[8] = p1_array_concat_8221_comb[8];
  assign p1_array_concat_8227_comb[9] = p1_array_concat_8221_comb[9];
  assign p1_array_concat_8227_comb[10] = p1_array_concat_8221_comb[10];
  assign p1_array_concat_8227_comb[11] = p1_array_concat_8221_comb[11];
  assign p1_array_concat_8227_comb[12] = p1_array_concat_8221_comb[12];
  assign p1_array_concat_8227_comb[13] = p1_array_concat_8221_comb[13];
  assign p1_array_concat_8227_comb[14] = p1_array_concat_8221_comb[14];
  assign p1_array_concat_8227_comb[15] = p1_array_concat_8221_comb[15];
  assign p1_array_concat_8227_comb[16] = p1_array_concat_8221_comb[16];
  assign p1_array_concat_8227_comb[17] = p1_array_concat_8221_comb[17];
  assign p1_array_concat_8227_comb[18] = p1_array_concat_8221_comb[18];
  assign p1_array_concat_8227_comb[19] = p1_array_concat_8221_comb[19];
  assign p1_array_concat_8227_comb[20] = p1_array_concat_8221_comb[20];
  assign p1_array_concat_8227_comb[21] = p1_array_concat_8221_comb[21];
  assign p1_array_concat_8227_comb[22] = p1_array_concat_8221_comb[22];
  assign p1_array_concat_8227_comb[23] = p1_array_concat_8221_comb[23];
  assign p1_array_concat_8227_comb[24] = p1_array_concat_8221_comb[24];
  assign p1_array_concat_8227_comb[25] = p1_array_concat_8221_comb[25];
  assign p1_array_concat_8227_comb[26] = p1_array_concat_8221_comb[26];
  assign p1_array_concat_8227_comb[27] = p1_array_concat_8221_comb[27];
  assign p1_array_concat_8227_comb[28] = p1_array_concat_8221_comb[28];
  assign p1_array_concat_8227_comb[29] = p1_array_concat_8221_comb[29];
  assign p1_array_concat_8227_comb[30] = p1_array_concat_8221_comb[30];
  assign p1_array_concat_8227_comb[31] = p1_array_concat_8221_comb[31];
  assign p1_array_concat_8227_comb[32] = p1_array_concat_8221_comb[32];
  assign p1_array_concat_8227_comb[33] = p1_array_concat_8221_comb[33];
  assign p1_array_concat_8227_comb[34] = p1_array_concat_8221_comb[34];
  assign p1_array_concat_8227_comb[35] = p1_array_concat_8221_comb[35];
  assign p1_array_concat_8227_comb[36] = p1_array_concat_8221_comb[36];
  assign p1_array_concat_8227_comb[37] = p1_array_concat_8221_comb[37];
  assign p1_array_concat_8227_comb[38] = p1_array_concat_8221_comb[38];
  assign p1_array_concat_8227_comb[39] = p1_array_concat_8221_comb[39];
  assign p1_array_concat_8227_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_8227_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_8227_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_8227_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_8227_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_8227_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_8227_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_8227_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[p1_idx_u8__6_squeezed_comb][0];
  assign p1_row6_comb[1] = p0_matrix[p1_idx_u8__6_squeezed_comb][1];
  assign p1_row6_comb[2] = p0_matrix[p1_idx_u8__6_squeezed_comb][2];
  assign p1_row6_comb[3] = p0_matrix[p1_idx_u8__6_squeezed_comb][3];
  assign p1_row6_comb[4] = p0_matrix[p1_idx_u8__6_squeezed_comb][4];
  assign p1_row6_comb[5] = p0_matrix[p1_idx_u8__6_squeezed_comb][5];
  assign p1_row6_comb[6] = p0_matrix[p1_idx_u8__6_squeezed_comb][6];
  assign p1_row6_comb[7] = p0_matrix[p1_idx_u8__6_squeezed_comb][7];
  assign p1_idx_u8__7_squeezed_comb = 3'h7;
  assign p1_add_8230_comb = p0_start_pix[7:1] + 7'h07;
  assign p1_actual_index__13_comb = p0_start_pix + p1_idx_u8__13_comb;
  assign p1_array_concat_8234_comb[0] = p1_array_concat_8227_comb[0];
  assign p1_array_concat_8234_comb[1] = p1_array_concat_8227_comb[1];
  assign p1_array_concat_8234_comb[2] = p1_array_concat_8227_comb[2];
  assign p1_array_concat_8234_comb[3] = p1_array_concat_8227_comb[3];
  assign p1_array_concat_8234_comb[4] = p1_array_concat_8227_comb[4];
  assign p1_array_concat_8234_comb[5] = p1_array_concat_8227_comb[5];
  assign p1_array_concat_8234_comb[6] = p1_array_concat_8227_comb[6];
  assign p1_array_concat_8234_comb[7] = p1_array_concat_8227_comb[7];
  assign p1_array_concat_8234_comb[8] = p1_array_concat_8227_comb[8];
  assign p1_array_concat_8234_comb[9] = p1_array_concat_8227_comb[9];
  assign p1_array_concat_8234_comb[10] = p1_array_concat_8227_comb[10];
  assign p1_array_concat_8234_comb[11] = p1_array_concat_8227_comb[11];
  assign p1_array_concat_8234_comb[12] = p1_array_concat_8227_comb[12];
  assign p1_array_concat_8234_comb[13] = p1_array_concat_8227_comb[13];
  assign p1_array_concat_8234_comb[14] = p1_array_concat_8227_comb[14];
  assign p1_array_concat_8234_comb[15] = p1_array_concat_8227_comb[15];
  assign p1_array_concat_8234_comb[16] = p1_array_concat_8227_comb[16];
  assign p1_array_concat_8234_comb[17] = p1_array_concat_8227_comb[17];
  assign p1_array_concat_8234_comb[18] = p1_array_concat_8227_comb[18];
  assign p1_array_concat_8234_comb[19] = p1_array_concat_8227_comb[19];
  assign p1_array_concat_8234_comb[20] = p1_array_concat_8227_comb[20];
  assign p1_array_concat_8234_comb[21] = p1_array_concat_8227_comb[21];
  assign p1_array_concat_8234_comb[22] = p1_array_concat_8227_comb[22];
  assign p1_array_concat_8234_comb[23] = p1_array_concat_8227_comb[23];
  assign p1_array_concat_8234_comb[24] = p1_array_concat_8227_comb[24];
  assign p1_array_concat_8234_comb[25] = p1_array_concat_8227_comb[25];
  assign p1_array_concat_8234_comb[26] = p1_array_concat_8227_comb[26];
  assign p1_array_concat_8234_comb[27] = p1_array_concat_8227_comb[27];
  assign p1_array_concat_8234_comb[28] = p1_array_concat_8227_comb[28];
  assign p1_array_concat_8234_comb[29] = p1_array_concat_8227_comb[29];
  assign p1_array_concat_8234_comb[30] = p1_array_concat_8227_comb[30];
  assign p1_array_concat_8234_comb[31] = p1_array_concat_8227_comb[31];
  assign p1_array_concat_8234_comb[32] = p1_array_concat_8227_comb[32];
  assign p1_array_concat_8234_comb[33] = p1_array_concat_8227_comb[33];
  assign p1_array_concat_8234_comb[34] = p1_array_concat_8227_comb[34];
  assign p1_array_concat_8234_comb[35] = p1_array_concat_8227_comb[35];
  assign p1_array_concat_8234_comb[36] = p1_array_concat_8227_comb[36];
  assign p1_array_concat_8234_comb[37] = p1_array_concat_8227_comb[37];
  assign p1_array_concat_8234_comb[38] = p1_array_concat_8227_comb[38];
  assign p1_array_concat_8234_comb[39] = p1_array_concat_8227_comb[39];
  assign p1_array_concat_8234_comb[40] = p1_array_concat_8227_comb[40];
  assign p1_array_concat_8234_comb[41] = p1_array_concat_8227_comb[41];
  assign p1_array_concat_8234_comb[42] = p1_array_concat_8227_comb[42];
  assign p1_array_concat_8234_comb[43] = p1_array_concat_8227_comb[43];
  assign p1_array_concat_8234_comb[44] = p1_array_concat_8227_comb[44];
  assign p1_array_concat_8234_comb[45] = p1_array_concat_8227_comb[45];
  assign p1_array_concat_8234_comb[46] = p1_array_concat_8227_comb[46];
  assign p1_array_concat_8234_comb[47] = p1_array_concat_8227_comb[47];
  assign p1_array_concat_8234_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_8234_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_8234_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_8234_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_8234_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_8234_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_8234_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_8234_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[p1_idx_u8__7_squeezed_comb][0];
  assign p1_row7_comb[1] = p0_matrix[p1_idx_u8__7_squeezed_comb][1];
  assign p1_row7_comb[2] = p0_matrix[p1_idx_u8__7_squeezed_comb][2];
  assign p1_row7_comb[3] = p0_matrix[p1_idx_u8__7_squeezed_comb][3];
  assign p1_row7_comb[4] = p0_matrix[p1_idx_u8__7_squeezed_comb][4];
  assign p1_row7_comb[5] = p0_matrix[p1_idx_u8__7_squeezed_comb][5];
  assign p1_row7_comb[6] = p0_matrix[p1_idx_u8__7_squeezed_comb][6];
  assign p1_row7_comb[7] = p0_matrix[p1_idx_u8__7_squeezed_comb][7];
  assign p1_add_8239_comb = p0_start_pix[7:2] + 6'h03;
  assign p1_flat_comb[0] = p1_array_concat_8234_comb[0];
  assign p1_flat_comb[1] = p1_array_concat_8234_comb[1];
  assign p1_flat_comb[2] = p1_array_concat_8234_comb[2];
  assign p1_flat_comb[3] = p1_array_concat_8234_comb[3];
  assign p1_flat_comb[4] = p1_array_concat_8234_comb[4];
  assign p1_flat_comb[5] = p1_array_concat_8234_comb[5];
  assign p1_flat_comb[6] = p1_array_concat_8234_comb[6];
  assign p1_flat_comb[7] = p1_array_concat_8234_comb[7];
  assign p1_flat_comb[8] = p1_array_concat_8234_comb[8];
  assign p1_flat_comb[9] = p1_array_concat_8234_comb[9];
  assign p1_flat_comb[10] = p1_array_concat_8234_comb[10];
  assign p1_flat_comb[11] = p1_array_concat_8234_comb[11];
  assign p1_flat_comb[12] = p1_array_concat_8234_comb[12];
  assign p1_flat_comb[13] = p1_array_concat_8234_comb[13];
  assign p1_flat_comb[14] = p1_array_concat_8234_comb[14];
  assign p1_flat_comb[15] = p1_array_concat_8234_comb[15];
  assign p1_flat_comb[16] = p1_array_concat_8234_comb[16];
  assign p1_flat_comb[17] = p1_array_concat_8234_comb[17];
  assign p1_flat_comb[18] = p1_array_concat_8234_comb[18];
  assign p1_flat_comb[19] = p1_array_concat_8234_comb[19];
  assign p1_flat_comb[20] = p1_array_concat_8234_comb[20];
  assign p1_flat_comb[21] = p1_array_concat_8234_comb[21];
  assign p1_flat_comb[22] = p1_array_concat_8234_comb[22];
  assign p1_flat_comb[23] = p1_array_concat_8234_comb[23];
  assign p1_flat_comb[24] = p1_array_concat_8234_comb[24];
  assign p1_flat_comb[25] = p1_array_concat_8234_comb[25];
  assign p1_flat_comb[26] = p1_array_concat_8234_comb[26];
  assign p1_flat_comb[27] = p1_array_concat_8234_comb[27];
  assign p1_flat_comb[28] = p1_array_concat_8234_comb[28];
  assign p1_flat_comb[29] = p1_array_concat_8234_comb[29];
  assign p1_flat_comb[30] = p1_array_concat_8234_comb[30];
  assign p1_flat_comb[31] = p1_array_concat_8234_comb[31];
  assign p1_flat_comb[32] = p1_array_concat_8234_comb[32];
  assign p1_flat_comb[33] = p1_array_concat_8234_comb[33];
  assign p1_flat_comb[34] = p1_array_concat_8234_comb[34];
  assign p1_flat_comb[35] = p1_array_concat_8234_comb[35];
  assign p1_flat_comb[36] = p1_array_concat_8234_comb[36];
  assign p1_flat_comb[37] = p1_array_concat_8234_comb[37];
  assign p1_flat_comb[38] = p1_array_concat_8234_comb[38];
  assign p1_flat_comb[39] = p1_array_concat_8234_comb[39];
  assign p1_flat_comb[40] = p1_array_concat_8234_comb[40];
  assign p1_flat_comb[41] = p1_array_concat_8234_comb[41];
  assign p1_flat_comb[42] = p1_array_concat_8234_comb[42];
  assign p1_flat_comb[43] = p1_array_concat_8234_comb[43];
  assign p1_flat_comb[44] = p1_array_concat_8234_comb[44];
  assign p1_flat_comb[45] = p1_array_concat_8234_comb[45];
  assign p1_flat_comb[46] = p1_array_concat_8234_comb[46];
  assign p1_flat_comb[47] = p1_array_concat_8234_comb[47];
  assign p1_flat_comb[48] = p1_array_concat_8234_comb[48];
  assign p1_flat_comb[49] = p1_array_concat_8234_comb[49];
  assign p1_flat_comb[50] = p1_array_concat_8234_comb[50];
  assign p1_flat_comb[51] = p1_array_concat_8234_comb[51];
  assign p1_flat_comb[52] = p1_array_concat_8234_comb[52];
  assign p1_flat_comb[53] = p1_array_concat_8234_comb[53];
  assign p1_flat_comb[54] = p1_array_concat_8234_comb[54];
  assign p1_flat_comb[55] = p1_array_concat_8234_comb[55];
  assign p1_flat_comb[56] = p1_row7_comb[0];
  assign p1_flat_comb[57] = p1_row7_comb[1];
  assign p1_flat_comb[58] = p1_row7_comb[2];
  assign p1_flat_comb[59] = p1_row7_comb[3];
  assign p1_flat_comb[60] = p1_row7_comb[4];
  assign p1_flat_comb[61] = p1_row7_comb[5];
  assign p1_flat_comb[62] = p1_row7_comb[6];
  assign p1_flat_comb[63] = p1_row7_comb[7];
  assign p1_actual_index__14_comb = {p1_add_8230_comb, p0_start_pix[0]};
  assign p1_idx_u8__1_comb = 8'h01;
  assign p1_idx_u8__3_comb = 8'h03;
  assign p1_idx_u8__5_comb = 8'h05;
  assign p1_idx_u8__7_comb = 8'h07;
  assign p1_idx_u8__9_comb = 8'h09;
  assign p1_idx_u8__11_comb = 8'h0b;
  assign p1_actual_index__12_comb = {p1_add_8239_comb, p0_start_pix[1:0]};
  assign p1_actual_index__1_comb = p0_start_pix + p1_idx_u8__1_comb;
  assign p1_add_8350_comb = p0_start_pix[7:1] + 7'h01;
  assign p1_actual_index__3_comb = p0_start_pix + p1_idx_u8__3_comb;
  assign p1_add_8333_comb = p0_start_pix[7:2] + 6'h01;
  assign p1_actual_index__5_comb = p0_start_pix + p1_idx_u8__5_comb;
  assign p1_add_8316_comb = p0_start_pix[7:1] + 7'h03;
  assign p1_actual_index__7_comb = p0_start_pix + p1_idx_u8__7_comb;
  assign p1_actual_index__9_comb = p0_start_pix + p1_idx_u8__9_comb;
  assign p1_add_8263_comb = p0_start_pix[7:1] + 7'h05;
  assign p1_actual_index__11_comb = p0_start_pix + p1_idx_u8__11_comb;
  assign p1_idx_u8__15_comb = 8'h0f;
  assign p1_idx_u8__17_comb = 8'h11;
  assign p1_idx_u8__19_comb = 8'h13;
  assign p1_idx_u8__21_comb = 8'h15;
  assign p1_idx_u8__23_comb = 8'h17;
  assign p1_idx_u8__25_comb = 8'h19;
  assign p1_idx_u8__27_comb = 8'h1b;
  assign p1_idx_u8__29_comb = 8'h1d;
  assign p1_idx_u8__31_comb = 8'h1f;
  assign p1_idx_u8__33_comb = 8'h21;
  assign p1_idx_u8__35_comb = 8'h23;
  assign p1_idx_u8__37_comb = 8'h25;
  assign p1_idx_u8__39_comb = 8'h27;
  assign p1_idx_u8__41_comb = 8'h29;
  assign p1_idx_u8__43_comb = 8'h2b;
  assign p1_idx_u8__45_comb = 8'h2d;
  assign p1_idx_u8__47_comb = 8'h2f;
  assign p1_idx_u8__49_comb = 8'h31;
  assign p1_idx_u8__51_comb = 8'h33;
  assign p1_idx_u8__53_comb = 8'h35;
  assign p1_idx_u8__55_comb = 8'h37;
  assign p1_idx_u8__57_comb = 8'h39;
  assign p1_idx_u8__59_comb = 8'h3b;
  assign p1_idx_u8__61_comb = 8'h3d;
  assign p1_and_8258_comb = p1_flat_comb[p1_actual_index__14_comb > 8'h3f ? 6'h3f : p1_actual_index__14_comb[5:0]] & {8{~(p1_add_8230_comb[5] | p1_add_8230_comb[6])}};
  assign p1_add_8282_comb = p0_start_pix[7:3] + 5'h01;
  assign p1_actual_index__15_comb = p0_start_pix + p1_idx_u8__15_comb;
  assign p1_add_8453_comb = p0_start_pix[7:4] + 4'h1;
  assign p1_actual_index__17_comb = p0_start_pix + p1_idx_u8__17_comb;
  assign p1_add_8455_comb = p0_start_pix[7:1] + 7'h09;
  assign p1_actual_index__19_comb = p0_start_pix + p1_idx_u8__19_comb;
  assign p1_add_8457_comb = p0_start_pix[7:2] + 6'h05;
  assign p1_actual_index__21_comb = p0_start_pix + p1_idx_u8__21_comb;
  assign p1_add_8459_comb = p0_start_pix[7:1] + 7'h0b;
  assign p1_actual_index__23_comb = p0_start_pix + p1_idx_u8__23_comb;
  assign p1_add_8461_comb = p0_start_pix[7:3] + 5'h03;
  assign p1_actual_index__25_comb = p0_start_pix + p1_idx_u8__25_comb;
  assign p1_add_8463_comb = p0_start_pix[7:1] + 7'h0d;
  assign p1_actual_index__27_comb = p0_start_pix + p1_idx_u8__27_comb;
  assign p1_add_8465_comb = p0_start_pix[7:2] + 6'h07;
  assign p1_actual_index__29_comb = p0_start_pix + p1_idx_u8__29_comb;
  assign p1_add_8467_comb = p0_start_pix[7:1] + 7'h0f;
  assign p1_actual_index__31_comb = p0_start_pix + p1_idx_u8__31_comb;
  assign p1_add_8469_comb = p0_start_pix[7:5] + 3'h1;
  assign p1_actual_index__33_comb = p0_start_pix + p1_idx_u8__33_comb;
  assign p1_add_8471_comb = p0_start_pix[7:1] + 7'h11;
  assign p1_actual_index__35_comb = p0_start_pix + p1_idx_u8__35_comb;
  assign p1_add_8473_comb = p0_start_pix[7:2] + 6'h09;
  assign p1_actual_index__37_comb = p0_start_pix + p1_idx_u8__37_comb;
  assign p1_add_8475_comb = p0_start_pix[7:1] + 7'h13;
  assign p1_actual_index__39_comb = p0_start_pix + p1_idx_u8__39_comb;
  assign p1_add_8477_comb = p0_start_pix[7:3] + 5'h05;
  assign p1_actual_index__41_comb = p0_start_pix + p1_idx_u8__41_comb;
  assign p1_add_8479_comb = p0_start_pix[7:1] + 7'h15;
  assign p1_actual_index__43_comb = p0_start_pix + p1_idx_u8__43_comb;
  assign p1_add_8481_comb = p0_start_pix[7:2] + 6'h0b;
  assign p1_actual_index__45_comb = p0_start_pix + p1_idx_u8__45_comb;
  assign p1_add_8483_comb = p0_start_pix[7:1] + 7'h17;
  assign p1_actual_index__47_comb = p0_start_pix + p1_idx_u8__47_comb;
  assign p1_add_8485_comb = p0_start_pix[7:4] + 4'h3;
  assign p1_actual_index__49_comb = p0_start_pix + p1_idx_u8__49_comb;
  assign p1_add_8487_comb = p0_start_pix[7:1] + 7'h19;
  assign p1_actual_index__51_comb = p0_start_pix + p1_idx_u8__51_comb;
  assign p1_add_8489_comb = p0_start_pix[7:2] + 6'h0d;
  assign p1_actual_index__53_comb = p0_start_pix + p1_idx_u8__53_comb;
  assign p1_add_8491_comb = p0_start_pix[7:1] + 7'h1b;
  assign p1_actual_index__55_comb = p0_start_pix + p1_idx_u8__55_comb;
  assign p1_add_8493_comb = p0_start_pix[7:3] + 5'h07;
  assign p1_actual_index__57_comb = p0_start_pix + p1_idx_u8__57_comb;
  assign p1_add_8495_comb = p0_start_pix[7:1] + 7'h1d;
  assign p1_actual_index__59_comb = p0_start_pix + p1_idx_u8__59_comb;
  assign p1_add_8497_comb = p0_start_pix[7:2] + 6'h0f;
  assign p1_actual_index__61_comb = p0_start_pix + p1_idx_u8__61_comb;
  assign p1_add_8499_comb = p0_start_pix[7:1] + 7'h1f;
  assign p1_and_8266_comb = p1_flat_comb[p1_actual_index__13_comb > 8'h3f ? 6'h3f : p1_actual_index__13_comb[5:0]] & {8{~(p1_actual_index__13_comb[6] | p1_actual_index__13_comb[7])}};
  assign p1_eq_8269_comb = p1_and_8258_comb == 8'h00;
  assign p1_and_8270_comb = p1_flat_comb[p1_actual_index__12_comb > 8'h3f ? 6'h3f : p1_actual_index__12_comb[5:0]] & {8{~(p1_add_8239_comb[4] | p1_add_8239_comb[5])}};
  assign p1_actual_index__2_comb = {p1_add_8350_comb, p0_start_pix[0]};
  assign p1_actual_index__4_comb = {p1_add_8333_comb, p0_start_pix[1:0]};
  assign p1_actual_index__6_comb = {p1_add_8316_comb, p0_start_pix[0]};
  assign p1_actual_index__10_comb = {p1_add_8263_comb, p0_start_pix[0]};
  assign p1_ne_8278_comb = p1_and_8266_comb != 8'h00;
  assign p1_idx_u8__1_squeezed_comb = 2'h1;
  assign p1_eq_8281_comb = p1_and_8270_comb == 8'h00;
  assign p1_actual_index__8_comb = {p1_add_8282_comb, p0_start_pix[2:0]};
  assign p1_actual_index__16_comb = {p1_add_8453_comb, p0_start_pix[3:0]};
  assign p1_actual_index__18_comb = {p1_add_8455_comb, p0_start_pix[0]};
  assign p1_actual_index__20_comb = {p1_add_8457_comb, p0_start_pix[1:0]};
  assign p1_actual_index__22_comb = {p1_add_8459_comb, p0_start_pix[0]};
  assign p1_actual_index__24_comb = {p1_add_8461_comb, p0_start_pix[2:0]};
  assign p1_actual_index__26_comb = {p1_add_8463_comb, p0_start_pix[0]};
  assign p1_actual_index__28_comb = {p1_add_8465_comb, p0_start_pix[1:0]};
  assign p1_actual_index__30_comb = {p1_add_8467_comb, p0_start_pix[0]};
  assign p1_actual_index__32_comb = {p1_add_8469_comb, p0_start_pix[4:0]};
  assign p1_actual_index__34_comb = {p1_add_8471_comb, p0_start_pix[0]};
  assign p1_actual_index__36_comb = {p1_add_8473_comb, p0_start_pix[1:0]};
  assign p1_actual_index__38_comb = {p1_add_8475_comb, p0_start_pix[0]};
  assign p1_actual_index__40_comb = {p1_add_8477_comb, p0_start_pix[2:0]};
  assign p1_actual_index__42_comb = {p1_add_8479_comb, p0_start_pix[0]};
  assign p1_actual_index__44_comb = {p1_add_8481_comb, p0_start_pix[1:0]};
  assign p1_actual_index__46_comb = {p1_add_8483_comb, p0_start_pix[0]};
  assign p1_actual_index__48_comb = {p1_add_8485_comb, p0_start_pix[3:0]};
  assign p1_actual_index__50_comb = {p1_add_8487_comb, p0_start_pix[0]};
  assign p1_actual_index__52_comb = {p1_add_8489_comb, p0_start_pix[1:0]};
  assign p1_actual_index__54_comb = {p1_add_8491_comb, p0_start_pix[0]};
  assign p1_actual_index__56_comb = {p1_add_8493_comb, p0_start_pix[2:0]};
  assign p1_actual_index__58_comb = {p1_add_8495_comb, p0_start_pix[0]};
  assign p1_actual_index__60_comb = {p1_add_8497_comb, p0_start_pix[1:0]};
  assign p1_actual_index__62_comb = {p1_add_8499_comb, p0_start_pix[0]};
  assign p1_and_8394_comb = p1_flat_comb[p0_start_pix > 8'h3f ? 6'h3f : p0_start_pix[5:0]] & {8{~(p0_start_pix[6] | p0_start_pix[7])}};
  assign p1_and_8396_comb = p1_flat_comb[p1_actual_index__1_comb > 8'h3f ? 6'h3f : p1_actual_index__1_comb[5:0]] & {8{~(p1_actual_index__1_comb[6] | p1_actual_index__1_comb[7])}};
  assign p1_and_8391_comb = p1_flat_comb[p1_actual_index__2_comb > 8'h3f ? 6'h3f : p1_actual_index__2_comb[5:0]] & {8{~(p1_add_8350_comb[5] | p1_add_8350_comb[6])}};
  assign p1_and_8384_comb = p1_flat_comb[p1_actual_index__3_comb > 8'h3f ? 6'h3f : p1_actual_index__3_comb[5:0]] & {8{~(p1_actual_index__3_comb[6] | p1_actual_index__3_comb[7])}};
  assign p1_and_8377_comb = p1_flat_comb[p1_actual_index__4_comb > 8'h3f ? 6'h3f : p1_actual_index__4_comb[5:0]] & {8{~(p1_add_8333_comb[4] | p1_add_8333_comb[5])}};
  assign p1_and_8366_comb = p1_flat_comb[p1_actual_index__5_comb > 8'h3f ? 6'h3f : p1_actual_index__5_comb[5:0]] & {8{~(p1_actual_index__5_comb[6] | p1_actual_index__5_comb[7])}};
  assign p1_and_8357_comb = p1_flat_comb[p1_actual_index__6_comb > 8'h3f ? 6'h3f : p1_actual_index__6_comb[5:0]] & {8{~(p1_add_8316_comb[5] | p1_add_8316_comb[6])}};
  assign p1_and_8347_comb = p1_flat_comb[p1_actual_index__7_comb > 8'h3f ? 6'h3f : p1_actual_index__7_comb[5:0]] & {8{~(p1_actual_index__7_comb[6] | p1_actual_index__7_comb[7])}};
  assign p1_and_8319_comb = p1_flat_comb[p1_actual_index__9_comb > 8'h3f ? 6'h3f : p1_actual_index__9_comb[5:0]] & {8{~(p1_actual_index__9_comb[6] | p1_actual_index__9_comb[7])}};
  assign p1_and_8308_comb = p1_flat_comb[p1_actual_index__10_comb > 8'h3f ? 6'h3f : p1_actual_index__10_comb[5:0]] & {8{~(p1_add_8263_comb[5] | p1_add_8263_comb[6])}};
  assign p1_and_8298_comb = p1_flat_comb[p1_actual_index__11_comb > 8'h3f ? 6'h3f : p1_actual_index__11_comb[5:0]] & {8{~(p1_actual_index__11_comb[6] | p1_actual_index__11_comb[7])}};
  assign p1_ne_8399_comb = p1_and_8394_comb != 8'h00;
  assign p1_ne_8400_comb = p1_and_8396_comb != 8'h00;
  assign p1_ne_8398_comb = p1_and_8391_comb != 8'h00;
  assign p1_ne_8393_comb = p1_and_8384_comb != 8'h00;
  assign p1_ne_8386_comb = p1_and_8377_comb != 8'h00;
  assign p1_ne_8379_comb = p1_and_8366_comb != 8'h00;
  assign p1_ne_8368_comb = p1_and_8357_comb != 8'h00;
  assign p1_ne_8359_comb = p1_and_8347_comb != 8'h00;
  assign p1_and_8323_comb = p1_flat_comb[p1_actual_index__8_comb > 8'h3f ? 6'h3f : p1_actual_index__8_comb[5:0]] & {8{~(p1_add_8282_comb[3] | p1_add_8282_comb[4])}};
  assign p1_ne_8330_comb = p1_and_8319_comb != 8'h00;
  assign p1_ne_8321_comb = p1_and_8308_comb != 8'h00;
  assign p1_ne_8310_comb = p1_and_8298_comb != 8'h00;
  assign p1_not_8401_comb = ~p1_ne_8399_comb;
  assign p1_eq_8331_comb = p1_and_8323_comb == 8'h00;
  assign p1_sel_8322_comb = p1_ne_8310_comb ? 3'h3 : {1'h1, (p1_ne_8278_comb ? p1_idx_u8__1_squeezed_comb : {1'h1, p1_eq_8269_comb}) & {2{p1_eq_8281_comb}}};
  assign p1_and_8921_comb = p1_not_8401_comb & ~p1_ne_8400_comb & ~p1_ne_8398_comb & ~p1_ne_8393_comb & ~p1_ne_8386_comb & ~p1_ne_8379_comb & ~p1_ne_8368_comb & ~p1_ne_8359_comb & p1_eq_8331_comb & ~p1_ne_8330_comb & ~p1_ne_8321_comb & ~p1_ne_8310_comb & p1_eq_8281_comb & ~p1_ne_8278_comb & p1_eq_8269_comb & (p1_flat_comb[p1_actual_index__15_comb > 8'h3f ? 6'h3f : p1_actual_index__15_comb[5:0]] & {8{~(p1_actual_index__15_comb[6] | p1_actual_index__15_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__16_comb > 8'h3f ? 6'h3f : p1_actual_index__16_comb[5:0]] & {8{~(p1_add_8453_comb[2] | p1_add_8453_comb[3])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__17_comb > 8'h3f ? 6'h3f : p1_actual_index__17_comb[5:0]] & {8{~(p1_actual_index__17_comb[6] | p1_actual_index__17_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__18_comb > 8'h3f ? 6'h3f : p1_actual_index__18_comb[5:0]] & {8{~(p1_add_8455_comb[5] | p1_add_8455_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__19_comb > 8'h3f ? 6'h3f : p1_actual_index__19_comb[5:0]] & {8{~(p1_actual_index__19_comb[6] | p1_actual_index__19_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__20_comb > 8'h3f ? 6'h3f : p1_actual_index__20_comb[5:0]] & {8{~(p1_add_8457_comb[4] | p1_add_8457_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__21_comb > 8'h3f ? 6'h3f : p1_actual_index__21_comb[5:0]] & {8{~(p1_actual_index__21_comb[6] | p1_actual_index__21_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__22_comb > 8'h3f ? 6'h3f : p1_actual_index__22_comb[5:0]] & {8{~(p1_add_8459_comb[5] | p1_add_8459_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__23_comb > 8'h3f ? 6'h3f : p1_actual_index__23_comb[5:0]] & {8{~(p1_actual_index__23_comb[6] | p1_actual_index__23_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__24_comb > 8'h3f ? 6'h3f : p1_actual_index__24_comb[5:0]] & {8{~(p1_add_8461_comb[3] | p1_add_8461_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__25_comb > 8'h3f ? 6'h3f : p1_actual_index__25_comb[5:0]] & {8{~(p1_actual_index__25_comb[6] | p1_actual_index__25_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__26_comb > 8'h3f ? 6'h3f : p1_actual_index__26_comb[5:0]] & {8{~(p1_add_8463_comb[5] | p1_add_8463_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__27_comb > 8'h3f ? 6'h3f : p1_actual_index__27_comb[5:0]] & {8{~(p1_actual_index__27_comb[6] | p1_actual_index__27_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__28_comb > 8'h3f ? 6'h3f : p1_actual_index__28_comb[5:0]] & {8{~(p1_add_8465_comb[4] | p1_add_8465_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__29_comb > 8'h3f ? 6'h3f : p1_actual_index__29_comb[5:0]] & {8{~(p1_actual_index__29_comb[6] | p1_actual_index__29_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__30_comb > 8'h3f ? 6'h3f : p1_actual_index__30_comb[5:0]] & {8{~(p1_add_8467_comb[5] | p1_add_8467_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__31_comb > 8'h3f ? 6'h3f : p1_actual_index__31_comb[5:0]] & {8{~(p1_actual_index__31_comb[6] | p1_actual_index__31_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__32_comb > 8'h3f ? 6'h3f : p1_actual_index__32_comb[5:0]] & {8{~(p1_add_8469_comb[1] | p1_add_8469_comb[2])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__33_comb > 8'h3f ? 6'h3f : p1_actual_index__33_comb[5:0]] & {8{~(p1_actual_index__33_comb[6] | p1_actual_index__33_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__34_comb > 8'h3f ? 6'h3f : p1_actual_index__34_comb[5:0]] & {8{~(p1_add_8471_comb[5] | p1_add_8471_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__35_comb > 8'h3f ? 6'h3f : p1_actual_index__35_comb[5:0]] & {8{~(p1_actual_index__35_comb[6] | p1_actual_index__35_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__36_comb > 8'h3f ? 6'h3f : p1_actual_index__36_comb[5:0]] & {8{~(p1_add_8473_comb[4] | p1_add_8473_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__37_comb > 8'h3f ? 6'h3f : p1_actual_index__37_comb[5:0]] & {8{~(p1_actual_index__37_comb[6] | p1_actual_index__37_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__38_comb > 8'h3f ? 6'h3f : p1_actual_index__38_comb[5:0]] & {8{~(p1_add_8475_comb[5] | p1_add_8475_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__39_comb > 8'h3f ? 6'h3f : p1_actual_index__39_comb[5:0]] & {8{~(p1_actual_index__39_comb[6] | p1_actual_index__39_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__40_comb > 8'h3f ? 6'h3f : p1_actual_index__40_comb[5:0]] & {8{~(p1_add_8477_comb[3] | p1_add_8477_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__41_comb > 8'h3f ? 6'h3f : p1_actual_index__41_comb[5:0]] & {8{~(p1_actual_index__41_comb[6] | p1_actual_index__41_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__42_comb > 8'h3f ? 6'h3f : p1_actual_index__42_comb[5:0]] & {8{~(p1_add_8479_comb[5] | p1_add_8479_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__43_comb > 8'h3f ? 6'h3f : p1_actual_index__43_comb[5:0]] & {8{~(p1_actual_index__43_comb[6] | p1_actual_index__43_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__44_comb > 8'h3f ? 6'h3f : p1_actual_index__44_comb[5:0]] & {8{~(p1_add_8481_comb[4] | p1_add_8481_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__45_comb > 8'h3f ? 6'h3f : p1_actual_index__45_comb[5:0]] & {8{~(p1_actual_index__45_comb[6] | p1_actual_index__45_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__46_comb > 8'h3f ? 6'h3f : p1_actual_index__46_comb[5:0]] & {8{~(p1_add_8483_comb[5] | p1_add_8483_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__47_comb > 8'h3f ? 6'h3f : p1_actual_index__47_comb[5:0]] & {8{~(p1_actual_index__47_comb[6] | p1_actual_index__47_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__48_comb > 8'h3f ? 6'h3f : p1_actual_index__48_comb[5:0]] & {8{~(p1_add_8485_comb[2] | p1_add_8485_comb[3])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__49_comb > 8'h3f ? 6'h3f : p1_actual_index__49_comb[5:0]] & {8{~(p1_actual_index__49_comb[6] | p1_actual_index__49_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__50_comb > 8'h3f ? 6'h3f : p1_actual_index__50_comb[5:0]] & {8{~(p1_add_8487_comb[5] | p1_add_8487_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__51_comb > 8'h3f ? 6'h3f : p1_actual_index__51_comb[5:0]] & {8{~(p1_actual_index__51_comb[6] | p1_actual_index__51_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__52_comb > 8'h3f ? 6'h3f : p1_actual_index__52_comb[5:0]] & {8{~(p1_add_8489_comb[4] | p1_add_8489_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__53_comb > 8'h3f ? 6'h3f : p1_actual_index__53_comb[5:0]] & {8{~(p1_actual_index__53_comb[6] | p1_actual_index__53_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__54_comb > 8'h3f ? 6'h3f : p1_actual_index__54_comb[5:0]] & {8{~(p1_add_8491_comb[5] | p1_add_8491_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__55_comb > 8'h3f ? 6'h3f : p1_actual_index__55_comb[5:0]] & {8{~(p1_actual_index__55_comb[6] | p1_actual_index__55_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__56_comb > 8'h3f ? 6'h3f : p1_actual_index__56_comb[5:0]] & {8{~(p1_add_8493_comb[3] | p1_add_8493_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__57_comb > 8'h3f ? 6'h3f : p1_actual_index__57_comb[5:0]] & {8{~(p1_actual_index__57_comb[6] | p1_actual_index__57_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__58_comb > 8'h3f ? 6'h3f : p1_actual_index__58_comb[5:0]] & {8{~(p1_add_8495_comb[5] | p1_add_8495_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__59_comb > 8'h3f ? 6'h3f : p1_actual_index__59_comb[5:0]] & {8{~(p1_actual_index__59_comb[6] | p1_actual_index__59_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__60_comb > 8'h3f ? 6'h3f : p1_actual_index__60_comb[5:0]] & {8{~(p1_add_8497_comb[4] | p1_add_8497_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__61_comb > 8'h3f ? 6'h3f : p1_actual_index__61_comb[5:0]] & {8{~(p1_actual_index__61_comb[6] | p1_actual_index__61_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__62_comb > 8'h3f ? 6'h3f : p1_actual_index__62_comb[5:0]] & {8{~(p1_add_8499_comb[5] | p1_add_8499_comb[6])}}) == 8'h00;
  assign p1_value_comb = p0_matrix[3'h0][3'h0];

  // Registers for pipe stage 1:
  reg p1_is_luminance;
  reg [7:0] p1_and_8258;
  reg [7:0] p1_and_8266;
  reg [7:0] p1_and_8270;
  reg [7:0] p1_and_8298;
  reg [7:0] p1_and_8308;
  reg [7:0] p1_and_8319;
  reg p1_ne_8321;
  reg [2:0] p1_sel_8322;
  reg [7:0] p1_and_8323;
  reg p1_ne_8330;
  reg p1_eq_8331;
  reg [7:0] p1_and_8347;
  reg [7:0] p1_and_8357;
  reg p1_ne_8359;
  reg [7:0] p1_and_8366;
  reg p1_ne_8368;
  reg [7:0] p1_and_8377;
  reg p1_ne_8379;
  reg [7:0] p1_and_8384;
  reg p1_ne_8386;
  reg [7:0] p1_and_8391;
  reg p1_ne_8393;
  reg [7:0] p1_and_8394;
  reg [7:0] p1_and_8396;
  reg p1_ne_8398;
  reg p1_ne_8399;
  reg p1_ne_8400;
  reg p1_not_8401;
  reg p1_and_8921;
  reg [7:0] p1_value;
  always @ (posedge clk) begin
    p1_is_luminance <= p0_is_luminance;
    p1_and_8258 <= p1_and_8258_comb;
    p1_and_8266 <= p1_and_8266_comb;
    p1_and_8270 <= p1_and_8270_comb;
    p1_and_8298 <= p1_and_8298_comb;
    p1_and_8308 <= p1_and_8308_comb;
    p1_and_8319 <= p1_and_8319_comb;
    p1_ne_8321 <= p1_ne_8321_comb;
    p1_sel_8322 <= p1_sel_8322_comb;
    p1_and_8323 <= p1_and_8323_comb;
    p1_ne_8330 <= p1_ne_8330_comb;
    p1_eq_8331 <= p1_eq_8331_comb;
    p1_and_8347 <= p1_and_8347_comb;
    p1_and_8357 <= p1_and_8357_comb;
    p1_ne_8359 <= p1_ne_8359_comb;
    p1_and_8366 <= p1_and_8366_comb;
    p1_ne_8368 <= p1_ne_8368_comb;
    p1_and_8377 <= p1_and_8377_comb;
    p1_ne_8379 <= p1_ne_8379_comb;
    p1_and_8384 <= p1_and_8384_comb;
    p1_ne_8386 <= p1_ne_8386_comb;
    p1_and_8391 <= p1_and_8391_comb;
    p1_ne_8393 <= p1_ne_8393_comb;
    p1_and_8394 <= p1_and_8394_comb;
    p1_and_8396 <= p1_and_8396_comb;
    p1_ne_8398 <= p1_ne_8398_comb;
    p1_ne_8399 <= p1_ne_8399_comb;
    p1_ne_8400 <= p1_ne_8400_comb;
    p1_not_8401 <= p1_not_8401_comb;
    p1_and_8921 <= p1_and_8921_comb;
    p1_value <= p1_value_comb;
  end

  // ===== Pipe stage 2:
  wire [3:0] p2_sel_8996_comb;
  wire [3:0] p2_sel_9004_comb;
  wire [3:0] p2_sel_9008_comb;
  wire [3:0] p2_run_comb;
  wire [7:0] p2_value__1_comb;
  wire p2_eq_9026_comb;
  wire [1:0] p2_idx_u8__1_squeezed__1_comb;
  wire [1:0] p2_idx_u8__2_squeezed_comb;
  wire [3:0] p2_add_9023_comb;
  wire p2_or_reduce_9018_comb;
  wire [1:0] p2_sel_9019_comb;
  wire [3:0] p2_run_u8__1_comb;
  wire [3:0] p2_and_9029_comb;
  assign p2_sel_8996_comb = p1_ne_8359 ? 4'h7 : {1'h1, (p1_ne_8330 ? 3'h1 : (p1_ne_8321 ? 3'h2 : p1_sel_8322)) & {3{p1_eq_8331}}};
  assign p2_sel_9004_comb = p1_ne_8393 ? 4'h3 : (p1_ne_8386 ? 4'h4 : (p1_ne_8379 ? 4'h5 : (p1_ne_8368 ? 4'h6 : p2_sel_8996_comb)));
  assign p2_sel_9008_comb = p1_ne_8400 ? 4'h1 : (p1_ne_8398 ? 4'h2 : p2_sel_9004_comb);
  assign p2_run_comb = p2_sel_9008_comb & {4{p1_not_8401}};
  assign p2_value__1_comb = p2_run_comb == 4'h0 ? p1_and_8394 : (p2_run_comb == 4'h1 ? p1_and_8396 : (p2_run_comb == 4'h2 ? p1_and_8391 : (p2_run_comb == 4'h3 ? p1_and_8384 : (p2_run_comb == 4'h4 ? p1_and_8377 : (p2_run_comb == 4'h5 ? p1_and_8366 : (p2_run_comb == 4'h6 ? p1_and_8357 : (p2_run_comb == 4'h7 ? p1_and_8347 : (p2_run_comb == 4'h8 ? p1_and_8323 : (p2_run_comb == 4'h9 ? p1_and_8319 : (p2_run_comb == 4'ha ? p1_and_8308 : (p2_run_comb == 4'hb ? p1_and_8298 : (p2_run_comb == 4'hc ? p1_and_8270 : (p2_run_comb == 4'hd ? p1_and_8266 : (p2_run_comb == 4'he ? p1_and_8258 : 8'h00))))))))))))));
  assign p2_eq_9026_comb = p2_run_comb == 4'hf;
  assign p2_idx_u8__1_squeezed__1_comb = 2'h1;
  assign p2_idx_u8__2_squeezed_comb = 2'h2;
  assign p2_add_9023_comb = p2_sel_9004_comb + 4'h7;
  assign p2_or_reduce_9018_comb = |p2_value__1_comb[7:2];
  assign p2_sel_9019_comb = |p2_value__1_comb[7:1] ? p2_idx_u8__2_squeezed_comb : p2_idx_u8__1_squeezed__1_comb;
  assign p2_run_u8__1_comb = p2_run_comb < 4'ha ? p2_run_comb : p2_add_9023_comb;
  assign p2_and_9029_comb = p2_sel_9008_comb & {4{~(p2_eq_9026_comb | p1_ne_8399)}};

  // Registers for pipe stage 2:
  reg p2_is_luminance;
  reg [7:0] p2_value__1;
  reg p2_or_reduce_9018;
  reg [1:0] p2_sel_9019;
  reg [3:0] p2_run_u8__1;
  reg p2_and_8921;
  reg p2_eq_9026;
  reg [7:0] p2_value;
  reg [3:0] p2_and_9029;
  always @ (posedge clk) begin
    p2_is_luminance <= p1_is_luminance;
    p2_value__1 <= p2_value__1_comb;
    p2_or_reduce_9018 <= p2_or_reduce_9018_comb;
    p2_sel_9019 <= p2_sel_9019_comb;
    p2_run_u8__1 <= p2_run_u8__1_comb;
    p2_and_8921 <= p1_and_8921;
    p2_eq_9026 <= p2_eq_9026_comb;
    p2_value <= p1_value;
    p2_and_9029 <= p2_and_9029_comb;
  end

  // ===== Pipe stage 3:
  wire [1:0] p3_idx_u8__3_squeezed_comb;
  wire [2:0] p3_idx_u8__4_squeezed__1_comb;
  wire [2:0] p3_idx_u8__5_squeezed__1_comb;
  wire [2:0] p3_idx_u8__6_squeezed__1_comb;
  wire [2:0] p3_idx_u8__7_squeezed__1_comb;
  wire [2:0] p3_sel_9068_comb;
  wire [3:0] p3_idx_u8__8_squeezed_comb;
  wire p3_eq_9073_comb;
  wire [7:0] p3_size__1_comb;
  wire [7:0] p3_idx_u8__48_comb;
  wire [7:0] p3_run_size_str_u8_comb;
  wire p3_or_9088_comb;
  wire [7:0] p3_flipped__1_comb;
  wire [4:0] p3_huffman_length_squeezed_comb;
  wire [4:0] p3_idx_u8__2_squeezed__1_comb;
  wire [7:0] p3_code_list__1_comb;
  wire [15:0] p3_huffman_code_full_comb;
  wire [35:0] p3_tuple_9110_comb;
  assign p3_idx_u8__3_squeezed_comb = 2'h3;
  assign p3_idx_u8__4_squeezed__1_comb = 3'h4;
  assign p3_idx_u8__5_squeezed__1_comb = 3'h5;
  assign p3_idx_u8__6_squeezed__1_comb = 3'h6;
  assign p3_idx_u8__7_squeezed__1_comb = 3'h7;
  assign p3_sel_9068_comb = |p2_value__1[7:6] ? p3_idx_u8__7_squeezed__1_comb : (|p2_value__1[7:5] ? p3_idx_u8__6_squeezed__1_comb : (|p2_value__1[7:4] ? p3_idx_u8__5_squeezed__1_comb : (|p2_value__1[7:3] ? p3_idx_u8__4_squeezed__1_comb : {1'h0, p2_or_reduce_9018 ? p3_idx_u8__3_squeezed_comb : p2_sel_9019})));
  assign p3_idx_u8__8_squeezed_comb = 4'h8;
  assign p3_eq_9073_comb = p2_value__1 == 8'h00;
  assign p3_size__1_comb = {4'h0, p2_value__1[7] ? p3_idx_u8__8_squeezed_comb : {1'h0, p3_sel_9068_comb}} & {8{~p3_eq_9073_comb}};
  assign p3_idx_u8__48_comb = 8'h30;
  assign p3_run_size_str_u8_comb = {p2_run_u8__1, 4'h0} | p3_size__1_comb | p3_idx_u8__48_comb;
  assign p3_or_9088_comb = p2_and_8921 | p2_eq_9026;
  assign p3_flipped__1_comb = 8'hff;
  assign p3_huffman_length_squeezed_comb = p2_is_luminance ? literal_9085[p3_run_size_str_u8_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8_comb] : literal_9083[p3_run_size_str_u8_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8_comb];
  assign p3_idx_u8__2_squeezed__1_comb = 5'h02;
  assign p3_code_list__1_comb = p3_eq_9073_comb ? p3_flipped__1_comb : p2_value__1;
  assign p3_huffman_code_full_comb = p2_is_luminance ? literal_9087[p3_run_size_str_u8_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8_comb] : literal_9086[p3_run_size_str_u8_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8_comb];
  assign p3_tuple_9110_comb = {p3_huffman_code_full_comb & {16{~p3_or_9088_comb}}, {3'h0, p3_or_9088_comb ? p3_idx_u8__2_squeezed__1_comb : p3_huffman_length_squeezed_comb}, p2_and_8921 ? p2_value : p3_code_list__1_comb & {8{~p2_eq_9026}}, p2_and_8921 ? 4'hf : p2_and_9029};

  // Registers for pipe stage 3:
  reg [35:0] p3_tuple_9110;
  always @ (posedge clk) begin
    p3_tuple_9110 <= p3_tuple_9110_comb;
  end
  assign out = p3_tuple_9110;
endmodule
