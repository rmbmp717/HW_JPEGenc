module Huffman_ACenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire [7:0] start_pix,
  input wire [7:0] pre_start_pix,
  input wire is_luminance,
  output wire [57:0] out
);
  wire [4:0] literal_11466[0:251];
  assign literal_11466[0] = 5'h02;
  assign literal_11466[1] = 5'h02;
  assign literal_11466[2] = 5'h03;
  assign literal_11466[3] = 5'h04;
  assign literal_11466[4] = 5'h05;
  assign literal_11466[5] = 5'h07;
  assign literal_11466[6] = 5'h08;
  assign literal_11466[7] = 5'h0e;
  assign literal_11466[8] = 5'h10;
  assign literal_11466[9] = 5'h10;
  assign literal_11466[10] = 5'h10;
  assign literal_11466[11] = 5'h00;
  assign literal_11466[12] = 5'h00;
  assign literal_11466[13] = 5'h00;
  assign literal_11466[14] = 5'h00;
  assign literal_11466[15] = 5'h00;
  assign literal_11466[16] = 5'h00;
  assign literal_11466[17] = 5'h03;
  assign literal_11466[18] = 5'h06;
  assign literal_11466[19] = 5'h07;
  assign literal_11466[20] = 5'h09;
  assign literal_11466[21] = 5'h0b;
  assign literal_11466[22] = 5'h0d;
  assign literal_11466[23] = 5'h10;
  assign literal_11466[24] = 5'h10;
  assign literal_11466[25] = 5'h10;
  assign literal_11466[26] = 5'h10;
  assign literal_11466[27] = 5'h00;
  assign literal_11466[28] = 5'h00;
  assign literal_11466[29] = 5'h00;
  assign literal_11466[30] = 5'h00;
  assign literal_11466[31] = 5'h00;
  assign literal_11466[32] = 5'h00;
  assign literal_11466[33] = 5'h05;
  assign literal_11466[34] = 5'h07;
  assign literal_11466[35] = 5'h0a;
  assign literal_11466[36] = 5'h0c;
  assign literal_11466[37] = 5'h0d;
  assign literal_11466[38] = 5'h10;
  assign literal_11466[39] = 5'h10;
  assign literal_11466[40] = 5'h10;
  assign literal_11466[41] = 5'h10;
  assign literal_11466[42] = 5'h10;
  assign literal_11466[43] = 5'h00;
  assign literal_11466[44] = 5'h00;
  assign literal_11466[45] = 5'h00;
  assign literal_11466[46] = 5'h00;
  assign literal_11466[47] = 5'h00;
  assign literal_11466[48] = 5'h00;
  assign literal_11466[49] = 5'h06;
  assign literal_11466[50] = 5'h08;
  assign literal_11466[51] = 5'h0b;
  assign literal_11466[52] = 5'h0c;
  assign literal_11466[53] = 5'h0f;
  assign literal_11466[54] = 5'h10;
  assign literal_11466[55] = 5'h10;
  assign literal_11466[56] = 5'h10;
  assign literal_11466[57] = 5'h10;
  assign literal_11466[58] = 5'h10;
  assign literal_11466[59] = 5'h00;
  assign literal_11466[60] = 5'h00;
  assign literal_11466[61] = 5'h00;
  assign literal_11466[62] = 5'h00;
  assign literal_11466[63] = 5'h00;
  assign literal_11466[64] = 5'h00;
  assign literal_11466[65] = 5'h06;
  assign literal_11466[66] = 5'h0a;
  assign literal_11466[67] = 5'h0c;
  assign literal_11466[68] = 5'h0f;
  assign literal_11466[69] = 5'h10;
  assign literal_11466[70] = 5'h10;
  assign literal_11466[71] = 5'h10;
  assign literal_11466[72] = 5'h10;
  assign literal_11466[73] = 5'h10;
  assign literal_11466[74] = 5'h10;
  assign literal_11466[75] = 5'h00;
  assign literal_11466[76] = 5'h00;
  assign literal_11466[77] = 5'h00;
  assign literal_11466[78] = 5'h00;
  assign literal_11466[79] = 5'h00;
  assign literal_11466[80] = 5'h00;
  assign literal_11466[81] = 5'h07;
  assign literal_11466[82] = 5'h0b;
  assign literal_11466[83] = 5'h0d;
  assign literal_11466[84] = 5'h10;
  assign literal_11466[85] = 5'h10;
  assign literal_11466[86] = 5'h10;
  assign literal_11466[87] = 5'h10;
  assign literal_11466[88] = 5'h10;
  assign literal_11466[89] = 5'h10;
  assign literal_11466[90] = 5'h10;
  assign literal_11466[91] = 5'h00;
  assign literal_11466[92] = 5'h00;
  assign literal_11466[93] = 5'h00;
  assign literal_11466[94] = 5'h00;
  assign literal_11466[95] = 5'h00;
  assign literal_11466[96] = 5'h00;
  assign literal_11466[97] = 5'h07;
  assign literal_11466[98] = 5'h0b;
  assign literal_11466[99] = 5'h0d;
  assign literal_11466[100] = 5'h10;
  assign literal_11466[101] = 5'h10;
  assign literal_11466[102] = 5'h10;
  assign literal_11466[103] = 5'h10;
  assign literal_11466[104] = 5'h10;
  assign literal_11466[105] = 5'h10;
  assign literal_11466[106] = 5'h10;
  assign literal_11466[107] = 5'h00;
  assign literal_11466[108] = 5'h00;
  assign literal_11466[109] = 5'h00;
  assign literal_11466[110] = 5'h00;
  assign literal_11466[111] = 5'h00;
  assign literal_11466[112] = 5'h00;
  assign literal_11466[113] = 5'h08;
  assign literal_11466[114] = 5'h0b;
  assign literal_11466[115] = 5'h0e;
  assign literal_11466[116] = 5'h10;
  assign literal_11466[117] = 5'h10;
  assign literal_11466[118] = 5'h10;
  assign literal_11466[119] = 5'h10;
  assign literal_11466[120] = 5'h10;
  assign literal_11466[121] = 5'h10;
  assign literal_11466[122] = 5'h10;
  assign literal_11466[123] = 5'h00;
  assign literal_11466[124] = 5'h00;
  assign literal_11466[125] = 5'h00;
  assign literal_11466[126] = 5'h00;
  assign literal_11466[127] = 5'h00;
  assign literal_11466[128] = 5'h00;
  assign literal_11466[129] = 5'h08;
  assign literal_11466[130] = 5'h0c;
  assign literal_11466[131] = 5'h10;
  assign literal_11466[132] = 5'h10;
  assign literal_11466[133] = 5'h10;
  assign literal_11466[134] = 5'h10;
  assign literal_11466[135] = 5'h10;
  assign literal_11466[136] = 5'h10;
  assign literal_11466[137] = 5'h10;
  assign literal_11466[138] = 5'h10;
  assign literal_11466[139] = 5'h00;
  assign literal_11466[140] = 5'h00;
  assign literal_11466[141] = 5'h00;
  assign literal_11466[142] = 5'h00;
  assign literal_11466[143] = 5'h00;
  assign literal_11466[144] = 5'h00;
  assign literal_11466[145] = 5'h08;
  assign literal_11466[146] = 5'h0d;
  assign literal_11466[147] = 5'h10;
  assign literal_11466[148] = 5'h10;
  assign literal_11466[149] = 5'h10;
  assign literal_11466[150] = 5'h10;
  assign literal_11466[151] = 5'h10;
  assign literal_11466[152] = 5'h10;
  assign literal_11466[153] = 5'h10;
  assign literal_11466[154] = 5'h10;
  assign literal_11466[155] = 5'h00;
  assign literal_11466[156] = 5'h00;
  assign literal_11466[157] = 5'h00;
  assign literal_11466[158] = 5'h00;
  assign literal_11466[159] = 5'h00;
  assign literal_11466[160] = 5'h00;
  assign literal_11466[161] = 5'h09;
  assign literal_11466[162] = 5'h0d;
  assign literal_11466[163] = 5'h10;
  assign literal_11466[164] = 5'h10;
  assign literal_11466[165] = 5'h10;
  assign literal_11466[166] = 5'h10;
  assign literal_11466[167] = 5'h10;
  assign literal_11466[168] = 5'h10;
  assign literal_11466[169] = 5'h10;
  assign literal_11466[170] = 5'h10;
  assign literal_11466[171] = 5'h00;
  assign literal_11466[172] = 5'h00;
  assign literal_11466[173] = 5'h00;
  assign literal_11466[174] = 5'h00;
  assign literal_11466[175] = 5'h00;
  assign literal_11466[176] = 5'h00;
  assign literal_11466[177] = 5'h09;
  assign literal_11466[178] = 5'h0d;
  assign literal_11466[179] = 5'h10;
  assign literal_11466[180] = 5'h10;
  assign literal_11466[181] = 5'h10;
  assign literal_11466[182] = 5'h10;
  assign literal_11466[183] = 5'h10;
  assign literal_11466[184] = 5'h10;
  assign literal_11466[185] = 5'h10;
  assign literal_11466[186] = 5'h10;
  assign literal_11466[187] = 5'h00;
  assign literal_11466[188] = 5'h00;
  assign literal_11466[189] = 5'h00;
  assign literal_11466[190] = 5'h00;
  assign literal_11466[191] = 5'h00;
  assign literal_11466[192] = 5'h00;
  assign literal_11466[193] = 5'h0a;
  assign literal_11466[194] = 5'h0d;
  assign literal_11466[195] = 5'h10;
  assign literal_11466[196] = 5'h10;
  assign literal_11466[197] = 5'h10;
  assign literal_11466[198] = 5'h10;
  assign literal_11466[199] = 5'h10;
  assign literal_11466[200] = 5'h10;
  assign literal_11466[201] = 5'h10;
  assign literal_11466[202] = 5'h10;
  assign literal_11466[203] = 5'h00;
  assign literal_11466[204] = 5'h00;
  assign literal_11466[205] = 5'h00;
  assign literal_11466[206] = 5'h00;
  assign literal_11466[207] = 5'h00;
  assign literal_11466[208] = 5'h00;
  assign literal_11466[209] = 5'h0a;
  assign literal_11466[210] = 5'h0e;
  assign literal_11466[211] = 5'h10;
  assign literal_11466[212] = 5'h10;
  assign literal_11466[213] = 5'h10;
  assign literal_11466[214] = 5'h10;
  assign literal_11466[215] = 5'h10;
  assign literal_11466[216] = 5'h10;
  assign literal_11466[217] = 5'h10;
  assign literal_11466[218] = 5'h10;
  assign literal_11466[219] = 5'h00;
  assign literal_11466[220] = 5'h00;
  assign literal_11466[221] = 5'h00;
  assign literal_11466[222] = 5'h00;
  assign literal_11466[223] = 5'h00;
  assign literal_11466[224] = 5'h00;
  assign literal_11466[225] = 5'h0a;
  assign literal_11466[226] = 5'h0f;
  assign literal_11466[227] = 5'h10;
  assign literal_11466[228] = 5'h10;
  assign literal_11466[229] = 5'h10;
  assign literal_11466[230] = 5'h10;
  assign literal_11466[231] = 5'h10;
  assign literal_11466[232] = 5'h10;
  assign literal_11466[233] = 5'h10;
  assign literal_11466[234] = 5'h10;
  assign literal_11466[235] = 5'h00;
  assign literal_11466[236] = 5'h00;
  assign literal_11466[237] = 5'h00;
  assign literal_11466[238] = 5'h00;
  assign literal_11466[239] = 5'h00;
  assign literal_11466[240] = 5'h09;
  assign literal_11466[241] = 5'h0b;
  assign literal_11466[242] = 5'h10;
  assign literal_11466[243] = 5'h10;
  assign literal_11466[244] = 5'h10;
  assign literal_11466[245] = 5'h10;
  assign literal_11466[246] = 5'h10;
  assign literal_11466[247] = 5'h10;
  assign literal_11466[248] = 5'h10;
  assign literal_11466[249] = 5'h10;
  assign literal_11466[250] = 5'h10;
  assign literal_11466[251] = 5'h00;
  wire [4:0] literal_11468[0:251];
  assign literal_11468[0] = 5'h04;
  assign literal_11468[1] = 5'h02;
  assign literal_11468[2] = 5'h02;
  assign literal_11468[3] = 5'h03;
  assign literal_11468[4] = 5'h04;
  assign literal_11468[5] = 5'h05;
  assign literal_11468[6] = 5'h07;
  assign literal_11468[7] = 5'h09;
  assign literal_11468[8] = 5'h10;
  assign literal_11468[9] = 5'h10;
  assign literal_11468[10] = 5'h10;
  assign literal_11468[11] = 5'h00;
  assign literal_11468[12] = 5'h00;
  assign literal_11468[13] = 5'h00;
  assign literal_11468[14] = 5'h00;
  assign literal_11468[15] = 5'h00;
  assign literal_11468[16] = 5'h00;
  assign literal_11468[17] = 5'h04;
  assign literal_11468[18] = 5'h05;
  assign literal_11468[19] = 5'h07;
  assign literal_11468[20] = 5'h09;
  assign literal_11468[21] = 5'h0a;
  assign literal_11468[22] = 5'h0b;
  assign literal_11468[23] = 5'h10;
  assign literal_11468[24] = 5'h10;
  assign literal_11468[25] = 5'h10;
  assign literal_11468[26] = 5'h10;
  assign literal_11468[27] = 5'h00;
  assign literal_11468[28] = 5'h00;
  assign literal_11468[29] = 5'h00;
  assign literal_11468[30] = 5'h00;
  assign literal_11468[31] = 5'h00;
  assign literal_11468[32] = 5'h00;
  assign literal_11468[33] = 5'h05;
  assign literal_11468[34] = 5'h08;
  assign literal_11468[35] = 5'h0a;
  assign literal_11468[36] = 5'h0c;
  assign literal_11468[37] = 5'h0e;
  assign literal_11468[38] = 5'h10;
  assign literal_11468[39] = 5'h10;
  assign literal_11468[40] = 5'h10;
  assign literal_11468[41] = 5'h10;
  assign literal_11468[42] = 5'h10;
  assign literal_11468[43] = 5'h00;
  assign literal_11468[44] = 5'h00;
  assign literal_11468[45] = 5'h00;
  assign literal_11468[46] = 5'h00;
  assign literal_11468[47] = 5'h00;
  assign literal_11468[48] = 5'h00;
  assign literal_11468[49] = 5'h06;
  assign literal_11468[50] = 5'h09;
  assign literal_11468[51] = 5'h0b;
  assign literal_11468[52] = 5'h0e;
  assign literal_11468[53] = 5'h10;
  assign literal_11468[54] = 5'h10;
  assign literal_11468[55] = 5'h10;
  assign literal_11468[56] = 5'h10;
  assign literal_11468[57] = 5'h10;
  assign literal_11468[58] = 5'h10;
  assign literal_11468[59] = 5'h00;
  assign literal_11468[60] = 5'h00;
  assign literal_11468[61] = 5'h00;
  assign literal_11468[62] = 5'h00;
  assign literal_11468[63] = 5'h00;
  assign literal_11468[64] = 5'h00;
  assign literal_11468[65] = 5'h06;
  assign literal_11468[66] = 5'h0a;
  assign literal_11468[67] = 5'h0e;
  assign literal_11468[68] = 5'h10;
  assign literal_11468[69] = 5'h10;
  assign literal_11468[70] = 5'h10;
  assign literal_11468[71] = 5'h10;
  assign literal_11468[72] = 5'h10;
  assign literal_11468[73] = 5'h10;
  assign literal_11468[74] = 5'h10;
  assign literal_11468[75] = 5'h00;
  assign literal_11468[76] = 5'h00;
  assign literal_11468[77] = 5'h00;
  assign literal_11468[78] = 5'h00;
  assign literal_11468[79] = 5'h00;
  assign literal_11468[80] = 5'h00;
  assign literal_11468[81] = 5'h07;
  assign literal_11468[82] = 5'h0a;
  assign literal_11468[83] = 5'h0e;
  assign literal_11468[84] = 5'h10;
  assign literal_11468[85] = 5'h10;
  assign literal_11468[86] = 5'h10;
  assign literal_11468[87] = 5'h10;
  assign literal_11468[88] = 5'h10;
  assign literal_11468[89] = 5'h10;
  assign literal_11468[90] = 5'h10;
  assign literal_11468[91] = 5'h00;
  assign literal_11468[92] = 5'h00;
  assign literal_11468[93] = 5'h00;
  assign literal_11468[94] = 5'h00;
  assign literal_11468[95] = 5'h00;
  assign literal_11468[96] = 5'h00;
  assign literal_11468[97] = 5'h07;
  assign literal_11468[98] = 5'h0c;
  assign literal_11468[99] = 5'h0f;
  assign literal_11468[100] = 5'h10;
  assign literal_11468[101] = 5'h10;
  assign literal_11468[102] = 5'h10;
  assign literal_11468[103] = 5'h10;
  assign literal_11468[104] = 5'h10;
  assign literal_11468[105] = 5'h10;
  assign literal_11468[106] = 5'h10;
  assign literal_11468[107] = 5'h00;
  assign literal_11468[108] = 5'h00;
  assign literal_11468[109] = 5'h00;
  assign literal_11468[110] = 5'h00;
  assign literal_11468[111] = 5'h00;
  assign literal_11468[112] = 5'h00;
  assign literal_11468[113] = 5'h08;
  assign literal_11468[114] = 5'h0c;
  assign literal_11468[115] = 5'h10;
  assign literal_11468[116] = 5'h10;
  assign literal_11468[117] = 5'h10;
  assign literal_11468[118] = 5'h10;
  assign literal_11468[119] = 5'h10;
  assign literal_11468[120] = 5'h10;
  assign literal_11468[121] = 5'h10;
  assign literal_11468[122] = 5'h10;
  assign literal_11468[123] = 5'h00;
  assign literal_11468[124] = 5'h00;
  assign literal_11468[125] = 5'h00;
  assign literal_11468[126] = 5'h00;
  assign literal_11468[127] = 5'h00;
  assign literal_11468[128] = 5'h00;
  assign literal_11468[129] = 5'h09;
  assign literal_11468[130] = 5'h0d;
  assign literal_11468[131] = 5'h10;
  assign literal_11468[132] = 5'h10;
  assign literal_11468[133] = 5'h10;
  assign literal_11468[134] = 5'h10;
  assign literal_11468[135] = 5'h10;
  assign literal_11468[136] = 5'h10;
  assign literal_11468[137] = 5'h10;
  assign literal_11468[138] = 5'h10;
  assign literal_11468[139] = 5'h00;
  assign literal_11468[140] = 5'h00;
  assign literal_11468[141] = 5'h00;
  assign literal_11468[142] = 5'h00;
  assign literal_11468[143] = 5'h00;
  assign literal_11468[144] = 5'h00;
  assign literal_11468[145] = 5'h09;
  assign literal_11468[146] = 5'h0e;
  assign literal_11468[147] = 5'h10;
  assign literal_11468[148] = 5'h10;
  assign literal_11468[149] = 5'h10;
  assign literal_11468[150] = 5'h10;
  assign literal_11468[151] = 5'h10;
  assign literal_11468[152] = 5'h10;
  assign literal_11468[153] = 5'h10;
  assign literal_11468[154] = 5'h10;
  assign literal_11468[155] = 5'h00;
  assign literal_11468[156] = 5'h00;
  assign literal_11468[157] = 5'h00;
  assign literal_11468[158] = 5'h00;
  assign literal_11468[159] = 5'h00;
  assign literal_11468[160] = 5'h00;
  assign literal_11468[161] = 5'h09;
  assign literal_11468[162] = 5'h0e;
  assign literal_11468[163] = 5'h10;
  assign literal_11468[164] = 5'h10;
  assign literal_11468[165] = 5'h10;
  assign literal_11468[166] = 5'h10;
  assign literal_11468[167] = 5'h10;
  assign literal_11468[168] = 5'h10;
  assign literal_11468[169] = 5'h10;
  assign literal_11468[170] = 5'h10;
  assign literal_11468[171] = 5'h00;
  assign literal_11468[172] = 5'h00;
  assign literal_11468[173] = 5'h00;
  assign literal_11468[174] = 5'h00;
  assign literal_11468[175] = 5'h00;
  assign literal_11468[176] = 5'h00;
  assign literal_11468[177] = 5'h0a;
  assign literal_11468[178] = 5'h0f;
  assign literal_11468[179] = 5'h10;
  assign literal_11468[180] = 5'h10;
  assign literal_11468[181] = 5'h10;
  assign literal_11468[182] = 5'h10;
  assign literal_11468[183] = 5'h10;
  assign literal_11468[184] = 5'h10;
  assign literal_11468[185] = 5'h10;
  assign literal_11468[186] = 5'h10;
  assign literal_11468[187] = 5'h00;
  assign literal_11468[188] = 5'h00;
  assign literal_11468[189] = 5'h00;
  assign literal_11468[190] = 5'h00;
  assign literal_11468[191] = 5'h00;
  assign literal_11468[192] = 5'h00;
  assign literal_11468[193] = 5'h0a;
  assign literal_11468[194] = 5'h10;
  assign literal_11468[195] = 5'h10;
  assign literal_11468[196] = 5'h10;
  assign literal_11468[197] = 5'h10;
  assign literal_11468[198] = 5'h10;
  assign literal_11468[199] = 5'h10;
  assign literal_11468[200] = 5'h10;
  assign literal_11468[201] = 5'h10;
  assign literal_11468[202] = 5'h10;
  assign literal_11468[203] = 5'h00;
  assign literal_11468[204] = 5'h00;
  assign literal_11468[205] = 5'h00;
  assign literal_11468[206] = 5'h00;
  assign literal_11468[207] = 5'h00;
  assign literal_11468[208] = 5'h00;
  assign literal_11468[209] = 5'h0a;
  assign literal_11468[210] = 5'h10;
  assign literal_11468[211] = 5'h10;
  assign literal_11468[212] = 5'h10;
  assign literal_11468[213] = 5'h10;
  assign literal_11468[214] = 5'h10;
  assign literal_11468[215] = 5'h10;
  assign literal_11468[216] = 5'h10;
  assign literal_11468[217] = 5'h10;
  assign literal_11468[218] = 5'h10;
  assign literal_11468[219] = 5'h00;
  assign literal_11468[220] = 5'h00;
  assign literal_11468[221] = 5'h00;
  assign literal_11468[222] = 5'h00;
  assign literal_11468[223] = 5'h00;
  assign literal_11468[224] = 5'h00;
  assign literal_11468[225] = 5'h0b;
  assign literal_11468[226] = 5'h10;
  assign literal_11468[227] = 5'h10;
  assign literal_11468[228] = 5'h10;
  assign literal_11468[229] = 5'h10;
  assign literal_11468[230] = 5'h10;
  assign literal_11468[231] = 5'h10;
  assign literal_11468[232] = 5'h10;
  assign literal_11468[233] = 5'h10;
  assign literal_11468[234] = 5'h10;
  assign literal_11468[235] = 5'h00;
  assign literal_11468[236] = 5'h00;
  assign literal_11468[237] = 5'h00;
  assign literal_11468[238] = 5'h00;
  assign literal_11468[239] = 5'h00;
  assign literal_11468[240] = 5'h0c;
  assign literal_11468[241] = 5'h0d;
  assign literal_11468[242] = 5'h10;
  assign literal_11468[243] = 5'h10;
  assign literal_11468[244] = 5'h10;
  assign literal_11468[245] = 5'h10;
  assign literal_11468[246] = 5'h10;
  assign literal_11468[247] = 5'h10;
  assign literal_11468[248] = 5'h10;
  assign literal_11468[249] = 5'h10;
  assign literal_11468[250] = 5'h10;
  assign literal_11468[251] = 5'h00;
  wire [15:0] literal_11472[0:251];
  assign literal_11472[0] = 16'h0001;
  assign literal_11472[1] = 16'h0000;
  assign literal_11472[2] = 16'h0004;
  assign literal_11472[3] = 16'h000c;
  assign literal_11472[4] = 16'h001a;
  assign literal_11472[5] = 16'h0076;
  assign literal_11472[6] = 16'h00f6;
  assign literal_11472[7] = 16'h3fe0;
  assign literal_11472[8] = 16'hff96;
  assign literal_11472[9] = 16'hff97;
  assign literal_11472[10] = 16'hff98;
  assign literal_11472[11] = 16'h0000;
  assign literal_11472[12] = 16'h0000;
  assign literal_11472[13] = 16'h0000;
  assign literal_11472[14] = 16'h0000;
  assign literal_11472[15] = 16'h0000;
  assign literal_11472[16] = 16'h0000;
  assign literal_11472[17] = 16'h0005;
  assign literal_11472[18] = 16'h0038;
  assign literal_11472[19] = 16'h0078;
  assign literal_11472[20] = 16'h01f9;
  assign literal_11472[21] = 16'h07f2;
  assign literal_11472[22] = 16'h1fe8;
  assign literal_11472[23] = 16'hff93;
  assign literal_11472[24] = 16'hff99;
  assign literal_11472[25] = 16'hff9a;
  assign literal_11472[26] = 16'hff9e;
  assign literal_11472[27] = 16'h0000;
  assign literal_11472[28] = 16'h0000;
  assign literal_11472[29] = 16'h0000;
  assign literal_11472[30] = 16'h0000;
  assign literal_11472[31] = 16'h0000;
  assign literal_11472[32] = 16'h0000;
  assign literal_11472[33] = 16'h001b;
  assign literal_11472[34] = 16'h007a;
  assign literal_11472[35] = 16'h03f7;
  assign literal_11472[36] = 16'h0ff0;
  assign literal_11472[37] = 16'h1feb;
  assign literal_11472[38] = 16'hff9b;
  assign literal_11472[39] = 16'hff9f;
  assign literal_11472[40] = 16'hffa8;
  assign literal_11472[41] = 16'hffa9;
  assign literal_11472[42] = 16'hfff1;
  assign literal_11472[43] = 16'h0000;
  assign literal_11472[44] = 16'h0000;
  assign literal_11472[45] = 16'h0000;
  assign literal_11472[46] = 16'h0000;
  assign literal_11472[47] = 16'h0000;
  assign literal_11472[48] = 16'h0000;
  assign literal_11472[49] = 16'h0039;
  assign literal_11472[50] = 16'h00fa;
  assign literal_11472[51] = 16'h07f7;
  assign literal_11472[52] = 16'h0ff1;
  assign literal_11472[53] = 16'h7fc6;
  assign literal_11472[54] = 16'hff9c;
  assign literal_11472[55] = 16'hffa3;
  assign literal_11472[56] = 16'hffd7;
  assign literal_11472[57] = 16'hffe4;
  assign literal_11472[58] = 16'hfff2;
  assign literal_11472[59] = 16'h0000;
  assign literal_11472[60] = 16'h0000;
  assign literal_11472[61] = 16'h0000;
  assign literal_11472[62] = 16'h0000;
  assign literal_11472[63] = 16'h0000;
  assign literal_11472[64] = 16'h0000;
  assign literal_11472[65] = 16'h003a;
  assign literal_11472[66] = 16'h03f8;
  assign literal_11472[67] = 16'h0ff2;
  assign literal_11472[68] = 16'h7fc8;
  assign literal_11472[69] = 16'hff9d;
  assign literal_11472[70] = 16'hffbf;
  assign literal_11472[71] = 16'hffcb;
  assign literal_11472[72] = 16'hffd8;
  assign literal_11472[73] = 16'hffe5;
  assign literal_11472[74] = 16'hfff3;
  assign literal_11472[75] = 16'h0000;
  assign literal_11472[76] = 16'h0000;
  assign literal_11472[77] = 16'h0000;
  assign literal_11472[78] = 16'h0000;
  assign literal_11472[79] = 16'h0000;
  assign literal_11472[80] = 16'h0000;
  assign literal_11472[81] = 16'h0077;
  assign literal_11472[82] = 16'h07f3;
  assign literal_11472[83] = 16'h1fea;
  assign literal_11472[84] = 16'hff94;
  assign literal_11472[85] = 16'hffa2;
  assign literal_11472[86] = 16'hffc0;
  assign literal_11472[87] = 16'hffcc;
  assign literal_11472[88] = 16'hffd9;
  assign literal_11472[89] = 16'hffe6;
  assign literal_11472[90] = 16'hfff4;
  assign literal_11472[91] = 16'h0000;
  assign literal_11472[92] = 16'h0000;
  assign literal_11472[93] = 16'h0000;
  assign literal_11472[94] = 16'h0000;
  assign literal_11472[95] = 16'h0000;
  assign literal_11472[96] = 16'h0000;
  assign literal_11472[97] = 16'h0079;
  assign literal_11472[98] = 16'h07f4;
  assign literal_11472[99] = 16'h1fed;
  assign literal_11472[100] = 16'hffa0;
  assign literal_11472[101] = 16'hffb5;
  assign literal_11472[102] = 16'hffc1;
  assign literal_11472[103] = 16'hffcd;
  assign literal_11472[104] = 16'hffda;
  assign literal_11472[105] = 16'hffe7;
  assign literal_11472[106] = 16'hfff5;
  assign literal_11472[107] = 16'h0000;
  assign literal_11472[108] = 16'h0000;
  assign literal_11472[109] = 16'h0000;
  assign literal_11472[110] = 16'h0000;
  assign literal_11472[111] = 16'h0000;
  assign literal_11472[112] = 16'h0000;
  assign literal_11472[113] = 16'h00f7;
  assign literal_11472[114] = 16'h07f5;
  assign literal_11472[115] = 16'h3fe1;
  assign literal_11472[116] = 16'hffa1;
  assign literal_11472[117] = 16'hffb6;
  assign literal_11472[118] = 16'hffc2;
  assign literal_11472[119] = 16'hffce;
  assign literal_11472[120] = 16'hffdb;
  assign literal_11472[121] = 16'hffe8;
  assign literal_11472[122] = 16'hfff6;
  assign literal_11472[123] = 16'h0000;
  assign literal_11472[124] = 16'h0000;
  assign literal_11472[125] = 16'h0000;
  assign literal_11472[126] = 16'h0000;
  assign literal_11472[127] = 16'h0000;
  assign literal_11472[128] = 16'h0000;
  assign literal_11472[129] = 16'h00f8;
  assign literal_11472[130] = 16'h0ff3;
  assign literal_11472[131] = 16'hff92;
  assign literal_11472[132] = 16'hffad;
  assign literal_11472[133] = 16'hffb7;
  assign literal_11472[134] = 16'hffc3;
  assign literal_11472[135] = 16'hffcf;
  assign literal_11472[136] = 16'hffdc;
  assign literal_11472[137] = 16'hffe9;
  assign literal_11472[138] = 16'hfff7;
  assign literal_11472[139] = 16'h0000;
  assign literal_11472[140] = 16'h0000;
  assign literal_11472[141] = 16'h0000;
  assign literal_11472[142] = 16'h0000;
  assign literal_11472[143] = 16'h0000;
  assign literal_11472[144] = 16'h0000;
  assign literal_11472[145] = 16'h00f9;
  assign literal_11472[146] = 16'h1fe9;
  assign literal_11472[147] = 16'hff95;
  assign literal_11472[148] = 16'hffae;
  assign literal_11472[149] = 16'hffb8;
  assign literal_11472[150] = 16'hffc4;
  assign literal_11472[151] = 16'hffd0;
  assign literal_11472[152] = 16'hffdd;
  assign literal_11472[153] = 16'hffea;
  assign literal_11472[154] = 16'hfff8;
  assign literal_11472[155] = 16'h0000;
  assign literal_11472[156] = 16'h0000;
  assign literal_11472[157] = 16'h0000;
  assign literal_11472[158] = 16'h0000;
  assign literal_11472[159] = 16'h0000;
  assign literal_11472[160] = 16'h0000;
  assign literal_11472[161] = 16'h01f6;
  assign literal_11472[162] = 16'h1fec;
  assign literal_11472[163] = 16'hffa5;
  assign literal_11472[164] = 16'hffaf;
  assign literal_11472[165] = 16'hffb9;
  assign literal_11472[166] = 16'hffc5;
  assign literal_11472[167] = 16'hffd1;
  assign literal_11472[168] = 16'hffde;
  assign literal_11472[169] = 16'hffeb;
  assign literal_11472[170] = 16'hfff9;
  assign literal_11472[171] = 16'h0000;
  assign literal_11472[172] = 16'h0000;
  assign literal_11472[173] = 16'h0000;
  assign literal_11472[174] = 16'h0000;
  assign literal_11472[175] = 16'h0000;
  assign literal_11472[176] = 16'h0000;
  assign literal_11472[177] = 16'h01f7;
  assign literal_11472[178] = 16'h1fee;
  assign literal_11472[179] = 16'hffa6;
  assign literal_11472[180] = 16'hffb0;
  assign literal_11472[181] = 16'hffba;
  assign literal_11472[182] = 16'hffc6;
  assign literal_11472[183] = 16'hffd2;
  assign literal_11472[184] = 16'hffdf;
  assign literal_11472[185] = 16'hffec;
  assign literal_11472[186] = 16'hfffa;
  assign literal_11472[187] = 16'h0000;
  assign literal_11472[188] = 16'h0000;
  assign literal_11472[189] = 16'h0000;
  assign literal_11472[190] = 16'h0000;
  assign literal_11472[191] = 16'h0000;
  assign literal_11472[192] = 16'h0000;
  assign literal_11472[193] = 16'h03f4;
  assign literal_11472[194] = 16'h1fef;
  assign literal_11472[195] = 16'hffa7;
  assign literal_11472[196] = 16'hffb1;
  assign literal_11472[197] = 16'hffbb;
  assign literal_11472[198] = 16'hffc7;
  assign literal_11472[199] = 16'hffd3;
  assign literal_11472[200] = 16'hffe0;
  assign literal_11472[201] = 16'hffed;
  assign literal_11472[202] = 16'hfffb;
  assign literal_11472[203] = 16'h0000;
  assign literal_11472[204] = 16'h0000;
  assign literal_11472[205] = 16'h0000;
  assign literal_11472[206] = 16'h0000;
  assign literal_11472[207] = 16'h0000;
  assign literal_11472[208] = 16'h0000;
  assign literal_11472[209] = 16'h03f5;
  assign literal_11472[210] = 16'h3fe2;
  assign literal_11472[211] = 16'hffaa;
  assign literal_11472[212] = 16'hffb2;
  assign literal_11472[213] = 16'hffbc;
  assign literal_11472[214] = 16'hffc8;
  assign literal_11472[215] = 16'hffd4;
  assign literal_11472[216] = 16'hffe1;
  assign literal_11472[217] = 16'hffee;
  assign literal_11472[218] = 16'hfffc;
  assign literal_11472[219] = 16'h0000;
  assign literal_11472[220] = 16'h0000;
  assign literal_11472[221] = 16'h0000;
  assign literal_11472[222] = 16'h0000;
  assign literal_11472[223] = 16'h0000;
  assign literal_11472[224] = 16'h0000;
  assign literal_11472[225] = 16'h03f6;
  assign literal_11472[226] = 16'h7fc7;
  assign literal_11472[227] = 16'hffab;
  assign literal_11472[228] = 16'hffb3;
  assign literal_11472[229] = 16'hffbd;
  assign literal_11472[230] = 16'hffc9;
  assign literal_11472[231] = 16'hffd5;
  assign literal_11472[232] = 16'hffe2;
  assign literal_11472[233] = 16'hffef;
  assign literal_11472[234] = 16'hfffd;
  assign literal_11472[235] = 16'h0000;
  assign literal_11472[236] = 16'h0000;
  assign literal_11472[237] = 16'h0000;
  assign literal_11472[238] = 16'h0000;
  assign literal_11472[239] = 16'h0000;
  assign literal_11472[240] = 16'h01f8;
  assign literal_11472[241] = 16'h07f6;
  assign literal_11472[242] = 16'hffa4;
  assign literal_11472[243] = 16'hffac;
  assign literal_11472[244] = 16'hffb4;
  assign literal_11472[245] = 16'hffbe;
  assign literal_11472[246] = 16'hffca;
  assign literal_11472[247] = 16'hffd6;
  assign literal_11472[248] = 16'hffe3;
  assign literal_11472[249] = 16'hfff0;
  assign literal_11472[250] = 16'hfffe;
  assign literal_11472[251] = 16'h0000;
  wire [15:0] literal_11473[0:251];
  assign literal_11473[0] = 16'h000c;
  assign literal_11473[1] = 16'h0000;
  assign literal_11473[2] = 16'h0001;
  assign literal_11473[3] = 16'h0004;
  assign literal_11473[4] = 16'h000b;
  assign literal_11473[5] = 16'h001a;
  assign literal_11473[6] = 16'h0079;
  assign literal_11473[7] = 16'h01f9;
  assign literal_11473[8] = 16'hff9c;
  assign literal_11473[9] = 16'hff9f;
  assign literal_11473[10] = 16'hffa0;
  assign literal_11473[11] = 16'h0000;
  assign literal_11473[12] = 16'h0000;
  assign literal_11473[13] = 16'h0000;
  assign literal_11473[14] = 16'h0000;
  assign literal_11473[15] = 16'h0000;
  assign literal_11473[16] = 16'h0000;
  assign literal_11473[17] = 16'h000a;
  assign literal_11473[18] = 16'h001c;
  assign literal_11473[19] = 16'h007a;
  assign literal_11473[20] = 16'h01f5;
  assign literal_11473[21] = 16'h03f4;
  assign literal_11473[22] = 16'h07f8;
  assign literal_11473[23] = 16'hff95;
  assign literal_11473[24] = 16'hffa1;
  assign literal_11473[25] = 16'hffa2;
  assign literal_11473[26] = 16'hffad;
  assign literal_11473[27] = 16'h0000;
  assign literal_11473[28] = 16'h0000;
  assign literal_11473[29] = 16'h0000;
  assign literal_11473[30] = 16'h0000;
  assign literal_11473[31] = 16'h0000;
  assign literal_11473[32] = 16'h0000;
  assign literal_11473[33] = 16'h001b;
  assign literal_11473[34] = 16'h00f8;
  assign literal_11473[35] = 16'h03f7;
  assign literal_11473[36] = 16'h0ff4;
  assign literal_11473[37] = 16'h3fdc;
  assign literal_11473[38] = 16'hff9d;
  assign literal_11473[39] = 16'hff90;
  assign literal_11473[40] = 16'hffac;
  assign literal_11473[41] = 16'hffe3;
  assign literal_11473[42] = 16'hfff1;
  assign literal_11473[43] = 16'h0000;
  assign literal_11473[44] = 16'h0000;
  assign literal_11473[45] = 16'h0000;
  assign literal_11473[46] = 16'h0000;
  assign literal_11473[47] = 16'h0000;
  assign literal_11473[48] = 16'h0000;
  assign literal_11473[49] = 16'h003a;
  assign literal_11473[50] = 16'h01f6;
  assign literal_11473[51] = 16'h07f7;
  assign literal_11473[52] = 16'h3fde;
  assign literal_11473[53] = 16'hff8e;
  assign literal_11473[54] = 16'hff94;
  assign literal_11473[55] = 16'hffc9;
  assign literal_11473[56] = 16'hffd6;
  assign literal_11473[57] = 16'hffe4;
  assign literal_11473[58] = 16'hfff2;
  assign literal_11473[59] = 16'h0000;
  assign literal_11473[60] = 16'h0000;
  assign literal_11473[61] = 16'h0000;
  assign literal_11473[62] = 16'h0000;
  assign literal_11473[63] = 16'h0000;
  assign literal_11473[64] = 16'h0000;
  assign literal_11473[65] = 16'h003b;
  assign literal_11473[66] = 16'h03f6;
  assign literal_11473[67] = 16'h3fdd;
  assign literal_11473[68] = 16'hff8f;
  assign literal_11473[69] = 16'hffa5;
  assign literal_11473[70] = 16'hffa6;
  assign literal_11473[71] = 16'hffca;
  assign literal_11473[72] = 16'hffd7;
  assign literal_11473[73] = 16'hffe5;
  assign literal_11473[74] = 16'hfff3;
  assign literal_11473[75] = 16'h0000;
  assign literal_11473[76] = 16'h0000;
  assign literal_11473[77] = 16'h0000;
  assign literal_11473[78] = 16'h0000;
  assign literal_11473[79] = 16'h0000;
  assign literal_11473[80] = 16'h0000;
  assign literal_11473[81] = 16'h0078;
  assign literal_11473[82] = 16'h03f9;
  assign literal_11473[83] = 16'h3fdf;
  assign literal_11473[84] = 16'hff96;
  assign literal_11473[85] = 16'hffab;
  assign literal_11473[86] = 16'hffa9;
  assign literal_11473[87] = 16'hffcb;
  assign literal_11473[88] = 16'hffd8;
  assign literal_11473[89] = 16'hffe6;
  assign literal_11473[90] = 16'hfff4;
  assign literal_11473[91] = 16'h0000;
  assign literal_11473[92] = 16'h0000;
  assign literal_11473[93] = 16'h0000;
  assign literal_11473[94] = 16'h0000;
  assign literal_11473[95] = 16'h0000;
  assign literal_11473[96] = 16'h0000;
  assign literal_11473[97] = 16'h007b;
  assign literal_11473[98] = 16'h0ff2;
  assign literal_11473[99] = 16'h7fc5;
  assign literal_11473[100] = 16'hff97;
  assign literal_11473[101] = 16'hffb5;
  assign literal_11473[102] = 16'hffbf;
  assign literal_11473[103] = 16'hffcc;
  assign literal_11473[104] = 16'hffd9;
  assign literal_11473[105] = 16'hffe7;
  assign literal_11473[106] = 16'hfff5;
  assign literal_11473[107] = 16'h0000;
  assign literal_11473[108] = 16'h0000;
  assign literal_11473[109] = 16'h0000;
  assign literal_11473[110] = 16'h0000;
  assign literal_11473[111] = 16'h0000;
  assign literal_11473[112] = 16'h0000;
  assign literal_11473[113] = 16'h00f9;
  assign literal_11473[114] = 16'h0ff5;
  assign literal_11473[115] = 16'hff8c;
  assign literal_11473[116] = 16'hff98;
  assign literal_11473[117] = 16'hffb6;
  assign literal_11473[118] = 16'hffc0;
  assign literal_11473[119] = 16'hffcd;
  assign literal_11473[120] = 16'hffda;
  assign literal_11473[121] = 16'hffe8;
  assign literal_11473[122] = 16'hfff6;
  assign literal_11473[123] = 16'h0000;
  assign literal_11473[124] = 16'h0000;
  assign literal_11473[125] = 16'h0000;
  assign literal_11473[126] = 16'h0000;
  assign literal_11473[127] = 16'h0000;
  assign literal_11473[128] = 16'h0000;
  assign literal_11473[129] = 16'h01f4;
  assign literal_11473[130] = 16'h1fec;
  assign literal_11473[131] = 16'hff9e;
  assign literal_11473[132] = 16'hffa3;
  assign literal_11473[133] = 16'hffb7;
  assign literal_11473[134] = 16'hffc1;
  assign literal_11473[135] = 16'hffce;
  assign literal_11473[136] = 16'hffdb;
  assign literal_11473[137] = 16'hffe9;
  assign literal_11473[138] = 16'hfff7;
  assign literal_11473[139] = 16'h0000;
  assign literal_11473[140] = 16'h0000;
  assign literal_11473[141] = 16'h0000;
  assign literal_11473[142] = 16'h0000;
  assign literal_11473[143] = 16'h0000;
  assign literal_11473[144] = 16'h0000;
  assign literal_11473[145] = 16'h01f7;
  assign literal_11473[146] = 16'h3fe0;
  assign literal_11473[147] = 16'hff91;
  assign literal_11473[148] = 16'hffa4;
  assign literal_11473[149] = 16'hffb8;
  assign literal_11473[150] = 16'hffc2;
  assign literal_11473[151] = 16'hffcf;
  assign literal_11473[152] = 16'hffdc;
  assign literal_11473[153] = 16'hffea;
  assign literal_11473[154] = 16'hfff8;
  assign literal_11473[155] = 16'h0000;
  assign literal_11473[156] = 16'h0000;
  assign literal_11473[157] = 16'h0000;
  assign literal_11473[158] = 16'h0000;
  assign literal_11473[159] = 16'h0000;
  assign literal_11473[160] = 16'h0000;
  assign literal_11473[161] = 16'h01f8;
  assign literal_11473[162] = 16'h3fe1;
  assign literal_11473[163] = 16'hff92;
  assign literal_11473[164] = 16'hffa7;
  assign literal_11473[165] = 16'hffb9;
  assign literal_11473[166] = 16'hffc3;
  assign literal_11473[167] = 16'hffd0;
  assign literal_11473[168] = 16'hffdd;
  assign literal_11473[169] = 16'hffeb;
  assign literal_11473[170] = 16'hfff9;
  assign literal_11473[171] = 16'h0000;
  assign literal_11473[172] = 16'h0000;
  assign literal_11473[173] = 16'h0000;
  assign literal_11473[174] = 16'h0000;
  assign literal_11473[175] = 16'h0000;
  assign literal_11473[176] = 16'h0000;
  assign literal_11473[177] = 16'h03f5;
  assign literal_11473[178] = 16'h7fc4;
  assign literal_11473[179] = 16'hff93;
  assign literal_11473[180] = 16'hffa8;
  assign literal_11473[181] = 16'hffba;
  assign literal_11473[182] = 16'hffc4;
  assign literal_11473[183] = 16'hffd1;
  assign literal_11473[184] = 16'hffde;
  assign literal_11473[185] = 16'hffec;
  assign literal_11473[186] = 16'hfffa;
  assign literal_11473[187] = 16'h0000;
  assign literal_11473[188] = 16'h0000;
  assign literal_11473[189] = 16'h0000;
  assign literal_11473[190] = 16'h0000;
  assign literal_11473[191] = 16'h0000;
  assign literal_11473[192] = 16'h0000;
  assign literal_11473[193] = 16'h03f8;
  assign literal_11473[194] = 16'hff8d;
  assign literal_11473[195] = 16'hff99;
  assign literal_11473[196] = 16'hffb1;
  assign literal_11473[197] = 16'hffbb;
  assign literal_11473[198] = 16'hffc5;
  assign literal_11473[199] = 16'hffd2;
  assign literal_11473[200] = 16'hffdf;
  assign literal_11473[201] = 16'hffed;
  assign literal_11473[202] = 16'hfffb;
  assign literal_11473[203] = 16'h0000;
  assign literal_11473[204] = 16'h0000;
  assign literal_11473[205] = 16'h0000;
  assign literal_11473[206] = 16'h0000;
  assign literal_11473[207] = 16'h0000;
  assign literal_11473[208] = 16'h0000;
  assign literal_11473[209] = 16'h03fa;
  assign literal_11473[210] = 16'hff9a;
  assign literal_11473[211] = 16'hffaa;
  assign literal_11473[212] = 16'hffb2;
  assign literal_11473[213] = 16'hffbc;
  assign literal_11473[214] = 16'hffc6;
  assign literal_11473[215] = 16'hffd3;
  assign literal_11473[216] = 16'hffe0;
  assign literal_11473[217] = 16'hffee;
  assign literal_11473[218] = 16'hfffc;
  assign literal_11473[219] = 16'h0000;
  assign literal_11473[220] = 16'h0000;
  assign literal_11473[221] = 16'h0000;
  assign literal_11473[222] = 16'h0000;
  assign literal_11473[223] = 16'h0000;
  assign literal_11473[224] = 16'h0000;
  assign literal_11473[225] = 16'h07f6;
  assign literal_11473[226] = 16'hff9b;
  assign literal_11473[227] = 16'hffaf;
  assign literal_11473[228] = 16'hffb3;
  assign literal_11473[229] = 16'hffbd;
  assign literal_11473[230] = 16'hffc7;
  assign literal_11473[231] = 16'hffd4;
  assign literal_11473[232] = 16'hffe1;
  assign literal_11473[233] = 16'hffef;
  assign literal_11473[234] = 16'hfffd;
  assign literal_11473[235] = 16'h0000;
  assign literal_11473[236] = 16'h0000;
  assign literal_11473[237] = 16'h0000;
  assign literal_11473[238] = 16'h0000;
  assign literal_11473[239] = 16'h0000;
  assign literal_11473[240] = 16'h0ff3;
  assign literal_11473[241] = 16'h1fed;
  assign literal_11473[242] = 16'hffae;
  assign literal_11473[243] = 16'hffb0;
  assign literal_11473[244] = 16'hffb4;
  assign literal_11473[245] = 16'hffbe;
  assign literal_11473[246] = 16'hffc8;
  assign literal_11473[247] = 16'hffd5;
  assign literal_11473[248] = 16'hffe2;
  assign literal_11473[249] = 16'hfff0;
  assign literal_11473[250] = 16'hfffe;
  assign literal_11473[251] = 16'h0000;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [2:0] p1_huff_length_squeezed_const_msb_bits_comb;
  wire [9:0] p1_row0_comb[0:7];
  wire [9:0] p1_row1_comb[0:7];
  wire [9:0] p1_array_concat_10453_comb[0:15];
  wire [9:0] p1_row2_comb[0:7];
  wire [9:0] p1_array_concat_10456_comb[0:23];
  wire [9:0] p1_row3_comb[0:7];
  wire [9:0] p1_array_concat_10459_comb[0:31];
  wire [9:0] p1_row4_comb[0:7];
  wire [9:0] p1_array_concat_10462_comb[0:39];
  wire [9:0] p1_row5_comb[0:7];
  wire p1_run__1_squeezed_const_msb_bits__6_comb;
  wire p1_run__1_squeezed_const_msb_bits_comb;
  wire [9:0] p1_array_concat_10468_comb[0:47];
  wire [9:0] p1_row6_comb[0:7];
  wire [7:0] p1_concat_10471_comb;
  wire [8:0] p1_concat_10473_comb;
  wire [9:0] p1_array_concat_10475_comb[0:55];
  wire [9:0] p1_row7_comb[0:7];
  wire [7:0] p1_add_10477_comb;
  wire [8:0] p1_add_10479_comb;
  wire [9:0] p1_flat_ac_comb[0:63];
  wire p1_run__1_squeezed_const_msb_bits__7_comb;
  wire p1_run__1_squeezed_const_msb_bits__8_comb;
  wire [8:0] p1_concat_10484_comb;
  wire [8:0] p1_add_10488_comb;
  wire [6:0] p1_concat_10489_comb;
  wire [6:0] p1_add_10499_comb;
  wire [7:0] p1_add_10514_comb;
  wire [5:0] p1_add_10543_comb;
  wire [7:0] p1_add_10555_comb;
  wire [6:0] p1_add_10568_comb;
  wire [7:0] p1_add_10585_comb;
  wire [8:0] p1_concat_10509_comb;
  wire [8:0] p1_add_10515_comb;
  wire [8:0] p1_concat_10524_comb;
  wire [8:0] p1_add_10531_comb;
  wire [8:0] p1_concat_10552_comb;
  wire [8:0] p1_add_10556_comb;
  wire [8:0] p1_concat_10562_comb;
  wire [8:0] p1_add_10569_comb;
  wire [8:0] p1_concat_10578_comb;
  wire [8:0] p1_add_10586_comb;
  wire [8:0] p1_concat_10593_comb;
  wire [8:0] p1_add_10607_comb;
  wire [1:0] p1_and_10530_comb;
  wire p1_or_10539_comb;
  wire p1_or_10547_comb;
  wire p1_or_10553_comb;
  wire p1_nor_10554_comb;
  wire p1_or_10575_comb;
  wire p1_or_10584_comb;
  wire p1_or_10592_comb;
  wire p1_or_10599_comb;
  wire p1_or_10606_comb;
  wire p1_or_10610_comb;
  wire p1_or_10614_comb;
  wire p1_nor_10617_comb;
  assign p1_huff_length_squeezed_const_msb_bits_comb = 3'h0;
  assign p1_row0_comb[0] = p0_matrix[p1_huff_length_squeezed_const_msb_bits_comb][0];
  assign p1_row0_comb[1] = p0_matrix[p1_huff_length_squeezed_const_msb_bits_comb][1];
  assign p1_row0_comb[2] = p0_matrix[p1_huff_length_squeezed_const_msb_bits_comb][2];
  assign p1_row0_comb[3] = p0_matrix[p1_huff_length_squeezed_const_msb_bits_comb][3];
  assign p1_row0_comb[4] = p0_matrix[p1_huff_length_squeezed_const_msb_bits_comb][4];
  assign p1_row0_comb[5] = p0_matrix[p1_huff_length_squeezed_const_msb_bits_comb][5];
  assign p1_row0_comb[6] = p0_matrix[p1_huff_length_squeezed_const_msb_bits_comb][6];
  assign p1_row0_comb[7] = p0_matrix[p1_huff_length_squeezed_const_msb_bits_comb][7];
  assign p1_row1_comb[0] = p0_matrix[3'h1][0];
  assign p1_row1_comb[1] = p0_matrix[3'h1][1];
  assign p1_row1_comb[2] = p0_matrix[3'h1][2];
  assign p1_row1_comb[3] = p0_matrix[3'h1][3];
  assign p1_row1_comb[4] = p0_matrix[3'h1][4];
  assign p1_row1_comb[5] = p0_matrix[3'h1][5];
  assign p1_row1_comb[6] = p0_matrix[3'h1][6];
  assign p1_row1_comb[7] = p0_matrix[3'h1][7];
  assign p1_array_concat_10453_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_10453_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_10453_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_10453_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_10453_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_10453_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_10453_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_10453_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_10453_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_10453_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_10453_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_10453_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_10453_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_10453_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_10453_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_10453_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_10456_comb[0] = p1_array_concat_10453_comb[0];
  assign p1_array_concat_10456_comb[1] = p1_array_concat_10453_comb[1];
  assign p1_array_concat_10456_comb[2] = p1_array_concat_10453_comb[2];
  assign p1_array_concat_10456_comb[3] = p1_array_concat_10453_comb[3];
  assign p1_array_concat_10456_comb[4] = p1_array_concat_10453_comb[4];
  assign p1_array_concat_10456_comb[5] = p1_array_concat_10453_comb[5];
  assign p1_array_concat_10456_comb[6] = p1_array_concat_10453_comb[6];
  assign p1_array_concat_10456_comb[7] = p1_array_concat_10453_comb[7];
  assign p1_array_concat_10456_comb[8] = p1_array_concat_10453_comb[8];
  assign p1_array_concat_10456_comb[9] = p1_array_concat_10453_comb[9];
  assign p1_array_concat_10456_comb[10] = p1_array_concat_10453_comb[10];
  assign p1_array_concat_10456_comb[11] = p1_array_concat_10453_comb[11];
  assign p1_array_concat_10456_comb[12] = p1_array_concat_10453_comb[12];
  assign p1_array_concat_10456_comb[13] = p1_array_concat_10453_comb[13];
  assign p1_array_concat_10456_comb[14] = p1_array_concat_10453_comb[14];
  assign p1_array_concat_10456_comb[15] = p1_array_concat_10453_comb[15];
  assign p1_array_concat_10456_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_10456_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_10456_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_10456_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_10456_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_10456_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_10456_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_10456_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_array_concat_10459_comb[0] = p1_array_concat_10456_comb[0];
  assign p1_array_concat_10459_comb[1] = p1_array_concat_10456_comb[1];
  assign p1_array_concat_10459_comb[2] = p1_array_concat_10456_comb[2];
  assign p1_array_concat_10459_comb[3] = p1_array_concat_10456_comb[3];
  assign p1_array_concat_10459_comb[4] = p1_array_concat_10456_comb[4];
  assign p1_array_concat_10459_comb[5] = p1_array_concat_10456_comb[5];
  assign p1_array_concat_10459_comb[6] = p1_array_concat_10456_comb[6];
  assign p1_array_concat_10459_comb[7] = p1_array_concat_10456_comb[7];
  assign p1_array_concat_10459_comb[8] = p1_array_concat_10456_comb[8];
  assign p1_array_concat_10459_comb[9] = p1_array_concat_10456_comb[9];
  assign p1_array_concat_10459_comb[10] = p1_array_concat_10456_comb[10];
  assign p1_array_concat_10459_comb[11] = p1_array_concat_10456_comb[11];
  assign p1_array_concat_10459_comb[12] = p1_array_concat_10456_comb[12];
  assign p1_array_concat_10459_comb[13] = p1_array_concat_10456_comb[13];
  assign p1_array_concat_10459_comb[14] = p1_array_concat_10456_comb[14];
  assign p1_array_concat_10459_comb[15] = p1_array_concat_10456_comb[15];
  assign p1_array_concat_10459_comb[16] = p1_array_concat_10456_comb[16];
  assign p1_array_concat_10459_comb[17] = p1_array_concat_10456_comb[17];
  assign p1_array_concat_10459_comb[18] = p1_array_concat_10456_comb[18];
  assign p1_array_concat_10459_comb[19] = p1_array_concat_10456_comb[19];
  assign p1_array_concat_10459_comb[20] = p1_array_concat_10456_comb[20];
  assign p1_array_concat_10459_comb[21] = p1_array_concat_10456_comb[21];
  assign p1_array_concat_10459_comb[22] = p1_array_concat_10456_comb[22];
  assign p1_array_concat_10459_comb[23] = p1_array_concat_10456_comb[23];
  assign p1_array_concat_10459_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_10459_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_10459_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_10459_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_10459_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_10459_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_10459_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_10459_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[3'h4][0];
  assign p1_row4_comb[1] = p0_matrix[3'h4][1];
  assign p1_row4_comb[2] = p0_matrix[3'h4][2];
  assign p1_row4_comb[3] = p0_matrix[3'h4][3];
  assign p1_row4_comb[4] = p0_matrix[3'h4][4];
  assign p1_row4_comb[5] = p0_matrix[3'h4][5];
  assign p1_row4_comb[6] = p0_matrix[3'h4][6];
  assign p1_row4_comb[7] = p0_matrix[3'h4][7];
  assign p1_array_concat_10462_comb[0] = p1_array_concat_10459_comb[0];
  assign p1_array_concat_10462_comb[1] = p1_array_concat_10459_comb[1];
  assign p1_array_concat_10462_comb[2] = p1_array_concat_10459_comb[2];
  assign p1_array_concat_10462_comb[3] = p1_array_concat_10459_comb[3];
  assign p1_array_concat_10462_comb[4] = p1_array_concat_10459_comb[4];
  assign p1_array_concat_10462_comb[5] = p1_array_concat_10459_comb[5];
  assign p1_array_concat_10462_comb[6] = p1_array_concat_10459_comb[6];
  assign p1_array_concat_10462_comb[7] = p1_array_concat_10459_comb[7];
  assign p1_array_concat_10462_comb[8] = p1_array_concat_10459_comb[8];
  assign p1_array_concat_10462_comb[9] = p1_array_concat_10459_comb[9];
  assign p1_array_concat_10462_comb[10] = p1_array_concat_10459_comb[10];
  assign p1_array_concat_10462_comb[11] = p1_array_concat_10459_comb[11];
  assign p1_array_concat_10462_comb[12] = p1_array_concat_10459_comb[12];
  assign p1_array_concat_10462_comb[13] = p1_array_concat_10459_comb[13];
  assign p1_array_concat_10462_comb[14] = p1_array_concat_10459_comb[14];
  assign p1_array_concat_10462_comb[15] = p1_array_concat_10459_comb[15];
  assign p1_array_concat_10462_comb[16] = p1_array_concat_10459_comb[16];
  assign p1_array_concat_10462_comb[17] = p1_array_concat_10459_comb[17];
  assign p1_array_concat_10462_comb[18] = p1_array_concat_10459_comb[18];
  assign p1_array_concat_10462_comb[19] = p1_array_concat_10459_comb[19];
  assign p1_array_concat_10462_comb[20] = p1_array_concat_10459_comb[20];
  assign p1_array_concat_10462_comb[21] = p1_array_concat_10459_comb[21];
  assign p1_array_concat_10462_comb[22] = p1_array_concat_10459_comb[22];
  assign p1_array_concat_10462_comb[23] = p1_array_concat_10459_comb[23];
  assign p1_array_concat_10462_comb[24] = p1_array_concat_10459_comb[24];
  assign p1_array_concat_10462_comb[25] = p1_array_concat_10459_comb[25];
  assign p1_array_concat_10462_comb[26] = p1_array_concat_10459_comb[26];
  assign p1_array_concat_10462_comb[27] = p1_array_concat_10459_comb[27];
  assign p1_array_concat_10462_comb[28] = p1_array_concat_10459_comb[28];
  assign p1_array_concat_10462_comb[29] = p1_array_concat_10459_comb[29];
  assign p1_array_concat_10462_comb[30] = p1_array_concat_10459_comb[30];
  assign p1_array_concat_10462_comb[31] = p1_array_concat_10459_comb[31];
  assign p1_array_concat_10462_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_10462_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_10462_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_10462_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_10462_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_10462_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_10462_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_10462_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[3'h5][0];
  assign p1_row5_comb[1] = p0_matrix[3'h5][1];
  assign p1_row5_comb[2] = p0_matrix[3'h5][2];
  assign p1_row5_comb[3] = p0_matrix[3'h5][3];
  assign p1_row5_comb[4] = p0_matrix[3'h5][4];
  assign p1_row5_comb[5] = p0_matrix[3'h5][5];
  assign p1_row5_comb[6] = p0_matrix[3'h5][6];
  assign p1_row5_comb[7] = p0_matrix[3'h5][7];
  assign p1_run__1_squeezed_const_msb_bits__6_comb = 1'h0;
  assign p1_run__1_squeezed_const_msb_bits_comb = 1'h0;
  assign p1_array_concat_10468_comb[0] = p1_array_concat_10462_comb[0];
  assign p1_array_concat_10468_comb[1] = p1_array_concat_10462_comb[1];
  assign p1_array_concat_10468_comb[2] = p1_array_concat_10462_comb[2];
  assign p1_array_concat_10468_comb[3] = p1_array_concat_10462_comb[3];
  assign p1_array_concat_10468_comb[4] = p1_array_concat_10462_comb[4];
  assign p1_array_concat_10468_comb[5] = p1_array_concat_10462_comb[5];
  assign p1_array_concat_10468_comb[6] = p1_array_concat_10462_comb[6];
  assign p1_array_concat_10468_comb[7] = p1_array_concat_10462_comb[7];
  assign p1_array_concat_10468_comb[8] = p1_array_concat_10462_comb[8];
  assign p1_array_concat_10468_comb[9] = p1_array_concat_10462_comb[9];
  assign p1_array_concat_10468_comb[10] = p1_array_concat_10462_comb[10];
  assign p1_array_concat_10468_comb[11] = p1_array_concat_10462_comb[11];
  assign p1_array_concat_10468_comb[12] = p1_array_concat_10462_comb[12];
  assign p1_array_concat_10468_comb[13] = p1_array_concat_10462_comb[13];
  assign p1_array_concat_10468_comb[14] = p1_array_concat_10462_comb[14];
  assign p1_array_concat_10468_comb[15] = p1_array_concat_10462_comb[15];
  assign p1_array_concat_10468_comb[16] = p1_array_concat_10462_comb[16];
  assign p1_array_concat_10468_comb[17] = p1_array_concat_10462_comb[17];
  assign p1_array_concat_10468_comb[18] = p1_array_concat_10462_comb[18];
  assign p1_array_concat_10468_comb[19] = p1_array_concat_10462_comb[19];
  assign p1_array_concat_10468_comb[20] = p1_array_concat_10462_comb[20];
  assign p1_array_concat_10468_comb[21] = p1_array_concat_10462_comb[21];
  assign p1_array_concat_10468_comb[22] = p1_array_concat_10462_comb[22];
  assign p1_array_concat_10468_comb[23] = p1_array_concat_10462_comb[23];
  assign p1_array_concat_10468_comb[24] = p1_array_concat_10462_comb[24];
  assign p1_array_concat_10468_comb[25] = p1_array_concat_10462_comb[25];
  assign p1_array_concat_10468_comb[26] = p1_array_concat_10462_comb[26];
  assign p1_array_concat_10468_comb[27] = p1_array_concat_10462_comb[27];
  assign p1_array_concat_10468_comb[28] = p1_array_concat_10462_comb[28];
  assign p1_array_concat_10468_comb[29] = p1_array_concat_10462_comb[29];
  assign p1_array_concat_10468_comb[30] = p1_array_concat_10462_comb[30];
  assign p1_array_concat_10468_comb[31] = p1_array_concat_10462_comb[31];
  assign p1_array_concat_10468_comb[32] = p1_array_concat_10462_comb[32];
  assign p1_array_concat_10468_comb[33] = p1_array_concat_10462_comb[33];
  assign p1_array_concat_10468_comb[34] = p1_array_concat_10462_comb[34];
  assign p1_array_concat_10468_comb[35] = p1_array_concat_10462_comb[35];
  assign p1_array_concat_10468_comb[36] = p1_array_concat_10462_comb[36];
  assign p1_array_concat_10468_comb[37] = p1_array_concat_10462_comb[37];
  assign p1_array_concat_10468_comb[38] = p1_array_concat_10462_comb[38];
  assign p1_array_concat_10468_comb[39] = p1_array_concat_10462_comb[39];
  assign p1_array_concat_10468_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_10468_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_10468_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_10468_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_10468_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_10468_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_10468_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_10468_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[3'h6][0];
  assign p1_row6_comb[1] = p0_matrix[3'h6][1];
  assign p1_row6_comb[2] = p0_matrix[3'h6][2];
  assign p1_row6_comb[3] = p0_matrix[3'h6][3];
  assign p1_row6_comb[4] = p0_matrix[3'h6][4];
  assign p1_row6_comb[5] = p0_matrix[3'h6][5];
  assign p1_row6_comb[6] = p0_matrix[3'h6][6];
  assign p1_row6_comb[7] = p0_matrix[3'h6][7];
  assign p1_concat_10471_comb = {p1_run__1_squeezed_const_msb_bits__6_comb, p0_start_pix[7:1]};
  assign p1_concat_10473_comb = {p1_run__1_squeezed_const_msb_bits_comb, p0_start_pix};
  assign p1_array_concat_10475_comb[0] = p1_array_concat_10468_comb[0];
  assign p1_array_concat_10475_comb[1] = p1_array_concat_10468_comb[1];
  assign p1_array_concat_10475_comb[2] = p1_array_concat_10468_comb[2];
  assign p1_array_concat_10475_comb[3] = p1_array_concat_10468_comb[3];
  assign p1_array_concat_10475_comb[4] = p1_array_concat_10468_comb[4];
  assign p1_array_concat_10475_comb[5] = p1_array_concat_10468_comb[5];
  assign p1_array_concat_10475_comb[6] = p1_array_concat_10468_comb[6];
  assign p1_array_concat_10475_comb[7] = p1_array_concat_10468_comb[7];
  assign p1_array_concat_10475_comb[8] = p1_array_concat_10468_comb[8];
  assign p1_array_concat_10475_comb[9] = p1_array_concat_10468_comb[9];
  assign p1_array_concat_10475_comb[10] = p1_array_concat_10468_comb[10];
  assign p1_array_concat_10475_comb[11] = p1_array_concat_10468_comb[11];
  assign p1_array_concat_10475_comb[12] = p1_array_concat_10468_comb[12];
  assign p1_array_concat_10475_comb[13] = p1_array_concat_10468_comb[13];
  assign p1_array_concat_10475_comb[14] = p1_array_concat_10468_comb[14];
  assign p1_array_concat_10475_comb[15] = p1_array_concat_10468_comb[15];
  assign p1_array_concat_10475_comb[16] = p1_array_concat_10468_comb[16];
  assign p1_array_concat_10475_comb[17] = p1_array_concat_10468_comb[17];
  assign p1_array_concat_10475_comb[18] = p1_array_concat_10468_comb[18];
  assign p1_array_concat_10475_comb[19] = p1_array_concat_10468_comb[19];
  assign p1_array_concat_10475_comb[20] = p1_array_concat_10468_comb[20];
  assign p1_array_concat_10475_comb[21] = p1_array_concat_10468_comb[21];
  assign p1_array_concat_10475_comb[22] = p1_array_concat_10468_comb[22];
  assign p1_array_concat_10475_comb[23] = p1_array_concat_10468_comb[23];
  assign p1_array_concat_10475_comb[24] = p1_array_concat_10468_comb[24];
  assign p1_array_concat_10475_comb[25] = p1_array_concat_10468_comb[25];
  assign p1_array_concat_10475_comb[26] = p1_array_concat_10468_comb[26];
  assign p1_array_concat_10475_comb[27] = p1_array_concat_10468_comb[27];
  assign p1_array_concat_10475_comb[28] = p1_array_concat_10468_comb[28];
  assign p1_array_concat_10475_comb[29] = p1_array_concat_10468_comb[29];
  assign p1_array_concat_10475_comb[30] = p1_array_concat_10468_comb[30];
  assign p1_array_concat_10475_comb[31] = p1_array_concat_10468_comb[31];
  assign p1_array_concat_10475_comb[32] = p1_array_concat_10468_comb[32];
  assign p1_array_concat_10475_comb[33] = p1_array_concat_10468_comb[33];
  assign p1_array_concat_10475_comb[34] = p1_array_concat_10468_comb[34];
  assign p1_array_concat_10475_comb[35] = p1_array_concat_10468_comb[35];
  assign p1_array_concat_10475_comb[36] = p1_array_concat_10468_comb[36];
  assign p1_array_concat_10475_comb[37] = p1_array_concat_10468_comb[37];
  assign p1_array_concat_10475_comb[38] = p1_array_concat_10468_comb[38];
  assign p1_array_concat_10475_comb[39] = p1_array_concat_10468_comb[39];
  assign p1_array_concat_10475_comb[40] = p1_array_concat_10468_comb[40];
  assign p1_array_concat_10475_comb[41] = p1_array_concat_10468_comb[41];
  assign p1_array_concat_10475_comb[42] = p1_array_concat_10468_comb[42];
  assign p1_array_concat_10475_comb[43] = p1_array_concat_10468_comb[43];
  assign p1_array_concat_10475_comb[44] = p1_array_concat_10468_comb[44];
  assign p1_array_concat_10475_comb[45] = p1_array_concat_10468_comb[45];
  assign p1_array_concat_10475_comb[46] = p1_array_concat_10468_comb[46];
  assign p1_array_concat_10475_comb[47] = p1_array_concat_10468_comb[47];
  assign p1_array_concat_10475_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_10475_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_10475_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_10475_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_10475_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_10475_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_10475_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_10475_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[3'h7][0];
  assign p1_row7_comb[1] = p0_matrix[3'h7][1];
  assign p1_row7_comb[2] = p0_matrix[3'h7][2];
  assign p1_row7_comb[3] = p0_matrix[3'h7][3];
  assign p1_row7_comb[4] = p0_matrix[3'h7][4];
  assign p1_row7_comb[5] = p0_matrix[3'h7][5];
  assign p1_row7_comb[6] = p0_matrix[3'h7][6];
  assign p1_row7_comb[7] = p0_matrix[3'h7][7];
  assign p1_add_10477_comb = p1_concat_10471_comb + 8'h07;
  assign p1_add_10479_comb = p1_concat_10473_comb + 9'h00f;
  assign p1_flat_ac_comb[0] = p1_array_concat_10475_comb[0];
  assign p1_flat_ac_comb[1] = p1_array_concat_10475_comb[1];
  assign p1_flat_ac_comb[2] = p1_array_concat_10475_comb[2];
  assign p1_flat_ac_comb[3] = p1_array_concat_10475_comb[3];
  assign p1_flat_ac_comb[4] = p1_array_concat_10475_comb[4];
  assign p1_flat_ac_comb[5] = p1_array_concat_10475_comb[5];
  assign p1_flat_ac_comb[6] = p1_array_concat_10475_comb[6];
  assign p1_flat_ac_comb[7] = p1_array_concat_10475_comb[7];
  assign p1_flat_ac_comb[8] = p1_array_concat_10475_comb[8];
  assign p1_flat_ac_comb[9] = p1_array_concat_10475_comb[9];
  assign p1_flat_ac_comb[10] = p1_array_concat_10475_comb[10];
  assign p1_flat_ac_comb[11] = p1_array_concat_10475_comb[11];
  assign p1_flat_ac_comb[12] = p1_array_concat_10475_comb[12];
  assign p1_flat_ac_comb[13] = p1_array_concat_10475_comb[13];
  assign p1_flat_ac_comb[14] = p1_array_concat_10475_comb[14];
  assign p1_flat_ac_comb[15] = p1_array_concat_10475_comb[15];
  assign p1_flat_ac_comb[16] = p1_array_concat_10475_comb[16];
  assign p1_flat_ac_comb[17] = p1_array_concat_10475_comb[17];
  assign p1_flat_ac_comb[18] = p1_array_concat_10475_comb[18];
  assign p1_flat_ac_comb[19] = p1_array_concat_10475_comb[19];
  assign p1_flat_ac_comb[20] = p1_array_concat_10475_comb[20];
  assign p1_flat_ac_comb[21] = p1_array_concat_10475_comb[21];
  assign p1_flat_ac_comb[22] = p1_array_concat_10475_comb[22];
  assign p1_flat_ac_comb[23] = p1_array_concat_10475_comb[23];
  assign p1_flat_ac_comb[24] = p1_array_concat_10475_comb[24];
  assign p1_flat_ac_comb[25] = p1_array_concat_10475_comb[25];
  assign p1_flat_ac_comb[26] = p1_array_concat_10475_comb[26];
  assign p1_flat_ac_comb[27] = p1_array_concat_10475_comb[27];
  assign p1_flat_ac_comb[28] = p1_array_concat_10475_comb[28];
  assign p1_flat_ac_comb[29] = p1_array_concat_10475_comb[29];
  assign p1_flat_ac_comb[30] = p1_array_concat_10475_comb[30];
  assign p1_flat_ac_comb[31] = p1_array_concat_10475_comb[31];
  assign p1_flat_ac_comb[32] = p1_array_concat_10475_comb[32];
  assign p1_flat_ac_comb[33] = p1_array_concat_10475_comb[33];
  assign p1_flat_ac_comb[34] = p1_array_concat_10475_comb[34];
  assign p1_flat_ac_comb[35] = p1_array_concat_10475_comb[35];
  assign p1_flat_ac_comb[36] = p1_array_concat_10475_comb[36];
  assign p1_flat_ac_comb[37] = p1_array_concat_10475_comb[37];
  assign p1_flat_ac_comb[38] = p1_array_concat_10475_comb[38];
  assign p1_flat_ac_comb[39] = p1_array_concat_10475_comb[39];
  assign p1_flat_ac_comb[40] = p1_array_concat_10475_comb[40];
  assign p1_flat_ac_comb[41] = p1_array_concat_10475_comb[41];
  assign p1_flat_ac_comb[42] = p1_array_concat_10475_comb[42];
  assign p1_flat_ac_comb[43] = p1_array_concat_10475_comb[43];
  assign p1_flat_ac_comb[44] = p1_array_concat_10475_comb[44];
  assign p1_flat_ac_comb[45] = p1_array_concat_10475_comb[45];
  assign p1_flat_ac_comb[46] = p1_array_concat_10475_comb[46];
  assign p1_flat_ac_comb[47] = p1_array_concat_10475_comb[47];
  assign p1_flat_ac_comb[48] = p1_array_concat_10475_comb[48];
  assign p1_flat_ac_comb[49] = p1_array_concat_10475_comb[49];
  assign p1_flat_ac_comb[50] = p1_array_concat_10475_comb[50];
  assign p1_flat_ac_comb[51] = p1_array_concat_10475_comb[51];
  assign p1_flat_ac_comb[52] = p1_array_concat_10475_comb[52];
  assign p1_flat_ac_comb[53] = p1_array_concat_10475_comb[53];
  assign p1_flat_ac_comb[54] = p1_array_concat_10475_comb[54];
  assign p1_flat_ac_comb[55] = p1_array_concat_10475_comb[55];
  assign p1_flat_ac_comb[56] = p1_row7_comb[0];
  assign p1_flat_ac_comb[57] = p1_row7_comb[1];
  assign p1_flat_ac_comb[58] = p1_row7_comb[2];
  assign p1_flat_ac_comb[59] = p1_row7_comb[3];
  assign p1_flat_ac_comb[60] = p1_row7_comb[4];
  assign p1_flat_ac_comb[61] = p1_row7_comb[5];
  assign p1_flat_ac_comb[62] = p1_row7_comb[6];
  assign p1_flat_ac_comb[63] = p1_row7_comb[7];
  assign p1_run__1_squeezed_const_msb_bits__7_comb = 1'h0;
  assign p1_run__1_squeezed_const_msb_bits__8_comb = 1'h0;
  assign p1_concat_10484_comb = {p1_add_10477_comb, p0_start_pix[0]};
  assign p1_add_10488_comb = p1_concat_10473_comb + 9'h00d;
  assign p1_concat_10489_comb = {p1_run__1_squeezed_const_msb_bits__7_comb, p0_start_pix[7:2]};
  assign p1_add_10499_comb = p1_concat_10489_comb + 7'h03;
  assign p1_add_10514_comb = p1_concat_10471_comb + 8'h05;
  assign p1_add_10543_comb = {p1_run__1_squeezed_const_msb_bits__8_comb, p0_start_pix[7:3]} + 6'h01;
  assign p1_add_10555_comb = p1_concat_10471_comb + 8'h03;
  assign p1_add_10568_comb = p1_concat_10489_comb + 7'h01;
  assign p1_add_10585_comb = p1_concat_10471_comb + 8'h01;
  assign p1_concat_10509_comb = {p1_add_10499_comb, p0_start_pix[1:0]};
  assign p1_add_10515_comb = p1_concat_10473_comb + 9'h00b;
  assign p1_concat_10524_comb = {p1_add_10514_comb, p0_start_pix[0]};
  assign p1_add_10531_comb = p1_concat_10473_comb + 9'h009;
  assign p1_concat_10552_comb = {p1_add_10543_comb, p0_start_pix[2:0]};
  assign p1_add_10556_comb = p1_concat_10473_comb + 9'h007;
  assign p1_concat_10562_comb = {p1_add_10555_comb, p0_start_pix[0]};
  assign p1_add_10569_comb = p1_concat_10473_comb + 9'h005;
  assign p1_concat_10578_comb = {p1_add_10568_comb, p0_start_pix[1:0]};
  assign p1_add_10586_comb = p1_concat_10473_comb + 9'h003;
  assign p1_concat_10593_comb = {p1_add_10585_comb, p0_start_pix[0]};
  assign p1_add_10607_comb = p1_concat_10473_comb + 9'h001;
  assign p1_and_10530_comb = ((|p1_add_10477_comb[7:5]) | p1_flat_ac_comb[p1_concat_10484_comb > 9'h03f ? 6'h3f : p1_concat_10484_comb[5:0]] != 10'h000 ? 2'h1 : {1'h1, ~((|p1_add_10479_comb[8:6]) | p1_flat_ac_comb[p1_add_10479_comb > 9'h03f ? 6'h3f : p1_add_10479_comb[5:0]] != 10'h000)}) & {2{~((|p1_add_10488_comb[8:6]) | p1_flat_ac_comb[p1_add_10488_comb > 9'h03f ? 6'h3f : p1_add_10488_comb[5:0]] != 10'h000)}};
  assign p1_or_10539_comb = (|p1_add_10499_comb[6:4]) | p1_flat_ac_comb[p1_concat_10509_comb > 9'h03f ? 6'h3f : p1_concat_10509_comb[5:0]] != 10'h000;
  assign p1_or_10547_comb = (|p1_add_10515_comb[8:6]) | p1_flat_ac_comb[p1_add_10515_comb > 9'h03f ? 6'h3f : p1_add_10515_comb[5:0]] != 10'h000;
  assign p1_or_10553_comb = (|p1_add_10514_comb[7:5]) | p1_flat_ac_comb[p1_concat_10524_comb > 9'h03f ? 6'h3f : p1_concat_10524_comb[5:0]] != 10'h000;
  assign p1_nor_10554_comb = ~((|p1_add_10531_comb[8:6]) | p1_flat_ac_comb[p1_add_10531_comb > 9'h03f ? 6'h3f : p1_add_10531_comb[5:0]] != 10'h000);
  assign p1_or_10575_comb = (|p1_add_10543_comb[5:3]) | p1_flat_ac_comb[p1_concat_10552_comb > 9'h03f ? 6'h3f : p1_concat_10552_comb[5:0]] != 10'h000;
  assign p1_or_10584_comb = (|p1_add_10556_comb[8:6]) | p1_flat_ac_comb[p1_add_10556_comb > 9'h03f ? 6'h3f : p1_add_10556_comb[5:0]] != 10'h000;
  assign p1_or_10592_comb = (|p1_add_10555_comb[7:5]) | p1_flat_ac_comb[p1_concat_10562_comb > 9'h03f ? 6'h3f : p1_concat_10562_comb[5:0]] != 10'h000;
  assign p1_or_10599_comb = (|p1_add_10569_comb[8:6]) | p1_flat_ac_comb[p1_add_10569_comb > 9'h03f ? 6'h3f : p1_add_10569_comb[5:0]] != 10'h000;
  assign p1_or_10606_comb = (|p1_add_10568_comb[6:4]) | p1_flat_ac_comb[p1_concat_10578_comb > 9'h03f ? 6'h3f : p1_concat_10578_comb[5:0]] != 10'h000;
  assign p1_or_10610_comb = (|p1_add_10586_comb[8:6]) | p1_flat_ac_comb[p1_add_10586_comb > 9'h03f ? 6'h3f : p1_add_10586_comb[5:0]] != 10'h000;
  assign p1_or_10614_comb = (|p1_add_10585_comb[7:5]) | p1_flat_ac_comb[p1_concat_10593_comb > 9'h03f ? 6'h3f : p1_concat_10593_comb[5:0]] != 10'h000;
  assign p1_nor_10617_comb = ~(p1_add_10607_comb > 9'h03e | p1_flat_ac_comb[p1_add_10607_comb > 9'h03f ? 6'h3f : p1_add_10607_comb[5:0]] != 10'h000);

  // Registers for pipe stage 1:
  reg [7:0] p1_start_pix;
  reg p1_is_luminance;
  reg [9:0] p1_flat_ac[0:63];
  reg [1:0] p1_and_10530;
  reg p1_or_10539;
  reg p1_or_10547;
  reg p1_or_10553;
  reg p1_nor_10554;
  reg p1_or_10575;
  reg p1_or_10584;
  reg p1_or_10592;
  reg p1_or_10599;
  reg p1_or_10606;
  reg p1_or_10610;
  reg p1_or_10614;
  reg p1_nor_10617;
  always @ (posedge clk) begin
    p1_start_pix <= p0_start_pix;
    p1_is_luminance <= p0_is_luminance;
    p1_flat_ac[0] <= p1_flat_ac_comb[0];
    p1_flat_ac[1] <= p1_flat_ac_comb[1];
    p1_flat_ac[2] <= p1_flat_ac_comb[2];
    p1_flat_ac[3] <= p1_flat_ac_comb[3];
    p1_flat_ac[4] <= p1_flat_ac_comb[4];
    p1_flat_ac[5] <= p1_flat_ac_comb[5];
    p1_flat_ac[6] <= p1_flat_ac_comb[6];
    p1_flat_ac[7] <= p1_flat_ac_comb[7];
    p1_flat_ac[8] <= p1_flat_ac_comb[8];
    p1_flat_ac[9] <= p1_flat_ac_comb[9];
    p1_flat_ac[10] <= p1_flat_ac_comb[10];
    p1_flat_ac[11] <= p1_flat_ac_comb[11];
    p1_flat_ac[12] <= p1_flat_ac_comb[12];
    p1_flat_ac[13] <= p1_flat_ac_comb[13];
    p1_flat_ac[14] <= p1_flat_ac_comb[14];
    p1_flat_ac[15] <= p1_flat_ac_comb[15];
    p1_flat_ac[16] <= p1_flat_ac_comb[16];
    p1_flat_ac[17] <= p1_flat_ac_comb[17];
    p1_flat_ac[18] <= p1_flat_ac_comb[18];
    p1_flat_ac[19] <= p1_flat_ac_comb[19];
    p1_flat_ac[20] <= p1_flat_ac_comb[20];
    p1_flat_ac[21] <= p1_flat_ac_comb[21];
    p1_flat_ac[22] <= p1_flat_ac_comb[22];
    p1_flat_ac[23] <= p1_flat_ac_comb[23];
    p1_flat_ac[24] <= p1_flat_ac_comb[24];
    p1_flat_ac[25] <= p1_flat_ac_comb[25];
    p1_flat_ac[26] <= p1_flat_ac_comb[26];
    p1_flat_ac[27] <= p1_flat_ac_comb[27];
    p1_flat_ac[28] <= p1_flat_ac_comb[28];
    p1_flat_ac[29] <= p1_flat_ac_comb[29];
    p1_flat_ac[30] <= p1_flat_ac_comb[30];
    p1_flat_ac[31] <= p1_flat_ac_comb[31];
    p1_flat_ac[32] <= p1_flat_ac_comb[32];
    p1_flat_ac[33] <= p1_flat_ac_comb[33];
    p1_flat_ac[34] <= p1_flat_ac_comb[34];
    p1_flat_ac[35] <= p1_flat_ac_comb[35];
    p1_flat_ac[36] <= p1_flat_ac_comb[36];
    p1_flat_ac[37] <= p1_flat_ac_comb[37];
    p1_flat_ac[38] <= p1_flat_ac_comb[38];
    p1_flat_ac[39] <= p1_flat_ac_comb[39];
    p1_flat_ac[40] <= p1_flat_ac_comb[40];
    p1_flat_ac[41] <= p1_flat_ac_comb[41];
    p1_flat_ac[42] <= p1_flat_ac_comb[42];
    p1_flat_ac[43] <= p1_flat_ac_comb[43];
    p1_flat_ac[44] <= p1_flat_ac_comb[44];
    p1_flat_ac[45] <= p1_flat_ac_comb[45];
    p1_flat_ac[46] <= p1_flat_ac_comb[46];
    p1_flat_ac[47] <= p1_flat_ac_comb[47];
    p1_flat_ac[48] <= p1_flat_ac_comb[48];
    p1_flat_ac[49] <= p1_flat_ac_comb[49];
    p1_flat_ac[50] <= p1_flat_ac_comb[50];
    p1_flat_ac[51] <= p1_flat_ac_comb[51];
    p1_flat_ac[52] <= p1_flat_ac_comb[52];
    p1_flat_ac[53] <= p1_flat_ac_comb[53];
    p1_flat_ac[54] <= p1_flat_ac_comb[54];
    p1_flat_ac[55] <= p1_flat_ac_comb[55];
    p1_flat_ac[56] <= p1_flat_ac_comb[56];
    p1_flat_ac[57] <= p1_flat_ac_comb[57];
    p1_flat_ac[58] <= p1_flat_ac_comb[58];
    p1_flat_ac[59] <= p1_flat_ac_comb[59];
    p1_flat_ac[60] <= p1_flat_ac_comb[60];
    p1_flat_ac[61] <= p1_flat_ac_comb[61];
    p1_flat_ac[62] <= p1_flat_ac_comb[62];
    p1_flat_ac[63] <= p1_flat_ac_comb[63];
    p1_and_10530 <= p1_and_10530_comb;
    p1_or_10539 <= p1_or_10539_comb;
    p1_or_10547 <= p1_or_10547_comb;
    p1_or_10553 <= p1_or_10553_comb;
    p1_nor_10554 <= p1_nor_10554_comb;
    p1_or_10575 <= p1_or_10575_comb;
    p1_or_10584 <= p1_or_10584_comb;
    p1_or_10592 <= p1_or_10592_comb;
    p1_or_10599 <= p1_or_10599_comb;
    p1_or_10606 <= p1_or_10606_comb;
    p1_or_10610 <= p1_or_10610_comb;
    p1_or_10614 <= p1_or_10614_comb;
    p1_nor_10617 <= p1_nor_10617_comb;
  end

  // ===== Pipe stage 2:
  wire [2:0] p2_and_10660_comb;
  wire [3:0] p2_sel_10669_comb;
  wire p2_run__1_squeezed_const_msb_bits__4_comb;
  wire [4:0] p2_concat_10677_comb;
  wire [4:0] p2_sign_ext_10678_comb;
  assign p2_and_10660_comb = (p1_or_10553 ? 3'h1 : (p1_or_10547 ? 3'h2 : (p1_or_10539 ? 3'h3 : {1'h1, p1_and_10530}))) & {3{p1_nor_10554}};
  assign p2_sel_10669_comb = p1_or_10599 ? 4'h4 : (p1_or_10592 ? 4'h5 : (p1_or_10584 ? 4'h6 : (p1_or_10575 ? 4'h7 : {1'h1, p2_and_10660_comb})));
  assign p2_run__1_squeezed_const_msb_bits__4_comb = 1'h0;
  assign p2_concat_10677_comb = {p2_run__1_squeezed_const_msb_bits__4_comb, p1_or_10614 ? 4'h1 : (p1_or_10610 ? 4'h2 : (p1_or_10606 ? 4'h3 : p2_sel_10669_comb))};
  assign p2_sign_ext_10678_comb = {5{p1_nor_10617}};

  // Registers for pipe stage 2:
  reg [7:0] p2_start_pix;
  reg p2_is_luminance;
  reg [9:0] p2_flat_ac[0:63];
  reg [4:0] p2_concat_10677;
  reg [4:0] p2_sign_ext_10678;
  always @ (posedge clk) begin
    p2_start_pix <= p1_start_pix;
    p2_is_luminance <= p1_is_luminance;
    p2_flat_ac[0] <= p1_flat_ac[0];
    p2_flat_ac[1] <= p1_flat_ac[1];
    p2_flat_ac[2] <= p1_flat_ac[2];
    p2_flat_ac[3] <= p1_flat_ac[3];
    p2_flat_ac[4] <= p1_flat_ac[4];
    p2_flat_ac[5] <= p1_flat_ac[5];
    p2_flat_ac[6] <= p1_flat_ac[6];
    p2_flat_ac[7] <= p1_flat_ac[7];
    p2_flat_ac[8] <= p1_flat_ac[8];
    p2_flat_ac[9] <= p1_flat_ac[9];
    p2_flat_ac[10] <= p1_flat_ac[10];
    p2_flat_ac[11] <= p1_flat_ac[11];
    p2_flat_ac[12] <= p1_flat_ac[12];
    p2_flat_ac[13] <= p1_flat_ac[13];
    p2_flat_ac[14] <= p1_flat_ac[14];
    p2_flat_ac[15] <= p1_flat_ac[15];
    p2_flat_ac[16] <= p1_flat_ac[16];
    p2_flat_ac[17] <= p1_flat_ac[17];
    p2_flat_ac[18] <= p1_flat_ac[18];
    p2_flat_ac[19] <= p1_flat_ac[19];
    p2_flat_ac[20] <= p1_flat_ac[20];
    p2_flat_ac[21] <= p1_flat_ac[21];
    p2_flat_ac[22] <= p1_flat_ac[22];
    p2_flat_ac[23] <= p1_flat_ac[23];
    p2_flat_ac[24] <= p1_flat_ac[24];
    p2_flat_ac[25] <= p1_flat_ac[25];
    p2_flat_ac[26] <= p1_flat_ac[26];
    p2_flat_ac[27] <= p1_flat_ac[27];
    p2_flat_ac[28] <= p1_flat_ac[28];
    p2_flat_ac[29] <= p1_flat_ac[29];
    p2_flat_ac[30] <= p1_flat_ac[30];
    p2_flat_ac[31] <= p1_flat_ac[31];
    p2_flat_ac[32] <= p1_flat_ac[32];
    p2_flat_ac[33] <= p1_flat_ac[33];
    p2_flat_ac[34] <= p1_flat_ac[34];
    p2_flat_ac[35] <= p1_flat_ac[35];
    p2_flat_ac[36] <= p1_flat_ac[36];
    p2_flat_ac[37] <= p1_flat_ac[37];
    p2_flat_ac[38] <= p1_flat_ac[38];
    p2_flat_ac[39] <= p1_flat_ac[39];
    p2_flat_ac[40] <= p1_flat_ac[40];
    p2_flat_ac[41] <= p1_flat_ac[41];
    p2_flat_ac[42] <= p1_flat_ac[42];
    p2_flat_ac[43] <= p1_flat_ac[43];
    p2_flat_ac[44] <= p1_flat_ac[44];
    p2_flat_ac[45] <= p1_flat_ac[45];
    p2_flat_ac[46] <= p1_flat_ac[46];
    p2_flat_ac[47] <= p1_flat_ac[47];
    p2_flat_ac[48] <= p1_flat_ac[48];
    p2_flat_ac[49] <= p1_flat_ac[49];
    p2_flat_ac[50] <= p1_flat_ac[50];
    p2_flat_ac[51] <= p1_flat_ac[51];
    p2_flat_ac[52] <= p1_flat_ac[52];
    p2_flat_ac[53] <= p1_flat_ac[53];
    p2_flat_ac[54] <= p1_flat_ac[54];
    p2_flat_ac[55] <= p1_flat_ac[55];
    p2_flat_ac[56] <= p1_flat_ac[56];
    p2_flat_ac[57] <= p1_flat_ac[57];
    p2_flat_ac[58] <= p1_flat_ac[58];
    p2_flat_ac[59] <= p1_flat_ac[59];
    p2_flat_ac[60] <= p1_flat_ac[60];
    p2_flat_ac[61] <= p1_flat_ac[61];
    p2_flat_ac[62] <= p1_flat_ac[62];
    p2_flat_ac[63] <= p1_flat_ac[63];
    p2_concat_10677 <= p2_concat_10677_comb;
    p2_sign_ext_10678 <= p2_sign_ext_10678_comb;
  end

  // ===== Pipe stage 3:
  wire [4:0] p3_zero_num__1_comb;
  wire [9:0] p3_value_comb;
  wire [2:0] p3_huff_length_squeezed_const_msb_bits__1_comb;
  wire [4:0] p3_add_10694_comb;
  wire [7:0] p3_start_pix_1__1_comb;
  wire [7:0] p3_value_pix_num_comb;
  wire [7:0] p3_add_10699_comb;
  wire [7:0] p3_actual_index__65_comb;
  wire [6:0] p3_add_10797_comb;
  wire [7:0] p3_actual_index__67_comb;
  wire [5:0] p3_add_10799_comb;
  wire [7:0] p3_actual_index__69_comb;
  wire [6:0] p3_add_10801_comb;
  wire [7:0] p3_actual_index__71_comb;
  wire [4:0] p3_add_10803_comb;
  wire [7:0] p3_actual_index__73_comb;
  wire [6:0] p3_add_10805_comb;
  wire [7:0] p3_actual_index__75_comb;
  wire [5:0] p3_add_10807_comb;
  wire [7:0] p3_actual_index__77_comb;
  wire [6:0] p3_add_10809_comb;
  wire [7:0] p3_actual_index__79_comb;
  wire [3:0] p3_add_10811_comb;
  wire [7:0] p3_actual_index__81_comb;
  wire [6:0] p3_add_10813_comb;
  wire [7:0] p3_actual_index__83_comb;
  wire [5:0] p3_add_10815_comb;
  wire [7:0] p3_actual_index__85_comb;
  wire [6:0] p3_add_10817_comb;
  wire [7:0] p3_actual_index__87_comb;
  wire [4:0] p3_add_10819_comb;
  wire [7:0] p3_actual_index__89_comb;
  wire [6:0] p3_add_10821_comb;
  wire [7:0] p3_actual_index__91_comb;
  wire [5:0] p3_add_10823_comb;
  wire [7:0] p3_actual_index__93_comb;
  wire [6:0] p3_add_10825_comb;
  wire [7:0] p3_actual_index__95_comb;
  wire [2:0] p3_add_10827_comb;
  wire [7:0] p3_actual_index__97_comb;
  wire [6:0] p3_add_10829_comb;
  wire [7:0] p3_actual_index__99_comb;
  wire [5:0] p3_add_10831_comb;
  wire [7:0] p3_actual_index__101_comb;
  wire [6:0] p3_add_10833_comb;
  wire [7:0] p3_actual_index__103_comb;
  wire [4:0] p3_add_10835_comb;
  wire [7:0] p3_actual_index__105_comb;
  wire [6:0] p3_add_10837_comb;
  wire [7:0] p3_actual_index__107_comb;
  wire [5:0] p3_add_10839_comb;
  wire [7:0] p3_actual_index__109_comb;
  wire [6:0] p3_add_10841_comb;
  wire [7:0] p3_actual_index__111_comb;
  wire [3:0] p3_add_10843_comb;
  wire [7:0] p3_actual_index__113_comb;
  wire [6:0] p3_add_10845_comb;
  wire [7:0] p3_actual_index__115_comb;
  wire [5:0] p3_add_10847_comb;
  wire [7:0] p3_actual_index__117_comb;
  wire [6:0] p3_add_10849_comb;
  wire [7:0] p3_actual_index__119_comb;
  wire [4:0] p3_add_10851_comb;
  wire [7:0] p3_actual_index__121_comb;
  wire [6:0] p3_add_10853_comb;
  wire [7:0] p3_actual_index__123_comb;
  wire [5:0] p3_add_10855_comb;
  wire [7:0] p3_actual_index__125_comb;
  wire [6:0] p3_add_10857_comb;
  wire [7:0] p3_actual_index__127_comb;
  wire [9:0] p3_value__1_comb;
  wire [7:0] p3_bin_value__1_comb;
  wire [7:0] p3_actual_index__66_comb;
  wire [7:0] p3_actual_index__68_comb;
  wire [7:0] p3_actual_index__70_comb;
  wire [7:0] p3_actual_index__72_comb;
  wire [7:0] p3_actual_index__74_comb;
  wire [7:0] p3_actual_index__76_comb;
  wire [7:0] p3_actual_index__78_comb;
  wire [7:0] p3_actual_index__80_comb;
  wire [7:0] p3_actual_index__82_comb;
  wire [7:0] p3_actual_index__84_comb;
  wire [7:0] p3_actual_index__86_comb;
  wire [7:0] p3_actual_index__88_comb;
  wire [7:0] p3_actual_index__90_comb;
  wire [7:0] p3_actual_index__92_comb;
  wire [7:0] p3_actual_index__94_comb;
  wire [7:0] p3_actual_index__96_comb;
  wire [7:0] p3_actual_index__98_comb;
  wire [7:0] p3_actual_index__100_comb;
  wire [7:0] p3_actual_index__102_comb;
  wire [7:0] p3_actual_index__104_comb;
  wire [7:0] p3_actual_index__106_comb;
  wire [7:0] p3_actual_index__108_comb;
  wire [7:0] p3_actual_index__110_comb;
  wire [7:0] p3_actual_index__112_comb;
  wire [7:0] p3_actual_index__114_comb;
  wire [7:0] p3_actual_index__116_comb;
  wire [7:0] p3_actual_index__118_comb;
  wire [7:0] p3_actual_index__120_comb;
  wire [7:0] p3_actual_index__122_comb;
  wire [7:0] p3_actual_index__124_comb;
  wire [7:0] p3_actual_index__126_comb;
  wire [7:0] p3_bin_value_comb;
  wire [7:0] p3_value_abs_comb;
  wire p3_and_11412_comb;
  wire [7:0] p3_flipped_comb;
  wire p3_run__1_squeezed_const_msb_bits__1_comb;
  wire [7:0] p3_Code_list_comb;
  wire p3_or_reduce_10718_comb;
  wire [2:0] p3_concat_10719_comb;
  wire p3_or_reduce_10723_comb;
  wire p3_or_reduce_10726_comb;
  wire p3_or_reduce_10795_comb;
  wire p3_bit_slice_10995_comb;
  wire p3_eq_10996_comb;
  wire [4:0] p3_run__1_squeezed_comb;
  wire [7:0] p3_code_list_comb;
  assign p3_zero_num__1_comb = p2_concat_10677 & p2_sign_ext_10678;
  assign p3_value_comb = p2_flat_ac[p2_start_pix > 8'h3f ? 6'h3f : p2_start_pix[5:0]];
  assign p3_huff_length_squeezed_const_msb_bits__1_comb = 3'h0;
  assign p3_add_10694_comb = p3_zero_num__1_comb + 5'h01;
  assign p3_start_pix_1__1_comb = p2_start_pix > 8'h40 ? 8'h40 : p2_start_pix;
  assign p3_value_pix_num_comb = {p3_huff_length_squeezed_const_msb_bits__1_comb, p3_add_10694_comb} & {8{p3_value_comb == 10'h000}};
  assign p3_add_10699_comb = p2_start_pix + p3_value_pix_num_comb;
  assign p3_actual_index__65_comb = p3_start_pix_1__1_comb + 8'h01;
  assign p3_add_10797_comb = p3_start_pix_1__1_comb[7:1] + 7'h01;
  assign p3_actual_index__67_comb = p3_start_pix_1__1_comb + 8'h03;
  assign p3_add_10799_comb = p3_start_pix_1__1_comb[7:2] + 6'h01;
  assign p3_actual_index__69_comb = p3_start_pix_1__1_comb + 8'h05;
  assign p3_add_10801_comb = p3_start_pix_1__1_comb[7:1] + 7'h03;
  assign p3_actual_index__71_comb = p3_start_pix_1__1_comb + 8'h07;
  assign p3_add_10803_comb = p3_start_pix_1__1_comb[7:3] + 5'h01;
  assign p3_actual_index__73_comb = p3_start_pix_1__1_comb + 8'h09;
  assign p3_add_10805_comb = p3_start_pix_1__1_comb[7:1] + 7'h05;
  assign p3_actual_index__75_comb = p3_start_pix_1__1_comb + 8'h0b;
  assign p3_add_10807_comb = p3_start_pix_1__1_comb[7:2] + 6'h03;
  assign p3_actual_index__77_comb = p3_start_pix_1__1_comb + 8'h0d;
  assign p3_add_10809_comb = p3_start_pix_1__1_comb[7:1] + 7'h07;
  assign p3_actual_index__79_comb = p3_start_pix_1__1_comb + 8'h0f;
  assign p3_add_10811_comb = p3_start_pix_1__1_comb[7:4] + 4'h1;
  assign p3_actual_index__81_comb = p3_start_pix_1__1_comb + 8'h11;
  assign p3_add_10813_comb = p3_start_pix_1__1_comb[7:1] + 7'h09;
  assign p3_actual_index__83_comb = p3_start_pix_1__1_comb + 8'h13;
  assign p3_add_10815_comb = p3_start_pix_1__1_comb[7:2] + 6'h05;
  assign p3_actual_index__85_comb = p3_start_pix_1__1_comb + 8'h15;
  assign p3_add_10817_comb = p3_start_pix_1__1_comb[7:1] + 7'h0b;
  assign p3_actual_index__87_comb = p3_start_pix_1__1_comb + 8'h17;
  assign p3_add_10819_comb = p3_start_pix_1__1_comb[7:3] + 5'h03;
  assign p3_actual_index__89_comb = p3_start_pix_1__1_comb + 8'h19;
  assign p3_add_10821_comb = p3_start_pix_1__1_comb[7:1] + 7'h0d;
  assign p3_actual_index__91_comb = p3_start_pix_1__1_comb + 8'h1b;
  assign p3_add_10823_comb = p3_start_pix_1__1_comb[7:2] + 6'h07;
  assign p3_actual_index__93_comb = p3_start_pix_1__1_comb + 8'h1d;
  assign p3_add_10825_comb = p3_start_pix_1__1_comb[7:1] + 7'h0f;
  assign p3_actual_index__95_comb = p3_start_pix_1__1_comb + 8'h1f;
  assign p3_add_10827_comb = p3_start_pix_1__1_comb[7:5] + 3'h1;
  assign p3_actual_index__97_comb = p3_start_pix_1__1_comb + 8'h21;
  assign p3_add_10829_comb = p3_start_pix_1__1_comb[7:1] + 7'h11;
  assign p3_actual_index__99_comb = p3_start_pix_1__1_comb + 8'h23;
  assign p3_add_10831_comb = p3_start_pix_1__1_comb[7:2] + 6'h09;
  assign p3_actual_index__101_comb = p3_start_pix_1__1_comb + 8'h25;
  assign p3_add_10833_comb = p3_start_pix_1__1_comb[7:1] + 7'h13;
  assign p3_actual_index__103_comb = p3_start_pix_1__1_comb + 8'h27;
  assign p3_add_10835_comb = p3_start_pix_1__1_comb[7:3] + 5'h05;
  assign p3_actual_index__105_comb = p3_start_pix_1__1_comb + 8'h29;
  assign p3_add_10837_comb = p3_start_pix_1__1_comb[7:1] + 7'h15;
  assign p3_actual_index__107_comb = p3_start_pix_1__1_comb + 8'h2b;
  assign p3_add_10839_comb = p3_start_pix_1__1_comb[7:2] + 6'h0b;
  assign p3_actual_index__109_comb = p3_start_pix_1__1_comb + 8'h2d;
  assign p3_add_10841_comb = p3_start_pix_1__1_comb[7:1] + 7'h17;
  assign p3_actual_index__111_comb = p3_start_pix_1__1_comb + 8'h2f;
  assign p3_add_10843_comb = p3_start_pix_1__1_comb[7:4] + 4'h3;
  assign p3_actual_index__113_comb = p3_start_pix_1__1_comb + 8'h31;
  assign p3_add_10845_comb = p3_start_pix_1__1_comb[7:1] + 7'h19;
  assign p3_actual_index__115_comb = p3_start_pix_1__1_comb + 8'h33;
  assign p3_add_10847_comb = p3_start_pix_1__1_comb[7:2] + 6'h0d;
  assign p3_actual_index__117_comb = p3_start_pix_1__1_comb + 8'h35;
  assign p3_add_10849_comb = p3_start_pix_1__1_comb[7:1] + 7'h1b;
  assign p3_actual_index__119_comb = p3_start_pix_1__1_comb + 8'h37;
  assign p3_add_10851_comb = p3_start_pix_1__1_comb[7:3] + 5'h07;
  assign p3_actual_index__121_comb = p3_start_pix_1__1_comb + 8'h39;
  assign p3_add_10853_comb = p3_start_pix_1__1_comb[7:1] + 7'h1d;
  assign p3_actual_index__123_comb = p3_start_pix_1__1_comb + 8'h3b;
  assign p3_add_10855_comb = p3_start_pix_1__1_comb[7:2] + 6'h0f;
  assign p3_actual_index__125_comb = p3_start_pix_1__1_comb + 8'h3d;
  assign p3_add_10857_comb = p3_start_pix_1__1_comb[7:1] + 7'h1f;
  assign p3_actual_index__127_comb = p3_start_pix_1__1_comb + 8'h3f;
  assign p3_value__1_comb = p2_flat_ac[p3_add_10699_comb > 8'h3f ? 6'h3f : p3_add_10699_comb[5:0]];
  assign p3_bin_value__1_comb = p3_value__1_comb[7:0];
  assign p3_actual_index__66_comb = {p3_add_10797_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__68_comb = {p3_add_10799_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__70_comb = {p3_add_10801_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__72_comb = {p3_add_10803_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__74_comb = {p3_add_10805_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__76_comb = {p3_add_10807_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__78_comb = {p3_add_10809_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__80_comb = {p3_add_10811_comb, p3_start_pix_1__1_comb[3:0]};
  assign p3_actual_index__82_comb = {p3_add_10813_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__84_comb = {p3_add_10815_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__86_comb = {p3_add_10817_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__88_comb = {p3_add_10819_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__90_comb = {p3_add_10821_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__92_comb = {p3_add_10823_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__94_comb = {p3_add_10825_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__96_comb = {p3_add_10827_comb, p3_start_pix_1__1_comb[4:0]};
  assign p3_actual_index__98_comb = {p3_add_10829_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__100_comb = {p3_add_10831_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__102_comb = {p3_add_10833_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__104_comb = {p3_add_10835_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__106_comb = {p3_add_10837_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__108_comb = {p3_add_10839_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__110_comb = {p3_add_10841_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__112_comb = {p3_add_10843_comb, p3_start_pix_1__1_comb[3:0]};
  assign p3_actual_index__114_comb = {p3_add_10845_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__116_comb = {p3_add_10847_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__118_comb = {p3_add_10849_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__120_comb = {p3_add_10851_comb, p3_start_pix_1__1_comb[2:0]};
  assign p3_actual_index__122_comb = {p3_add_10853_comb, p3_start_pix_1__1_comb[0]};
  assign p3_actual_index__124_comb = {p3_add_10855_comb, p3_start_pix_1__1_comb[1:0]};
  assign p3_actual_index__126_comb = {p3_add_10857_comb, p3_start_pix_1__1_comb[0]};
  assign p3_bin_value_comb = -p3_bin_value__1_comb;
  assign p3_value_abs_comb = p3_value__1_comb[9] ? p3_bin_value_comb : p3_bin_value__1_comb;
  assign p3_and_11412_comb = (p3_value_comb & {10{~p3_start_pix_1__1_comb[6]}}) == 10'h000 & (p2_flat_ac[p3_actual_index__65_comb > 8'h3f ? 6'h3f : p3_actual_index__65_comb[5:0]] & {10{~(p3_actual_index__65_comb[6] | p3_actual_index__65_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__66_comb > 8'h3f ? 6'h3f : p3_actual_index__66_comb[5:0]] & {10{~(p3_add_10797_comb[5] | p3_add_10797_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__67_comb > 8'h3f ? 6'h3f : p3_actual_index__67_comb[5:0]] & {10{~(p3_actual_index__67_comb[6] | p3_actual_index__67_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__68_comb > 8'h3f ? 6'h3f : p3_actual_index__68_comb[5:0]] & {10{~(p3_add_10799_comb[4] | p3_add_10799_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__69_comb > 8'h3f ? 6'h3f : p3_actual_index__69_comb[5:0]] & {10{~(p3_actual_index__69_comb[6] | p3_actual_index__69_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__70_comb > 8'h3f ? 6'h3f : p3_actual_index__70_comb[5:0]] & {10{~(p3_add_10801_comb[5] | p3_add_10801_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__71_comb > 8'h3f ? 6'h3f : p3_actual_index__71_comb[5:0]] & {10{~(p3_actual_index__71_comb[6] | p3_actual_index__71_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__72_comb > 8'h3f ? 6'h3f : p3_actual_index__72_comb[5:0]] & {10{~(p3_add_10803_comb[3] | p3_add_10803_comb[4])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__73_comb > 8'h3f ? 6'h3f : p3_actual_index__73_comb[5:0]] & {10{~(p3_actual_index__73_comb[6] | p3_actual_index__73_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__74_comb > 8'h3f ? 6'h3f : p3_actual_index__74_comb[5:0]] & {10{~(p3_add_10805_comb[5] | p3_add_10805_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__75_comb > 8'h3f ? 6'h3f : p3_actual_index__75_comb[5:0]] & {10{~(p3_actual_index__75_comb[6] | p3_actual_index__75_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__76_comb > 8'h3f ? 6'h3f : p3_actual_index__76_comb[5:0]] & {10{~(p3_add_10807_comb[4] | p3_add_10807_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__77_comb > 8'h3f ? 6'h3f : p3_actual_index__77_comb[5:0]] & {10{~(p3_actual_index__77_comb[6] | p3_actual_index__77_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__78_comb > 8'h3f ? 6'h3f : p3_actual_index__78_comb[5:0]] & {10{~(p3_add_10809_comb[5] | p3_add_10809_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__79_comb > 8'h3f ? 6'h3f : p3_actual_index__79_comb[5:0]] & {10{~(p3_actual_index__79_comb[6] | p3_actual_index__79_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__80_comb > 8'h3f ? 6'h3f : p3_actual_index__80_comb[5:0]] & {10{~(p3_add_10811_comb[2] | p3_add_10811_comb[3])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__81_comb > 8'h3f ? 6'h3f : p3_actual_index__81_comb[5:0]] & {10{~(p3_actual_index__81_comb[6] | p3_actual_index__81_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__82_comb > 8'h3f ? 6'h3f : p3_actual_index__82_comb[5:0]] & {10{~(p3_add_10813_comb[5] | p3_add_10813_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__83_comb > 8'h3f ? 6'h3f : p3_actual_index__83_comb[5:0]] & {10{~(p3_actual_index__83_comb[6] | p3_actual_index__83_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__84_comb > 8'h3f ? 6'h3f : p3_actual_index__84_comb[5:0]] & {10{~(p3_add_10815_comb[4] | p3_add_10815_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__85_comb > 8'h3f ? 6'h3f : p3_actual_index__85_comb[5:0]] & {10{~(p3_actual_index__85_comb[6] | p3_actual_index__85_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__86_comb > 8'h3f ? 6'h3f : p3_actual_index__86_comb[5:0]] & {10{~(p3_add_10817_comb[5] | p3_add_10817_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__87_comb > 8'h3f ? 6'h3f : p3_actual_index__87_comb[5:0]] & {10{~(p3_actual_index__87_comb[6] | p3_actual_index__87_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__88_comb > 8'h3f ? 6'h3f : p3_actual_index__88_comb[5:0]] & {10{~(p3_add_10819_comb[3] | p3_add_10819_comb[4])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__89_comb > 8'h3f ? 6'h3f : p3_actual_index__89_comb[5:0]] & {10{~(p3_actual_index__89_comb[6] | p3_actual_index__89_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__90_comb > 8'h3f ? 6'h3f : p3_actual_index__90_comb[5:0]] & {10{~(p3_add_10821_comb[5] | p3_add_10821_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__91_comb > 8'h3f ? 6'h3f : p3_actual_index__91_comb[5:0]] & {10{~(p3_actual_index__91_comb[6] | p3_actual_index__91_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__92_comb > 8'h3f ? 6'h3f : p3_actual_index__92_comb[5:0]] & {10{~(p3_add_10823_comb[4] | p3_add_10823_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__93_comb > 8'h3f ? 6'h3f : p3_actual_index__93_comb[5:0]] & {10{~(p3_actual_index__93_comb[6] | p3_actual_index__93_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__94_comb > 8'h3f ? 6'h3f : p3_actual_index__94_comb[5:0]] & {10{~(p3_add_10825_comb[5] | p3_add_10825_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__95_comb > 8'h3f ? 6'h3f : p3_actual_index__95_comb[5:0]] & {10{~(p3_actual_index__95_comb[6] | p3_actual_index__95_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__96_comb > 8'h3f ? 6'h3f : p3_actual_index__96_comb[5:0]] & {10{~(p3_add_10827_comb[1] | p3_add_10827_comb[2])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__97_comb > 8'h3f ? 6'h3f : p3_actual_index__97_comb[5:0]] & {10{~(p3_actual_index__97_comb[6] | p3_actual_index__97_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__98_comb > 8'h3f ? 6'h3f : p3_actual_index__98_comb[5:0]] & {10{~(p3_add_10829_comb[5] | p3_add_10829_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__99_comb > 8'h3f ? 6'h3f : p3_actual_index__99_comb[5:0]] & {10{~(p3_actual_index__99_comb[6] | p3_actual_index__99_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__100_comb > 8'h3f ? 6'h3f : p3_actual_index__100_comb[5:0]] & {10{~(p3_add_10831_comb[4] | p3_add_10831_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__101_comb > 8'h3f ? 6'h3f : p3_actual_index__101_comb[5:0]] & {10{~(p3_actual_index__101_comb[6] | p3_actual_index__101_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__102_comb > 8'h3f ? 6'h3f : p3_actual_index__102_comb[5:0]] & {10{~(p3_add_10833_comb[5] | p3_add_10833_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__103_comb > 8'h3f ? 6'h3f : p3_actual_index__103_comb[5:0]] & {10{~(p3_actual_index__103_comb[6] | p3_actual_index__103_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__104_comb > 8'h3f ? 6'h3f : p3_actual_index__104_comb[5:0]] & {10{~(p3_add_10835_comb[3] | p3_add_10835_comb[4])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__105_comb > 8'h3f ? 6'h3f : p3_actual_index__105_comb[5:0]] & {10{~(p3_actual_index__105_comb[6] | p3_actual_index__105_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__106_comb > 8'h3f ? 6'h3f : p3_actual_index__106_comb[5:0]] & {10{~(p3_add_10837_comb[5] | p3_add_10837_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__107_comb > 8'h3f ? 6'h3f : p3_actual_index__107_comb[5:0]] & {10{~(p3_actual_index__107_comb[6] | p3_actual_index__107_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__108_comb > 8'h3f ? 6'h3f : p3_actual_index__108_comb[5:0]] & {10{~(p3_add_10839_comb[4] | p3_add_10839_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__109_comb > 8'h3f ? 6'h3f : p3_actual_index__109_comb[5:0]] & {10{~(p3_actual_index__109_comb[6] | p3_actual_index__109_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__110_comb > 8'h3f ? 6'h3f : p3_actual_index__110_comb[5:0]] & {10{~(p3_add_10841_comb[5] | p3_add_10841_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__111_comb > 8'h3f ? 6'h3f : p3_actual_index__111_comb[5:0]] & {10{~(p3_actual_index__111_comb[6] | p3_actual_index__111_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__112_comb > 8'h3f ? 6'h3f : p3_actual_index__112_comb[5:0]] & {10{~(p3_add_10843_comb[2] | p3_add_10843_comb[3])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__113_comb > 8'h3f ? 6'h3f : p3_actual_index__113_comb[5:0]] & {10{~(p3_actual_index__113_comb[6] | p3_actual_index__113_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__114_comb > 8'h3f ? 6'h3f : p3_actual_index__114_comb[5:0]] & {10{~(p3_add_10845_comb[5] | p3_add_10845_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__115_comb > 8'h3f ? 6'h3f : p3_actual_index__115_comb[5:0]] & {10{~(p3_actual_index__115_comb[6] | p3_actual_index__115_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__116_comb > 8'h3f ? 6'h3f : p3_actual_index__116_comb[5:0]] & {10{~(p3_add_10847_comb[4] | p3_add_10847_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__117_comb > 8'h3f ? 6'h3f : p3_actual_index__117_comb[5:0]] & {10{~(p3_actual_index__117_comb[6] | p3_actual_index__117_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__118_comb > 8'h3f ? 6'h3f : p3_actual_index__118_comb[5:0]] & {10{~(p3_add_10849_comb[5] | p3_add_10849_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__119_comb > 8'h3f ? 6'h3f : p3_actual_index__119_comb[5:0]] & {10{~(p3_actual_index__119_comb[6] | p3_actual_index__119_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__120_comb > 8'h3f ? 6'h3f : p3_actual_index__120_comb[5:0]] & {10{~(p3_add_10851_comb[3] | p3_add_10851_comb[4])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__121_comb > 8'h3f ? 6'h3f : p3_actual_index__121_comb[5:0]] & {10{~(p3_actual_index__121_comb[6] | p3_actual_index__121_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__122_comb > 8'h3f ? 6'h3f : p3_actual_index__122_comb[5:0]] & {10{~(p3_add_10853_comb[5] | p3_add_10853_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__123_comb > 8'h3f ? 6'h3f : p3_actual_index__123_comb[5:0]] & {10{~(p3_actual_index__123_comb[6] | p3_actual_index__123_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__124_comb > 8'h3f ? 6'h3f : p3_actual_index__124_comb[5:0]] & {10{~(p3_add_10855_comb[4] | p3_add_10855_comb[5])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__125_comb > 8'h3f ? 6'h3f : p3_actual_index__125_comb[5:0]] & {10{~(p3_actual_index__125_comb[6] | p3_actual_index__125_comb[7])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__126_comb > 8'h3f ? 6'h3f : p3_actual_index__126_comb[5:0]] & {10{~(p3_add_10857_comb[5] | p3_add_10857_comb[6])}}) == 10'h000 & (p2_flat_ac[p3_actual_index__127_comb > 8'h3f ? 6'h3f : p3_actual_index__127_comb[5:0]] & {10{~(p3_actual_index__127_comb[6] | p3_actual_index__127_comb[7])}}) == 10'h000;
  assign p3_flipped_comb = ~p3_bin_value_comb;
  assign p3_run__1_squeezed_const_msb_bits__1_comb = 1'h0;
  assign p3_Code_list_comb = $signed(p3_value__1_comb) <= $signed(10'h000) ? p3_flipped_comb : p3_bin_value__1_comb;
  assign p3_or_reduce_10718_comb = |p3_value_abs_comb[7:3];
  assign p3_concat_10719_comb = {p3_run__1_squeezed_const_msb_bits__1_comb, |p3_value_abs_comb[7:2] ? 2'h3 : (|p3_value_abs_comb[7:1] ? 2'h2 : 2'h1)};
  assign p3_or_reduce_10723_comb = |p3_value_abs_comb[7:4];
  assign p3_or_reduce_10726_comb = |p3_value_abs_comb[7:5];
  assign p3_or_reduce_10795_comb = |p3_value_abs_comb[7:6];
  assign p3_bit_slice_10995_comb = p3_value_abs_comb[7];
  assign p3_eq_10996_comb = p3_value_abs_comb == 8'h00;
  assign p3_run__1_squeezed_comb = p3_value_pix_num_comb[4] ? 5'h0f : p3_value_pix_num_comb[4:0];
  assign p3_code_list_comb = p3_Code_list_comb & {8{~p3_and_11412_comb}};

  // Registers for pipe stage 3:
  reg p3_is_luminance;
  reg [9:0] p3_value;
  reg p3_or_reduce_10718;
  reg [2:0] p3_concat_10719;
  reg p3_or_reduce_10723;
  reg p3_or_reduce_10726;
  reg p3_or_reduce_10795;
  reg p3_bit_slice_10995;
  reg p3_eq_10996;
  reg [4:0] p3_run__1_squeezed;
  reg p3_and_11412;
  reg [7:0] p3_code_list;
  always @ (posedge clk) begin
    p3_is_luminance <= p2_is_luminance;
    p3_value <= p3_value_comb;
    p3_or_reduce_10718 <= p3_or_reduce_10718_comb;
    p3_concat_10719 <= p3_concat_10719_comb;
    p3_or_reduce_10723 <= p3_or_reduce_10723_comb;
    p3_or_reduce_10726 <= p3_or_reduce_10726_comb;
    p3_or_reduce_10795 <= p3_or_reduce_10795_comb;
    p3_bit_slice_10995 <= p3_bit_slice_10995_comb;
    p3_eq_10996 <= p3_eq_10996_comb;
    p3_run__1_squeezed <= p3_run__1_squeezed_comb;
    p3_and_11412 <= p3_and_11412_comb;
    p3_code_list <= p3_code_list_comb;
  end

  // ===== Pipe stage 4:
  wire p4_run__1_squeezed_const_msb_bits__2_comb;
  wire [3:0] p4_concat_11453_comb;
  wire [7:0] p4_concat_11460_comb;
  wire [7:0] p4_Code_size_comb;
  wire [7:0] p4_run_size_str_u8_comb;
  wire p4_run__1_squeezed_const_msb_bits__5_comb;
  wire [2:0] p4_sel_11474_comb;
  wire [1:0] p4_next_pix_squeezed_const_msb_bits_comb;
  wire p4_run__1_squeezed_const_msb_bits__3_comb;
  wire [5:0] p4_run__1_comb;
  wire [4:0] p4_Huffman_length_squeezed_comb;
  wire [5:0] p4_next_pix__1_squeezed_comb;
  wire [15:0] p4_Huffman_code_full_comb;
  wire [2:0] p4_huff_length_squeezed_const_msb_bits__2_comb;
  wire [4:0] p4_huff_length_squeezed_comb;
  wire [1:0] p4_next_pix_squeezed_const_msb_bits__1_comb;
  wire [5:0] p4_next_pix_squeezed_comb;
  wire [15:0] p4_huff_code_comb;
  wire [7:0] p4_huff_length_comb;
  wire [7:0] p4_code_size_comb;
  wire [7:0] p4_next_pix_comb;
  wire [57:0] p4_tuple_11503_comb;
  assign p4_run__1_squeezed_const_msb_bits__2_comb = 1'h0;
  assign p4_concat_11453_comb = {p4_run__1_squeezed_const_msb_bits__2_comb, p3_or_reduce_10795 ? 3'h7 : (p3_or_reduce_10726 ? 3'h6 : (p3_or_reduce_10723 ? 3'h5 : (p3_or_reduce_10718 ? 3'h4 : p3_concat_10719)))};
  assign p4_concat_11460_comb = {4'h0, p3_bit_slice_10995 ? 4'h8 : p4_concat_11453_comb};
  assign p4_Code_size_comb = p4_concat_11460_comb & {8{~p3_eq_10996}};
  assign p4_run_size_str_u8_comb = {p3_run__1_squeezed[3:0], 4'h0} | p4_Code_size_comb;
  assign p4_run__1_squeezed_const_msb_bits__5_comb = 1'h0;
  assign p4_sel_11474_comb = p3_is_luminance ? 3'h4 : 3'h1;
  assign p4_next_pix_squeezed_const_msb_bits_comb = 2'h0;
  assign p4_run__1_squeezed_const_msb_bits__3_comb = 1'h0;
  assign p4_run__1_comb = {p4_run__1_squeezed_const_msb_bits__5_comb, p3_run__1_squeezed};
  assign p4_Huffman_length_squeezed_comb = p3_is_luminance ? literal_11468[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_11466[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_next_pix__1_squeezed_comb = p4_run__1_comb + 6'h01;
  assign p4_Huffman_code_full_comb = p3_is_luminance ? literal_11473[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_11472[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_huff_length_squeezed_const_msb_bits__2_comb = 3'h0;
  assign p4_huff_length_squeezed_comb = p3_and_11412 ? {p4_next_pix_squeezed_const_msb_bits_comb, p3_is_luminance ? 2'h2 : 2'h1, p4_run__1_squeezed_const_msb_bits__3_comb} : p4_Huffman_length_squeezed_comb;
  assign p4_next_pix_squeezed_const_msb_bits__1_comb = 2'h0;
  assign p4_next_pix_squeezed_comb = p3_and_11412 ? 6'h3f : p4_next_pix__1_squeezed_comb;
  assign p4_huff_code_comb = p3_and_11412 ? {12'h000, {{1{p4_sel_11474_comb[2]}}, p4_sel_11474_comb}} : p4_Huffman_code_full_comb;
  assign p4_huff_length_comb = {p4_huff_length_squeezed_const_msb_bits__2_comb, p4_huff_length_squeezed_comb};
  assign p4_code_size_comb = p4_concat_11460_comb & {8{~(p3_and_11412 | p3_eq_10996)}};
  assign p4_next_pix_comb = {p4_next_pix_squeezed_const_msb_bits__1_comb, p4_next_pix_squeezed_comb};
  assign p4_tuple_11503_comb = {p4_huff_code_comb, p4_huff_length_comb, p3_code_list, p4_code_size_comb, p4_next_pix_comb, p3_value};

  // Registers for pipe stage 4:
  reg [57:0] p4_tuple_11503;
  always @ (posedge clk) begin
    p4_tuple_11503 <= p4_tuple_11503_comb;
  end
  assign out = p4_tuple_11503;
endmodule
