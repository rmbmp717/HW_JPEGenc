module Huffman_DCenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire is_luminance,
  output wire [23:0] out
);
  wire [3:0] literal_815[0:12];
  assign literal_815[0] = 4'h2;
  assign literal_815[1] = 4'h2;
  assign literal_815[2] = 4'h3;
  assign literal_815[3] = 4'h3;
  assign literal_815[4] = 4'h4;
  assign literal_815[5] = 4'h4;
  assign literal_815[6] = 4'h4;
  assign literal_815[7] = 4'h5;
  assign literal_815[8] = 4'h6;
  assign literal_815[9] = 4'h7;
  assign literal_815[10] = 4'h8;
  assign literal_815[11] = 4'h9;
  assign literal_815[12] = 4'h0;
  wire [3:0] literal_817[0:12];
  assign literal_817[0] = 4'h3;
  assign literal_817[1] = 4'h3;
  assign literal_817[2] = 4'h3;
  assign literal_817[3] = 4'h3;
  assign literal_817[4] = 4'h3;
  assign literal_817[5] = 4'h3;
  assign literal_817[6] = 4'h3;
  assign literal_817[7] = 4'h4;
  assign literal_817[8] = 4'h5;
  assign literal_817[9] = 4'h6;
  assign literal_817[10] = 4'h7;
  assign literal_817[11] = 4'h8;
  assign literal_817[12] = 4'h0;
  wire [6:0] literal_818[0:12];
  assign literal_818[0] = 7'h60;
  assign literal_818[1] = 7'h50;
  assign literal_818[2] = 7'h30;
  assign literal_818[3] = 7'h20;
  assign literal_818[4] = 7'h00;
  assign literal_818[5] = 7'h10;
  assign literal_818[6] = 7'h40;
  assign literal_818[7] = 7'h70;
  assign literal_818[8] = 7'h78;
  assign literal_818[9] = 7'h7c;
  assign literal_818[10] = 7'h7e;
  assign literal_818[11] = 7'h7f;
  assign literal_818[12] = 7'h00;
  wire [7:0] literal_821[0:12];
  assign literal_821[0] = 8'h02;
  assign literal_821[1] = 8'h00;
  assign literal_821[2] = 8'h20;
  assign literal_821[3] = 8'h28;
  assign literal_821[4] = 8'h60;
  assign literal_821[5] = 8'h68;
  assign literal_821[6] = 8'h70;
  assign literal_821[7] = 8'h78;
  assign literal_821[8] = 8'h7c;
  assign literal_821[9] = 8'h7e;
  assign literal_821[10] = 8'h7f;
  assign literal_821[11] = 8'hfe;
  assign literal_821[12] = 8'h00;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [9:0] p1_dc_comb;
  wire [7:0] p1_bin_value_comb;
  wire [7:0] p1_dc_abs_comb;
  wire [2:0] p1_sel_797_comb;
  wire [3:0] p1_concat_810_comb;
  wire [3:0] p1_size__1_comb;
  wire [2:0] p1_length_squeezed_squeezed_comb;
  wire [7:0] p1_flipped_comb;
  wire [7:0] p1_BoolList_comb;
  wire [7:0] p1_length_comb;
  wire [7:0] p1_code_list_comb;
  wire [23:0] p1_tuple_836_comb;
  assign p1_dc_comb = p0_matrix[3'h0][3'h0];
  assign p1_bin_value_comb = p1_dc_comb[7:0];
  assign p1_dc_abs_comb = p1_dc_comb[9] ? -p1_bin_value_comb : p1_bin_value_comb;
  assign p1_sel_797_comb = |p1_dc_abs_comb[7:3] ? 3'h4 : {1'h0, |p1_dc_abs_comb[7:2] ? 2'h3 : (|p1_dc_abs_comb[7:1] ? 2'h2 : 2'h1)};
  assign p1_concat_810_comb = {1'h0, |p1_dc_abs_comb[7:6] ? 3'h7 : (|p1_dc_abs_comb[7:5] ? 3'h6 : (|p1_dc_abs_comb[7:4] ? 3'h5 : p1_sel_797_comb))};
  assign p1_size__1_comb = (p1_dc_abs_comb[7] ? 4'h8 : p1_concat_810_comb) & {4{p1_dc_abs_comb != 8'h00}};
  assign p1_length_squeezed_squeezed_comb = p0_is_luminance ? literal_817[p1_size__1_comb > 4'hc ? 4'hc : p1_size__1_comb][2:0] : literal_815[p1_size__1_comb > 4'hc ? 4'hc : p1_size__1_comb][2:0];
  assign p1_flipped_comb = ~p1_bin_value_comb;
  assign p1_BoolList_comb = p0_is_luminance ? {literal_818[p1_size__1_comb > 4'hc ? 4'hc : p1_size__1_comb], 1'h0} : literal_821[p1_size__1_comb];
  assign p1_length_comb = {5'h00, p1_length_squeezed_squeezed_comb};
  assign p1_code_list_comb = $signed(p1_dc_comb) <= $signed(10'h000) ? p1_flipped_comb : p1_bin_value_comb;
  assign p1_tuple_836_comb = {p1_BoolList_comb, p1_length_comb, p1_code_list_comb};

  // Registers for pipe stage 1:
  reg [23:0] p1_tuple_836;
  always @ (posedge clk) begin
    p1_tuple_836 <= p1_tuple_836_comb;
  end
  assign out = p1_tuple_836;
endmodule
