module Huffman_ACenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [47:0] out
);
  wire [4:0] literal_10574[0:251];
  assign literal_10574[0] = 5'h02;
  assign literal_10574[1] = 5'h02;
  assign literal_10574[2] = 5'h03;
  assign literal_10574[3] = 5'h04;
  assign literal_10574[4] = 5'h05;
  assign literal_10574[5] = 5'h07;
  assign literal_10574[6] = 5'h08;
  assign literal_10574[7] = 5'h0e;
  assign literal_10574[8] = 5'h10;
  assign literal_10574[9] = 5'h10;
  assign literal_10574[10] = 5'h10;
  assign literal_10574[11] = 5'h00;
  assign literal_10574[12] = 5'h00;
  assign literal_10574[13] = 5'h00;
  assign literal_10574[14] = 5'h00;
  assign literal_10574[15] = 5'h00;
  assign literal_10574[16] = 5'h00;
  assign literal_10574[17] = 5'h03;
  assign literal_10574[18] = 5'h06;
  assign literal_10574[19] = 5'h07;
  assign literal_10574[20] = 5'h09;
  assign literal_10574[21] = 5'h0b;
  assign literal_10574[22] = 5'h0d;
  assign literal_10574[23] = 5'h10;
  assign literal_10574[24] = 5'h10;
  assign literal_10574[25] = 5'h10;
  assign literal_10574[26] = 5'h10;
  assign literal_10574[27] = 5'h00;
  assign literal_10574[28] = 5'h00;
  assign literal_10574[29] = 5'h00;
  assign literal_10574[30] = 5'h00;
  assign literal_10574[31] = 5'h00;
  assign literal_10574[32] = 5'h00;
  assign literal_10574[33] = 5'h05;
  assign literal_10574[34] = 5'h07;
  assign literal_10574[35] = 5'h0a;
  assign literal_10574[36] = 5'h0c;
  assign literal_10574[37] = 5'h0d;
  assign literal_10574[38] = 5'h10;
  assign literal_10574[39] = 5'h10;
  assign literal_10574[40] = 5'h10;
  assign literal_10574[41] = 5'h10;
  assign literal_10574[42] = 5'h10;
  assign literal_10574[43] = 5'h00;
  assign literal_10574[44] = 5'h00;
  assign literal_10574[45] = 5'h00;
  assign literal_10574[46] = 5'h00;
  assign literal_10574[47] = 5'h00;
  assign literal_10574[48] = 5'h00;
  assign literal_10574[49] = 5'h06;
  assign literal_10574[50] = 5'h08;
  assign literal_10574[51] = 5'h0b;
  assign literal_10574[52] = 5'h0c;
  assign literal_10574[53] = 5'h0f;
  assign literal_10574[54] = 5'h10;
  assign literal_10574[55] = 5'h10;
  assign literal_10574[56] = 5'h10;
  assign literal_10574[57] = 5'h10;
  assign literal_10574[58] = 5'h10;
  assign literal_10574[59] = 5'h00;
  assign literal_10574[60] = 5'h00;
  assign literal_10574[61] = 5'h00;
  assign literal_10574[62] = 5'h00;
  assign literal_10574[63] = 5'h00;
  assign literal_10574[64] = 5'h00;
  assign literal_10574[65] = 5'h06;
  assign literal_10574[66] = 5'h0a;
  assign literal_10574[67] = 5'h0c;
  assign literal_10574[68] = 5'h0f;
  assign literal_10574[69] = 5'h10;
  assign literal_10574[70] = 5'h10;
  assign literal_10574[71] = 5'h10;
  assign literal_10574[72] = 5'h10;
  assign literal_10574[73] = 5'h10;
  assign literal_10574[74] = 5'h10;
  assign literal_10574[75] = 5'h00;
  assign literal_10574[76] = 5'h00;
  assign literal_10574[77] = 5'h00;
  assign literal_10574[78] = 5'h00;
  assign literal_10574[79] = 5'h00;
  assign literal_10574[80] = 5'h00;
  assign literal_10574[81] = 5'h07;
  assign literal_10574[82] = 5'h0b;
  assign literal_10574[83] = 5'h0d;
  assign literal_10574[84] = 5'h10;
  assign literal_10574[85] = 5'h10;
  assign literal_10574[86] = 5'h10;
  assign literal_10574[87] = 5'h10;
  assign literal_10574[88] = 5'h10;
  assign literal_10574[89] = 5'h10;
  assign literal_10574[90] = 5'h10;
  assign literal_10574[91] = 5'h00;
  assign literal_10574[92] = 5'h00;
  assign literal_10574[93] = 5'h00;
  assign literal_10574[94] = 5'h00;
  assign literal_10574[95] = 5'h00;
  assign literal_10574[96] = 5'h00;
  assign literal_10574[97] = 5'h07;
  assign literal_10574[98] = 5'h0b;
  assign literal_10574[99] = 5'h0d;
  assign literal_10574[100] = 5'h10;
  assign literal_10574[101] = 5'h10;
  assign literal_10574[102] = 5'h10;
  assign literal_10574[103] = 5'h10;
  assign literal_10574[104] = 5'h10;
  assign literal_10574[105] = 5'h10;
  assign literal_10574[106] = 5'h10;
  assign literal_10574[107] = 5'h00;
  assign literal_10574[108] = 5'h00;
  assign literal_10574[109] = 5'h00;
  assign literal_10574[110] = 5'h00;
  assign literal_10574[111] = 5'h00;
  assign literal_10574[112] = 5'h00;
  assign literal_10574[113] = 5'h08;
  assign literal_10574[114] = 5'h0b;
  assign literal_10574[115] = 5'h0e;
  assign literal_10574[116] = 5'h10;
  assign literal_10574[117] = 5'h10;
  assign literal_10574[118] = 5'h10;
  assign literal_10574[119] = 5'h10;
  assign literal_10574[120] = 5'h10;
  assign literal_10574[121] = 5'h10;
  assign literal_10574[122] = 5'h10;
  assign literal_10574[123] = 5'h00;
  assign literal_10574[124] = 5'h00;
  assign literal_10574[125] = 5'h00;
  assign literal_10574[126] = 5'h00;
  assign literal_10574[127] = 5'h00;
  assign literal_10574[128] = 5'h00;
  assign literal_10574[129] = 5'h08;
  assign literal_10574[130] = 5'h0c;
  assign literal_10574[131] = 5'h10;
  assign literal_10574[132] = 5'h10;
  assign literal_10574[133] = 5'h10;
  assign literal_10574[134] = 5'h10;
  assign literal_10574[135] = 5'h10;
  assign literal_10574[136] = 5'h10;
  assign literal_10574[137] = 5'h10;
  assign literal_10574[138] = 5'h10;
  assign literal_10574[139] = 5'h00;
  assign literal_10574[140] = 5'h00;
  assign literal_10574[141] = 5'h00;
  assign literal_10574[142] = 5'h00;
  assign literal_10574[143] = 5'h00;
  assign literal_10574[144] = 5'h00;
  assign literal_10574[145] = 5'h08;
  assign literal_10574[146] = 5'h0d;
  assign literal_10574[147] = 5'h10;
  assign literal_10574[148] = 5'h10;
  assign literal_10574[149] = 5'h10;
  assign literal_10574[150] = 5'h10;
  assign literal_10574[151] = 5'h10;
  assign literal_10574[152] = 5'h10;
  assign literal_10574[153] = 5'h10;
  assign literal_10574[154] = 5'h10;
  assign literal_10574[155] = 5'h00;
  assign literal_10574[156] = 5'h00;
  assign literal_10574[157] = 5'h00;
  assign literal_10574[158] = 5'h00;
  assign literal_10574[159] = 5'h00;
  assign literal_10574[160] = 5'h00;
  assign literal_10574[161] = 5'h09;
  assign literal_10574[162] = 5'h0d;
  assign literal_10574[163] = 5'h10;
  assign literal_10574[164] = 5'h10;
  assign literal_10574[165] = 5'h10;
  assign literal_10574[166] = 5'h10;
  assign literal_10574[167] = 5'h10;
  assign literal_10574[168] = 5'h10;
  assign literal_10574[169] = 5'h10;
  assign literal_10574[170] = 5'h10;
  assign literal_10574[171] = 5'h00;
  assign literal_10574[172] = 5'h00;
  assign literal_10574[173] = 5'h00;
  assign literal_10574[174] = 5'h00;
  assign literal_10574[175] = 5'h00;
  assign literal_10574[176] = 5'h00;
  assign literal_10574[177] = 5'h09;
  assign literal_10574[178] = 5'h0d;
  assign literal_10574[179] = 5'h10;
  assign literal_10574[180] = 5'h10;
  assign literal_10574[181] = 5'h10;
  assign literal_10574[182] = 5'h10;
  assign literal_10574[183] = 5'h10;
  assign literal_10574[184] = 5'h10;
  assign literal_10574[185] = 5'h10;
  assign literal_10574[186] = 5'h10;
  assign literal_10574[187] = 5'h00;
  assign literal_10574[188] = 5'h00;
  assign literal_10574[189] = 5'h00;
  assign literal_10574[190] = 5'h00;
  assign literal_10574[191] = 5'h00;
  assign literal_10574[192] = 5'h00;
  assign literal_10574[193] = 5'h0a;
  assign literal_10574[194] = 5'h0d;
  assign literal_10574[195] = 5'h10;
  assign literal_10574[196] = 5'h10;
  assign literal_10574[197] = 5'h10;
  assign literal_10574[198] = 5'h10;
  assign literal_10574[199] = 5'h10;
  assign literal_10574[200] = 5'h10;
  assign literal_10574[201] = 5'h10;
  assign literal_10574[202] = 5'h10;
  assign literal_10574[203] = 5'h00;
  assign literal_10574[204] = 5'h00;
  assign literal_10574[205] = 5'h00;
  assign literal_10574[206] = 5'h00;
  assign literal_10574[207] = 5'h00;
  assign literal_10574[208] = 5'h00;
  assign literal_10574[209] = 5'h0a;
  assign literal_10574[210] = 5'h0e;
  assign literal_10574[211] = 5'h10;
  assign literal_10574[212] = 5'h10;
  assign literal_10574[213] = 5'h10;
  assign literal_10574[214] = 5'h10;
  assign literal_10574[215] = 5'h10;
  assign literal_10574[216] = 5'h10;
  assign literal_10574[217] = 5'h10;
  assign literal_10574[218] = 5'h10;
  assign literal_10574[219] = 5'h00;
  assign literal_10574[220] = 5'h00;
  assign literal_10574[221] = 5'h00;
  assign literal_10574[222] = 5'h00;
  assign literal_10574[223] = 5'h00;
  assign literal_10574[224] = 5'h00;
  assign literal_10574[225] = 5'h0a;
  assign literal_10574[226] = 5'h0f;
  assign literal_10574[227] = 5'h10;
  assign literal_10574[228] = 5'h10;
  assign literal_10574[229] = 5'h10;
  assign literal_10574[230] = 5'h10;
  assign literal_10574[231] = 5'h10;
  assign literal_10574[232] = 5'h10;
  assign literal_10574[233] = 5'h10;
  assign literal_10574[234] = 5'h10;
  assign literal_10574[235] = 5'h00;
  assign literal_10574[236] = 5'h00;
  assign literal_10574[237] = 5'h00;
  assign literal_10574[238] = 5'h00;
  assign literal_10574[239] = 5'h00;
  assign literal_10574[240] = 5'h09;
  assign literal_10574[241] = 5'h0b;
  assign literal_10574[242] = 5'h10;
  assign literal_10574[243] = 5'h10;
  assign literal_10574[244] = 5'h10;
  assign literal_10574[245] = 5'h10;
  assign literal_10574[246] = 5'h10;
  assign literal_10574[247] = 5'h10;
  assign literal_10574[248] = 5'h10;
  assign literal_10574[249] = 5'h10;
  assign literal_10574[250] = 5'h10;
  assign literal_10574[251] = 5'h00;
  wire [4:0] literal_10576[0:251];
  assign literal_10576[0] = 5'h04;
  assign literal_10576[1] = 5'h02;
  assign literal_10576[2] = 5'h02;
  assign literal_10576[3] = 5'h03;
  assign literal_10576[4] = 5'h04;
  assign literal_10576[5] = 5'h05;
  assign literal_10576[6] = 5'h07;
  assign literal_10576[7] = 5'h09;
  assign literal_10576[8] = 5'h10;
  assign literal_10576[9] = 5'h10;
  assign literal_10576[10] = 5'h10;
  assign literal_10576[11] = 5'h00;
  assign literal_10576[12] = 5'h00;
  assign literal_10576[13] = 5'h00;
  assign literal_10576[14] = 5'h00;
  assign literal_10576[15] = 5'h00;
  assign literal_10576[16] = 5'h00;
  assign literal_10576[17] = 5'h04;
  assign literal_10576[18] = 5'h05;
  assign literal_10576[19] = 5'h07;
  assign literal_10576[20] = 5'h09;
  assign literal_10576[21] = 5'h0a;
  assign literal_10576[22] = 5'h0b;
  assign literal_10576[23] = 5'h10;
  assign literal_10576[24] = 5'h10;
  assign literal_10576[25] = 5'h10;
  assign literal_10576[26] = 5'h10;
  assign literal_10576[27] = 5'h00;
  assign literal_10576[28] = 5'h00;
  assign literal_10576[29] = 5'h00;
  assign literal_10576[30] = 5'h00;
  assign literal_10576[31] = 5'h00;
  assign literal_10576[32] = 5'h00;
  assign literal_10576[33] = 5'h05;
  assign literal_10576[34] = 5'h08;
  assign literal_10576[35] = 5'h0a;
  assign literal_10576[36] = 5'h0c;
  assign literal_10576[37] = 5'h0e;
  assign literal_10576[38] = 5'h10;
  assign literal_10576[39] = 5'h10;
  assign literal_10576[40] = 5'h10;
  assign literal_10576[41] = 5'h10;
  assign literal_10576[42] = 5'h10;
  assign literal_10576[43] = 5'h00;
  assign literal_10576[44] = 5'h00;
  assign literal_10576[45] = 5'h00;
  assign literal_10576[46] = 5'h00;
  assign literal_10576[47] = 5'h00;
  assign literal_10576[48] = 5'h00;
  assign literal_10576[49] = 5'h06;
  assign literal_10576[50] = 5'h09;
  assign literal_10576[51] = 5'h0b;
  assign literal_10576[52] = 5'h0e;
  assign literal_10576[53] = 5'h10;
  assign literal_10576[54] = 5'h10;
  assign literal_10576[55] = 5'h10;
  assign literal_10576[56] = 5'h10;
  assign literal_10576[57] = 5'h10;
  assign literal_10576[58] = 5'h10;
  assign literal_10576[59] = 5'h00;
  assign literal_10576[60] = 5'h00;
  assign literal_10576[61] = 5'h00;
  assign literal_10576[62] = 5'h00;
  assign literal_10576[63] = 5'h00;
  assign literal_10576[64] = 5'h00;
  assign literal_10576[65] = 5'h06;
  assign literal_10576[66] = 5'h0a;
  assign literal_10576[67] = 5'h0e;
  assign literal_10576[68] = 5'h10;
  assign literal_10576[69] = 5'h10;
  assign literal_10576[70] = 5'h10;
  assign literal_10576[71] = 5'h10;
  assign literal_10576[72] = 5'h10;
  assign literal_10576[73] = 5'h10;
  assign literal_10576[74] = 5'h10;
  assign literal_10576[75] = 5'h00;
  assign literal_10576[76] = 5'h00;
  assign literal_10576[77] = 5'h00;
  assign literal_10576[78] = 5'h00;
  assign literal_10576[79] = 5'h00;
  assign literal_10576[80] = 5'h00;
  assign literal_10576[81] = 5'h07;
  assign literal_10576[82] = 5'h0a;
  assign literal_10576[83] = 5'h0e;
  assign literal_10576[84] = 5'h10;
  assign literal_10576[85] = 5'h10;
  assign literal_10576[86] = 5'h10;
  assign literal_10576[87] = 5'h10;
  assign literal_10576[88] = 5'h10;
  assign literal_10576[89] = 5'h10;
  assign literal_10576[90] = 5'h10;
  assign literal_10576[91] = 5'h00;
  assign literal_10576[92] = 5'h00;
  assign literal_10576[93] = 5'h00;
  assign literal_10576[94] = 5'h00;
  assign literal_10576[95] = 5'h00;
  assign literal_10576[96] = 5'h00;
  assign literal_10576[97] = 5'h07;
  assign literal_10576[98] = 5'h0c;
  assign literal_10576[99] = 5'h0f;
  assign literal_10576[100] = 5'h10;
  assign literal_10576[101] = 5'h10;
  assign literal_10576[102] = 5'h10;
  assign literal_10576[103] = 5'h10;
  assign literal_10576[104] = 5'h10;
  assign literal_10576[105] = 5'h10;
  assign literal_10576[106] = 5'h10;
  assign literal_10576[107] = 5'h00;
  assign literal_10576[108] = 5'h00;
  assign literal_10576[109] = 5'h00;
  assign literal_10576[110] = 5'h00;
  assign literal_10576[111] = 5'h00;
  assign literal_10576[112] = 5'h00;
  assign literal_10576[113] = 5'h08;
  assign literal_10576[114] = 5'h0c;
  assign literal_10576[115] = 5'h10;
  assign literal_10576[116] = 5'h10;
  assign literal_10576[117] = 5'h10;
  assign literal_10576[118] = 5'h10;
  assign literal_10576[119] = 5'h10;
  assign literal_10576[120] = 5'h10;
  assign literal_10576[121] = 5'h10;
  assign literal_10576[122] = 5'h10;
  assign literal_10576[123] = 5'h00;
  assign literal_10576[124] = 5'h00;
  assign literal_10576[125] = 5'h00;
  assign literal_10576[126] = 5'h00;
  assign literal_10576[127] = 5'h00;
  assign literal_10576[128] = 5'h00;
  assign literal_10576[129] = 5'h09;
  assign literal_10576[130] = 5'h0d;
  assign literal_10576[131] = 5'h10;
  assign literal_10576[132] = 5'h10;
  assign literal_10576[133] = 5'h10;
  assign literal_10576[134] = 5'h10;
  assign literal_10576[135] = 5'h10;
  assign literal_10576[136] = 5'h10;
  assign literal_10576[137] = 5'h10;
  assign literal_10576[138] = 5'h10;
  assign literal_10576[139] = 5'h00;
  assign literal_10576[140] = 5'h00;
  assign literal_10576[141] = 5'h00;
  assign literal_10576[142] = 5'h00;
  assign literal_10576[143] = 5'h00;
  assign literal_10576[144] = 5'h00;
  assign literal_10576[145] = 5'h09;
  assign literal_10576[146] = 5'h0e;
  assign literal_10576[147] = 5'h10;
  assign literal_10576[148] = 5'h10;
  assign literal_10576[149] = 5'h10;
  assign literal_10576[150] = 5'h10;
  assign literal_10576[151] = 5'h10;
  assign literal_10576[152] = 5'h10;
  assign literal_10576[153] = 5'h10;
  assign literal_10576[154] = 5'h10;
  assign literal_10576[155] = 5'h00;
  assign literal_10576[156] = 5'h00;
  assign literal_10576[157] = 5'h00;
  assign literal_10576[158] = 5'h00;
  assign literal_10576[159] = 5'h00;
  assign literal_10576[160] = 5'h00;
  assign literal_10576[161] = 5'h09;
  assign literal_10576[162] = 5'h0e;
  assign literal_10576[163] = 5'h10;
  assign literal_10576[164] = 5'h10;
  assign literal_10576[165] = 5'h10;
  assign literal_10576[166] = 5'h10;
  assign literal_10576[167] = 5'h10;
  assign literal_10576[168] = 5'h10;
  assign literal_10576[169] = 5'h10;
  assign literal_10576[170] = 5'h10;
  assign literal_10576[171] = 5'h00;
  assign literal_10576[172] = 5'h00;
  assign literal_10576[173] = 5'h00;
  assign literal_10576[174] = 5'h00;
  assign literal_10576[175] = 5'h00;
  assign literal_10576[176] = 5'h00;
  assign literal_10576[177] = 5'h0a;
  assign literal_10576[178] = 5'h0f;
  assign literal_10576[179] = 5'h10;
  assign literal_10576[180] = 5'h10;
  assign literal_10576[181] = 5'h10;
  assign literal_10576[182] = 5'h10;
  assign literal_10576[183] = 5'h10;
  assign literal_10576[184] = 5'h10;
  assign literal_10576[185] = 5'h10;
  assign literal_10576[186] = 5'h10;
  assign literal_10576[187] = 5'h00;
  assign literal_10576[188] = 5'h00;
  assign literal_10576[189] = 5'h00;
  assign literal_10576[190] = 5'h00;
  assign literal_10576[191] = 5'h00;
  assign literal_10576[192] = 5'h00;
  assign literal_10576[193] = 5'h0a;
  assign literal_10576[194] = 5'h10;
  assign literal_10576[195] = 5'h10;
  assign literal_10576[196] = 5'h10;
  assign literal_10576[197] = 5'h10;
  assign literal_10576[198] = 5'h10;
  assign literal_10576[199] = 5'h10;
  assign literal_10576[200] = 5'h10;
  assign literal_10576[201] = 5'h10;
  assign literal_10576[202] = 5'h10;
  assign literal_10576[203] = 5'h00;
  assign literal_10576[204] = 5'h00;
  assign literal_10576[205] = 5'h00;
  assign literal_10576[206] = 5'h00;
  assign literal_10576[207] = 5'h00;
  assign literal_10576[208] = 5'h00;
  assign literal_10576[209] = 5'h0a;
  assign literal_10576[210] = 5'h10;
  assign literal_10576[211] = 5'h10;
  assign literal_10576[212] = 5'h10;
  assign literal_10576[213] = 5'h10;
  assign literal_10576[214] = 5'h10;
  assign literal_10576[215] = 5'h10;
  assign literal_10576[216] = 5'h10;
  assign literal_10576[217] = 5'h10;
  assign literal_10576[218] = 5'h10;
  assign literal_10576[219] = 5'h00;
  assign literal_10576[220] = 5'h00;
  assign literal_10576[221] = 5'h00;
  assign literal_10576[222] = 5'h00;
  assign literal_10576[223] = 5'h00;
  assign literal_10576[224] = 5'h00;
  assign literal_10576[225] = 5'h0b;
  assign literal_10576[226] = 5'h10;
  assign literal_10576[227] = 5'h10;
  assign literal_10576[228] = 5'h10;
  assign literal_10576[229] = 5'h10;
  assign literal_10576[230] = 5'h10;
  assign literal_10576[231] = 5'h10;
  assign literal_10576[232] = 5'h10;
  assign literal_10576[233] = 5'h10;
  assign literal_10576[234] = 5'h10;
  assign literal_10576[235] = 5'h00;
  assign literal_10576[236] = 5'h00;
  assign literal_10576[237] = 5'h00;
  assign literal_10576[238] = 5'h00;
  assign literal_10576[239] = 5'h00;
  assign literal_10576[240] = 5'h0c;
  assign literal_10576[241] = 5'h0d;
  assign literal_10576[242] = 5'h10;
  assign literal_10576[243] = 5'h10;
  assign literal_10576[244] = 5'h10;
  assign literal_10576[245] = 5'h10;
  assign literal_10576[246] = 5'h10;
  assign literal_10576[247] = 5'h10;
  assign literal_10576[248] = 5'h10;
  assign literal_10576[249] = 5'h10;
  assign literal_10576[250] = 5'h10;
  assign literal_10576[251] = 5'h00;
  wire [15:0] literal_10580[0:251];
  assign literal_10580[0] = 16'h0001;
  assign literal_10580[1] = 16'h0000;
  assign literal_10580[2] = 16'h0004;
  assign literal_10580[3] = 16'h000c;
  assign literal_10580[4] = 16'h001a;
  assign literal_10580[5] = 16'h0076;
  assign literal_10580[6] = 16'h00f6;
  assign literal_10580[7] = 16'h3fe0;
  assign literal_10580[8] = 16'hff96;
  assign literal_10580[9] = 16'hff97;
  assign literal_10580[10] = 16'hff98;
  assign literal_10580[11] = 16'h0000;
  assign literal_10580[12] = 16'h0000;
  assign literal_10580[13] = 16'h0000;
  assign literal_10580[14] = 16'h0000;
  assign literal_10580[15] = 16'h0000;
  assign literal_10580[16] = 16'h0000;
  assign literal_10580[17] = 16'h0005;
  assign literal_10580[18] = 16'h0038;
  assign literal_10580[19] = 16'h0078;
  assign literal_10580[20] = 16'h01f9;
  assign literal_10580[21] = 16'h07f2;
  assign literal_10580[22] = 16'h1fe8;
  assign literal_10580[23] = 16'hff93;
  assign literal_10580[24] = 16'hff99;
  assign literal_10580[25] = 16'hff9a;
  assign literal_10580[26] = 16'hff9e;
  assign literal_10580[27] = 16'h0000;
  assign literal_10580[28] = 16'h0000;
  assign literal_10580[29] = 16'h0000;
  assign literal_10580[30] = 16'h0000;
  assign literal_10580[31] = 16'h0000;
  assign literal_10580[32] = 16'h0000;
  assign literal_10580[33] = 16'h001b;
  assign literal_10580[34] = 16'h007a;
  assign literal_10580[35] = 16'h03f7;
  assign literal_10580[36] = 16'h0ff0;
  assign literal_10580[37] = 16'h1feb;
  assign literal_10580[38] = 16'hff9b;
  assign literal_10580[39] = 16'hff9f;
  assign literal_10580[40] = 16'hffa8;
  assign literal_10580[41] = 16'hffa9;
  assign literal_10580[42] = 16'hfff1;
  assign literal_10580[43] = 16'h0000;
  assign literal_10580[44] = 16'h0000;
  assign literal_10580[45] = 16'h0000;
  assign literal_10580[46] = 16'h0000;
  assign literal_10580[47] = 16'h0000;
  assign literal_10580[48] = 16'h0000;
  assign literal_10580[49] = 16'h0039;
  assign literal_10580[50] = 16'h00fa;
  assign literal_10580[51] = 16'h07f7;
  assign literal_10580[52] = 16'h0ff1;
  assign literal_10580[53] = 16'h7fc6;
  assign literal_10580[54] = 16'hff9c;
  assign literal_10580[55] = 16'hffa3;
  assign literal_10580[56] = 16'hffd7;
  assign literal_10580[57] = 16'hffe4;
  assign literal_10580[58] = 16'hfff2;
  assign literal_10580[59] = 16'h0000;
  assign literal_10580[60] = 16'h0000;
  assign literal_10580[61] = 16'h0000;
  assign literal_10580[62] = 16'h0000;
  assign literal_10580[63] = 16'h0000;
  assign literal_10580[64] = 16'h0000;
  assign literal_10580[65] = 16'h003a;
  assign literal_10580[66] = 16'h03f8;
  assign literal_10580[67] = 16'h0ff2;
  assign literal_10580[68] = 16'h7fc8;
  assign literal_10580[69] = 16'hff9d;
  assign literal_10580[70] = 16'hffbf;
  assign literal_10580[71] = 16'hffcb;
  assign literal_10580[72] = 16'hffd8;
  assign literal_10580[73] = 16'hffe5;
  assign literal_10580[74] = 16'hfff3;
  assign literal_10580[75] = 16'h0000;
  assign literal_10580[76] = 16'h0000;
  assign literal_10580[77] = 16'h0000;
  assign literal_10580[78] = 16'h0000;
  assign literal_10580[79] = 16'h0000;
  assign literal_10580[80] = 16'h0000;
  assign literal_10580[81] = 16'h0077;
  assign literal_10580[82] = 16'h07f3;
  assign literal_10580[83] = 16'h1fea;
  assign literal_10580[84] = 16'hff94;
  assign literal_10580[85] = 16'hffa2;
  assign literal_10580[86] = 16'hffc0;
  assign literal_10580[87] = 16'hffcc;
  assign literal_10580[88] = 16'hffd9;
  assign literal_10580[89] = 16'hffe6;
  assign literal_10580[90] = 16'hfff4;
  assign literal_10580[91] = 16'h0000;
  assign literal_10580[92] = 16'h0000;
  assign literal_10580[93] = 16'h0000;
  assign literal_10580[94] = 16'h0000;
  assign literal_10580[95] = 16'h0000;
  assign literal_10580[96] = 16'h0000;
  assign literal_10580[97] = 16'h0079;
  assign literal_10580[98] = 16'h07f4;
  assign literal_10580[99] = 16'h1fed;
  assign literal_10580[100] = 16'hffa0;
  assign literal_10580[101] = 16'hffb5;
  assign literal_10580[102] = 16'hffc1;
  assign literal_10580[103] = 16'hffcd;
  assign literal_10580[104] = 16'hffda;
  assign literal_10580[105] = 16'hffe7;
  assign literal_10580[106] = 16'hfff5;
  assign literal_10580[107] = 16'h0000;
  assign literal_10580[108] = 16'h0000;
  assign literal_10580[109] = 16'h0000;
  assign literal_10580[110] = 16'h0000;
  assign literal_10580[111] = 16'h0000;
  assign literal_10580[112] = 16'h0000;
  assign literal_10580[113] = 16'h00f7;
  assign literal_10580[114] = 16'h07f5;
  assign literal_10580[115] = 16'h3fe1;
  assign literal_10580[116] = 16'hffa1;
  assign literal_10580[117] = 16'hffb6;
  assign literal_10580[118] = 16'hffc2;
  assign literal_10580[119] = 16'hffce;
  assign literal_10580[120] = 16'hffdb;
  assign literal_10580[121] = 16'hffe8;
  assign literal_10580[122] = 16'hfff6;
  assign literal_10580[123] = 16'h0000;
  assign literal_10580[124] = 16'h0000;
  assign literal_10580[125] = 16'h0000;
  assign literal_10580[126] = 16'h0000;
  assign literal_10580[127] = 16'h0000;
  assign literal_10580[128] = 16'h0000;
  assign literal_10580[129] = 16'h00f8;
  assign literal_10580[130] = 16'h0ff3;
  assign literal_10580[131] = 16'hff92;
  assign literal_10580[132] = 16'hffad;
  assign literal_10580[133] = 16'hffb7;
  assign literal_10580[134] = 16'hffc3;
  assign literal_10580[135] = 16'hffcf;
  assign literal_10580[136] = 16'hffdc;
  assign literal_10580[137] = 16'hffe9;
  assign literal_10580[138] = 16'hfff7;
  assign literal_10580[139] = 16'h0000;
  assign literal_10580[140] = 16'h0000;
  assign literal_10580[141] = 16'h0000;
  assign literal_10580[142] = 16'h0000;
  assign literal_10580[143] = 16'h0000;
  assign literal_10580[144] = 16'h0000;
  assign literal_10580[145] = 16'h00f9;
  assign literal_10580[146] = 16'h1fe9;
  assign literal_10580[147] = 16'hff95;
  assign literal_10580[148] = 16'hffae;
  assign literal_10580[149] = 16'hffb8;
  assign literal_10580[150] = 16'hffc4;
  assign literal_10580[151] = 16'hffd0;
  assign literal_10580[152] = 16'hffdd;
  assign literal_10580[153] = 16'hffea;
  assign literal_10580[154] = 16'hfff8;
  assign literal_10580[155] = 16'h0000;
  assign literal_10580[156] = 16'h0000;
  assign literal_10580[157] = 16'h0000;
  assign literal_10580[158] = 16'h0000;
  assign literal_10580[159] = 16'h0000;
  assign literal_10580[160] = 16'h0000;
  assign literal_10580[161] = 16'h01f6;
  assign literal_10580[162] = 16'h1fec;
  assign literal_10580[163] = 16'hffa5;
  assign literal_10580[164] = 16'hffaf;
  assign literal_10580[165] = 16'hffb9;
  assign literal_10580[166] = 16'hffc5;
  assign literal_10580[167] = 16'hffd1;
  assign literal_10580[168] = 16'hffde;
  assign literal_10580[169] = 16'hffeb;
  assign literal_10580[170] = 16'hfff9;
  assign literal_10580[171] = 16'h0000;
  assign literal_10580[172] = 16'h0000;
  assign literal_10580[173] = 16'h0000;
  assign literal_10580[174] = 16'h0000;
  assign literal_10580[175] = 16'h0000;
  assign literal_10580[176] = 16'h0000;
  assign literal_10580[177] = 16'h01f7;
  assign literal_10580[178] = 16'h1fee;
  assign literal_10580[179] = 16'hffa6;
  assign literal_10580[180] = 16'hffb0;
  assign literal_10580[181] = 16'hffba;
  assign literal_10580[182] = 16'hffc6;
  assign literal_10580[183] = 16'hffd2;
  assign literal_10580[184] = 16'hffdf;
  assign literal_10580[185] = 16'hffec;
  assign literal_10580[186] = 16'hfffa;
  assign literal_10580[187] = 16'h0000;
  assign literal_10580[188] = 16'h0000;
  assign literal_10580[189] = 16'h0000;
  assign literal_10580[190] = 16'h0000;
  assign literal_10580[191] = 16'h0000;
  assign literal_10580[192] = 16'h0000;
  assign literal_10580[193] = 16'h03f4;
  assign literal_10580[194] = 16'h1fef;
  assign literal_10580[195] = 16'hffa7;
  assign literal_10580[196] = 16'hffb1;
  assign literal_10580[197] = 16'hffbb;
  assign literal_10580[198] = 16'hffc7;
  assign literal_10580[199] = 16'hffd3;
  assign literal_10580[200] = 16'hffe0;
  assign literal_10580[201] = 16'hffed;
  assign literal_10580[202] = 16'hfffb;
  assign literal_10580[203] = 16'h0000;
  assign literal_10580[204] = 16'h0000;
  assign literal_10580[205] = 16'h0000;
  assign literal_10580[206] = 16'h0000;
  assign literal_10580[207] = 16'h0000;
  assign literal_10580[208] = 16'h0000;
  assign literal_10580[209] = 16'h03f5;
  assign literal_10580[210] = 16'h3fe2;
  assign literal_10580[211] = 16'hffaa;
  assign literal_10580[212] = 16'hffb2;
  assign literal_10580[213] = 16'hffbc;
  assign literal_10580[214] = 16'hffc8;
  assign literal_10580[215] = 16'hffd4;
  assign literal_10580[216] = 16'hffe1;
  assign literal_10580[217] = 16'hffee;
  assign literal_10580[218] = 16'hfffc;
  assign literal_10580[219] = 16'h0000;
  assign literal_10580[220] = 16'h0000;
  assign literal_10580[221] = 16'h0000;
  assign literal_10580[222] = 16'h0000;
  assign literal_10580[223] = 16'h0000;
  assign literal_10580[224] = 16'h0000;
  assign literal_10580[225] = 16'h03f6;
  assign literal_10580[226] = 16'h7fc7;
  assign literal_10580[227] = 16'hffab;
  assign literal_10580[228] = 16'hffb3;
  assign literal_10580[229] = 16'hffbd;
  assign literal_10580[230] = 16'hffc9;
  assign literal_10580[231] = 16'hffd5;
  assign literal_10580[232] = 16'hffe2;
  assign literal_10580[233] = 16'hffef;
  assign literal_10580[234] = 16'hfffd;
  assign literal_10580[235] = 16'h0000;
  assign literal_10580[236] = 16'h0000;
  assign literal_10580[237] = 16'h0000;
  assign literal_10580[238] = 16'h0000;
  assign literal_10580[239] = 16'h0000;
  assign literal_10580[240] = 16'h01f8;
  assign literal_10580[241] = 16'h07f6;
  assign literal_10580[242] = 16'hffa4;
  assign literal_10580[243] = 16'hffac;
  assign literal_10580[244] = 16'hffb4;
  assign literal_10580[245] = 16'hffbe;
  assign literal_10580[246] = 16'hffca;
  assign literal_10580[247] = 16'hffd6;
  assign literal_10580[248] = 16'hffe3;
  assign literal_10580[249] = 16'hfff0;
  assign literal_10580[250] = 16'hfffe;
  assign literal_10580[251] = 16'h0000;
  wire [15:0] literal_10581[0:251];
  assign literal_10581[0] = 16'h000c;
  assign literal_10581[1] = 16'h0000;
  assign literal_10581[2] = 16'h0001;
  assign literal_10581[3] = 16'h0004;
  assign literal_10581[4] = 16'h000b;
  assign literal_10581[5] = 16'h001a;
  assign literal_10581[6] = 16'h0079;
  assign literal_10581[7] = 16'h01f9;
  assign literal_10581[8] = 16'hff9c;
  assign literal_10581[9] = 16'hff9f;
  assign literal_10581[10] = 16'hffa0;
  assign literal_10581[11] = 16'h0000;
  assign literal_10581[12] = 16'h0000;
  assign literal_10581[13] = 16'h0000;
  assign literal_10581[14] = 16'h0000;
  assign literal_10581[15] = 16'h0000;
  assign literal_10581[16] = 16'h0000;
  assign literal_10581[17] = 16'h000a;
  assign literal_10581[18] = 16'h001c;
  assign literal_10581[19] = 16'h007a;
  assign literal_10581[20] = 16'h01f5;
  assign literal_10581[21] = 16'h03f4;
  assign literal_10581[22] = 16'h07f8;
  assign literal_10581[23] = 16'hff95;
  assign literal_10581[24] = 16'hffa1;
  assign literal_10581[25] = 16'hffa2;
  assign literal_10581[26] = 16'hffad;
  assign literal_10581[27] = 16'h0000;
  assign literal_10581[28] = 16'h0000;
  assign literal_10581[29] = 16'h0000;
  assign literal_10581[30] = 16'h0000;
  assign literal_10581[31] = 16'h0000;
  assign literal_10581[32] = 16'h0000;
  assign literal_10581[33] = 16'h001b;
  assign literal_10581[34] = 16'h00f8;
  assign literal_10581[35] = 16'h03f7;
  assign literal_10581[36] = 16'h0ff4;
  assign literal_10581[37] = 16'h3fdc;
  assign literal_10581[38] = 16'hff9d;
  assign literal_10581[39] = 16'hff90;
  assign literal_10581[40] = 16'hffac;
  assign literal_10581[41] = 16'hffe3;
  assign literal_10581[42] = 16'hfff1;
  assign literal_10581[43] = 16'h0000;
  assign literal_10581[44] = 16'h0000;
  assign literal_10581[45] = 16'h0000;
  assign literal_10581[46] = 16'h0000;
  assign literal_10581[47] = 16'h0000;
  assign literal_10581[48] = 16'h0000;
  assign literal_10581[49] = 16'h003a;
  assign literal_10581[50] = 16'h01f6;
  assign literal_10581[51] = 16'h07f7;
  assign literal_10581[52] = 16'h3fde;
  assign literal_10581[53] = 16'hff8e;
  assign literal_10581[54] = 16'hff94;
  assign literal_10581[55] = 16'hffc9;
  assign literal_10581[56] = 16'hffd6;
  assign literal_10581[57] = 16'hffe4;
  assign literal_10581[58] = 16'hfff2;
  assign literal_10581[59] = 16'h0000;
  assign literal_10581[60] = 16'h0000;
  assign literal_10581[61] = 16'h0000;
  assign literal_10581[62] = 16'h0000;
  assign literal_10581[63] = 16'h0000;
  assign literal_10581[64] = 16'h0000;
  assign literal_10581[65] = 16'h003b;
  assign literal_10581[66] = 16'h03f6;
  assign literal_10581[67] = 16'h3fdd;
  assign literal_10581[68] = 16'hff8f;
  assign literal_10581[69] = 16'hffa5;
  assign literal_10581[70] = 16'hffa6;
  assign literal_10581[71] = 16'hffca;
  assign literal_10581[72] = 16'hffd7;
  assign literal_10581[73] = 16'hffe5;
  assign literal_10581[74] = 16'hfff3;
  assign literal_10581[75] = 16'h0000;
  assign literal_10581[76] = 16'h0000;
  assign literal_10581[77] = 16'h0000;
  assign literal_10581[78] = 16'h0000;
  assign literal_10581[79] = 16'h0000;
  assign literal_10581[80] = 16'h0000;
  assign literal_10581[81] = 16'h0078;
  assign literal_10581[82] = 16'h03f9;
  assign literal_10581[83] = 16'h3fdf;
  assign literal_10581[84] = 16'hff96;
  assign literal_10581[85] = 16'hffab;
  assign literal_10581[86] = 16'hffa9;
  assign literal_10581[87] = 16'hffcb;
  assign literal_10581[88] = 16'hffd8;
  assign literal_10581[89] = 16'hffe6;
  assign literal_10581[90] = 16'hfff4;
  assign literal_10581[91] = 16'h0000;
  assign literal_10581[92] = 16'h0000;
  assign literal_10581[93] = 16'h0000;
  assign literal_10581[94] = 16'h0000;
  assign literal_10581[95] = 16'h0000;
  assign literal_10581[96] = 16'h0000;
  assign literal_10581[97] = 16'h007b;
  assign literal_10581[98] = 16'h0ff2;
  assign literal_10581[99] = 16'h7fc5;
  assign literal_10581[100] = 16'hff97;
  assign literal_10581[101] = 16'hffb5;
  assign literal_10581[102] = 16'hffbf;
  assign literal_10581[103] = 16'hffcc;
  assign literal_10581[104] = 16'hffd9;
  assign literal_10581[105] = 16'hffe7;
  assign literal_10581[106] = 16'hfff5;
  assign literal_10581[107] = 16'h0000;
  assign literal_10581[108] = 16'h0000;
  assign literal_10581[109] = 16'h0000;
  assign literal_10581[110] = 16'h0000;
  assign literal_10581[111] = 16'h0000;
  assign literal_10581[112] = 16'h0000;
  assign literal_10581[113] = 16'h00f9;
  assign literal_10581[114] = 16'h0ff5;
  assign literal_10581[115] = 16'hff8c;
  assign literal_10581[116] = 16'hff98;
  assign literal_10581[117] = 16'hffb6;
  assign literal_10581[118] = 16'hffc0;
  assign literal_10581[119] = 16'hffcd;
  assign literal_10581[120] = 16'hffda;
  assign literal_10581[121] = 16'hffe8;
  assign literal_10581[122] = 16'hfff6;
  assign literal_10581[123] = 16'h0000;
  assign literal_10581[124] = 16'h0000;
  assign literal_10581[125] = 16'h0000;
  assign literal_10581[126] = 16'h0000;
  assign literal_10581[127] = 16'h0000;
  assign literal_10581[128] = 16'h0000;
  assign literal_10581[129] = 16'h01f4;
  assign literal_10581[130] = 16'h1fec;
  assign literal_10581[131] = 16'hff9e;
  assign literal_10581[132] = 16'hffa3;
  assign literal_10581[133] = 16'hffb7;
  assign literal_10581[134] = 16'hffc1;
  assign literal_10581[135] = 16'hffce;
  assign literal_10581[136] = 16'hffdb;
  assign literal_10581[137] = 16'hffe9;
  assign literal_10581[138] = 16'hfff7;
  assign literal_10581[139] = 16'h0000;
  assign literal_10581[140] = 16'h0000;
  assign literal_10581[141] = 16'h0000;
  assign literal_10581[142] = 16'h0000;
  assign literal_10581[143] = 16'h0000;
  assign literal_10581[144] = 16'h0000;
  assign literal_10581[145] = 16'h01f7;
  assign literal_10581[146] = 16'h3fe0;
  assign literal_10581[147] = 16'hff91;
  assign literal_10581[148] = 16'hffa4;
  assign literal_10581[149] = 16'hffb8;
  assign literal_10581[150] = 16'hffc2;
  assign literal_10581[151] = 16'hffcf;
  assign literal_10581[152] = 16'hffdc;
  assign literal_10581[153] = 16'hffea;
  assign literal_10581[154] = 16'hfff8;
  assign literal_10581[155] = 16'h0000;
  assign literal_10581[156] = 16'h0000;
  assign literal_10581[157] = 16'h0000;
  assign literal_10581[158] = 16'h0000;
  assign literal_10581[159] = 16'h0000;
  assign literal_10581[160] = 16'h0000;
  assign literal_10581[161] = 16'h01f8;
  assign literal_10581[162] = 16'h3fe1;
  assign literal_10581[163] = 16'hff92;
  assign literal_10581[164] = 16'hffa7;
  assign literal_10581[165] = 16'hffb9;
  assign literal_10581[166] = 16'hffc3;
  assign literal_10581[167] = 16'hffd0;
  assign literal_10581[168] = 16'hffdd;
  assign literal_10581[169] = 16'hffeb;
  assign literal_10581[170] = 16'hfff9;
  assign literal_10581[171] = 16'h0000;
  assign literal_10581[172] = 16'h0000;
  assign literal_10581[173] = 16'h0000;
  assign literal_10581[174] = 16'h0000;
  assign literal_10581[175] = 16'h0000;
  assign literal_10581[176] = 16'h0000;
  assign literal_10581[177] = 16'h03f5;
  assign literal_10581[178] = 16'h7fc4;
  assign literal_10581[179] = 16'hff93;
  assign literal_10581[180] = 16'hffa8;
  assign literal_10581[181] = 16'hffba;
  assign literal_10581[182] = 16'hffc4;
  assign literal_10581[183] = 16'hffd1;
  assign literal_10581[184] = 16'hffde;
  assign literal_10581[185] = 16'hffec;
  assign literal_10581[186] = 16'hfffa;
  assign literal_10581[187] = 16'h0000;
  assign literal_10581[188] = 16'h0000;
  assign literal_10581[189] = 16'h0000;
  assign literal_10581[190] = 16'h0000;
  assign literal_10581[191] = 16'h0000;
  assign literal_10581[192] = 16'h0000;
  assign literal_10581[193] = 16'h03f8;
  assign literal_10581[194] = 16'hff8d;
  assign literal_10581[195] = 16'hff99;
  assign literal_10581[196] = 16'hffb1;
  assign literal_10581[197] = 16'hffbb;
  assign literal_10581[198] = 16'hffc5;
  assign literal_10581[199] = 16'hffd2;
  assign literal_10581[200] = 16'hffdf;
  assign literal_10581[201] = 16'hffed;
  assign literal_10581[202] = 16'hfffb;
  assign literal_10581[203] = 16'h0000;
  assign literal_10581[204] = 16'h0000;
  assign literal_10581[205] = 16'h0000;
  assign literal_10581[206] = 16'h0000;
  assign literal_10581[207] = 16'h0000;
  assign literal_10581[208] = 16'h0000;
  assign literal_10581[209] = 16'h03fa;
  assign literal_10581[210] = 16'hff9a;
  assign literal_10581[211] = 16'hffaa;
  assign literal_10581[212] = 16'hffb2;
  assign literal_10581[213] = 16'hffbc;
  assign literal_10581[214] = 16'hffc6;
  assign literal_10581[215] = 16'hffd3;
  assign literal_10581[216] = 16'hffe0;
  assign literal_10581[217] = 16'hffee;
  assign literal_10581[218] = 16'hfffc;
  assign literal_10581[219] = 16'h0000;
  assign literal_10581[220] = 16'h0000;
  assign literal_10581[221] = 16'h0000;
  assign literal_10581[222] = 16'h0000;
  assign literal_10581[223] = 16'h0000;
  assign literal_10581[224] = 16'h0000;
  assign literal_10581[225] = 16'h07f6;
  assign literal_10581[226] = 16'hff9b;
  assign literal_10581[227] = 16'hffaf;
  assign literal_10581[228] = 16'hffb3;
  assign literal_10581[229] = 16'hffbd;
  assign literal_10581[230] = 16'hffc7;
  assign literal_10581[231] = 16'hffd4;
  assign literal_10581[232] = 16'hffe1;
  assign literal_10581[233] = 16'hffef;
  assign literal_10581[234] = 16'hfffd;
  assign literal_10581[235] = 16'h0000;
  assign literal_10581[236] = 16'h0000;
  assign literal_10581[237] = 16'h0000;
  assign literal_10581[238] = 16'h0000;
  assign literal_10581[239] = 16'h0000;
  assign literal_10581[240] = 16'h0ff3;
  assign literal_10581[241] = 16'h1fed;
  assign literal_10581[242] = 16'hffae;
  assign literal_10581[243] = 16'hffb0;
  assign literal_10581[244] = 16'hffb4;
  assign literal_10581[245] = 16'hffbe;
  assign literal_10581[246] = 16'hffc8;
  assign literal_10581[247] = 16'hffd5;
  assign literal_10581[248] = 16'hffe2;
  assign literal_10581[249] = 16'hfff0;
  assign literal_10581[250] = 16'hfffe;
  assign literal_10581[251] = 16'h0000;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [8:0] p1_concat_9678_comb;
  wire [7:0] p1_concat_9676_comb;
  wire [6:0] p1_concat_9878_comb;
  wire [8:0] p1_add_9898_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed_comb;
  wire [2:0] p1_huff_length_squeezed_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__1_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__2_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__3_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__4_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__5_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__6_comb;
  wire [2:0] p1_huff_length_squeezed__1_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__7_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__8_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__9_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__10_comb;
  wire [2:0] p1_huff_length_squeezed__3_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__11_comb;
  wire [2:0] p1_huff_length_squeezed__4_comb;
  wire [2:0] p1_huff_length_squeezed__5_comb;
  wire [2:0] p1_huff_length_squeezed__6_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__12_comb;
  wire [2:0] p1_huff_length_squeezed__7_comb;
  wire [2:0] p1_huff_length_squeezed__8_comb;
  wire [2:0] p1_huff_length_squeezed__9_comb;
  wire [2:0] p1_huff_length_squeezed__10_comb;
  wire [2:0] p1_huff_length_squeezed__11_comb;
  wire [2:0] p1_huff_length_squeezed__12_comb;
  wire [2:0] p1_huff_length_squeezed__13_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__13_comb;
  wire [2:0] p1_huff_length_squeezed__14_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__14_comb;
  wire [2:0] p1_huff_length_squeezed__15_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__15_comb;
  wire [2:0] p1_huff_length_squeezed__16_comb;
  wire [5:0] p1_concat_9943_comb;
  wire [7:0] p1_flipped__2_comb;
  wire [7:0] p1_add_9680_comb;
  wire [6:0] p1_add_9886_comb;
  wire [7:0] p1_add_9909_comb;
  wire [9:0] p1_array_index_9814_comb;
  wire [9:0] p1_array_index_9815_comb;
  wire [9:0] p1_array_index_9816_comb;
  wire [9:0] p1_array_index_9817_comb;
  wire [9:0] p1_array_index_9818_comb;
  wire [9:0] p1_array_index_9819_comb;
  wire [9:0] p1_array_index_9820_comb;
  wire [9:0] p1_array_index_9821_comb;
  wire [9:0] p1_array_index_9822_comb;
  wire [9:0] p1_array_index_9823_comb;
  wire [9:0] p1_array_index_9824_comb;
  wire [9:0] p1_array_index_9825_comb;
  wire [9:0] p1_array_index_9826_comb;
  wire [9:0] p1_array_index_9827_comb;
  wire [9:0] p1_array_index_9828_comb;
  wire [9:0] p1_array_index_9829_comb;
  wire [9:0] p1_array_index_9830_comb;
  wire [9:0] p1_array_index_9831_comb;
  wire [9:0] p1_array_index_9832_comb;
  wire [9:0] p1_array_index_9833_comb;
  wire [9:0] p1_array_index_9834_comb;
  wire [9:0] p1_array_index_9835_comb;
  wire [9:0] p1_array_index_9836_comb;
  wire [9:0] p1_array_index_9837_comb;
  wire [9:0] p1_array_index_9838_comb;
  wire [9:0] p1_array_index_9839_comb;
  wire [9:0] p1_array_index_9840_comb;
  wire [9:0] p1_array_index_9841_comb;
  wire [9:0] p1_array_index_9842_comb;
  wire [9:0] p1_array_index_9843_comb;
  wire [9:0] p1_array_index_9844_comb;
  wire [9:0] p1_array_index_9845_comb;
  wire [9:0] p1_array_index_9846_comb;
  wire [9:0] p1_array_index_9847_comb;
  wire [9:0] p1_array_index_9848_comb;
  wire [9:0] p1_array_index_9849_comb;
  wire [9:0] p1_array_index_9850_comb;
  wire [9:0] p1_array_index_9851_comb;
  wire [9:0] p1_array_index_9852_comb;
  wire [9:0] p1_array_index_9853_comb;
  wire [9:0] p1_array_index_9854_comb;
  wire [9:0] p1_array_index_9855_comb;
  wire [9:0] p1_array_index_9856_comb;
  wire [9:0] p1_array_index_9857_comb;
  wire [9:0] p1_array_index_9858_comb;
  wire [9:0] p1_array_index_9859_comb;
  wire [9:0] p1_array_index_9860_comb;
  wire [9:0] p1_array_index_9861_comb;
  wire [9:0] p1_array_index_9862_comb;
  wire [9:0] p1_array_index_9863_comb;
  wire [9:0] p1_array_index_9864_comb;
  wire [9:0] p1_array_index_9865_comb;
  wire [9:0] p1_array_index_9866_comb;
  wire [9:0] p1_array_index_9867_comb;
  wire [9:0] p1_array_index_9868_comb;
  wire [9:0] p1_array_index_9869_comb;
  wire [9:0] p1_array_index_9870_comb;
  wire [9:0] p1_array_index_9871_comb;
  wire [9:0] p1_array_index_9872_comb;
  wire [9:0] p1_array_index_9873_comb;
  wire [9:0] p1_array_index_9874_comb;
  wire [9:0] p1_array_index_9875_comb;
  wire [9:0] p1_array_index_9876_comb;
  wire [8:0] p1_add_9912_comb;
  wire [7:0] p1_add_9913_comb;
  wire [5:0] p1_add_9961_comb;
  wire [7:0] p1_add_10000_comb;
  wire [6:0] p1_add_10030_comb;
  wire [7:0] p1_add_10062_comb;
  wire [8:0] p1_add_9682_comb;
  wire [8:0] p1_concat_9812_comb;
  wire [8:0] p1_add_9877_comb;
  wire [8:0] p1_concat_9902_comb;
  wire [8:0] p1_add_9914_comb;
  wire [8:0] p1_concat_9926_comb;
  wire [8:0] p1_add_9931_comb;
  wire [6:0] p1_add_9954_comb;
  wire [8:0] p1_add_9974_comb;
  wire [8:0] p1_concat_9983_comb;
  wire [7:0] p1_add_9990_comb;
  wire [8:0] p1_add_9999_comb;
  wire [8:0] p1_add_10001_comb;
  wire [8:0] p1_concat_10014_comb;
  wire [8:0] p1_add_10031_comb;
  wire [5:0] p1_add_10040_comb;
  wire [8:0] p1_concat_10048_comb;
  wire [8:0] p1_add_10058_comb;
  wire [8:0] p1_add_10063_comb;
  wire [7:0] p1_add_10074_comb;
  wire [8:0] p1_concat_10080_comb;
  wire [8:0] p1_add_10091_comb;
  wire [6:0] p1_add_10108_comb;
  wire [8:0] p1_add_10128_comb;
  wire [7:0] p1_add_10143_comb;
  wire [8:0] p1_add_10153_comb;
  wire [8:0] p1_add_10088_comb;
  wire [7:0] p1_huff_length_comb;
  wire [7:0] p1_huff_length__1_comb;
  wire [1:0] p1_concat_9977_comb;
  wire [1:0] p1_huff_length__1_squeezed__2_comb;
  wire p1_nor_9905_comb;
  wire p1_or_9916_comb;
  wire p1_nor_9917_comb;
  wire [9:0] p1_value__1_comb;
  wire p1_or_9968_comb;
  wire p1_or_9986_comb;
  wire [1:0] p1_sel_9996_comb;
  wire [1:0] p1_sign_ext_9997_comb;
  wire p1_or_10003_comb;
  wire p1_nor_10004_comb;
  wire p1_or_10026_comb;
  wire p1_or_10043_comb;
  wire p1_or_10055_comb;
  wire p1_or_10060_comb;
  wire p1_nor_10061_comb;
  wire p1_or_10070_comb;
  wire p1_or_10087_comb;
  wire p1_or_10104_comb;
  wire p1_or_10116_comb;
  wire p1_or_10122_comb;
  wire p1_or_10135_comb;
  wire p1_or_10139_comb;
  wire p1_eq_10140_comb;
  wire p1_ne_10141_comb;
  wire p1_or_10151_comb;
  wire p1_or_10154_comb;
  wire p1_or_10161_comb;
  wire p1_or_10169_comb;
  wire p1_or_10175_comb;
  wire p1_or_10241_comb;
  wire p1_nor_10242_comb;
  wire p1_and_10306_comb;
  assign p1_concat_9678_comb = {1'h0, p0_start_pix};
  assign p1_concat_9676_comb = {1'h0, p0_start_pix[7:1]};
  assign p1_concat_9878_comb = {1'h0, p0_start_pix[7:2]};
  assign p1_add_9898_comb = p1_concat_9678_comb + 9'h00f;
  assign p1_huff_code__1_squeezed_squeezed_comb = 3'h1;
  assign p1_huff_length_squeezed_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__1_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__2_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__3_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__4_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__5_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__6_comb = 3'h1;
  assign p1_huff_length_squeezed__1_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__7_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__8_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__9_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__10_comb = 3'h1;
  assign p1_huff_length_squeezed__3_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__11_comb = 3'h1;
  assign p1_huff_length_squeezed__4_comb = 3'h4;
  assign p1_huff_length_squeezed__5_comb = 3'h4;
  assign p1_huff_length_squeezed__6_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__12_comb = 3'h1;
  assign p1_huff_length_squeezed__7_comb = 3'h4;
  assign p1_huff_length_squeezed__8_comb = 3'h4;
  assign p1_huff_length_squeezed__9_comb = 3'h4;
  assign p1_huff_length_squeezed__10_comb = 3'h4;
  assign p1_huff_length_squeezed__11_comb = 3'h4;
  assign p1_huff_length_squeezed__12_comb = 3'h4;
  assign p1_huff_length_squeezed__13_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__13_comb = 3'h1;
  assign p1_huff_length_squeezed__14_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__14_comb = 3'h1;
  assign p1_huff_length_squeezed__15_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__15_comb = 3'h1;
  assign p1_huff_length_squeezed__16_comb = 3'h4;
  assign p1_concat_9943_comb = {1'h0, p0_start_pix[7:3]};
  assign p1_flipped__2_comb = 8'hff;
  assign p1_add_9680_comb = p1_concat_9676_comb + 8'hf9;
  assign p1_add_9886_comb = p1_concat_9878_comb + 7'h7d;
  assign p1_add_9909_comb = p1_concat_9676_comb + 8'h07;
  assign p1_array_index_9814_comb = p0_matrix[3'h0][3'h0];
  assign p1_array_index_9815_comb = p0_matrix[3'h0][p1_huff_code__1_squeezed_squeezed_comb];
  assign p1_array_index_9816_comb = p0_matrix[3'h0][3'h2];
  assign p1_array_index_9817_comb = p0_matrix[3'h0][3'h3];
  assign p1_array_index_9818_comb = p0_matrix[3'h0][p1_huff_length_squeezed_comb];
  assign p1_array_index_9819_comb = p0_matrix[3'h0][3'h5];
  assign p1_array_index_9820_comb = p0_matrix[3'h0][3'h6];
  assign p1_array_index_9821_comb = p0_matrix[3'h0][3'h7];
  assign p1_array_index_9822_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__1_comb][3'h0];
  assign p1_array_index_9823_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__2_comb][p1_huff_code__1_squeezed_squeezed__3_comb];
  assign p1_array_index_9824_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__4_comb][3'h2];
  assign p1_array_index_9825_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__5_comb][3'h3];
  assign p1_array_index_9826_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__6_comb][p1_huff_length_squeezed__1_comb];
  assign p1_array_index_9827_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__7_comb][3'h5];
  assign p1_array_index_9828_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__8_comb][3'h6];
  assign p1_array_index_9829_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__9_comb][3'h7];
  assign p1_array_index_9830_comb = p0_matrix[3'h2][3'h0];
  assign p1_array_index_9831_comb = p0_matrix[3'h2][p1_huff_code__1_squeezed_squeezed__10_comb];
  assign p1_array_index_9832_comb = p0_matrix[3'h2][3'h2];
  assign p1_array_index_9833_comb = p0_matrix[3'h2][3'h3];
  assign p1_array_index_9834_comb = p0_matrix[3'h2][p1_huff_length_squeezed__3_comb];
  assign p1_array_index_9835_comb = p0_matrix[3'h2][3'h5];
  assign p1_array_index_9836_comb = p0_matrix[3'h2][3'h6];
  assign p1_array_index_9837_comb = p0_matrix[3'h2][3'h7];
  assign p1_array_index_9838_comb = p0_matrix[3'h3][3'h0];
  assign p1_array_index_9839_comb = p0_matrix[3'h3][p1_huff_code__1_squeezed_squeezed__11_comb];
  assign p1_array_index_9840_comb = p0_matrix[3'h3][3'h2];
  assign p1_array_index_9841_comb = p0_matrix[3'h3][3'h3];
  assign p1_array_index_9842_comb = p0_matrix[3'h3][p1_huff_length_squeezed__4_comb];
  assign p1_array_index_9843_comb = p0_matrix[3'h3][3'h5];
  assign p1_array_index_9844_comb = p0_matrix[3'h3][3'h6];
  assign p1_array_index_9845_comb = p0_matrix[3'h3][3'h7];
  assign p1_array_index_9846_comb = p0_matrix[p1_huff_length_squeezed__5_comb][3'h0];
  assign p1_array_index_9847_comb = p0_matrix[p1_huff_length_squeezed__6_comb][p1_huff_code__1_squeezed_squeezed__12_comb];
  assign p1_array_index_9848_comb = p0_matrix[p1_huff_length_squeezed__7_comb][3'h2];
  assign p1_array_index_9849_comb = p0_matrix[p1_huff_length_squeezed__8_comb][3'h3];
  assign p1_array_index_9850_comb = p0_matrix[p1_huff_length_squeezed__9_comb][p1_huff_length_squeezed__10_comb];
  assign p1_array_index_9851_comb = p0_matrix[p1_huff_length_squeezed__11_comb][3'h5];
  assign p1_array_index_9852_comb = p0_matrix[p1_huff_length_squeezed__12_comb][3'h6];
  assign p1_array_index_9853_comb = p0_matrix[p1_huff_length_squeezed__13_comb][3'h7];
  assign p1_array_index_9854_comb = p0_matrix[3'h5][3'h0];
  assign p1_array_index_9855_comb = p0_matrix[3'h5][p1_huff_code__1_squeezed_squeezed__13_comb];
  assign p1_array_index_9856_comb = p0_matrix[3'h5][3'h2];
  assign p1_array_index_9857_comb = p0_matrix[3'h5][3'h3];
  assign p1_array_index_9858_comb = p0_matrix[3'h5][p1_huff_length_squeezed__14_comb];
  assign p1_array_index_9859_comb = p0_matrix[3'h5][3'h5];
  assign p1_array_index_9860_comb = p0_matrix[3'h5][3'h6];
  assign p1_array_index_9861_comb = p0_matrix[3'h5][3'h7];
  assign p1_array_index_9862_comb = p0_matrix[3'h6][3'h0];
  assign p1_array_index_9863_comb = p0_matrix[3'h6][p1_huff_code__1_squeezed_squeezed__14_comb];
  assign p1_array_index_9864_comb = p0_matrix[3'h6][3'h2];
  assign p1_array_index_9865_comb = p0_matrix[3'h6][3'h3];
  assign p1_array_index_9866_comb = p0_matrix[3'h6][p1_huff_length_squeezed__15_comb];
  assign p1_array_index_9867_comb = p0_matrix[3'h6][3'h5];
  assign p1_array_index_9868_comb = p0_matrix[3'h6][3'h6];
  assign p1_array_index_9869_comb = p0_matrix[3'h6][3'h7];
  assign p1_array_index_9870_comb = p0_matrix[3'h7][3'h0];
  assign p1_array_index_9871_comb = p0_matrix[3'h7][p1_huff_code__1_squeezed_squeezed__15_comb];
  assign p1_array_index_9872_comb = p0_matrix[3'h7][3'h2];
  assign p1_array_index_9873_comb = p0_matrix[3'h7][3'h3];
  assign p1_array_index_9874_comb = p0_matrix[3'h7][p1_huff_length_squeezed__16_comb];
  assign p1_array_index_9875_comb = p0_matrix[3'h7][3'h5];
  assign p1_array_index_9876_comb = p0_matrix[3'h7][3'h6];
  assign p1_add_9912_comb = p1_concat_9678_comb + 9'h00d;
  assign p1_add_9913_comb = p1_concat_9676_comb + 8'hfb;
  assign p1_add_9961_comb = p1_concat_9943_comb + 6'h3f;
  assign p1_add_10000_comb = p1_concat_9676_comb + 8'hfd;
  assign p1_add_10030_comb = p1_concat_9878_comb + 7'h7f;
  assign p1_add_10062_comb = p1_concat_9676_comb + p1_flipped__2_comb;
  assign p1_add_9682_comb = p1_concat_9678_comb + 9'h1f1;
  assign p1_concat_9812_comb = {p1_add_9680_comb, p0_start_pix[0]};
  assign p1_add_9877_comb = p1_concat_9678_comb + 9'h1f3;
  assign p1_concat_9902_comb = {p1_add_9886_comb, p0_start_pix[1:0]};
  assign p1_add_9914_comb = p1_concat_9678_comb + 9'h1f5;
  assign p1_concat_9926_comb = {p1_add_9913_comb, p0_start_pix[0]};
  assign p1_add_9931_comb = p1_concat_9678_comb + 9'h1f7;
  assign p1_add_9954_comb = p1_concat_9878_comb + 7'h03;
  assign p1_add_9974_comb = p1_concat_9678_comb + 9'h00b;
  assign p1_concat_9983_comb = {p1_add_9961_comb, p0_start_pix[2:0]};
  assign p1_add_9990_comb = p1_concat_9676_comb + 8'h05;
  assign p1_add_9999_comb = p1_concat_9678_comb + 9'h009;
  assign p1_add_10001_comb = p1_concat_9678_comb + 9'h1f9;
  assign p1_concat_10014_comb = {p1_add_10000_comb, p0_start_pix[0]};
  assign p1_add_10031_comb = p1_concat_9678_comb + 9'h1fb;
  assign p1_add_10040_comb = p1_concat_9943_comb + 6'h01;
  assign p1_concat_10048_comb = {p1_add_10030_comb, p0_start_pix[1:0]};
  assign p1_add_10058_comb = p1_concat_9678_comb + 9'h007;
  assign p1_add_10063_comb = p1_concat_9678_comb + 9'h1fd;
  assign p1_add_10074_comb = p1_concat_9676_comb + 8'h03;
  assign p1_concat_10080_comb = {p1_add_10062_comb, p0_start_pix[0]};
  assign p1_add_10091_comb = p1_concat_9678_comb + 9'h005;
  assign p1_add_10108_comb = p1_concat_9878_comb + 7'h01;
  assign p1_add_10128_comb = p1_concat_9678_comb + 9'h003;
  assign p1_add_10143_comb = p1_concat_9676_comb + 8'h01;
  assign p1_add_10153_comb = p1_concat_9678_comb + 9'h001;
  assign p1_add_10088_comb = p1_concat_9678_comb + 9'h1ff;
  assign p1_huff_length_comb = 8'h04;
  assign p1_huff_length__1_comb = 8'h02;
  assign p1_concat_9977_comb = {1'h1, ~(p1_add_9898_comb > 9'h03e | ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_9898_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000)};
  assign p1_huff_length__1_squeezed__2_comb = 2'h1;
  assign p1_nor_9905_comb = ~(p0_start_pix == 8'h0e | ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_add_9682_comb[8]}}, p1_add_9682_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000);
  assign p1_or_9916_comb = p0_start_pix == 8'h0d | ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_concat_9812_comb[8]}}, p1_concat_9812_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_nor_9917_comb = ~(p0_start_pix == 8'h0c | ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_add_9877_comb[8]}}, p1_add_9877_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000);
  assign p1_value__1_comb = p0_start_pix == 8'h00 ? p1_array_index_9814_comb : (p0_start_pix == 8'h01 ? p1_array_index_9815_comb : (p0_start_pix == 8'h02 ? p1_array_index_9816_comb : (p0_start_pix == 8'h03 ? p1_array_index_9817_comb : (p0_start_pix == 8'h04 ? p1_array_index_9818_comb : (p0_start_pix == 8'h05 ? p1_array_index_9819_comb : (p0_start_pix == 8'h06 ? p1_array_index_9820_comb : (p0_start_pix == 8'h07 ? p1_array_index_9821_comb : (p0_start_pix == 8'h08 ? p1_array_index_9822_comb : (p0_start_pix == 8'h09 ? p1_array_index_9823_comb : (p0_start_pix == 8'h0a ? p1_array_index_9824_comb : (p0_start_pix == 8'h0b ? p1_array_index_9825_comb : (p0_start_pix == 8'h0c ? p1_array_index_9826_comb : (p0_start_pix == 8'h0d ? p1_array_index_9827_comb : (p0_start_pix == 8'h0e ? p1_array_index_9828_comb : (p0_start_pix == 8'h0f ? p1_array_index_9829_comb : (p0_start_pix == 8'h10 ? p1_array_index_9830_comb : (p0_start_pix == 8'h11 ? p1_array_index_9831_comb : (p0_start_pix == 8'h12 ? p1_array_index_9832_comb : (p0_start_pix == 8'h13 ? p1_array_index_9833_comb : (p0_start_pix == 8'h14 ? p1_array_index_9834_comb : (p0_start_pix == 8'h15 ? p1_array_index_9835_comb : (p0_start_pix == 8'h16 ? p1_array_index_9836_comb : (p0_start_pix == 8'h17 ? p1_array_index_9837_comb : (p0_start_pix == 8'h18 ? p1_array_index_9838_comb : (p0_start_pix == 8'h19 ? p1_array_index_9839_comb : (p0_start_pix == 8'h1a ? p1_array_index_9840_comb : (p0_start_pix == 8'h1b ? p1_array_index_9841_comb : (p0_start_pix == 8'h1c ? p1_array_index_9842_comb : (p0_start_pix == 8'h1d ? p1_array_index_9843_comb : (p0_start_pix == 8'h1e ? p1_array_index_9844_comb : (p0_start_pix == 8'h1f ? p1_array_index_9845_comb : (p0_start_pix == 8'h20 ? p1_array_index_9846_comb : (p0_start_pix == 8'h21 ? p1_array_index_9847_comb : (p0_start_pix == 8'h22 ? p1_array_index_9848_comb : (p0_start_pix == 8'h23 ? p1_array_index_9849_comb : (p0_start_pix == 8'h24 ? p1_array_index_9850_comb : (p0_start_pix == 8'h25 ? p1_array_index_9851_comb : (p0_start_pix == 8'h26 ? p1_array_index_9852_comb : (p0_start_pix == 8'h27 ? p1_array_index_9853_comb : (p0_start_pix == 8'h28 ? p1_array_index_9854_comb : (p0_start_pix == 8'h29 ? p1_array_index_9855_comb : (p0_start_pix == 8'h2a ? p1_array_index_9856_comb : (p0_start_pix == 8'h2b ? p1_array_index_9857_comb : (p0_start_pix == 8'h2c ? p1_array_index_9858_comb : (p0_start_pix == 8'h2d ? p1_array_index_9859_comb : (p0_start_pix == 8'h2e ? p1_array_index_9860_comb : (p0_start_pix == 8'h2f ? p1_array_index_9861_comb : (p0_start_pix == 8'h30 ? p1_array_index_9862_comb : (p0_start_pix == 8'h31 ? p1_array_index_9863_comb : (p0_start_pix == 8'h32 ? p1_array_index_9864_comb : (p0_start_pix == 8'h33 ? p1_array_index_9865_comb : (p0_start_pix == 8'h34 ? p1_array_index_9866_comb : (p0_start_pix == 8'h35 ? p1_array_index_9867_comb : (p0_start_pix == 8'h36 ? p1_array_index_9868_comb : (p0_start_pix == 8'h37 ? p1_array_index_9869_comb : (p0_start_pix == 8'h38 ? p1_array_index_9870_comb : (p0_start_pix == 8'h39 ? p1_array_index_9871_comb : (p0_start_pix == 8'h3a ? p1_array_index_9872_comb : (p0_start_pix == 8'h3b ? p1_array_index_9873_comb : (p0_start_pix == 8'h3c ? p1_array_index_9874_comb : (p0_start_pix == 8'h3d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign p1_or_9968_comb = p0_start_pix == 8'h0b | ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_concat_9902_comb[8]}}, p1_concat_9902_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_9986_comb = p0_start_pix == 8'h0a | ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_add_9914_comb[8]}}, p1_add_9914_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_sel_9996_comb = {p1_add_9909_comb, p0_start_pix[0]} > 9'h03e | ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_9909_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000 ? p1_huff_length__1_squeezed__2_comb : p1_concat_9977_comb;
  assign p1_sign_ext_9997_comb = {2{~(p1_add_9912_comb > 9'h03e | ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_9912_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000)}};
  assign p1_or_10003_comb = p0_start_pix == 8'h09 | ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_concat_9926_comb[8]}}, p1_concat_9926_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_nor_10004_comb = ~(p0_start_pix == 8'h08 | ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_add_9931_comb[8]}}, p1_add_9931_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000);
  assign p1_or_10026_comb = {p1_add_9954_comb, p0_start_pix[1:0]} > 9'h03e | ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_9954_comb, p0_start_pix[1:0]} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10043_comb = p1_add_9974_comb > 9'h03e | ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_9974_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10055_comb = p0_start_pix == 8'h07 | ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_concat_9983_comb[8]}}, p1_concat_9983_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10060_comb = {p1_add_9990_comb, p0_start_pix[0]} > 9'h03e | ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_9990_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_nor_10061_comb = ~(p1_add_9999_comb > 9'h03e | ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_9999_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000);
  assign p1_or_10070_comb = p0_start_pix == 8'h06 | ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_add_10001_comb[8]}}, p1_add_10001_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10087_comb = p0_start_pix == 8'h05 | ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_concat_10014_comb[8]}}, p1_concat_10014_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10104_comb = p0_start_pix == p1_huff_length_comb | ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_add_10031_comb[8]}}, p1_add_10031_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10116_comb = {p1_add_10040_comb, p0_start_pix[2:0]} > 9'h03e | ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_10040_comb, p0_start_pix[2:0]} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10122_comb = p0_start_pix == 8'h03 | ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_concat_10048_comb[8]}}, p1_concat_10048_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10135_comb = p1_add_10058_comb > 9'h03e | ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_10058_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10139_comb = p0_start_pix == p1_huff_length__1_comb | ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_add_10063_comb[8]}}, p1_add_10063_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_eq_10140_comb = p0_start_pix == 8'h00;
  assign p1_ne_10141_comb = ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_add_10088_comb[8]}}, p1_add_10088_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10151_comb = {p1_add_10074_comb, p0_start_pix[0]} > 9'h03e | ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_10074_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10154_comb = p0_start_pix == 8'h01 | ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({{23{p1_concat_10080_comb[8]}}, p1_concat_10080_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10161_comb = p1_add_10091_comb > 9'h03e | ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_10091_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10169_comb = {p1_add_10108_comb, p0_start_pix[1:0]} > 9'h03e | ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_10108_comb, p0_start_pix[1:0]} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10175_comb = p1_add_10128_comb > 9'h03e | ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_10128_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10241_comb = {p1_add_10143_comb, p0_start_pix[0]} > 9'h03e | ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_10143_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_nor_10242_comb = ~(p1_add_10153_comb > 9'h03e | ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0000 ? p1_array_index_9814_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0001 ? p1_array_index_9815_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0002 ? p1_array_index_9816_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0003 ? p1_array_index_9817_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0004 ? p1_array_index_9818_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0005 ? p1_array_index_9819_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0006 ? p1_array_index_9820_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0007 ? p1_array_index_9821_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0008 ? p1_array_index_9822_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0009 ? p1_array_index_9823_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_000a ? p1_array_index_9824_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_000b ? p1_array_index_9825_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_000c ? p1_array_index_9826_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_000d ? p1_array_index_9827_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_000e ? p1_array_index_9828_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_000f ? p1_array_index_9829_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0010 ? p1_array_index_9830_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0011 ? p1_array_index_9831_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0012 ? p1_array_index_9832_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0013 ? p1_array_index_9833_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0014 ? p1_array_index_9834_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0015 ? p1_array_index_9835_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0016 ? p1_array_index_9836_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0017 ? p1_array_index_9837_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0018 ? p1_array_index_9838_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0019 ? p1_array_index_9839_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_001a ? p1_array_index_9840_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_001b ? p1_array_index_9841_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_001c ? p1_array_index_9842_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_001d ? p1_array_index_9843_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_001e ? p1_array_index_9844_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_001f ? p1_array_index_9845_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0020 ? p1_array_index_9846_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0021 ? p1_array_index_9847_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0022 ? p1_array_index_9848_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0023 ? p1_array_index_9849_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0024 ? p1_array_index_9850_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0025 ? p1_array_index_9851_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0026 ? p1_array_index_9852_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0027 ? p1_array_index_9853_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0028 ? p1_array_index_9854_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0029 ? p1_array_index_9855_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_002a ? p1_array_index_9856_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_002b ? p1_array_index_9857_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_002c ? p1_array_index_9858_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_002d ? p1_array_index_9859_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_002e ? p1_array_index_9860_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_002f ? p1_array_index_9861_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0030 ? p1_array_index_9862_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0031 ? p1_array_index_9863_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0032 ? p1_array_index_9864_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0033 ? p1_array_index_9865_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0034 ? p1_array_index_9866_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0035 ? p1_array_index_9867_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0036 ? p1_array_index_9868_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0037 ? p1_array_index_9869_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0038 ? p1_array_index_9870_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_0039 ? p1_array_index_9871_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_003a ? p1_array_index_9872_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_003b ? p1_array_index_9873_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_003c ? p1_array_index_9874_comb : ({23'h00_0000, p1_add_10153_comb} == 32'h0000_003d ? p1_array_index_9875_comb : p1_array_index_9876_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000);
  assign p1_and_10306_comb = p1_array_index_9814_comb == 10'h000 & p1_array_index_9815_comb == 10'h000 & p1_array_index_9816_comb == 10'h000 & p1_array_index_9817_comb == 10'h000 & p1_array_index_9818_comb == 10'h000 & p1_array_index_9819_comb == 10'h000 & p1_array_index_9820_comb == 10'h000 & p1_array_index_9821_comb == 10'h000 & p1_array_index_9822_comb == 10'h000 & p1_array_index_9823_comb == 10'h000 & p1_array_index_9824_comb == 10'h000 & p1_array_index_9825_comb == 10'h000 & p1_array_index_9826_comb == 10'h000 & p1_array_index_9827_comb == 10'h000 & p1_array_index_9828_comb == 10'h000 & p1_array_index_9829_comb == 10'h000 & p1_array_index_9830_comb == 10'h000 & p1_array_index_9831_comb == 10'h000 & p1_array_index_9832_comb == 10'h000 & p1_array_index_9833_comb == 10'h000 & p1_array_index_9834_comb == 10'h000 & p1_array_index_9835_comb == 10'h000 & p1_array_index_9836_comb == 10'h000 & p1_array_index_9837_comb == 10'h000 & p1_array_index_9838_comb == 10'h000 & p1_array_index_9839_comb == 10'h000 & p1_array_index_9840_comb == 10'h000 & p1_array_index_9841_comb == 10'h000 & p1_array_index_9842_comb == 10'h000 & p1_array_index_9843_comb == 10'h000 & p1_array_index_9844_comb == 10'h000 & p1_array_index_9845_comb == 10'h000 & p1_array_index_9846_comb == 10'h000 & p1_array_index_9847_comb == 10'h000 & p1_array_index_9848_comb == 10'h000 & p1_array_index_9849_comb == 10'h000 & p1_array_index_9850_comb == 10'h000 & p1_array_index_9851_comb == 10'h000 & p1_array_index_9852_comb == 10'h000 & p1_array_index_9853_comb == 10'h000 & p1_array_index_9854_comb == 10'h000 & p1_array_index_9855_comb == 10'h000 & p1_array_index_9856_comb == 10'h000 & p1_array_index_9857_comb == 10'h000 & p1_array_index_9858_comb == 10'h000 & p1_array_index_9859_comb == 10'h000 & p1_array_index_9860_comb == 10'h000 & p1_array_index_9861_comb == 10'h000 & p1_array_index_9862_comb == 10'h000 & p1_array_index_9863_comb == 10'h000 & p1_array_index_9864_comb == 10'h000 & p1_array_index_9865_comb == 10'h000 & p1_array_index_9866_comb == 10'h000 & p1_array_index_9867_comb == 10'h000 & p1_array_index_9868_comb == 10'h000 & p1_array_index_9869_comb == 10'h000 & p1_array_index_9870_comb == 10'h000 & p1_array_index_9871_comb == 10'h000 & p1_array_index_9872_comb == 10'h000 & p1_array_index_9873_comb == 10'h000 & p1_array_index_9874_comb == 10'h000 & p1_array_index_9875_comb == 10'h000 & p1_array_index_9876_comb == 10'h000;

  // Registers for pipe stage 1:
  reg p1_is_luminance;
  reg p1_nor_9905;
  reg p1_or_9916;
  reg p1_nor_9917;
  reg [9:0] p1_value__1;
  reg p1_or_9968;
  reg p1_or_9986;
  reg [1:0] p1_sel_9996;
  reg [1:0] p1_sign_ext_9997;
  reg p1_or_10003;
  reg p1_nor_10004;
  reg p1_or_10026;
  reg p1_or_10043;
  reg p1_or_10055;
  reg p1_or_10060;
  reg p1_nor_10061;
  reg p1_or_10070;
  reg p1_or_10087;
  reg p1_or_10104;
  reg p1_or_10116;
  reg p1_or_10122;
  reg p1_or_10135;
  reg p1_or_10139;
  reg p1_eq_10140;
  reg p1_ne_10141;
  reg p1_or_10151;
  reg p1_or_10154;
  reg p1_or_10161;
  reg p1_or_10169;
  reg p1_or_10175;
  reg p1_or_10241;
  reg p1_nor_10242;
  reg p1_and_10306;
  always @ (posedge clk) begin
    p1_is_luminance <= p0_is_luminance;
    p1_nor_9905 <= p1_nor_9905_comb;
    p1_or_9916 <= p1_or_9916_comb;
    p1_nor_9917 <= p1_nor_9917_comb;
    p1_value__1 <= p1_value__1_comb;
    p1_or_9968 <= p1_or_9968_comb;
    p1_or_9986 <= p1_or_9986_comb;
    p1_sel_9996 <= p1_sel_9996_comb;
    p1_sign_ext_9997 <= p1_sign_ext_9997_comb;
    p1_or_10003 <= p1_or_10003_comb;
    p1_nor_10004 <= p1_nor_10004_comb;
    p1_or_10026 <= p1_or_10026_comb;
    p1_or_10043 <= p1_or_10043_comb;
    p1_or_10055 <= p1_or_10055_comb;
    p1_or_10060 <= p1_or_10060_comb;
    p1_nor_10061 <= p1_nor_10061_comb;
    p1_or_10070 <= p1_or_10070_comb;
    p1_or_10087 <= p1_or_10087_comb;
    p1_or_10104 <= p1_or_10104_comb;
    p1_or_10116 <= p1_or_10116_comb;
    p1_or_10122 <= p1_or_10122_comb;
    p1_or_10135 <= p1_or_10135_comb;
    p1_or_10139 <= p1_or_10139_comb;
    p1_eq_10140 <= p1_eq_10140_comb;
    p1_ne_10141 <= p1_ne_10141_comb;
    p1_or_10151 <= p1_or_10151_comb;
    p1_or_10154 <= p1_or_10154_comb;
    p1_or_10161 <= p1_or_10161_comb;
    p1_or_10169 <= p1_or_10169_comb;
    p1_or_10175 <= p1_or_10175_comb;
    p1_or_10241 <= p1_or_10241_comb;
    p1_nor_10242 <= p1_nor_10242_comb;
    p1_and_10306 <= p1_and_10306_comb;
  end

  // ===== Pipe stage 2:
  wire [1:0] p2_huff_length__1_squeezed__1_comb;
  wire [7:0] p2_bin_value__2_comb;
  wire [7:0] p2_bin_value__3_comb;
  wire [7:0] p2_value_abs_comb;
  wire [2:0] p2_huff_code__1_squeezed_squeezed__17_comb;
  wire [2:0] p2_sel_10385_comb;
  wire [2:0] p2_huff_code__1_squeezed_squeezed__16_comb;
  wire [1:0] p2_huff_length__1_squeezed__3_comb;
  wire [1:0] p2_huff_length__1_squeezed_comb;
  wire [2:0] p2_and_10418_comb;
  wire [7:0] p2_flipped__1_comb;
  wire [7:0] p2_flipped_comb;
  wire [2:0] p2_and_10401_comb;
  wire [1:0] p2_sel_10408_comb;
  wire p2_or_reduce_10412_comb;
  wire p2_or_reduce_10416_comb;
  wire p2_or_reduce_10420_comb;
  wire p2_or_reduce_10423_comb;
  wire [3:0] p2_sel_10424_comb;
  wire p2_bit_slice_10425_comb;
  wire p2_ne_10427_comb;
  wire [7:0] p2_Code_list_comb;
  wire [7:0] p2_code_list_comb;
  assign p2_huff_length__1_squeezed__1_comb = 2'h1;
  assign p2_bin_value__2_comb = p1_value__1[7:0];
  assign p2_bin_value__3_comb = -p2_bin_value__2_comb;
  assign p2_value_abs_comb = p1_value__1[9] ? p2_bin_value__3_comb : p2_bin_value__2_comb;
  assign p2_huff_code__1_squeezed_squeezed__17_comb = 3'h1;
  assign p2_sel_10385_comb = p1_or_9968 ? 3'h3 : {1'h1, (p1_or_9916 ? p2_huff_length__1_squeezed__1_comb : {1'h1, p1_nor_9905}) & {2{p1_nor_9917}}};
  assign p2_huff_code__1_squeezed_squeezed__16_comb = 3'h1;
  assign p2_huff_length__1_squeezed__3_comb = 2'h1;
  assign p2_huff_length__1_squeezed_comb = 2'h2;
  assign p2_and_10418_comb = (p1_or_10060 ? p2_huff_code__1_squeezed_squeezed__17_comb : (p1_or_10043 ? 3'h2 : (p1_or_10026 ? 3'h3 : {1'h1, p1_sel_9996 & p1_sign_ext_9997}))) & {3{p1_nor_10061}};
  assign p2_flipped__1_comb = ~p2_bin_value__3_comb;
  assign p2_flipped_comb = 8'hff;
  assign p2_and_10401_comb = (p1_or_10003 ? p2_huff_code__1_squeezed_squeezed__16_comb : (p1_or_9986 ? 3'h2 : p2_sel_10385_comb)) & {3{p1_nor_10004}};
  assign p2_sel_10408_comb = |p2_value_abs_comb[7:2] ? 2'h3 : (|p2_value_abs_comb[7:1] ? p2_huff_length__1_squeezed_comb : p2_huff_length__1_squeezed__3_comb);
  assign p2_or_reduce_10412_comb = |p2_value_abs_comb[7:3];
  assign p2_or_reduce_10416_comb = |p2_value_abs_comb[7:4];
  assign p2_or_reduce_10420_comb = |p2_value_abs_comb[7:5];
  assign p2_or_reduce_10423_comb = |p2_value_abs_comb[7:6];
  assign p2_sel_10424_comb = p1_or_10116 ? 4'h7 : {1'h1, p2_and_10418_comb};
  assign p2_bit_slice_10425_comb = p2_value_abs_comb[7];
  assign p2_ne_10427_comb = p2_value_abs_comb != 8'h00;
  assign p2_Code_list_comb = $signed(p1_value__1) <= $signed(10'h000) ? p2_flipped__1_comb : p2_bin_value__2_comb;
  assign p2_code_list_comb = p1_value__1 == 10'h000 ? p2_flipped_comb : p2_bin_value__2_comb;

  // Registers for pipe stage 2:
  reg p2_is_luminance;
  reg [2:0] p2_and_10401;
  reg p2_or_10055;
  reg [1:0] p2_sel_10408;
  reg p2_or_10070;
  reg p2_or_reduce_10412;
  reg p2_or_10087;
  reg p2_or_reduce_10416;
  reg p2_or_10104;
  reg p2_or_reduce_10420;
  reg p2_or_10122;
  reg p2_or_reduce_10423;
  reg p2_or_10135;
  reg [3:0] p2_sel_10424;
  reg p2_or_10139;
  reg p2_eq_10140;
  reg p2_ne_10141;
  reg p2_or_10151;
  reg p2_or_10154;
  reg p2_bit_slice_10425;
  reg p2_or_10161;
  reg p2_ne_10427;
  reg p2_or_10169;
  reg p2_or_10175;
  reg p2_or_10241;
  reg p2_nor_10242;
  reg p2_and_10306;
  reg [7:0] p2_Code_list;
  reg [7:0] p2_code_list;
  always @ (posedge clk) begin
    p2_is_luminance <= p1_is_luminance;
    p2_and_10401 <= p2_and_10401_comb;
    p2_or_10055 <= p1_or_10055;
    p2_sel_10408 <= p2_sel_10408_comb;
    p2_or_10070 <= p1_or_10070;
    p2_or_reduce_10412 <= p2_or_reduce_10412_comb;
    p2_or_10087 <= p1_or_10087;
    p2_or_reduce_10416 <= p2_or_reduce_10416_comb;
    p2_or_10104 <= p1_or_10104;
    p2_or_reduce_10420 <= p2_or_reduce_10420_comb;
    p2_or_10122 <= p1_or_10122;
    p2_or_reduce_10423 <= p2_or_reduce_10423_comb;
    p2_or_10135 <= p1_or_10135;
    p2_sel_10424 <= p2_sel_10424_comb;
    p2_or_10139 <= p1_or_10139;
    p2_eq_10140 <= p1_eq_10140;
    p2_ne_10141 <= p1_ne_10141;
    p2_or_10151 <= p1_or_10151;
    p2_or_10154 <= p1_or_10154;
    p2_bit_slice_10425 <= p2_bit_slice_10425_comb;
    p2_or_10161 <= p1_or_10161;
    p2_ne_10427 <= p2_ne_10427_comb;
    p2_or_10169 <= p1_or_10169;
    p2_or_10175 <= p1_or_10175;
    p2_or_10241 <= p1_or_10241;
    p2_nor_10242 <= p1_nor_10242;
    p2_and_10306 <= p1_and_10306;
    p2_Code_list <= p2_Code_list_comb;
    p2_code_list <= p2_code_list_comb;
  end

  // ===== Pipe stage 3:
  wire [2:0] p3_huff_length_squeezed__17_comb;
  wire [3:0] p3_huff_length_squeezed__2_comb;
  wire [3:0] p3_huff_length_squeezed__19_comb;
  wire [3:0] p3_sel_10510_comb;
  wire [3:0] p3_sel_10535_comb;
  wire [3:0] p3_huff_code__1_squeezed_comb;
  wire [2:0] p3_sel_10518_comb;
  wire [3:0] p3_huff_code__1_squeezed__2_comb;
  wire [3:0] p3_huff_code__1_squeezed__1_comb;
  wire [3:0] p3_sel_10528_comb;
  wire [3:0] p3_sign_ext_10529_comb;
  wire [3:0] p3_sel_10530_comb;
  wire [3:0] p3_next_pix_comb;
  assign p3_huff_length_squeezed__17_comb = 3'h4;
  assign p3_huff_length_squeezed__2_comb = 4'h4;
  assign p3_huff_length_squeezed__19_comb = 4'h4;
  assign p3_sel_10510_comb = p2_or_10104 ? p3_huff_length_squeezed__19_comb : (p2_or_10087 ? 4'h5 : (p2_or_10070 ? 4'h6 : (p2_or_10055 ? 4'h7 : {1'h1, p2_and_10401})));
  assign p3_sel_10535_comb = p2_or_10175 ? 4'h2 : (p2_or_10169 ? 4'h3 : (p2_or_10161 ? p3_huff_length_squeezed__2_comb : (p2_or_10151 ? 4'h5 : (p2_or_10135 ? 4'h6 : p2_sel_10424))));
  assign p3_huff_code__1_squeezed_comb = 4'h1;
  assign p3_sel_10518_comb = p2_or_reduce_10423 ? 3'h7 : (p2_or_reduce_10420 ? 3'h6 : (p2_or_reduce_10416 ? 3'h5 : (p2_or_reduce_10412 ? p3_huff_length_squeezed__17_comb : {1'h0, p2_sel_10408})));
  assign p3_huff_code__1_squeezed__2_comb = 4'h1;
  assign p3_huff_code__1_squeezed__1_comb = 4'h1;
  assign p3_sel_10528_comb = p2_or_10154 ? p3_huff_code__1_squeezed__2_comb : (p2_or_10139 ? 4'h2 : (p2_or_10122 ? 4'h3 : p3_sel_10510_comb));
  assign p3_sign_ext_10529_comb = {4{~(p2_eq_10140 | p2_ne_10141)}};
  assign p3_sel_10530_comb = p2_bit_slice_10425 ? 4'h8 : {1'h0, p3_sel_10518_comb};
  assign p3_next_pix_comb = ((p2_or_10241 ? p3_huff_code__1_squeezed_comb : p3_sel_10535_comb) & {4{p2_nor_10242}}) + p3_huff_code__1_squeezed__1_comb;

  // Registers for pipe stage 3:
  reg p3_is_luminance;
  reg p3_eq_10140;
  reg p3_ne_10141;
  reg [3:0] p3_sel_10528;
  reg [3:0] p3_sign_ext_10529;
  reg [3:0] p3_sel_10530;
  reg p3_ne_10427;
  reg p3_and_10306;
  reg [7:0] p3_Code_list;
  reg [3:0] p3_next_pix;
  reg [7:0] p3_code_list;
  always @ (posedge clk) begin
    p3_is_luminance <= p2_is_luminance;
    p3_eq_10140 <= p2_eq_10140;
    p3_ne_10141 <= p2_ne_10141;
    p3_sel_10528 <= p3_sel_10528_comb;
    p3_sign_ext_10529 <= p3_sign_ext_10529_comb;
    p3_sel_10530 <= p3_sel_10530_comb;
    p3_ne_10427 <= p2_ne_10427;
    p3_and_10306 <= p2_and_10306;
    p3_Code_list <= p2_Code_list;
    p3_next_pix <= p3_next_pix_comb;
    p3_code_list <= p2_code_list;
  end

  // ===== Pipe stage 4:
  wire [3:0] p4_run_comb;
  wire [7:0] p4_Code_size_comb;
  wire [2:0] p4_huff_code__1_squeezed_squeezed__18_comb;
  wire [2:0] p4_huff_length_squeezed__18_comb;
  wire [7:0] p4_run_size_str_u8_comb;
  wire [1:0] p4_huff_length__1_squeezed__4_comb;
  wire [1:0] p4_huff_length__1_squeezed__5_comb;
  wire p4_eq_10579_comb;
  wire [2:0] p4_sel_10582_comb;
  wire [3:0] p4_Code_size_squeezed_comb;
  wire [3:0] p4_huff_length_squeezed__20_comb;
  wire p4_or_10596_comb;
  wire [4:0] p4_Huffman_length_squeezed_comb;
  wire [15:0] p4_Huffman_code_full_comb;
  wire [47:0] p4_tuple_10622_comb;
  assign p4_run_comb = p3_sel_10528 & p3_sign_ext_10529;
  assign p4_Code_size_comb = {4'h0, p3_sel_10530} & {8{p3_ne_10427}};
  assign p4_huff_code__1_squeezed_squeezed__18_comb = 3'h1;
  assign p4_huff_length_squeezed__18_comb = 3'h4;
  assign p4_run_size_str_u8_comb = {p4_run_comb, 4'h0} | p4_Code_size_comb;
  assign p4_huff_length__1_squeezed__4_comb = 2'h1;
  assign p4_huff_length__1_squeezed__5_comb = 2'h2;
  assign p4_eq_10579_comb = p4_run_comb == 4'hf;
  assign p4_sel_10582_comb = p3_is_luminance ? p4_huff_length_squeezed__18_comb : p4_huff_code__1_squeezed_squeezed__18_comb;
  assign p4_Code_size_squeezed_comb = p4_Code_size_comb[3:0];
  assign p4_huff_length_squeezed__20_comb = 4'h4;
  assign p4_or_10596_comb = p3_and_10306 | p4_eq_10579_comb;
  assign p4_Huffman_length_squeezed_comb = p3_is_luminance ? literal_10576[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_10574[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_Huffman_code_full_comb = p3_is_luminance ? literal_10581[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_10580[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_tuple_10622_comb = {p4_or_10596_comb ? {12'h000, {{1{p4_sel_10582_comb[2]}}, p4_sel_10582_comb}} : p4_Huffman_code_full_comb, {3'h0, p4_or_10596_comb ? {2'h0, p3_is_luminance ? p4_huff_length__1_squeezed__5_comb : p4_huff_length__1_squeezed__4_comb, 1'h0} : p4_Huffman_length_squeezed_comb}, p3_and_10306 ? p3_code_list : p3_Code_list & {8{~p4_eq_10579_comb}}, {4'h0, p4_eq_10579_comb ? p4_huff_length_squeezed__20_comb : p4_Code_size_squeezed_comb} & {8{~p3_and_10306}}, p3_and_10306 ? 4'hf : p3_sel_10528 & {4{~(p4_eq_10579_comb | p3_eq_10140 | p3_ne_10141)}}, p3_and_10306 ? 4'hf : p3_next_pix & {4{~p4_eq_10579_comb}}};

  // Registers for pipe stage 4:
  reg [47:0] p4_tuple_10622;
  always @ (posedge clk) begin
    p4_tuple_10622 <= p4_tuple_10622_comb;
  end
  assign out = p4_tuple_10622;
endmodule
