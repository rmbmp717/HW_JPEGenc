module Data_flip64(
  input wire clk,
  input wire [639:0] data_in,
  input wire is_flip,
  output wire [639:0] out
);
  wire [9:0] data_in_unflattened[0:63];
  assign data_in_unflattened[0] = data_in[9:0];
  assign data_in_unflattened[1] = data_in[19:10];
  assign data_in_unflattened[2] = data_in[29:20];
  assign data_in_unflattened[3] = data_in[39:30];
  assign data_in_unflattened[4] = data_in[49:40];
  assign data_in_unflattened[5] = data_in[59:50];
  assign data_in_unflattened[6] = data_in[69:60];
  assign data_in_unflattened[7] = data_in[79:70];
  assign data_in_unflattened[8] = data_in[89:80];
  assign data_in_unflattened[9] = data_in[99:90];
  assign data_in_unflattened[10] = data_in[109:100];
  assign data_in_unflattened[11] = data_in[119:110];
  assign data_in_unflattened[12] = data_in[129:120];
  assign data_in_unflattened[13] = data_in[139:130];
  assign data_in_unflattened[14] = data_in[149:140];
  assign data_in_unflattened[15] = data_in[159:150];
  assign data_in_unflattened[16] = data_in[169:160];
  assign data_in_unflattened[17] = data_in[179:170];
  assign data_in_unflattened[18] = data_in[189:180];
  assign data_in_unflattened[19] = data_in[199:190];
  assign data_in_unflattened[20] = data_in[209:200];
  assign data_in_unflattened[21] = data_in[219:210];
  assign data_in_unflattened[22] = data_in[229:220];
  assign data_in_unflattened[23] = data_in[239:230];
  assign data_in_unflattened[24] = data_in[249:240];
  assign data_in_unflattened[25] = data_in[259:250];
  assign data_in_unflattened[26] = data_in[269:260];
  assign data_in_unflattened[27] = data_in[279:270];
  assign data_in_unflattened[28] = data_in[289:280];
  assign data_in_unflattened[29] = data_in[299:290];
  assign data_in_unflattened[30] = data_in[309:300];
  assign data_in_unflattened[31] = data_in[319:310];
  assign data_in_unflattened[32] = data_in[329:320];
  assign data_in_unflattened[33] = data_in[339:330];
  assign data_in_unflattened[34] = data_in[349:340];
  assign data_in_unflattened[35] = data_in[359:350];
  assign data_in_unflattened[36] = data_in[369:360];
  assign data_in_unflattened[37] = data_in[379:370];
  assign data_in_unflattened[38] = data_in[389:380];
  assign data_in_unflattened[39] = data_in[399:390];
  assign data_in_unflattened[40] = data_in[409:400];
  assign data_in_unflattened[41] = data_in[419:410];
  assign data_in_unflattened[42] = data_in[429:420];
  assign data_in_unflattened[43] = data_in[439:430];
  assign data_in_unflattened[44] = data_in[449:440];
  assign data_in_unflattened[45] = data_in[459:450];
  assign data_in_unflattened[46] = data_in[469:460];
  assign data_in_unflattened[47] = data_in[479:470];
  assign data_in_unflattened[48] = data_in[489:480];
  assign data_in_unflattened[49] = data_in[499:490];
  assign data_in_unflattened[50] = data_in[509:500];
  assign data_in_unflattened[51] = data_in[519:510];
  assign data_in_unflattened[52] = data_in[529:520];
  assign data_in_unflattened[53] = data_in[539:530];
  assign data_in_unflattened[54] = data_in[549:540];
  assign data_in_unflattened[55] = data_in[559:550];
  assign data_in_unflattened[56] = data_in[569:560];
  assign data_in_unflattened[57] = data_in[579:570];
  assign data_in_unflattened[58] = data_in[589:580];
  assign data_in_unflattened[59] = data_in[599:590];
  assign data_in_unflattened[60] = data_in[609:600];
  assign data_in_unflattened[61] = data_in[619:610];
  assign data_in_unflattened[62] = data_in[629:620];
  assign data_in_unflattened[63] = data_in[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_data_in[0:63];
  reg p0_is_flip;
  always @ (posedge clk) begin
    p0_data_in[0] <= data_in_unflattened[0];
    p0_data_in[1] <= data_in_unflattened[1];
    p0_data_in[2] <= data_in_unflattened[2];
    p0_data_in[3] <= data_in_unflattened[3];
    p0_data_in[4] <= data_in_unflattened[4];
    p0_data_in[5] <= data_in_unflattened[5];
    p0_data_in[6] <= data_in_unflattened[6];
    p0_data_in[7] <= data_in_unflattened[7];
    p0_data_in[8] <= data_in_unflattened[8];
    p0_data_in[9] <= data_in_unflattened[9];
    p0_data_in[10] <= data_in_unflattened[10];
    p0_data_in[11] <= data_in_unflattened[11];
    p0_data_in[12] <= data_in_unflattened[12];
    p0_data_in[13] <= data_in_unflattened[13];
    p0_data_in[14] <= data_in_unflattened[14];
    p0_data_in[15] <= data_in_unflattened[15];
    p0_data_in[16] <= data_in_unflattened[16];
    p0_data_in[17] <= data_in_unflattened[17];
    p0_data_in[18] <= data_in_unflattened[18];
    p0_data_in[19] <= data_in_unflattened[19];
    p0_data_in[20] <= data_in_unflattened[20];
    p0_data_in[21] <= data_in_unflattened[21];
    p0_data_in[22] <= data_in_unflattened[22];
    p0_data_in[23] <= data_in_unflattened[23];
    p0_data_in[24] <= data_in_unflattened[24];
    p0_data_in[25] <= data_in_unflattened[25];
    p0_data_in[26] <= data_in_unflattened[26];
    p0_data_in[27] <= data_in_unflattened[27];
    p0_data_in[28] <= data_in_unflattened[28];
    p0_data_in[29] <= data_in_unflattened[29];
    p0_data_in[30] <= data_in_unflattened[30];
    p0_data_in[31] <= data_in_unflattened[31];
    p0_data_in[32] <= data_in_unflattened[32];
    p0_data_in[33] <= data_in_unflattened[33];
    p0_data_in[34] <= data_in_unflattened[34];
    p0_data_in[35] <= data_in_unflattened[35];
    p0_data_in[36] <= data_in_unflattened[36];
    p0_data_in[37] <= data_in_unflattened[37];
    p0_data_in[38] <= data_in_unflattened[38];
    p0_data_in[39] <= data_in_unflattened[39];
    p0_data_in[40] <= data_in_unflattened[40];
    p0_data_in[41] <= data_in_unflattened[41];
    p0_data_in[42] <= data_in_unflattened[42];
    p0_data_in[43] <= data_in_unflattened[43];
    p0_data_in[44] <= data_in_unflattened[44];
    p0_data_in[45] <= data_in_unflattened[45];
    p0_data_in[46] <= data_in_unflattened[46];
    p0_data_in[47] <= data_in_unflattened[47];
    p0_data_in[48] <= data_in_unflattened[48];
    p0_data_in[49] <= data_in_unflattened[49];
    p0_data_in[50] <= data_in_unflattened[50];
    p0_data_in[51] <= data_in_unflattened[51];
    p0_data_in[52] <= data_in_unflattened[52];
    p0_data_in[53] <= data_in_unflattened[53];
    p0_data_in[54] <= data_in_unflattened[54];
    p0_data_in[55] <= data_in_unflattened[55];
    p0_data_in[56] <= data_in_unflattened[56];
    p0_data_in[57] <= data_in_unflattened[57];
    p0_data_in[58] <= data_in_unflattened[58];
    p0_data_in[59] <= data_in_unflattened[59];
    p0_data_in[60] <= data_in_unflattened[60];
    p0_data_in[61] <= data_in_unflattened[61];
    p0_data_in[62] <= data_in_unflattened[62];
    p0_data_in[63] <= data_in_unflattened[63];
    p0_is_flip <= is_flip;
  end

  // ===== Pipe stage 1:
  wire [1:0] p1_src_index__65_squeezed_comb;
  wire [2:0] p1_src_index__66_squeezed_comb;
  wire [2:0] p1_src_index__67_squeezed_comb;
  wire [3:0] p1_src_index__68_squeezed_comb;
  wire [3:0] p1_src_index__69_squeezed_comb;
  wire [3:0] p1_src_index__70_squeezed_comb;
  wire [3:0] p1_src_index__71_squeezed_comb;
  wire [4:0] p1_src_index__72_squeezed_comb;
  wire [4:0] p1_src_index__73_squeezed_comb;
  wire [4:0] p1_src_index__74_squeezed_comb;
  wire [4:0] p1_src_index__75_squeezed_comb;
  wire [4:0] p1_src_index__76_squeezed_comb;
  wire [4:0] p1_src_index__77_squeezed_comb;
  wire [4:0] p1_src_index__78_squeezed_comb;
  wire [4:0] p1_src_index__79_squeezed_comb;
  wire [4:0] p1_src_index__112_squeezed_comb;
  wire [4:0] p1_src_index__113_squeezed_comb;
  wire [4:0] p1_src_index__114_squeezed_comb;
  wire [4:0] p1_src_index__115_squeezed_comb;
  wire [4:0] p1_src_index__116_squeezed_comb;
  wire [4:0] p1_src_index__117_squeezed_comb;
  wire [4:0] p1_src_index__118_squeezed_comb;
  wire [4:0] p1_src_index__119_squeezed_comb;
  wire [3:0] p1_src_index__120_squeezed_comb;
  wire [3:0] p1_src_index__121_squeezed_comb;
  wire [3:0] p1_src_index__122_squeezed_comb;
  wire [3:0] p1_src_index__123_squeezed_comb;
  wire [2:0] p1_src_index__124_squeezed_comb;
  wire [2:0] p1_src_index__125_squeezed_comb;
  wire [1:0] p1_src_index__126_squeezed_comb;
  wire [5:0] p1_src_index__64_comb;
  wire [5:0] p1_src_index__65_comb;
  wire [5:0] p1_src_index__66_comb;
  wire [5:0] p1_src_index__67_comb;
  wire [5:0] p1_src_index__68_comb;
  wire [5:0] p1_src_index__69_comb;
  wire [5:0] p1_src_index__70_comb;
  wire [5:0] p1_src_index__71_comb;
  wire [5:0] p1_src_index__72_comb;
  wire [5:0] p1_src_index__73_comb;
  wire [5:0] p1_src_index__74_comb;
  wire [5:0] p1_src_index__75_comb;
  wire [5:0] p1_src_index__76_comb;
  wire [5:0] p1_src_index__77_comb;
  wire [5:0] p1_src_index__78_comb;
  wire [5:0] p1_src_index__79_comb;
  wire [5:0] p1_src_index__80_comb;
  wire [5:0] p1_src_index__81_comb;
  wire [5:0] p1_src_index__82_comb;
  wire [5:0] p1_src_index__83_comb;
  wire [5:0] p1_src_index__84_comb;
  wire [5:0] p1_src_index__85_comb;
  wire [5:0] p1_src_index__86_comb;
  wire [5:0] p1_src_index__87_comb;
  wire [5:0] p1_src_index__88_comb;
  wire [5:0] p1_src_index__89_comb;
  wire [5:0] p1_src_index__90_comb;
  wire [5:0] p1_src_index__91_comb;
  wire [5:0] p1_src_index__92_comb;
  wire [5:0] p1_src_index__93_comb;
  wire [5:0] p1_src_index__94_comb;
  wire [5:0] p1_src_index__95_comb;
  wire [5:0] p1_src_index__96_comb;
  wire [5:0] p1_src_index__97_comb;
  wire [5:0] p1_src_index__98_comb;
  wire [5:0] p1_src_index__99_comb;
  wire [5:0] p1_src_index__100_comb;
  wire [5:0] p1_src_index__101_comb;
  wire [5:0] p1_src_index__102_comb;
  wire [5:0] p1_src_index__103_comb;
  wire [5:0] p1_src_index__104_comb;
  wire [5:0] p1_src_index__105_comb;
  wire [5:0] p1_src_index__106_comb;
  wire [5:0] p1_src_index__107_comb;
  wire [5:0] p1_src_index__108_comb;
  wire [5:0] p1_src_index__109_comb;
  wire [5:0] p1_src_index__110_comb;
  wire [5:0] p1_src_index__111_comb;
  wire [5:0] p1_src_index__112_comb;
  wire [5:0] p1_src_index__113_comb;
  wire [5:0] p1_src_index__114_comb;
  wire [5:0] p1_src_index__115_comb;
  wire [5:0] p1_src_index__116_comb;
  wire [5:0] p1_src_index__117_comb;
  wire [5:0] p1_src_index__118_comb;
  wire [5:0] p1_src_index__119_comb;
  wire [5:0] p1_src_index__120_comb;
  wire [5:0] p1_src_index__121_comb;
  wire [5:0] p1_src_index__122_comb;
  wire [5:0] p1_src_index__123_comb;
  wire [5:0] p1_src_index__124_comb;
  wire [5:0] p1_src_index__125_comb;
  wire [5:0] p1_src_index__126_comb;
  wire [5:0] p1_src_index__127_comb;
  wire [9:0] p1_result_comb[0:63];
  assign p1_src_index__65_squeezed_comb = p0_is_flip ? 2'h2 : 2'h1;
  assign p1_src_index__66_squeezed_comb = p0_is_flip ? 3'h5 : 3'h2;
  assign p1_src_index__67_squeezed_comb = p0_is_flip ? 3'h4 : 3'h3;
  assign p1_src_index__68_squeezed_comb = p0_is_flip ? 4'hb : 4'h4;
  assign p1_src_index__69_squeezed_comb = p0_is_flip ? 4'ha : 4'h5;
  assign p1_src_index__70_squeezed_comb = p0_is_flip ? 4'h9 : 4'h6;
  assign p1_src_index__71_squeezed_comb = p0_is_flip ? 4'h8 : 4'h7;
  assign p1_src_index__72_squeezed_comb = p0_is_flip ? 5'h17 : 5'h08;
  assign p1_src_index__73_squeezed_comb = p0_is_flip ? 5'h16 : 5'h09;
  assign p1_src_index__74_squeezed_comb = p0_is_flip ? 5'h15 : 5'h0a;
  assign p1_src_index__75_squeezed_comb = p0_is_flip ? 5'h14 : 5'h0b;
  assign p1_src_index__76_squeezed_comb = p0_is_flip ? 5'h13 : 5'h0c;
  assign p1_src_index__77_squeezed_comb = p0_is_flip ? 5'h12 : 5'h0d;
  assign p1_src_index__78_squeezed_comb = p0_is_flip ? 5'h11 : 5'h0e;
  assign p1_src_index__79_squeezed_comb = p0_is_flip ? 5'h10 : 5'h0f;
  assign p1_src_index__112_squeezed_comb = p0_is_flip ? 5'h0f : 5'h10;
  assign p1_src_index__113_squeezed_comb = p0_is_flip ? 5'h0e : 5'h11;
  assign p1_src_index__114_squeezed_comb = p0_is_flip ? 5'h0d : 5'h12;
  assign p1_src_index__115_squeezed_comb = p0_is_flip ? 5'h0c : 5'h13;
  assign p1_src_index__116_squeezed_comb = p0_is_flip ? 5'h0b : 5'h14;
  assign p1_src_index__117_squeezed_comb = p0_is_flip ? 5'h0a : 5'h15;
  assign p1_src_index__118_squeezed_comb = p0_is_flip ? 5'h09 : 5'h16;
  assign p1_src_index__119_squeezed_comb = p0_is_flip ? 5'h08 : 5'h17;
  assign p1_src_index__120_squeezed_comb = p0_is_flip ? 4'h7 : 4'h8;
  assign p1_src_index__121_squeezed_comb = p0_is_flip ? 4'h6 : 4'h9;
  assign p1_src_index__122_squeezed_comb = p0_is_flip ? 4'h5 : 4'ha;
  assign p1_src_index__123_squeezed_comb = p0_is_flip ? 4'h4 : 4'hb;
  assign p1_src_index__124_squeezed_comb = p0_is_flip ? 3'h3 : 3'h4;
  assign p1_src_index__125_squeezed_comb = p0_is_flip ? 3'h2 : 3'h5;
  assign p1_src_index__126_squeezed_comb = p0_is_flip ? 2'h1 : 2'h2;
  assign p1_src_index__64_comb = {6{p0_is_flip}};
  assign p1_src_index__65_comb = {{4{p1_src_index__65_squeezed_comb[1]}}, p1_src_index__65_squeezed_comb};
  assign p1_src_index__66_comb = {{3{p1_src_index__66_squeezed_comb[2]}}, p1_src_index__66_squeezed_comb};
  assign p1_src_index__67_comb = {{3{p1_src_index__67_squeezed_comb[2]}}, p1_src_index__67_squeezed_comb};
  assign p1_src_index__68_comb = {{2{p1_src_index__68_squeezed_comb[3]}}, p1_src_index__68_squeezed_comb};
  assign p1_src_index__69_comb = {{2{p1_src_index__69_squeezed_comb[3]}}, p1_src_index__69_squeezed_comb};
  assign p1_src_index__70_comb = {{2{p1_src_index__70_squeezed_comb[3]}}, p1_src_index__70_squeezed_comb};
  assign p1_src_index__71_comb = {{2{p1_src_index__71_squeezed_comb[3]}}, p1_src_index__71_squeezed_comb};
  assign p1_src_index__72_comb = {{1{p1_src_index__72_squeezed_comb[4]}}, p1_src_index__72_squeezed_comb};
  assign p1_src_index__73_comb = {{1{p1_src_index__73_squeezed_comb[4]}}, p1_src_index__73_squeezed_comb};
  assign p1_src_index__74_comb = {{1{p1_src_index__74_squeezed_comb[4]}}, p1_src_index__74_squeezed_comb};
  assign p1_src_index__75_comb = {{1{p1_src_index__75_squeezed_comb[4]}}, p1_src_index__75_squeezed_comb};
  assign p1_src_index__76_comb = {{1{p1_src_index__76_squeezed_comb[4]}}, p1_src_index__76_squeezed_comb};
  assign p1_src_index__77_comb = {{1{p1_src_index__77_squeezed_comb[4]}}, p1_src_index__77_squeezed_comb};
  assign p1_src_index__78_comb = {{1{p1_src_index__78_squeezed_comb[4]}}, p1_src_index__78_squeezed_comb};
  assign p1_src_index__79_comb = {{1{p1_src_index__79_squeezed_comb[4]}}, p1_src_index__79_squeezed_comb};
  assign p1_src_index__80_comb = p0_is_flip ? 6'h2f : 6'h10;
  assign p1_src_index__81_comb = p0_is_flip ? 6'h2e : 6'h11;
  assign p1_src_index__82_comb = p0_is_flip ? 6'h2d : 6'h12;
  assign p1_src_index__83_comb = p0_is_flip ? 6'h2c : 6'h13;
  assign p1_src_index__84_comb = p0_is_flip ? 6'h2b : 6'h14;
  assign p1_src_index__85_comb = p0_is_flip ? 6'h2a : 6'h15;
  assign p1_src_index__86_comb = p0_is_flip ? 6'h29 : 6'h16;
  assign p1_src_index__87_comb = p0_is_flip ? 6'h28 : 6'h17;
  assign p1_src_index__88_comb = p0_is_flip ? 6'h27 : 6'h18;
  assign p1_src_index__89_comb = p0_is_flip ? 6'h26 : 6'h19;
  assign p1_src_index__90_comb = p0_is_flip ? 6'h25 : 6'h1a;
  assign p1_src_index__91_comb = p0_is_flip ? 6'h24 : 6'h1b;
  assign p1_src_index__92_comb = p0_is_flip ? 6'h23 : 6'h1c;
  assign p1_src_index__93_comb = p0_is_flip ? 6'h22 : 6'h1d;
  assign p1_src_index__94_comb = p0_is_flip ? 6'h21 : 6'h1e;
  assign p1_src_index__95_comb = p0_is_flip ? 6'h20 : 6'h1f;
  assign p1_src_index__96_comb = p0_is_flip ? 6'h1f : 6'h20;
  assign p1_src_index__97_comb = p0_is_flip ? 6'h1e : 6'h21;
  assign p1_src_index__98_comb = p0_is_flip ? 6'h1d : 6'h22;
  assign p1_src_index__99_comb = p0_is_flip ? 6'h1c : 6'h23;
  assign p1_src_index__100_comb = p0_is_flip ? 6'h1b : 6'h24;
  assign p1_src_index__101_comb = p0_is_flip ? 6'h1a : 6'h25;
  assign p1_src_index__102_comb = p0_is_flip ? 6'h19 : 6'h26;
  assign p1_src_index__103_comb = p0_is_flip ? 6'h18 : 6'h27;
  assign p1_src_index__104_comb = p0_is_flip ? 6'h17 : 6'h28;
  assign p1_src_index__105_comb = p0_is_flip ? 6'h16 : 6'h29;
  assign p1_src_index__106_comb = p0_is_flip ? 6'h15 : 6'h2a;
  assign p1_src_index__107_comb = p0_is_flip ? 6'h14 : 6'h2b;
  assign p1_src_index__108_comb = p0_is_flip ? 6'h13 : 6'h2c;
  assign p1_src_index__109_comb = p0_is_flip ? 6'h12 : 6'h2d;
  assign p1_src_index__110_comb = p0_is_flip ? 6'h11 : 6'h2e;
  assign p1_src_index__111_comb = p0_is_flip ? 6'h10 : 6'h2f;
  assign p1_src_index__112_comb = {{1{p1_src_index__112_squeezed_comb[4]}}, p1_src_index__112_squeezed_comb};
  assign p1_src_index__113_comb = {{1{p1_src_index__113_squeezed_comb[4]}}, p1_src_index__113_squeezed_comb};
  assign p1_src_index__114_comb = {{1{p1_src_index__114_squeezed_comb[4]}}, p1_src_index__114_squeezed_comb};
  assign p1_src_index__115_comb = {{1{p1_src_index__115_squeezed_comb[4]}}, p1_src_index__115_squeezed_comb};
  assign p1_src_index__116_comb = {{1{p1_src_index__116_squeezed_comb[4]}}, p1_src_index__116_squeezed_comb};
  assign p1_src_index__117_comb = {{1{p1_src_index__117_squeezed_comb[4]}}, p1_src_index__117_squeezed_comb};
  assign p1_src_index__118_comb = {{1{p1_src_index__118_squeezed_comb[4]}}, p1_src_index__118_squeezed_comb};
  assign p1_src_index__119_comb = {{1{p1_src_index__119_squeezed_comb[4]}}, p1_src_index__119_squeezed_comb};
  assign p1_src_index__120_comb = {{2{p1_src_index__120_squeezed_comb[3]}}, p1_src_index__120_squeezed_comb};
  assign p1_src_index__121_comb = {{2{p1_src_index__121_squeezed_comb[3]}}, p1_src_index__121_squeezed_comb};
  assign p1_src_index__122_comb = {{2{p1_src_index__122_squeezed_comb[3]}}, p1_src_index__122_squeezed_comb};
  assign p1_src_index__123_comb = {{2{p1_src_index__123_squeezed_comb[3]}}, p1_src_index__123_squeezed_comb};
  assign p1_src_index__124_comb = {{3{p1_src_index__124_squeezed_comb[2]}}, p1_src_index__124_squeezed_comb};
  assign p1_src_index__125_comb = {{3{p1_src_index__125_squeezed_comb[2]}}, p1_src_index__125_squeezed_comb};
  assign p1_src_index__126_comb = {{4{p1_src_index__126_squeezed_comb[1]}}, p1_src_index__126_squeezed_comb};
  assign p1_src_index__127_comb = {6{~p0_is_flip}};
  assign p1_result_comb[0] = p0_data_in[p1_src_index__64_comb];
  assign p1_result_comb[1] = p0_data_in[p1_src_index__65_comb];
  assign p1_result_comb[2] = p0_data_in[p1_src_index__66_comb];
  assign p1_result_comb[3] = p0_data_in[p1_src_index__67_comb];
  assign p1_result_comb[4] = p0_data_in[p1_src_index__68_comb];
  assign p1_result_comb[5] = p0_data_in[p1_src_index__69_comb];
  assign p1_result_comb[6] = p0_data_in[p1_src_index__70_comb];
  assign p1_result_comb[7] = p0_data_in[p1_src_index__71_comb];
  assign p1_result_comb[8] = p0_data_in[p1_src_index__72_comb];
  assign p1_result_comb[9] = p0_data_in[p1_src_index__73_comb];
  assign p1_result_comb[10] = p0_data_in[p1_src_index__74_comb];
  assign p1_result_comb[11] = p0_data_in[p1_src_index__75_comb];
  assign p1_result_comb[12] = p0_data_in[p1_src_index__76_comb];
  assign p1_result_comb[13] = p0_data_in[p1_src_index__77_comb];
  assign p1_result_comb[14] = p0_data_in[p1_src_index__78_comb];
  assign p1_result_comb[15] = p0_data_in[p1_src_index__79_comb];
  assign p1_result_comb[16] = p0_data_in[p1_src_index__80_comb];
  assign p1_result_comb[17] = p0_data_in[p1_src_index__81_comb];
  assign p1_result_comb[18] = p0_data_in[p1_src_index__82_comb];
  assign p1_result_comb[19] = p0_data_in[p1_src_index__83_comb];
  assign p1_result_comb[20] = p0_data_in[p1_src_index__84_comb];
  assign p1_result_comb[21] = p0_data_in[p1_src_index__85_comb];
  assign p1_result_comb[22] = p0_data_in[p1_src_index__86_comb];
  assign p1_result_comb[23] = p0_data_in[p1_src_index__87_comb];
  assign p1_result_comb[24] = p0_data_in[p1_src_index__88_comb];
  assign p1_result_comb[25] = p0_data_in[p1_src_index__89_comb];
  assign p1_result_comb[26] = p0_data_in[p1_src_index__90_comb];
  assign p1_result_comb[27] = p0_data_in[p1_src_index__91_comb];
  assign p1_result_comb[28] = p0_data_in[p1_src_index__92_comb];
  assign p1_result_comb[29] = p0_data_in[p1_src_index__93_comb];
  assign p1_result_comb[30] = p0_data_in[p1_src_index__94_comb];
  assign p1_result_comb[31] = p0_data_in[p1_src_index__95_comb];
  assign p1_result_comb[32] = p0_data_in[p1_src_index__96_comb];
  assign p1_result_comb[33] = p0_data_in[p1_src_index__97_comb];
  assign p1_result_comb[34] = p0_data_in[p1_src_index__98_comb];
  assign p1_result_comb[35] = p0_data_in[p1_src_index__99_comb];
  assign p1_result_comb[36] = p0_data_in[p1_src_index__100_comb];
  assign p1_result_comb[37] = p0_data_in[p1_src_index__101_comb];
  assign p1_result_comb[38] = p0_data_in[p1_src_index__102_comb];
  assign p1_result_comb[39] = p0_data_in[p1_src_index__103_comb];
  assign p1_result_comb[40] = p0_data_in[p1_src_index__104_comb];
  assign p1_result_comb[41] = p0_data_in[p1_src_index__105_comb];
  assign p1_result_comb[42] = p0_data_in[p1_src_index__106_comb];
  assign p1_result_comb[43] = p0_data_in[p1_src_index__107_comb];
  assign p1_result_comb[44] = p0_data_in[p1_src_index__108_comb];
  assign p1_result_comb[45] = p0_data_in[p1_src_index__109_comb];
  assign p1_result_comb[46] = p0_data_in[p1_src_index__110_comb];
  assign p1_result_comb[47] = p0_data_in[p1_src_index__111_comb];
  assign p1_result_comb[48] = p0_data_in[p1_src_index__112_comb];
  assign p1_result_comb[49] = p0_data_in[p1_src_index__113_comb];
  assign p1_result_comb[50] = p0_data_in[p1_src_index__114_comb];
  assign p1_result_comb[51] = p0_data_in[p1_src_index__115_comb];
  assign p1_result_comb[52] = p0_data_in[p1_src_index__116_comb];
  assign p1_result_comb[53] = p0_data_in[p1_src_index__117_comb];
  assign p1_result_comb[54] = p0_data_in[p1_src_index__118_comb];
  assign p1_result_comb[55] = p0_data_in[p1_src_index__119_comb];
  assign p1_result_comb[56] = p0_data_in[p1_src_index__120_comb];
  assign p1_result_comb[57] = p0_data_in[p1_src_index__121_comb];
  assign p1_result_comb[58] = p0_data_in[p1_src_index__122_comb];
  assign p1_result_comb[59] = p0_data_in[p1_src_index__123_comb];
  assign p1_result_comb[60] = p0_data_in[p1_src_index__124_comb];
  assign p1_result_comb[61] = p0_data_in[p1_src_index__125_comb];
  assign p1_result_comb[62] = p0_data_in[p1_src_index__126_comb];
  assign p1_result_comb[63] = p0_data_in[p1_src_index__127_comb];

  // Registers for pipe stage 1:
  reg [9:0] p1_result[0:63];
  always @ (posedge clk) begin
    p1_result[0] <= p1_result_comb[0];
    p1_result[1] <= p1_result_comb[1];
    p1_result[2] <= p1_result_comb[2];
    p1_result[3] <= p1_result_comb[3];
    p1_result[4] <= p1_result_comb[4];
    p1_result[5] <= p1_result_comb[5];
    p1_result[6] <= p1_result_comb[6];
    p1_result[7] <= p1_result_comb[7];
    p1_result[8] <= p1_result_comb[8];
    p1_result[9] <= p1_result_comb[9];
    p1_result[10] <= p1_result_comb[10];
    p1_result[11] <= p1_result_comb[11];
    p1_result[12] <= p1_result_comb[12];
    p1_result[13] <= p1_result_comb[13];
    p1_result[14] <= p1_result_comb[14];
    p1_result[15] <= p1_result_comb[15];
    p1_result[16] <= p1_result_comb[16];
    p1_result[17] <= p1_result_comb[17];
    p1_result[18] <= p1_result_comb[18];
    p1_result[19] <= p1_result_comb[19];
    p1_result[20] <= p1_result_comb[20];
    p1_result[21] <= p1_result_comb[21];
    p1_result[22] <= p1_result_comb[22];
    p1_result[23] <= p1_result_comb[23];
    p1_result[24] <= p1_result_comb[24];
    p1_result[25] <= p1_result_comb[25];
    p1_result[26] <= p1_result_comb[26];
    p1_result[27] <= p1_result_comb[27];
    p1_result[28] <= p1_result_comb[28];
    p1_result[29] <= p1_result_comb[29];
    p1_result[30] <= p1_result_comb[30];
    p1_result[31] <= p1_result_comb[31];
    p1_result[32] <= p1_result_comb[32];
    p1_result[33] <= p1_result_comb[33];
    p1_result[34] <= p1_result_comb[34];
    p1_result[35] <= p1_result_comb[35];
    p1_result[36] <= p1_result_comb[36];
    p1_result[37] <= p1_result_comb[37];
    p1_result[38] <= p1_result_comb[38];
    p1_result[39] <= p1_result_comb[39];
    p1_result[40] <= p1_result_comb[40];
    p1_result[41] <= p1_result_comb[41];
    p1_result[42] <= p1_result_comb[42];
    p1_result[43] <= p1_result_comb[43];
    p1_result[44] <= p1_result_comb[44];
    p1_result[45] <= p1_result_comb[45];
    p1_result[46] <= p1_result_comb[46];
    p1_result[47] <= p1_result_comb[47];
    p1_result[48] <= p1_result_comb[48];
    p1_result[49] <= p1_result_comb[49];
    p1_result[50] <= p1_result_comb[50];
    p1_result[51] <= p1_result_comb[51];
    p1_result[52] <= p1_result_comb[52];
    p1_result[53] <= p1_result_comb[53];
    p1_result[54] <= p1_result_comb[54];
    p1_result[55] <= p1_result_comb[55];
    p1_result[56] <= p1_result_comb[56];
    p1_result[57] <= p1_result_comb[57];
    p1_result[58] <= p1_result_comb[58];
    p1_result[59] <= p1_result_comb[59];
    p1_result[60] <= p1_result_comb[60];
    p1_result[61] <= p1_result_comb[61];
    p1_result[62] <= p1_result_comb[62];
    p1_result[63] <= p1_result_comb[63];
  end
  assign out = {p1_result[63], p1_result[62], p1_result[61], p1_result[60], p1_result[59], p1_result[58], p1_result[57], p1_result[56], p1_result[55], p1_result[54], p1_result[53], p1_result[52], p1_result[51], p1_result[50], p1_result[49], p1_result[48], p1_result[47], p1_result[46], p1_result[45], p1_result[44], p1_result[43], p1_result[42], p1_result[41], p1_result[40], p1_result[39], p1_result[38], p1_result[37], p1_result[36], p1_result[35], p1_result[34], p1_result[33], p1_result[32], p1_result[31], p1_result[30], p1_result[29], p1_result[28], p1_result[27], p1_result[26], p1_result[25], p1_result[24], p1_result[23], p1_result[22], p1_result[21], p1_result[20], p1_result[19], p1_result[18], p1_result[17], p1_result[16], p1_result[15], p1_result[14], p1_result[13], p1_result[12], p1_result[11], p1_result[10], p1_result[9], p1_result[8], p1_result[7], p1_result[6], p1_result[5], p1_result[4], p1_result[3], p1_result[2], p1_result[1], p1_result[0]};
endmodule
