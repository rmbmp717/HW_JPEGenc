module dct_1d_u8(
  input wire clk,
  input wire [63:0] x,
  output wire [63:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [15:0] smul16b_8b_x_9b (input reg [7:0] lhs, input reg [8:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [8:0] signed_rhs;
    reg signed [15:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul16b_8b_x_9b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_6b (input reg [7:0] lhs, input reg [5:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [5:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_6b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [14:0] smul15b_8b_x_8b (input reg [7:0] lhs, input reg [7:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [7:0] signed_rhs;
    reg signed [14:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul15b_8b_x_8b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [13:0] smul14b_8b_x_7b (input reg [7:0] lhs, input reg [6:0] rhs);
    reg signed [7:0] signed_lhs;
    reg signed [6:0] signed_rhs;
    reg signed [13:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul14b_8b_x_7b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [23:0] umul24b_24b_x_7b (input reg [23:0] lhs, input reg [6:0] rhs);
    begin
      umul24b_24b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [7:0] x_unflattened[0:7];
  assign x_unflattened[0] = x[7:0];
  assign x_unflattened[1] = x[15:8];
  assign x_unflattened[2] = x[23:16];
  assign x_unflattened[3] = x[31:24];
  assign x_unflattened[4] = x[39:32];
  assign x_unflattened[5] = x[47:40];
  assign x_unflattened[6] = x[55:48];
  assign x_unflattened[7] = x[63:56];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_x[0:7];
  always @ (posedge clk) begin
    p0_x[0] <= x_unflattened[0];
    p0_x[1] <= x_unflattened[1];
    p0_x[2] <= x_unflattened[2];
    p0_x[3] <= x_unflattened[3];
    p0_x[4] <= x_unflattened[4];
    p0_x[5] <= x_unflattened[5];
    p0_x[6] <= x_unflattened[6];
    p0_x[7] <= x_unflattened[7];
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_array_index_5918_comb;
  wire [7:0] p1_array_index_5922_comb;
  wire [7:0] p1_array_index_5923_comb;
  wire [7:0] p1_array_index_5921_comb;
  wire [7:0] p1_array_index_5919_comb;
  wire [7:0] p1_array_index_5924_comb;
  wire [7:0] p1_array_index_5925_comb;
  wire [7:0] p1_array_index_5920_comb;
  wire [7:0] p1_concat_5950_comb;
  wire [7:0] p1_concat_5959_comb;
  wire [7:0] p1_concat_5961_comb;
  wire [7:0] p1_concat_5956_comb;
  wire [7:0] p1_concat_5952_comb;
  wire [7:0] p1_concat_5965_comb;
  wire [7:0] p1_concat_5967_comb;
  wire [7:0] p1_concat_5954_comb;
  wire [15:0] p1_smul_3287_NarrowedMult__comb;
  wire [15:0] p1_smul_3285_NarrowedMult__comb;
  wire [15:0] p1_smul_3282_NarrowedMult__comb;
  wire [15:0] p1_smul_3280_NarrowedMult__comb;
  wire [15:0] p1_smul_3270_NarrowedMult__comb;
  wire [15:0] p1_smul_3268_NarrowedMult__comb;
  wire [15:0] p1_smul_3267_NarrowedMult__comb;
  wire [15:0] p1_smul_3265_NarrowedMult__comb;
  wire [14:0] p1_smul_3294_NarrowedMult__comb;
  wire [14:0] p1_smul_3293_NarrowedMult__comb;
  wire [14:0] p1_smul_3290_NarrowedMult__comb;
  wire [14:0] p1_smul_3289_NarrowedMult__comb;
  wire [15:0] p1_smul_3279_NarrowedMult__comb;
  wire [15:0] p1_smul_3278_NarrowedMult__comb;
  wire [15:0] p1_smul_3277_NarrowedMult__comb;
  wire [15:0] p1_smul_3276_NarrowedMult__comb;
  wire [15:0] p1_smul_3275_NarrowedMult__comb;
  wire [15:0] p1_smul_3274_NarrowedMult__comb;
  wire [15:0] p1_smul_3273_NarrowedMult__comb;
  wire [15:0] p1_smul_3272_NarrowedMult__comb;
  wire [14:0] p1_smul_3263_NarrowedMult__comb;
  wire [14:0] p1_smul_3261_NarrowedMult__comb;
  wire [14:0] p1_smul_3258_NarrowedMult__comb;
  wire [14:0] p1_smul_3256_NarrowedMult__comb;
  wire [15:0] p1_smul_3303_NarrowedMult__comb;
  wire [15:0] p1_smul_3302_NarrowedMult__comb;
  wire [15:0] p1_smul_3297_NarrowedMult__comb;
  wire [15:0] p1_smul_3296_NarrowedMult__comb;
  wire [15:0] p1_smul_3253_NarrowedMult__comb;
  wire [15:0] p1_smul_3252_NarrowedMult__comb;
  wire [15:0] p1_smul_3251_NarrowedMult__comb;
  wire [15:0] p1_smul_3250_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6018_comb;
  wire [13:0] p1_smul_3378_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6020_comb;
  wire [14:0] p1_smul_3284_NarrowedMult__comb;
  wire [14:0] p1_smul_3283_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6023_comb;
  wire [13:0] p1_smul_3398_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6025_comb;
  wire [14:0] p1_smul_3271_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6035_comb;
  wire [13:0] p1_smul_3445_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6037_comb;
  wire [14:0] p1_bit_slice_6038_comb;
  wire [13:0] p1_smul_3455_NarrowedMult__comb;
  wire [14:0] p1_bit_slice_6040_comb;
  wire [14:0] p1_smul_3264_NarrowedMult__comb;
  wire [13:0] p1_smul_3295_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6111_comb;
  wire [13:0] p1_bit_slice_6112_comb;
  wire [13:0] p1_smul_3292_NarrowedMult__comb;
  wire [13:0] p1_smul_3291_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6115_comb;
  wire [13:0] p1_bit_slice_6116_comb;
  wire [13:0] p1_smul_3288_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6142_comb;
  wire [13:0] p1_smul_3262_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6144_comb;
  wire [13:0] p1_smul_3260_NarrowedMult__comb;
  wire [13:0] p1_smul_3259_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6147_comb;
  wire [13:0] p1_smul_3257_NarrowedMult__comb;
  wire [13:0] p1_bit_slice_6149_comb;
  wire [8:0] p1_add_6190_comb;
  wire [8:0] p1_add_6191_comb;
  wire [8:0] p1_add_6192_comb;
  wire [8:0] p1_add_6193_comb;
  wire [14:0] p1_smul_3301_NarrowedMult__comb;
  wire [13:0] p1_smul_3317_NarrowedMult__comb;
  wire [13:0] p1_smul_3319_NarrowedMult__comb;
  wire [14:0] p1_smul_3298_NarrowedMult__comb;
  wire [13:0] p1_smul_3506_NarrowedMult__comb;
  wire [14:0] p1_smul_3254_NarrowedMult__comb;
  wire [14:0] p1_smul_3249_NarrowedMult__comb;
  wire [13:0] p1_smul_3534_NarrowedMult__comb;
  wire [16:0] p1_add_6174_comb;
  wire [16:0] p1_add_6175_comb;
  wire [16:0] p1_add_6176_comb;
  wire [16:0] p1_add_6177_comb;
  wire [16:0] p1_add_6054_comb;
  wire [16:0] p1_add_6059_comb;
  wire [16:0] p1_add_6102_comb;
  wire [16:0] p1_add_6103_comb;
  wire [15:0] p1_add_6118_comb;
  wire [15:0] p1_add_6120_comb;
  wire [15:0] p1_add_6122_comb;
  wire [15:0] p1_add_6124_comb;
  wire [15:0] p1_add_6134_comb;
  wire [15:0] p1_add_6136_comb;
  wire [15:0] p1_add_6138_comb;
  wire [15:0] p1_add_6140_comb;
  wire [14:0] p1_add_6196_comb;
  wire [14:0] p1_add_6198_comb;
  wire [14:0] p1_add_6200_comb;
  wire [14:0] p1_add_6202_comb;
  wire [24:0] p1_sum__97_comb;
  wire [24:0] p1_sum__98_comb;
  wire [24:0] p1_sum__99_comb;
  wire [24:0] p1_sum__100_comb;
  wire [14:0] p1_add_6208_comb;
  wire [14:0] p1_add_6210_comb;
  wire [14:0] p1_add_6212_comb;
  wire [14:0] p1_add_6214_comb;
  wire [23:0] p1_add_6232_comb;
  wire [23:0] p1_add_6233_comb;
  wire [15:0] p1_bit_slice_6106_comb;
  wire [15:0] p1_add_6107_comb;
  wire [15:0] p1_add_6108_comb;
  wire [15:0] p1_bit_slice_6109_comb;
  wire [15:0] p1_add_6150_comb;
  wire [15:0] p1_bit_slice_6151_comb;
  wire [15:0] p1_bit_slice_6152_comb;
  wire [15:0] p1_add_6153_comb;
  wire [16:0] p1_concat_6170_comb;
  wire [16:0] p1_concat_6171_comb;
  wire [16:0] p1_concat_6172_comb;
  wire [16:0] p1_concat_6173_comb;
  wire [16:0] p1_concat_6178_comb;
  wire [16:0] p1_concat_6179_comb;
  wire [16:0] p1_concat_6180_comb;
  wire [16:0] p1_concat_6181_comb;
  wire p1_bit_slice_6194_comb;
  wire p1_bit_slice_6195_comb;
  wire p1_bit_slice_6216_comb;
  wire p1_bit_slice_6217_comb;
  wire [15:0] p1_concat_6222_comb;
  wire [15:0] p1_concat_6223_comb;
  wire [15:0] p1_concat_6224_comb;
  wire [15:0] p1_concat_6225_comb;
  wire [24:0] p1_sum__77_comb;
  wire [24:0] p1_sum__78_comb;
  wire [15:0] p1_concat_6228_comb;
  wire [15:0] p1_concat_6229_comb;
  wire [15:0] p1_concat_6230_comb;
  wire [15:0] p1_concat_6231_comb;
  wire [23:0] p1_add_6234_comb;
  assign p1_array_index_5918_comb = p0_x[3'h0];
  assign p1_array_index_5922_comb = p0_x[3'h2];
  assign p1_array_index_5923_comb = p0_x[3'h5];
  assign p1_array_index_5921_comb = p0_x[3'h7];
  assign p1_array_index_5919_comb = p0_x[3'h1];
  assign p1_array_index_5924_comb = p0_x[3'h3];
  assign p1_array_index_5925_comb = p0_x[3'h4];
  assign p1_array_index_5920_comb = p0_x[3'h6];
  assign p1_concat_5950_comb = {~p1_array_index_5918_comb[7], p1_array_index_5918_comb[6:0]};
  assign p1_concat_5959_comb = {~p1_array_index_5922_comb[7], p1_array_index_5922_comb[6:0]};
  assign p1_concat_5961_comb = {~p1_array_index_5923_comb[7], p1_array_index_5923_comb[6:0]};
  assign p1_concat_5956_comb = {~p1_array_index_5921_comb[7], p1_array_index_5921_comb[6:0]};
  assign p1_concat_5952_comb = {~p1_array_index_5919_comb[7], p1_array_index_5919_comb[6:0]};
  assign p1_concat_5965_comb = {~p1_array_index_5924_comb[7], p1_array_index_5924_comb[6:0]};
  assign p1_concat_5967_comb = {~p1_array_index_5925_comb[7], p1_array_index_5925_comb[6:0]};
  assign p1_concat_5954_comb = {~p1_array_index_5920_comb[7], p1_array_index_5920_comb[6:0]};
  assign p1_smul_3287_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5950_comb, 9'h0d5);
  assign p1_smul_3285_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5959_comb, 9'h105);
  assign p1_smul_3282_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5961_comb, 9'h0fb);
  assign p1_smul_3280_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5956_comb, 9'h12b);
  assign p1_smul_3270_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5952_comb, 9'h105);
  assign p1_smul_3268_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5965_comb, 9'h0d5);
  assign p1_smul_3267_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5967_comb, 9'h0d5);
  assign p1_smul_3265_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5954_comb, 9'h105);
  assign p1_smul_3294_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5952_comb, 7'h31);
  assign p1_smul_3293_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5959_comb, 7'h4f);
  assign p1_smul_3290_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5961_comb, 7'h4f);
  assign p1_smul_3289_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5954_comb, 7'h31);
  assign p1_smul_3279_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5950_comb, 9'h0b5);
  assign p1_smul_3278_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5952_comb, 9'h14b);
  assign p1_smul_3277_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5959_comb, 9'h14b);
  assign p1_smul_3276_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5965_comb, 9'h0b5);
  assign p1_smul_3275_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5967_comb, 9'h0b5);
  assign p1_smul_3274_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5961_comb, 9'h14b);
  assign p1_smul_3273_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5954_comb, 9'h14b);
  assign p1_smul_3272_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5956_comb, 9'h0b5);
  assign p1_smul_3263_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5950_comb, 7'h31);
  assign p1_smul_3261_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5959_comb, 7'h31);
  assign p1_smul_3258_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5961_comb, 7'h31);
  assign p1_smul_3256_NarrowedMult__comb = smul15b_8b_x_7b(p1_concat_5956_comb, 7'h31);
  assign p1_smul_3303_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5950_comb, 9'h0fb);
  assign p1_smul_3302_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5952_comb, 9'h0d5);
  assign p1_smul_3297_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5954_comb, 9'h12b);
  assign p1_smul_3296_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5956_comb, 9'h105);
  assign p1_smul_3253_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5959_comb, 9'h0d5);
  assign p1_smul_3252_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5965_comb, 9'h105);
  assign p1_smul_3251_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5967_comb, 9'h105);
  assign p1_smul_3250_NarrowedMult__comb = smul16b_8b_x_9b(p1_concat_5961_comb, 9'h0d5);
  assign p1_bit_slice_6018_comb = p1_smul_3287_NarrowedMult__comb[15:1];
  assign p1_smul_3378_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5952_comb, 6'h27);
  assign p1_bit_slice_6020_comb = p1_smul_3285_NarrowedMult__comb[15:1];
  assign p1_smul_3284_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5965_comb, 8'hb9);
  assign p1_smul_3283_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5967_comb, 8'h47);
  assign p1_bit_slice_6023_comb = p1_smul_3282_NarrowedMult__comb[15:1];
  assign p1_smul_3398_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5954_comb, 6'h19);
  assign p1_bit_slice_6025_comb = p1_smul_3280_NarrowedMult__comb[15:1];
  assign p1_smul_3271_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5950_comb, 8'h47);
  assign p1_bit_slice_6035_comb = p1_smul_3270_NarrowedMult__comb[15:1];
  assign p1_smul_3445_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5959_comb, 6'h27);
  assign p1_bit_slice_6037_comb = p1_smul_3268_NarrowedMult__comb[15:1];
  assign p1_bit_slice_6038_comb = p1_smul_3267_NarrowedMult__comb[15:1];
  assign p1_smul_3455_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5961_comb, 6'h27);
  assign p1_bit_slice_6040_comb = p1_smul_3265_NarrowedMult__comb[15:1];
  assign p1_smul_3264_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5956_comb, 8'h47);
  assign p1_smul_3295_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5950_comb, 7'h3b);
  assign p1_bit_slice_6111_comb = p1_smul_3294_NarrowedMult__comb[14:1];
  assign p1_bit_slice_6112_comb = p1_smul_3293_NarrowedMult__comb[14:1];
  assign p1_smul_3292_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5965_comb, 7'h45);
  assign p1_smul_3291_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5967_comb, 7'h45);
  assign p1_bit_slice_6115_comb = p1_smul_3290_NarrowedMult__comb[14:1];
  assign p1_bit_slice_6116_comb = p1_smul_3289_NarrowedMult__comb[14:1];
  assign p1_smul_3288_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5956_comb, 7'h3b);
  assign p1_bit_slice_6142_comb = p1_smul_3263_NarrowedMult__comb[14:1];
  assign p1_smul_3262_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5952_comb, 7'h45);
  assign p1_bit_slice_6144_comb = p1_smul_3261_NarrowedMult__comb[14:1];
  assign p1_smul_3260_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5965_comb, 7'h3b);
  assign p1_smul_3259_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5967_comb, 7'h3b);
  assign p1_bit_slice_6147_comb = p1_smul_3258_NarrowedMult__comb[14:1];
  assign p1_smul_3257_NarrowedMult__comb = smul14b_8b_x_7b(p1_concat_5954_comb, 7'h45);
  assign p1_bit_slice_6149_comb = p1_smul_3256_NarrowedMult__comb[14:1];
  assign p1_add_6190_comb = {{1{p1_concat_5950_comb[7]}}, p1_concat_5950_comb} + {{1{p1_concat_5952_comb[7]}}, p1_concat_5952_comb};
  assign p1_add_6191_comb = {{1{p1_concat_5959_comb[7]}}, p1_concat_5959_comb} + {{1{p1_concat_5965_comb[7]}}, p1_concat_5965_comb};
  assign p1_add_6192_comb = {{1{p1_concat_5967_comb[7]}}, p1_concat_5967_comb} + {{1{p1_concat_5961_comb[7]}}, p1_concat_5961_comb};
  assign p1_add_6193_comb = {{1{p1_concat_5954_comb[7]}}, p1_concat_5954_comb} + {{1{p1_concat_5956_comb[7]}}, p1_concat_5956_comb};
  assign p1_smul_3301_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5959_comb, 8'h47);
  assign p1_smul_3317_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5965_comb, 6'h19);
  assign p1_smul_3319_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5967_comb, 6'h27);
  assign p1_smul_3298_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5961_comb, 8'hb9);
  assign p1_smul_3506_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5950_comb, 6'h19);
  assign p1_smul_3254_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5952_comb, 8'hb9);
  assign p1_smul_3249_NarrowedMult__comb = smul15b_8b_x_8b(p1_concat_5954_comb, 8'hb9);
  assign p1_smul_3534_NarrowedMult__comb = smul14b_8b_x_6b(p1_concat_5956_comb, 6'h19);
  assign p1_add_6174_comb = {{1{p1_smul_3279_NarrowedMult__comb[15]}}, p1_smul_3279_NarrowedMult__comb} + {{1{p1_smul_3278_NarrowedMult__comb[15]}}, p1_smul_3278_NarrowedMult__comb};
  assign p1_add_6175_comb = {{1{p1_smul_3277_NarrowedMult__comb[15]}}, p1_smul_3277_NarrowedMult__comb} + {{1{p1_smul_3276_NarrowedMult__comb[15]}}, p1_smul_3276_NarrowedMult__comb};
  assign p1_add_6176_comb = {{1{p1_smul_3275_NarrowedMult__comb[15]}}, p1_smul_3275_NarrowedMult__comb} + {{1{p1_smul_3274_NarrowedMult__comb[15]}}, p1_smul_3274_NarrowedMult__comb};
  assign p1_add_6177_comb = {{1{p1_smul_3273_NarrowedMult__comb[15]}}, p1_smul_3273_NarrowedMult__comb} + {{1{p1_smul_3272_NarrowedMult__comb[15]}}, p1_smul_3272_NarrowedMult__comb};
  assign p1_add_6054_comb = {{1{p1_smul_3303_NarrowedMult__comb[15]}}, p1_smul_3303_NarrowedMult__comb} + {{1{p1_smul_3302_NarrowedMult__comb[15]}}, p1_smul_3302_NarrowedMult__comb};
  assign p1_add_6059_comb = {{1{p1_smul_3297_NarrowedMult__comb[15]}}, p1_smul_3297_NarrowedMult__comb} + {{1{p1_smul_3296_NarrowedMult__comb[15]}}, p1_smul_3296_NarrowedMult__comb};
  assign p1_add_6102_comb = {{1{p1_smul_3253_NarrowedMult__comb[15]}}, p1_smul_3253_NarrowedMult__comb} + {{1{p1_smul_3252_NarrowedMult__comb[15]}}, p1_smul_3252_NarrowedMult__comb};
  assign p1_add_6103_comb = {{1{p1_smul_3251_NarrowedMult__comb[15]}}, p1_smul_3251_NarrowedMult__comb} + {{1{p1_smul_3250_NarrowedMult__comb[15]}}, p1_smul_3250_NarrowedMult__comb};
  assign p1_add_6118_comb = {{1{p1_bit_slice_6018_comb[14]}}, p1_bit_slice_6018_comb} + {{2{p1_smul_3378_NarrowedMult__comb[13]}}, p1_smul_3378_NarrowedMult__comb};
  assign p1_add_6120_comb = {{1{p1_bit_slice_6020_comb[14]}}, p1_bit_slice_6020_comb} + {{1{p1_smul_3284_NarrowedMult__comb[14]}}, p1_smul_3284_NarrowedMult__comb};
  assign p1_add_6122_comb = {{1{p1_smul_3283_NarrowedMult__comb[14]}}, p1_smul_3283_NarrowedMult__comb} + {{1{p1_bit_slice_6023_comb[14]}}, p1_bit_slice_6023_comb};
  assign p1_add_6124_comb = {{2{p1_smul_3398_NarrowedMult__comb[13]}}, p1_smul_3398_NarrowedMult__comb} + {{1{p1_bit_slice_6025_comb[14]}}, p1_bit_slice_6025_comb};
  assign p1_add_6134_comb = {{1{p1_smul_3271_NarrowedMult__comb[14]}}, p1_smul_3271_NarrowedMult__comb} + {{1{p1_bit_slice_6035_comb[14]}}, p1_bit_slice_6035_comb};
  assign p1_add_6136_comb = {{2{p1_smul_3445_NarrowedMult__comb[13]}}, p1_smul_3445_NarrowedMult__comb} + {{1{p1_bit_slice_6037_comb[14]}}, p1_bit_slice_6037_comb};
  assign p1_add_6138_comb = {{1{p1_bit_slice_6038_comb[14]}}, p1_bit_slice_6038_comb} + {{2{p1_smul_3455_NarrowedMult__comb[13]}}, p1_smul_3455_NarrowedMult__comb};
  assign p1_add_6140_comb = {{1{p1_bit_slice_6040_comb[14]}}, p1_bit_slice_6040_comb} + {{1{p1_smul_3264_NarrowedMult__comb[14]}}, p1_smul_3264_NarrowedMult__comb};
  assign p1_add_6196_comb = {{1{p1_smul_3295_NarrowedMult__comb[13]}}, p1_smul_3295_NarrowedMult__comb} + {{1{p1_bit_slice_6111_comb[13]}}, p1_bit_slice_6111_comb};
  assign p1_add_6198_comb = {{1{p1_bit_slice_6112_comb[13]}}, p1_bit_slice_6112_comb} + {{1{p1_smul_3292_NarrowedMult__comb[13]}}, p1_smul_3292_NarrowedMult__comb};
  assign p1_add_6200_comb = {{1{p1_smul_3291_NarrowedMult__comb[13]}}, p1_smul_3291_NarrowedMult__comb} + {{1{p1_bit_slice_6115_comb[13]}}, p1_bit_slice_6115_comb};
  assign p1_add_6202_comb = {{1{p1_bit_slice_6116_comb[13]}}, p1_bit_slice_6116_comb} + {{1{p1_smul_3288_NarrowedMult__comb[13]}}, p1_smul_3288_NarrowedMult__comb};
  assign p1_sum__97_comb = {{8{p1_add_6174_comb[16]}}, p1_add_6174_comb};
  assign p1_sum__98_comb = {{8{p1_add_6175_comb[16]}}, p1_add_6175_comb};
  assign p1_sum__99_comb = {{8{p1_add_6176_comb[16]}}, p1_add_6176_comb};
  assign p1_sum__100_comb = {{8{p1_add_6177_comb[16]}}, p1_add_6177_comb};
  assign p1_add_6208_comb = {{1{p1_bit_slice_6142_comb[13]}}, p1_bit_slice_6142_comb} + {{1{p1_smul_3262_NarrowedMult__comb[13]}}, p1_smul_3262_NarrowedMult__comb};
  assign p1_add_6210_comb = {{1{p1_bit_slice_6144_comb[13]}}, p1_bit_slice_6144_comb} + {{1{p1_smul_3260_NarrowedMult__comb[13]}}, p1_smul_3260_NarrowedMult__comb};
  assign p1_add_6212_comb = {{1{p1_smul_3259_NarrowedMult__comb[13]}}, p1_smul_3259_NarrowedMult__comb} + {{1{p1_bit_slice_6147_comb[13]}}, p1_bit_slice_6147_comb};
  assign p1_add_6214_comb = {{1{p1_smul_3257_NarrowedMult__comb[13]}}, p1_smul_3257_NarrowedMult__comb} + {{1{p1_bit_slice_6149_comb[13]}}, p1_bit_slice_6149_comb};
  assign p1_add_6232_comb = {{15{p1_add_6190_comb[8]}}, p1_add_6190_comb} + {{15{p1_add_6191_comb[8]}}, p1_add_6191_comb};
  assign p1_add_6233_comb = {{15{p1_add_6192_comb[8]}}, p1_add_6192_comb} + {{15{p1_add_6193_comb[8]}}, p1_add_6193_comb};
  assign p1_bit_slice_6106_comb = p1_add_6054_comb[16:1];
  assign p1_add_6107_comb = {{1{p1_smul_3301_NarrowedMult__comb[14]}}, p1_smul_3301_NarrowedMult__comb} + {{2{p1_smul_3317_NarrowedMult__comb[13]}}, p1_smul_3317_NarrowedMult__comb};
  assign p1_add_6108_comb = {{2{p1_smul_3319_NarrowedMult__comb[13]}}, p1_smul_3319_NarrowedMult__comb} + {{1{p1_smul_3298_NarrowedMult__comb[14]}}, p1_smul_3298_NarrowedMult__comb};
  assign p1_bit_slice_6109_comb = p1_add_6059_comb[16:1];
  assign p1_add_6150_comb = {{2{p1_smul_3506_NarrowedMult__comb[13]}}, p1_smul_3506_NarrowedMult__comb} + {{1{p1_smul_3254_NarrowedMult__comb[14]}}, p1_smul_3254_NarrowedMult__comb};
  assign p1_bit_slice_6151_comb = p1_add_6102_comb[16:1];
  assign p1_bit_slice_6152_comb = p1_add_6103_comb[16:1];
  assign p1_add_6153_comb = {{1{p1_smul_3249_NarrowedMult__comb[14]}}, p1_smul_3249_NarrowedMult__comb} + {{2{p1_smul_3534_NarrowedMult__comb[13]}}, p1_smul_3534_NarrowedMult__comb};
  assign p1_concat_6170_comb = {p1_add_6118_comb, p1_smul_3287_NarrowedMult__comb[0]};
  assign p1_concat_6171_comb = {p1_add_6120_comb, p1_smul_3285_NarrowedMult__comb[0]};
  assign p1_concat_6172_comb = {p1_add_6122_comb, p1_smul_3282_NarrowedMult__comb[0]};
  assign p1_concat_6173_comb = {p1_add_6124_comb, p1_smul_3280_NarrowedMult__comb[0]};
  assign p1_concat_6178_comb = {p1_add_6134_comb, p1_smul_3270_NarrowedMult__comb[0]};
  assign p1_concat_6179_comb = {p1_add_6136_comb, p1_smul_3268_NarrowedMult__comb[0]};
  assign p1_concat_6180_comb = {p1_add_6138_comb, p1_smul_3267_NarrowedMult__comb[0]};
  assign p1_concat_6181_comb = {p1_add_6140_comb, p1_smul_3265_NarrowedMult__comb[0]};
  assign p1_bit_slice_6194_comb = p1_add_6054_comb[0];
  assign p1_bit_slice_6195_comb = p1_add_6059_comb[0];
  assign p1_bit_slice_6216_comb = p1_add_6102_comb[0];
  assign p1_bit_slice_6217_comb = p1_add_6103_comb[0];
  assign p1_concat_6222_comb = {p1_add_6196_comb, p1_smul_3294_NarrowedMult__comb[0]};
  assign p1_concat_6223_comb = {p1_add_6198_comb, p1_smul_3293_NarrowedMult__comb[0]};
  assign p1_concat_6224_comb = {p1_add_6200_comb, p1_smul_3290_NarrowedMult__comb[0]};
  assign p1_concat_6225_comb = {p1_add_6202_comb, p1_smul_3289_NarrowedMult__comb[0]};
  assign p1_sum__77_comb = p1_sum__97_comb + p1_sum__98_comb;
  assign p1_sum__78_comb = p1_sum__99_comb + p1_sum__100_comb;
  assign p1_concat_6228_comb = {p1_add_6208_comb, p1_smul_3263_NarrowedMult__comb[0]};
  assign p1_concat_6229_comb = {p1_add_6210_comb, p1_smul_3261_NarrowedMult__comb[0]};
  assign p1_concat_6230_comb = {p1_add_6212_comb, p1_smul_3258_NarrowedMult__comb[0]};
  assign p1_concat_6231_comb = {p1_add_6214_comb, p1_smul_3256_NarrowedMult__comb[0]};
  assign p1_add_6234_comb = p1_add_6232_comb + p1_add_6233_comb;

  // Registers for pipe stage 1:
  reg [15:0] p1_bit_slice_6106;
  reg [15:0] p1_add_6107;
  reg [15:0] p1_add_6108;
  reg [15:0] p1_bit_slice_6109;
  reg [15:0] p1_add_6150;
  reg [15:0] p1_bit_slice_6151;
  reg [15:0] p1_bit_slice_6152;
  reg [15:0] p1_add_6153;
  reg [16:0] p1_concat_6170;
  reg [16:0] p1_concat_6171;
  reg [16:0] p1_concat_6172;
  reg [16:0] p1_concat_6173;
  reg [16:0] p1_concat_6178;
  reg [16:0] p1_concat_6179;
  reg [16:0] p1_concat_6180;
  reg [16:0] p1_concat_6181;
  reg p1_bit_slice_6194;
  reg p1_bit_slice_6195;
  reg p1_bit_slice_6216;
  reg p1_bit_slice_6217;
  reg [15:0] p1_concat_6222;
  reg [15:0] p1_concat_6223;
  reg [15:0] p1_concat_6224;
  reg [15:0] p1_concat_6225;
  reg [24:0] p1_sum__77;
  reg [24:0] p1_sum__78;
  reg [15:0] p1_concat_6228;
  reg [15:0] p1_concat_6229;
  reg [15:0] p1_concat_6230;
  reg [15:0] p1_concat_6231;
  reg [23:0] p1_add_6234;
  always @ (posedge clk) begin
    p1_bit_slice_6106 <= p1_bit_slice_6106_comb;
    p1_add_6107 <= p1_add_6107_comb;
    p1_add_6108 <= p1_add_6108_comb;
    p1_bit_slice_6109 <= p1_bit_slice_6109_comb;
    p1_add_6150 <= p1_add_6150_comb;
    p1_bit_slice_6151 <= p1_bit_slice_6151_comb;
    p1_bit_slice_6152 <= p1_bit_slice_6152_comb;
    p1_add_6153 <= p1_add_6153_comb;
    p1_concat_6170 <= p1_concat_6170_comb;
    p1_concat_6171 <= p1_concat_6171_comb;
    p1_concat_6172 <= p1_concat_6172_comb;
    p1_concat_6173 <= p1_concat_6173_comb;
    p1_concat_6178 <= p1_concat_6178_comb;
    p1_concat_6179 <= p1_concat_6179_comb;
    p1_concat_6180 <= p1_concat_6180_comb;
    p1_concat_6181 <= p1_concat_6181_comb;
    p1_bit_slice_6194 <= p1_bit_slice_6194_comb;
    p1_bit_slice_6195 <= p1_bit_slice_6195_comb;
    p1_bit_slice_6216 <= p1_bit_slice_6216_comb;
    p1_bit_slice_6217 <= p1_bit_slice_6217_comb;
    p1_concat_6222 <= p1_concat_6222_comb;
    p1_concat_6223 <= p1_concat_6223_comb;
    p1_concat_6224 <= p1_concat_6224_comb;
    p1_concat_6225 <= p1_concat_6225_comb;
    p1_sum__77 <= p1_sum__77_comb;
    p1_sum__78 <= p1_sum__78_comb;
    p1_concat_6228 <= p1_concat_6228_comb;
    p1_concat_6229 <= p1_concat_6229_comb;
    p1_concat_6230 <= p1_concat_6230_comb;
    p1_concat_6231 <= p1_concat_6231_comb;
    p1_add_6234 <= p1_add_6234_comb;
  end

  // ===== Pipe stage 2:
  wire [24:0] p2_sum__67_comb;
  wire [23:0] p2_add_6305_comb;
  wire [23:0] p2_add_6306_comb;
  wire [24:0] p2_sum__101_comb;
  wire [24:0] p2_sum__102_comb;
  wire [24:0] p2_sum__103_comb;
  wire [24:0] p2_sum__104_comb;
  wire [24:0] p2_sum__93_comb;
  wire [24:0] p2_sum__94_comb;
  wire [24:0] p2_sum__95_comb;
  wire [24:0] p2_sum__96_comb;
  wire [23:0] p2_add_6315_comb;
  wire [23:0] p2_add_6316_comb;
  wire [23:0] p2_add_6345_comb;
  wire [23:0] p2_add_6346_comb;
  wire [24:0] p2_add_6348_comb;
  wire [23:0] p2_add_6350_comb;
  wire [23:0] p2_add_6351_comb;
  wire [24:0] p2_sum__83_comb;
  wire [24:0] p2_sum__84_comb;
  wire [24:0] p2_sum__79_comb;
  wire [24:0] p2_sum__80_comb;
  wire [24:0] p2_sum__75_comb;
  wire [24:0] p2_sum__76_comb;
  wire [24:0] p2_sum__71_comb;
  wire [24:0] p2_sum__72_comb;
  wire [23:0] p2_umul_2792_NarrowedMult__comb;
  wire [23:0] p2_add_6357_comb;
  wire [23:0] p2_add_6365_comb;
  wire [24:0] p2_sum__70_comb;
  wire [24:0] p2_sum__68_comb;
  wire [24:0] p2_sum__66_comb;
  wire [24:0] p2_sum__64_comb;
  wire [24:0] p2_add_6344_comb;
  wire [24:0] p2_add_6347_comb;
  wire [24:0] p2_add_6349_comb;
  wire [24:0] p2_add_6352_comb;
  wire [8:0] p2_clipped__16_comb;
  wire [8:0] p2_clipped__18_comb;
  wire [8:0] p2_clipped__20_comb;
  wire [8:0] p2_clipped__22_comb;
  wire [9:0] p2_add_6441_comb;
  wire [9:0] p2_add_6442_comb;
  wire [9:0] p2_add_6443_comb;
  wire [9:0] p2_add_6444_comb;
  wire [8:0] p2_clipped__17_comb;
  wire [8:0] p2_clipped__19_comb;
  wire [8:0] p2_clipped__21_comb;
  wire [8:0] p2_clipped__23_comb;
  wire [1:0] p2_bit_slice_6445_comb;
  wire [1:0] p2_bit_slice_6446_comb;
  wire [1:0] p2_bit_slice_6447_comb;
  wire [1:0] p2_bit_slice_6448_comb;
  wire [6:0] p2_bit_slice_6449_comb;
  wire [6:0] p2_bit_slice_6450_comb;
  wire [6:0] p2_bit_slice_6451_comb;
  wire [6:0] p2_bit_slice_6452_comb;
  assign p2_sum__67_comb = p1_sum__77 + p1_sum__78;
  assign p2_add_6305_comb = {{8{p1_bit_slice_6106[15]}}, p1_bit_slice_6106} + {{8{p1_add_6107[15]}}, p1_add_6107};
  assign p2_add_6306_comb = {{8{p1_add_6108[15]}}, p1_add_6108} + {{8{p1_bit_slice_6109[15]}}, p1_bit_slice_6109};
  assign p2_sum__101_comb = {{8{p1_concat_6170[16]}}, p1_concat_6170};
  assign p2_sum__102_comb = {{8{p1_concat_6171[16]}}, p1_concat_6171};
  assign p2_sum__103_comb = {{8{p1_concat_6172[16]}}, p1_concat_6172};
  assign p2_sum__104_comb = {{8{p1_concat_6173[16]}}, p1_concat_6173};
  assign p2_sum__93_comb = {{8{p1_concat_6178[16]}}, p1_concat_6178};
  assign p2_sum__94_comb = {{8{p1_concat_6179[16]}}, p1_concat_6179};
  assign p2_sum__95_comb = {{8{p1_concat_6180[16]}}, p1_concat_6180};
  assign p2_sum__96_comb = {{8{p1_concat_6181[16]}}, p1_concat_6181};
  assign p2_add_6315_comb = {{8{p1_add_6150[15]}}, p1_add_6150} + {{8{p1_bit_slice_6151[15]}}, p1_bit_slice_6151};
  assign p2_add_6316_comb = {{8{p1_bit_slice_6152[15]}}, p1_bit_slice_6152} + {{8{p1_add_6153[15]}}, p1_add_6153};
  assign p2_add_6345_comb = {{8{p1_concat_6222[15]}}, p1_concat_6222} + {{8{p1_concat_6223[15]}}, p1_concat_6223};
  assign p2_add_6346_comb = {{8{p1_concat_6224[15]}}, p1_concat_6224} + {{8{p1_concat_6225[15]}}, p1_concat_6225};
  assign p2_add_6348_comb = p2_sum__67_comb + 25'h000_0001;
  assign p2_add_6350_comb = {{8{p1_concat_6228[15]}}, p1_concat_6228} + {{8{p1_concat_6229[15]}}, p1_concat_6229};
  assign p2_add_6351_comb = {{8{p1_concat_6230[15]}}, p1_concat_6230} + {{8{p1_concat_6231[15]}}, p1_concat_6231};
  assign p2_sum__83_comb = {p2_add_6305_comb, p1_bit_slice_6194};
  assign p2_sum__84_comb = {p2_add_6306_comb, p1_bit_slice_6195};
  assign p2_sum__79_comb = p2_sum__101_comb + p2_sum__102_comb;
  assign p2_sum__80_comb = p2_sum__103_comb + p2_sum__104_comb;
  assign p2_sum__75_comb = p2_sum__93_comb + p2_sum__94_comb;
  assign p2_sum__76_comb = p2_sum__95_comb + p2_sum__96_comb;
  assign p2_sum__71_comb = {p2_add_6315_comb, p1_bit_slice_6216};
  assign p2_sum__72_comb = {p2_add_6316_comb, p1_bit_slice_6217};
  assign p2_umul_2792_NarrowedMult__comb = umul24b_24b_x_7b(p1_add_6234, 7'h5b);
  assign p2_add_6357_comb = p2_add_6345_comb + p2_add_6346_comb;
  assign p2_add_6365_comb = p2_add_6350_comb + p2_add_6351_comb;
  assign p2_sum__70_comb = p2_sum__83_comb + p2_sum__84_comb;
  assign p2_sum__68_comb = p2_sum__79_comb + p2_sum__80_comb;
  assign p2_sum__66_comb = p2_sum__75_comb + p2_sum__76_comb;
  assign p2_sum__64_comb = p2_sum__71_comb + p2_sum__72_comb;
  assign p2_add_6344_comb = p2_sum__70_comb + 25'h000_0001;
  assign p2_add_6347_comb = p2_sum__68_comb + 25'h000_0001;
  assign p2_add_6349_comb = p2_sum__66_comb + 25'h000_0001;
  assign p2_add_6352_comb = p2_sum__64_comb + 25'h000_0001;
  assign p2_clipped__16_comb = $signed(p2_umul_2792_NarrowedMult__comb) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_umul_2792_NarrowedMult__comb) > $signed(24'h00_7fff) ? 9'h0ff : p2_umul_2792_NarrowedMult__comb[15:7]);
  assign p2_clipped__18_comb = $signed(p2_add_6357_comb) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6357_comb) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6357_comb[15:7]);
  assign p2_clipped__20_comb = $signed(p2_add_6348_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6348_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6348_comb[16:8]);
  assign p2_clipped__22_comb = $signed(p2_add_6365_comb) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6365_comb) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6365_comb[15:7]);
  assign p2_add_6441_comb = {{1{p2_clipped__16_comb[8]}}, p2_clipped__16_comb} + 10'h001;
  assign p2_add_6442_comb = {{1{p2_clipped__18_comb[8]}}, p2_clipped__18_comb} + 10'h001;
  assign p2_add_6443_comb = {{1{p2_clipped__20_comb[8]}}, p2_clipped__20_comb} + 10'h001;
  assign p2_add_6444_comb = {{1{p2_clipped__22_comb[8]}}, p2_clipped__22_comb} + 10'h001;
  assign p2_clipped__17_comb = $signed(p2_add_6344_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6344_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6344_comb[16:8]);
  assign p2_clipped__19_comb = $signed(p2_add_6347_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6347_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6347_comb[16:8]);
  assign p2_clipped__21_comb = $signed(p2_add_6349_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6349_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6349_comb[16:8]);
  assign p2_clipped__23_comb = $signed(p2_add_6352_comb[24:1]) < $signed(24'hff_8000) ? 9'h100 : ($signed(p2_add_6352_comb[24:1]) > $signed(24'h00_7fff) ? 9'h0ff : p2_add_6352_comb[16:8]);
  assign p2_bit_slice_6445_comb = p2_add_6441_comb[9:8];
  assign p2_bit_slice_6446_comb = p2_add_6442_comb[9:8];
  assign p2_bit_slice_6447_comb = p2_add_6443_comb[9:8];
  assign p2_bit_slice_6448_comb = p2_add_6444_comb[9:8];
  assign p2_bit_slice_6449_comb = p2_add_6441_comb[7:1];
  assign p2_bit_slice_6450_comb = p2_add_6442_comb[7:1];
  assign p2_bit_slice_6451_comb = p2_add_6443_comb[7:1];
  assign p2_bit_slice_6452_comb = p2_add_6444_comb[7:1];

  // Registers for pipe stage 2:
  reg [8:0] p2_clipped__17;
  reg [8:0] p2_clipped__19;
  reg [8:0] p2_clipped__21;
  reg [8:0] p2_clipped__23;
  reg [1:0] p2_bit_slice_6445;
  reg [1:0] p2_bit_slice_6446;
  reg [1:0] p2_bit_slice_6447;
  reg [1:0] p2_bit_slice_6448;
  reg [6:0] p2_bit_slice_6449;
  reg [6:0] p2_bit_slice_6450;
  reg [6:0] p2_bit_slice_6451;
  reg [6:0] p2_bit_slice_6452;
  always @ (posedge clk) begin
    p2_clipped__17 <= p2_clipped__17_comb;
    p2_clipped__19 <= p2_clipped__19_comb;
    p2_clipped__21 <= p2_clipped__21_comb;
    p2_clipped__23 <= p2_clipped__23_comb;
    p2_bit_slice_6445 <= p2_bit_slice_6445_comb;
    p2_bit_slice_6446 <= p2_bit_slice_6446_comb;
    p2_bit_slice_6447 <= p2_bit_slice_6447_comb;
    p2_bit_slice_6448 <= p2_bit_slice_6448_comb;
    p2_bit_slice_6449 <= p2_bit_slice_6449_comb;
    p2_bit_slice_6450 <= p2_bit_slice_6450_comb;
    p2_bit_slice_6451 <= p2_bit_slice_6451_comb;
    p2_bit_slice_6452 <= p2_bit_slice_6452_comb;
  end

  // ===== Pipe stage 3:
  wire [9:0] p3_add_6485_comb;
  wire [9:0] p3_add_6486_comb;
  wire [9:0] p3_add_6487_comb;
  wire [9:0] p3_add_6488_comb;
  wire [1:0] p3_bit_slice_6489_comb;
  wire [1:0] p3_bit_slice_6490_comb;
  wire [1:0] p3_bit_slice_6491_comb;
  wire [1:0] p3_bit_slice_6492_comb;
  wire [2:0] p3_add_6509_comb;
  wire [2:0] p3_add_6510_comb;
  wire [2:0] p3_add_6511_comb;
  wire [2:0] p3_add_6512_comb;
  wire [2:0] p3_add_6513_comb;
  wire [2:0] p3_add_6514_comb;
  wire [2:0] p3_add_6515_comb;
  wire [2:0] p3_add_6516_comb;
  wire [7:0] p3_clipped__8_comb;
  wire [7:0] p3_clipped__9_comb;
  wire [7:0] p3_clipped__10_comb;
  wire [7:0] p3_clipped__11_comb;
  wire [7:0] p3_clipped__12_comb;
  wire [7:0] p3_clipped__13_comb;
  wire [7:0] p3_clipped__14_comb;
  wire [7:0] p3_clipped__15_comb;
  wire [7:0] p3_result_comb[0:7];
  assign p3_add_6485_comb = {{1{p2_clipped__17[8]}}, p2_clipped__17} + 10'h001;
  assign p3_add_6486_comb = {{1{p2_clipped__19[8]}}, p2_clipped__19} + 10'h001;
  assign p3_add_6487_comb = {{1{p2_clipped__21[8]}}, p2_clipped__21} + 10'h001;
  assign p3_add_6488_comb = {{1{p2_clipped__23[8]}}, p2_clipped__23} + 10'h001;
  assign p3_bit_slice_6489_comb = p3_add_6485_comb[9:8];
  assign p3_bit_slice_6490_comb = p3_add_6486_comb[9:8];
  assign p3_bit_slice_6491_comb = p3_add_6487_comb[9:8];
  assign p3_bit_slice_6492_comb = p3_add_6488_comb[9:8];
  assign p3_add_6509_comb = {{1{p2_bit_slice_6445[1]}}, p2_bit_slice_6445} + 3'h1;
  assign p3_add_6510_comb = {{1{p3_bit_slice_6489_comb[1]}}, p3_bit_slice_6489_comb} + 3'h1;
  assign p3_add_6511_comb = {{1{p2_bit_slice_6446[1]}}, p2_bit_slice_6446} + 3'h1;
  assign p3_add_6512_comb = {{1{p3_bit_slice_6490_comb[1]}}, p3_bit_slice_6490_comb} + 3'h1;
  assign p3_add_6513_comb = {{1{p2_bit_slice_6447[1]}}, p2_bit_slice_6447} + 3'h1;
  assign p3_add_6514_comb = {{1{p3_bit_slice_6491_comb[1]}}, p3_bit_slice_6491_comb} + 3'h1;
  assign p3_add_6515_comb = {{1{p2_bit_slice_6448[1]}}, p2_bit_slice_6448} + 3'h1;
  assign p3_add_6516_comb = {{1{p3_bit_slice_6492_comb[1]}}, p3_bit_slice_6492_comb} + 3'h1;
  assign p3_clipped__8_comb = p3_add_6509_comb[1] ? 8'hff : {p3_add_6509_comb[0], p2_bit_slice_6449};
  assign p3_clipped__9_comb = p3_add_6510_comb[1] ? 8'hff : {p3_add_6510_comb[0], p3_add_6485_comb[7:1]};
  assign p3_clipped__10_comb = p3_add_6511_comb[1] ? 8'hff : {p3_add_6511_comb[0], p2_bit_slice_6450};
  assign p3_clipped__11_comb = p3_add_6512_comb[1] ? 8'hff : {p3_add_6512_comb[0], p3_add_6486_comb[7:1]};
  assign p3_clipped__12_comb = p3_add_6513_comb[1] ? 8'hff : {p3_add_6513_comb[0], p2_bit_slice_6451};
  assign p3_clipped__13_comb = p3_add_6514_comb[1] ? 8'hff : {p3_add_6514_comb[0], p3_add_6487_comb[7:1]};
  assign p3_clipped__14_comb = p3_add_6515_comb[1] ? 8'hff : {p3_add_6515_comb[0], p2_bit_slice_6452};
  assign p3_clipped__15_comb = p3_add_6516_comb[1] ? 8'hff : {p3_add_6516_comb[0], p3_add_6488_comb[7:1]};
  assign p3_result_comb[0] = p3_clipped__8_comb;
  assign p3_result_comb[1] = p3_clipped__9_comb;
  assign p3_result_comb[2] = p3_clipped__10_comb;
  assign p3_result_comb[3] = p3_clipped__11_comb;
  assign p3_result_comb[4] = p3_clipped__12_comb;
  assign p3_result_comb[5] = p3_clipped__13_comb;
  assign p3_result_comb[6] = p3_clipped__14_comb;
  assign p3_result_comb[7] = p3_clipped__15_comb;

  // Registers for pipe stage 3:
  reg [7:0] p3_result[0:7];
  always @ (posedge clk) begin
    p3_result[0] <= p3_result_comb[0];
    p3_result[1] <= p3_result_comb[1];
    p3_result[2] <= p3_result_comb[2];
    p3_result[3] <= p3_result_comb[3];
    p3_result[4] <= p3_result_comb[4];
    p3_result[5] <= p3_result_comb[5];
    p3_result[6] <= p3_result_comb[6];
    p3_result[7] <= p3_result_comb[7];
  end
  assign out = {p3_result[7], p3_result[6], p3_result[5], p3_result[4], p3_result[3], p3_result[2], p3_result[1], p3_result[0]};
endmodule
