module Quantize(
  input wire clk,
  input wire [767:0] dct_coeffs,
  input wire [7:0] matrix_row,
  input wire is_luminance,
  input wire quantize_off,
  output wire [79:0] out
);
  function automatic [31:0] sdiv_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    begin
      sdiv_32b = rhs == 32'h0000_0000 ? (lhs[31] ? 32'h8000_0000 : 32'h7fff_ffff) : (lhs == 32'h8000_0000 && rhs == 32'hffff_ffff ? 32'h8000_0000 : $unsigned($signed(lhs) / $signed(rhs)));
    end
  endfunction
  wire [15:0] CHROMINANCE_QUANT_TBL[0:7][0:7];
  assign CHROMINANCE_QUANT_TBL[0][0] = 16'h0002;
  assign CHROMINANCE_QUANT_TBL[0][1] = 16'h0002;
  assign CHROMINANCE_QUANT_TBL[0][2] = 16'h0002;
  assign CHROMINANCE_QUANT_TBL[0][3] = 16'h0005;
  assign CHROMINANCE_QUANT_TBL[0][4] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[0][5] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[0][6] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[0][7] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[1][0] = 16'h0002;
  assign CHROMINANCE_QUANT_TBL[1][1] = 16'h0002;
  assign CHROMINANCE_QUANT_TBL[1][2] = 16'h0003;
  assign CHROMINANCE_QUANT_TBL[1][3] = 16'h0007;
  assign CHROMINANCE_QUANT_TBL[1][4] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[1][5] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[1][6] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[1][7] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[2][0] = 16'h0002;
  assign CHROMINANCE_QUANT_TBL[2][1] = 16'h0003;
  assign CHROMINANCE_QUANT_TBL[2][2] = 16'h0006;
  assign CHROMINANCE_QUANT_TBL[2][3] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[2][4] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[2][5] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[2][6] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[2][7] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[3][0] = 16'h0005;
  assign CHROMINANCE_QUANT_TBL[3][1] = 16'h0007;
  assign CHROMINANCE_QUANT_TBL[3][2] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[3][3] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[3][4] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[3][5] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[3][6] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[3][7] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[4][0] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[4][1] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[4][2] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[4][3] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[4][4] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[4][5] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[4][6] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[4][7] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[5][0] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[5][1] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[5][2] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[5][3] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[5][4] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[5][5] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[5][6] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[5][7] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[6][0] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[6][1] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[6][2] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[6][3] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[6][4] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[6][5] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[6][6] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[6][7] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[7][0] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[7][1] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[7][2] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[7][3] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[7][4] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[7][5] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[7][6] = 16'h000a;
  assign CHROMINANCE_QUANT_TBL[7][7] = 16'h000a;
  wire [15:0] LUMINANCE_QUANT_TBL[0:7][0:7];
  assign LUMINANCE_QUANT_TBL[0][0] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[0][1] = 16'h0001;
  assign LUMINANCE_QUANT_TBL[0][2] = 16'h0001;
  assign LUMINANCE_QUANT_TBL[0][3] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[0][4] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[0][5] = 16'h0004;
  assign LUMINANCE_QUANT_TBL[0][6] = 16'h0005;
  assign LUMINANCE_QUANT_TBL[0][7] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[1][0] = 16'h0001;
  assign LUMINANCE_QUANT_TBL[1][1] = 16'h0001;
  assign LUMINANCE_QUANT_TBL[1][2] = 16'h0001;
  assign LUMINANCE_QUANT_TBL[1][3] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[1][4] = 16'h0003;
  assign LUMINANCE_QUANT_TBL[1][5] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[1][6] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[1][7] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[2][0] = 16'h0001;
  assign LUMINANCE_QUANT_TBL[2][1] = 16'h0001;
  assign LUMINANCE_QUANT_TBL[2][2] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[2][3] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[2][4] = 16'h0004;
  assign LUMINANCE_QUANT_TBL[2][5] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[2][6] = 16'h0007;
  assign LUMINANCE_QUANT_TBL[2][7] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[3][0] = 16'h0001;
  assign LUMINANCE_QUANT_TBL[3][1] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[3][2] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[3][3] = 16'h0003;
  assign LUMINANCE_QUANT_TBL[3][4] = 16'h0005;
  assign LUMINANCE_QUANT_TBL[3][5] = 16'h0009;
  assign LUMINANCE_QUANT_TBL[3][6] = 16'h0008;
  assign LUMINANCE_QUANT_TBL[3][7] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[4][0] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[4][1] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[4][2] = 16'h0004;
  assign LUMINANCE_QUANT_TBL[4][3] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[4][4] = 16'h0007;
  assign LUMINANCE_QUANT_TBL[4][5] = 16'h000b;
  assign LUMINANCE_QUANT_TBL[4][6] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[4][7] = 16'h0008;
  assign LUMINANCE_QUANT_TBL[5][0] = 16'h0002;
  assign LUMINANCE_QUANT_TBL[5][1] = 16'h0004;
  assign LUMINANCE_QUANT_TBL[5][2] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[5][3] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[5][4] = 16'h0008;
  assign LUMINANCE_QUANT_TBL[5][5] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[5][6] = 16'h000b;
  assign LUMINANCE_QUANT_TBL[5][7] = 16'h0009;
  assign LUMINANCE_QUANT_TBL[6][0] = 16'h0005;
  assign LUMINANCE_QUANT_TBL[6][1] = 16'h0006;
  assign LUMINANCE_QUANT_TBL[6][2] = 16'h0008;
  assign LUMINANCE_QUANT_TBL[6][3] = 16'h0009;
  assign LUMINANCE_QUANT_TBL[6][4] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[6][5] = 16'h000c;
  assign LUMINANCE_QUANT_TBL[6][6] = 16'h000c;
  assign LUMINANCE_QUANT_TBL[6][7] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[7][0] = 16'h0007;
  assign LUMINANCE_QUANT_TBL[7][1] = 16'h0009;
  assign LUMINANCE_QUANT_TBL[7][2] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[7][3] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[7][4] = 16'h000b;
  assign LUMINANCE_QUANT_TBL[7][5] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[7][6] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[7][7] = 16'h000a;
  wire [11:0] dct_coeffs_unflattened[0:7][0:7];
  assign dct_coeffs_unflattened[0][0] = dct_coeffs[11:0];
  assign dct_coeffs_unflattened[0][1] = dct_coeffs[23:12];
  assign dct_coeffs_unflattened[0][2] = dct_coeffs[35:24];
  assign dct_coeffs_unflattened[0][3] = dct_coeffs[47:36];
  assign dct_coeffs_unflattened[0][4] = dct_coeffs[59:48];
  assign dct_coeffs_unflattened[0][5] = dct_coeffs[71:60];
  assign dct_coeffs_unflattened[0][6] = dct_coeffs[83:72];
  assign dct_coeffs_unflattened[0][7] = dct_coeffs[95:84];
  assign dct_coeffs_unflattened[1][0] = dct_coeffs[107:96];
  assign dct_coeffs_unflattened[1][1] = dct_coeffs[119:108];
  assign dct_coeffs_unflattened[1][2] = dct_coeffs[131:120];
  assign dct_coeffs_unflattened[1][3] = dct_coeffs[143:132];
  assign dct_coeffs_unflattened[1][4] = dct_coeffs[155:144];
  assign dct_coeffs_unflattened[1][5] = dct_coeffs[167:156];
  assign dct_coeffs_unflattened[1][6] = dct_coeffs[179:168];
  assign dct_coeffs_unflattened[1][7] = dct_coeffs[191:180];
  assign dct_coeffs_unflattened[2][0] = dct_coeffs[203:192];
  assign dct_coeffs_unflattened[2][1] = dct_coeffs[215:204];
  assign dct_coeffs_unflattened[2][2] = dct_coeffs[227:216];
  assign dct_coeffs_unflattened[2][3] = dct_coeffs[239:228];
  assign dct_coeffs_unflattened[2][4] = dct_coeffs[251:240];
  assign dct_coeffs_unflattened[2][5] = dct_coeffs[263:252];
  assign dct_coeffs_unflattened[2][6] = dct_coeffs[275:264];
  assign dct_coeffs_unflattened[2][7] = dct_coeffs[287:276];
  assign dct_coeffs_unflattened[3][0] = dct_coeffs[299:288];
  assign dct_coeffs_unflattened[3][1] = dct_coeffs[311:300];
  assign dct_coeffs_unflattened[3][2] = dct_coeffs[323:312];
  assign dct_coeffs_unflattened[3][3] = dct_coeffs[335:324];
  assign dct_coeffs_unflattened[3][4] = dct_coeffs[347:336];
  assign dct_coeffs_unflattened[3][5] = dct_coeffs[359:348];
  assign dct_coeffs_unflattened[3][6] = dct_coeffs[371:360];
  assign dct_coeffs_unflattened[3][7] = dct_coeffs[383:372];
  assign dct_coeffs_unflattened[4][0] = dct_coeffs[395:384];
  assign dct_coeffs_unflattened[4][1] = dct_coeffs[407:396];
  assign dct_coeffs_unflattened[4][2] = dct_coeffs[419:408];
  assign dct_coeffs_unflattened[4][3] = dct_coeffs[431:420];
  assign dct_coeffs_unflattened[4][4] = dct_coeffs[443:432];
  assign dct_coeffs_unflattened[4][5] = dct_coeffs[455:444];
  assign dct_coeffs_unflattened[4][6] = dct_coeffs[467:456];
  assign dct_coeffs_unflattened[4][7] = dct_coeffs[479:468];
  assign dct_coeffs_unflattened[5][0] = dct_coeffs[491:480];
  assign dct_coeffs_unflattened[5][1] = dct_coeffs[503:492];
  assign dct_coeffs_unflattened[5][2] = dct_coeffs[515:504];
  assign dct_coeffs_unflattened[5][3] = dct_coeffs[527:516];
  assign dct_coeffs_unflattened[5][4] = dct_coeffs[539:528];
  assign dct_coeffs_unflattened[5][5] = dct_coeffs[551:540];
  assign dct_coeffs_unflattened[5][6] = dct_coeffs[563:552];
  assign dct_coeffs_unflattened[5][7] = dct_coeffs[575:564];
  assign dct_coeffs_unflattened[6][0] = dct_coeffs[587:576];
  assign dct_coeffs_unflattened[6][1] = dct_coeffs[599:588];
  assign dct_coeffs_unflattened[6][2] = dct_coeffs[611:600];
  assign dct_coeffs_unflattened[6][3] = dct_coeffs[623:612];
  assign dct_coeffs_unflattened[6][4] = dct_coeffs[635:624];
  assign dct_coeffs_unflattened[6][5] = dct_coeffs[647:636];
  assign dct_coeffs_unflattened[6][6] = dct_coeffs[659:648];
  assign dct_coeffs_unflattened[6][7] = dct_coeffs[671:660];
  assign dct_coeffs_unflattened[7][0] = dct_coeffs[683:672];
  assign dct_coeffs_unflattened[7][1] = dct_coeffs[695:684];
  assign dct_coeffs_unflattened[7][2] = dct_coeffs[707:696];
  assign dct_coeffs_unflattened[7][3] = dct_coeffs[719:708];
  assign dct_coeffs_unflattened[7][4] = dct_coeffs[731:720];
  assign dct_coeffs_unflattened[7][5] = dct_coeffs[743:732];
  assign dct_coeffs_unflattened[7][6] = dct_coeffs[755:744];
  assign dct_coeffs_unflattened[7][7] = dct_coeffs[767:756];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [11:0] p0_dct_coeffs[0:7][0:7];
  reg [7:0] p0_matrix_row;
  reg p0_is_luminance;
  reg p0_quantize_off;
  always @ (posedge clk) begin
    p0_dct_coeffs[0][0] <= dct_coeffs_unflattened[0][0];
    p0_dct_coeffs[0][1] <= dct_coeffs_unflattened[0][1];
    p0_dct_coeffs[0][2] <= dct_coeffs_unflattened[0][2];
    p0_dct_coeffs[0][3] <= dct_coeffs_unflattened[0][3];
    p0_dct_coeffs[0][4] <= dct_coeffs_unflattened[0][4];
    p0_dct_coeffs[0][5] <= dct_coeffs_unflattened[0][5];
    p0_dct_coeffs[0][6] <= dct_coeffs_unflattened[0][6];
    p0_dct_coeffs[0][7] <= dct_coeffs_unflattened[0][7];
    p0_dct_coeffs[1][0] <= dct_coeffs_unflattened[1][0];
    p0_dct_coeffs[1][1] <= dct_coeffs_unflattened[1][1];
    p0_dct_coeffs[1][2] <= dct_coeffs_unflattened[1][2];
    p0_dct_coeffs[1][3] <= dct_coeffs_unflattened[1][3];
    p0_dct_coeffs[1][4] <= dct_coeffs_unflattened[1][4];
    p0_dct_coeffs[1][5] <= dct_coeffs_unflattened[1][5];
    p0_dct_coeffs[1][6] <= dct_coeffs_unflattened[1][6];
    p0_dct_coeffs[1][7] <= dct_coeffs_unflattened[1][7];
    p0_dct_coeffs[2][0] <= dct_coeffs_unflattened[2][0];
    p0_dct_coeffs[2][1] <= dct_coeffs_unflattened[2][1];
    p0_dct_coeffs[2][2] <= dct_coeffs_unflattened[2][2];
    p0_dct_coeffs[2][3] <= dct_coeffs_unflattened[2][3];
    p0_dct_coeffs[2][4] <= dct_coeffs_unflattened[2][4];
    p0_dct_coeffs[2][5] <= dct_coeffs_unflattened[2][5];
    p0_dct_coeffs[2][6] <= dct_coeffs_unflattened[2][6];
    p0_dct_coeffs[2][7] <= dct_coeffs_unflattened[2][7];
    p0_dct_coeffs[3][0] <= dct_coeffs_unflattened[3][0];
    p0_dct_coeffs[3][1] <= dct_coeffs_unflattened[3][1];
    p0_dct_coeffs[3][2] <= dct_coeffs_unflattened[3][2];
    p0_dct_coeffs[3][3] <= dct_coeffs_unflattened[3][3];
    p0_dct_coeffs[3][4] <= dct_coeffs_unflattened[3][4];
    p0_dct_coeffs[3][5] <= dct_coeffs_unflattened[3][5];
    p0_dct_coeffs[3][6] <= dct_coeffs_unflattened[3][6];
    p0_dct_coeffs[3][7] <= dct_coeffs_unflattened[3][7];
    p0_dct_coeffs[4][0] <= dct_coeffs_unflattened[4][0];
    p0_dct_coeffs[4][1] <= dct_coeffs_unflattened[4][1];
    p0_dct_coeffs[4][2] <= dct_coeffs_unflattened[4][2];
    p0_dct_coeffs[4][3] <= dct_coeffs_unflattened[4][3];
    p0_dct_coeffs[4][4] <= dct_coeffs_unflattened[4][4];
    p0_dct_coeffs[4][5] <= dct_coeffs_unflattened[4][5];
    p0_dct_coeffs[4][6] <= dct_coeffs_unflattened[4][6];
    p0_dct_coeffs[4][7] <= dct_coeffs_unflattened[4][7];
    p0_dct_coeffs[5][0] <= dct_coeffs_unflattened[5][0];
    p0_dct_coeffs[5][1] <= dct_coeffs_unflattened[5][1];
    p0_dct_coeffs[5][2] <= dct_coeffs_unflattened[5][2];
    p0_dct_coeffs[5][3] <= dct_coeffs_unflattened[5][3];
    p0_dct_coeffs[5][4] <= dct_coeffs_unflattened[5][4];
    p0_dct_coeffs[5][5] <= dct_coeffs_unflattened[5][5];
    p0_dct_coeffs[5][6] <= dct_coeffs_unflattened[5][6];
    p0_dct_coeffs[5][7] <= dct_coeffs_unflattened[5][7];
    p0_dct_coeffs[6][0] <= dct_coeffs_unflattened[6][0];
    p0_dct_coeffs[6][1] <= dct_coeffs_unflattened[6][1];
    p0_dct_coeffs[6][2] <= dct_coeffs_unflattened[6][2];
    p0_dct_coeffs[6][3] <= dct_coeffs_unflattened[6][3];
    p0_dct_coeffs[6][4] <= dct_coeffs_unflattened[6][4];
    p0_dct_coeffs[6][5] <= dct_coeffs_unflattened[6][5];
    p0_dct_coeffs[6][6] <= dct_coeffs_unflattened[6][6];
    p0_dct_coeffs[6][7] <= dct_coeffs_unflattened[6][7];
    p0_dct_coeffs[7][0] <= dct_coeffs_unflattened[7][0];
    p0_dct_coeffs[7][1] <= dct_coeffs_unflattened[7][1];
    p0_dct_coeffs[7][2] <= dct_coeffs_unflattened[7][2];
    p0_dct_coeffs[7][3] <= dct_coeffs_unflattened[7][3];
    p0_dct_coeffs[7][4] <= dct_coeffs_unflattened[7][4];
    p0_dct_coeffs[7][5] <= dct_coeffs_unflattened[7][5];
    p0_dct_coeffs[7][6] <= dct_coeffs_unflattened[7][6];
    p0_dct_coeffs[7][7] <= dct_coeffs_unflattened[7][7];
    p0_matrix_row <= matrix_row;
    p0_is_luminance <= is_luminance;
    p0_quantize_off <= quantize_off;
  end

  // ===== Pipe stage 1:
  wire [11:0] p1_array_index_816_comb;
  wire [3:0] p1_q_value_squeezed_comb;
  wire [11:0] p1_array_index_819_comb;
  wire [3:0] p1_q_value__1_squeezed_comb;
  wire [11:0] p1_array_index_822_comb;
  wire [3:0] p1_q_value__2_squeezed_comb;
  wire [11:0] p1_array_index_825_comb;
  wire [3:0] p1_q_value__3_squeezed_comb;
  wire [11:0] p1_array_index_828_comb;
  wire [3:0] p1_q_value__4_squeezed_comb;
  wire [11:0] p1_array_index_831_comb;
  wire [3:0] p1_q_value__5_squeezed_comb;
  wire [11:0] p1_array_index_834_comb;
  wire [3:0] p1_q_value__6_squeezed_comb;
  wire [11:0] p1_array_index_837_comb;
  wire [3:0] p1_q_value__7_squeezed_comb;
  wire [31:0] p1_sdiv_856_comb;
  wire [31:0] p1_sdiv_857_comb;
  wire [31:0] p1_sdiv_858_comb;
  wire [31:0] p1_sdiv_859_comb;
  wire [31:0] p1_sdiv_860_comb;
  wire [31:0] p1_sdiv_861_comb;
  wire [31:0] p1_sdiv_862_comb;
  wire [31:0] p1_sdiv_863_comb;
  wire [11:0] p1_divided_squeezed_comb;
  wire [11:0] p1_divided__1_squeezed_comb;
  wire [11:0] p1_divided__2_squeezed_comb;
  wire [11:0] p1_divided__3_squeezed_comb;
  wire [11:0] p1_divided__4_squeezed_comb;
  wire [11:0] p1_divided__5_squeezed_comb;
  wire [11:0] p1_divided__6_squeezed_comb;
  wire [11:0] p1_divided__7_squeezed_comb;
  wire [9:0] p1_clipped_comb;
  wire [9:0] p1_clipped__1_comb;
  wire [9:0] p1_clipped__2_comb;
  wire [9:0] p1_clipped__3_comb;
  wire [9:0] p1_clipped__4_comb;
  wire [9:0] p1_clipped__5_comb;
  wire [9:0] p1_clipped__6_comb;
  wire [9:0] p1_clipped__7_comb;
  wire [9:0] p1_array_952_comb[0:7];
  assign p1_array_index_816_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h0];
  assign p1_q_value_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h0][3:0] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h0][3:0];
  assign p1_array_index_819_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h1];
  assign p1_q_value__1_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h1][3:0] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h1][3:0];
  assign p1_array_index_822_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h2];
  assign p1_q_value__2_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h2][3:0] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h2][3:0];
  assign p1_array_index_825_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h3];
  assign p1_q_value__3_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h3][3:0] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h3][3:0];
  assign p1_array_index_828_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h4];
  assign p1_q_value__4_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h4][3:0] : 4'ha;
  assign p1_array_index_831_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h5];
  assign p1_q_value__5_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h5][3:0] : 4'ha;
  assign p1_array_index_834_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h6];
  assign p1_q_value__6_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h6][3:0] : 4'ha;
  assign p1_array_index_837_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h7];
  assign p1_q_value__7_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h7][3:0] : 4'ha;
  assign p1_sdiv_856_comb = sdiv_32b({{20{p1_array_index_816_comb[11]}}, p1_array_index_816_comb}, {28'h000_0000, p1_q_value_squeezed_comb});
  assign p1_sdiv_857_comb = sdiv_32b({{20{p1_array_index_819_comb[11]}}, p1_array_index_819_comb}, {28'h000_0000, p1_q_value__1_squeezed_comb});
  assign p1_sdiv_858_comb = sdiv_32b({{20{p1_array_index_822_comb[11]}}, p1_array_index_822_comb}, {28'h000_0000, p1_q_value__2_squeezed_comb});
  assign p1_sdiv_859_comb = sdiv_32b({{20{p1_array_index_825_comb[11]}}, p1_array_index_825_comb}, {28'h000_0000, p1_q_value__3_squeezed_comb});
  assign p1_sdiv_860_comb = sdiv_32b({{20{p1_array_index_828_comb[11]}}, p1_array_index_828_comb}, {28'h000_0000, p1_q_value__4_squeezed_comb});
  assign p1_sdiv_861_comb = sdiv_32b({{20{p1_array_index_831_comb[11]}}, p1_array_index_831_comb}, {28'h000_0000, p1_q_value__5_squeezed_comb});
  assign p1_sdiv_862_comb = sdiv_32b({{20{p1_array_index_834_comb[11]}}, p1_array_index_834_comb}, {28'h000_0000, p1_q_value__6_squeezed_comb});
  assign p1_sdiv_863_comb = sdiv_32b({{20{p1_array_index_837_comb[11]}}, p1_array_index_837_comb}, {28'h000_0000, p1_q_value__7_squeezed_comb});
  assign p1_divided_squeezed_comb = p0_quantize_off ? p1_array_index_816_comb : p1_sdiv_856_comb[11:0];
  assign p1_divided__1_squeezed_comb = p0_quantize_off ? p1_array_index_819_comb : p1_sdiv_857_comb[11:0];
  assign p1_divided__2_squeezed_comb = p0_quantize_off ? p1_array_index_822_comb : p1_sdiv_858_comb[11:0];
  assign p1_divided__3_squeezed_comb = p0_quantize_off ? p1_array_index_825_comb : p1_sdiv_859_comb[11:0];
  assign p1_divided__4_squeezed_comb = p0_quantize_off ? p1_array_index_828_comb : p1_sdiv_860_comb[11:0];
  assign p1_divided__5_squeezed_comb = p0_quantize_off ? p1_array_index_831_comb : p1_sdiv_861_comb[11:0];
  assign p1_divided__6_squeezed_comb = p0_quantize_off ? p1_array_index_834_comb : p1_sdiv_862_comb[11:0];
  assign p1_divided__7_squeezed_comb = p0_quantize_off ? p1_array_index_837_comb : p1_sdiv_863_comb[11:0];
  assign p1_clipped_comb = $signed(p1_divided_squeezed_comb) > $signed(12'h0ff) ? 10'h0ff : ($signed(p1_divided_squeezed_comb) < $signed(12'hf01) ? 10'h301 : p1_divided_squeezed_comb[9:0]);
  assign p1_clipped__1_comb = $signed(p1_divided__1_squeezed_comb) > $signed(12'h0ff) ? 10'h0ff : ($signed(p1_divided__1_squeezed_comb) < $signed(12'hf01) ? 10'h301 : p1_divided__1_squeezed_comb[9:0]);
  assign p1_clipped__2_comb = $signed(p1_divided__2_squeezed_comb) > $signed(12'h0ff) ? 10'h0ff : ($signed(p1_divided__2_squeezed_comb) < $signed(12'hf01) ? 10'h301 : p1_divided__2_squeezed_comb[9:0]);
  assign p1_clipped__3_comb = $signed(p1_divided__3_squeezed_comb) > $signed(12'h0ff) ? 10'h0ff : ($signed(p1_divided__3_squeezed_comb) < $signed(12'hf01) ? 10'h301 : p1_divided__3_squeezed_comb[9:0]);
  assign p1_clipped__4_comb = $signed(p1_divided__4_squeezed_comb) > $signed(12'h0ff) ? 10'h0ff : ($signed(p1_divided__4_squeezed_comb) < $signed(12'hf01) ? 10'h301 : p1_divided__4_squeezed_comb[9:0]);
  assign p1_clipped__5_comb = $signed(p1_divided__5_squeezed_comb) > $signed(12'h0ff) ? 10'h0ff : ($signed(p1_divided__5_squeezed_comb) < $signed(12'hf01) ? 10'h301 : p1_divided__5_squeezed_comb[9:0]);
  assign p1_clipped__6_comb = $signed(p1_divided__6_squeezed_comb) > $signed(12'h0ff) ? 10'h0ff : ($signed(p1_divided__6_squeezed_comb) < $signed(12'hf01) ? 10'h301 : p1_divided__6_squeezed_comb[9:0]);
  assign p1_clipped__7_comb = $signed(p1_divided__7_squeezed_comb) > $signed(12'h0ff) ? 10'h0ff : ($signed(p1_divided__7_squeezed_comb) < $signed(12'hf01) ? 10'h301 : p1_divided__7_squeezed_comb[9:0]);
  assign p1_array_952_comb[0] = p1_clipped_comb;
  assign p1_array_952_comb[1] = p1_clipped__1_comb;
  assign p1_array_952_comb[2] = p1_clipped__2_comb;
  assign p1_array_952_comb[3] = p1_clipped__3_comb;
  assign p1_array_952_comb[4] = p1_clipped__4_comb;
  assign p1_array_952_comb[5] = p1_clipped__5_comb;
  assign p1_array_952_comb[6] = p1_clipped__6_comb;
  assign p1_array_952_comb[7] = p1_clipped__7_comb;

  // Registers for pipe stage 1:
  reg [9:0] p1_array_952[0:7];
  always @ (posedge clk) begin
    p1_array_952[0] <= p1_array_952_comb[0];
    p1_array_952[1] <= p1_array_952_comb[1];
    p1_array_952[2] <= p1_array_952_comb[2];
    p1_array_952[3] <= p1_array_952_comb[3];
    p1_array_952[4] <= p1_array_952_comb[4];
    p1_array_952[5] <= p1_array_952_comb[5];
    p1_array_952[6] <= p1_array_952_comb[6];
    p1_array_952[7] <= p1_array_952_comb[7];
  end
  assign out = {p1_array_952[7], p1_array_952[6], p1_array_952[5], p1_array_952[4], p1_array_952[3], p1_array_952[2], p1_array_952[1], p1_array_952[0]};
endmodule
