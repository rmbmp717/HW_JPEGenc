module Huffman_ACenc(
  input wire clk,
  input wire [511:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [35:0] out
);
  wire [4:0] literal_10818[0:251];
  assign literal_10818[0] = 5'h02;
  assign literal_10818[1] = 5'h02;
  assign literal_10818[2] = 5'h03;
  assign literal_10818[3] = 5'h04;
  assign literal_10818[4] = 5'h05;
  assign literal_10818[5] = 5'h07;
  assign literal_10818[6] = 5'h08;
  assign literal_10818[7] = 5'h0e;
  assign literal_10818[8] = 5'h10;
  assign literal_10818[9] = 5'h10;
  assign literal_10818[10] = 5'h10;
  assign literal_10818[11] = 5'h00;
  assign literal_10818[12] = 5'h00;
  assign literal_10818[13] = 5'h00;
  assign literal_10818[14] = 5'h00;
  assign literal_10818[15] = 5'h00;
  assign literal_10818[16] = 5'h00;
  assign literal_10818[17] = 5'h03;
  assign literal_10818[18] = 5'h06;
  assign literal_10818[19] = 5'h07;
  assign literal_10818[20] = 5'h09;
  assign literal_10818[21] = 5'h0b;
  assign literal_10818[22] = 5'h0d;
  assign literal_10818[23] = 5'h10;
  assign literal_10818[24] = 5'h10;
  assign literal_10818[25] = 5'h10;
  assign literal_10818[26] = 5'h10;
  assign literal_10818[27] = 5'h00;
  assign literal_10818[28] = 5'h00;
  assign literal_10818[29] = 5'h00;
  assign literal_10818[30] = 5'h00;
  assign literal_10818[31] = 5'h00;
  assign literal_10818[32] = 5'h00;
  assign literal_10818[33] = 5'h05;
  assign literal_10818[34] = 5'h07;
  assign literal_10818[35] = 5'h0a;
  assign literal_10818[36] = 5'h0c;
  assign literal_10818[37] = 5'h0d;
  assign literal_10818[38] = 5'h10;
  assign literal_10818[39] = 5'h10;
  assign literal_10818[40] = 5'h10;
  assign literal_10818[41] = 5'h10;
  assign literal_10818[42] = 5'h10;
  assign literal_10818[43] = 5'h00;
  assign literal_10818[44] = 5'h00;
  assign literal_10818[45] = 5'h00;
  assign literal_10818[46] = 5'h00;
  assign literal_10818[47] = 5'h00;
  assign literal_10818[48] = 5'h00;
  assign literal_10818[49] = 5'h06;
  assign literal_10818[50] = 5'h08;
  assign literal_10818[51] = 5'h0b;
  assign literal_10818[52] = 5'h0c;
  assign literal_10818[53] = 5'h0f;
  assign literal_10818[54] = 5'h10;
  assign literal_10818[55] = 5'h10;
  assign literal_10818[56] = 5'h10;
  assign literal_10818[57] = 5'h10;
  assign literal_10818[58] = 5'h10;
  assign literal_10818[59] = 5'h00;
  assign literal_10818[60] = 5'h00;
  assign literal_10818[61] = 5'h00;
  assign literal_10818[62] = 5'h00;
  assign literal_10818[63] = 5'h00;
  assign literal_10818[64] = 5'h00;
  assign literal_10818[65] = 5'h06;
  assign literal_10818[66] = 5'h0a;
  assign literal_10818[67] = 5'h0c;
  assign literal_10818[68] = 5'h0f;
  assign literal_10818[69] = 5'h10;
  assign literal_10818[70] = 5'h10;
  assign literal_10818[71] = 5'h10;
  assign literal_10818[72] = 5'h10;
  assign literal_10818[73] = 5'h10;
  assign literal_10818[74] = 5'h10;
  assign literal_10818[75] = 5'h00;
  assign literal_10818[76] = 5'h00;
  assign literal_10818[77] = 5'h00;
  assign literal_10818[78] = 5'h00;
  assign literal_10818[79] = 5'h00;
  assign literal_10818[80] = 5'h00;
  assign literal_10818[81] = 5'h07;
  assign literal_10818[82] = 5'h0b;
  assign literal_10818[83] = 5'h0d;
  assign literal_10818[84] = 5'h10;
  assign literal_10818[85] = 5'h10;
  assign literal_10818[86] = 5'h10;
  assign literal_10818[87] = 5'h10;
  assign literal_10818[88] = 5'h10;
  assign literal_10818[89] = 5'h10;
  assign literal_10818[90] = 5'h10;
  assign literal_10818[91] = 5'h00;
  assign literal_10818[92] = 5'h00;
  assign literal_10818[93] = 5'h00;
  assign literal_10818[94] = 5'h00;
  assign literal_10818[95] = 5'h00;
  assign literal_10818[96] = 5'h00;
  assign literal_10818[97] = 5'h07;
  assign literal_10818[98] = 5'h0b;
  assign literal_10818[99] = 5'h0d;
  assign literal_10818[100] = 5'h10;
  assign literal_10818[101] = 5'h10;
  assign literal_10818[102] = 5'h10;
  assign literal_10818[103] = 5'h10;
  assign literal_10818[104] = 5'h10;
  assign literal_10818[105] = 5'h10;
  assign literal_10818[106] = 5'h10;
  assign literal_10818[107] = 5'h00;
  assign literal_10818[108] = 5'h00;
  assign literal_10818[109] = 5'h00;
  assign literal_10818[110] = 5'h00;
  assign literal_10818[111] = 5'h00;
  assign literal_10818[112] = 5'h00;
  assign literal_10818[113] = 5'h08;
  assign literal_10818[114] = 5'h0b;
  assign literal_10818[115] = 5'h0e;
  assign literal_10818[116] = 5'h10;
  assign literal_10818[117] = 5'h10;
  assign literal_10818[118] = 5'h10;
  assign literal_10818[119] = 5'h10;
  assign literal_10818[120] = 5'h10;
  assign literal_10818[121] = 5'h10;
  assign literal_10818[122] = 5'h10;
  assign literal_10818[123] = 5'h00;
  assign literal_10818[124] = 5'h00;
  assign literal_10818[125] = 5'h00;
  assign literal_10818[126] = 5'h00;
  assign literal_10818[127] = 5'h00;
  assign literal_10818[128] = 5'h00;
  assign literal_10818[129] = 5'h08;
  assign literal_10818[130] = 5'h0c;
  assign literal_10818[131] = 5'h10;
  assign literal_10818[132] = 5'h10;
  assign literal_10818[133] = 5'h10;
  assign literal_10818[134] = 5'h10;
  assign literal_10818[135] = 5'h10;
  assign literal_10818[136] = 5'h10;
  assign literal_10818[137] = 5'h10;
  assign literal_10818[138] = 5'h10;
  assign literal_10818[139] = 5'h00;
  assign literal_10818[140] = 5'h00;
  assign literal_10818[141] = 5'h00;
  assign literal_10818[142] = 5'h00;
  assign literal_10818[143] = 5'h00;
  assign literal_10818[144] = 5'h00;
  assign literal_10818[145] = 5'h08;
  assign literal_10818[146] = 5'h0d;
  assign literal_10818[147] = 5'h10;
  assign literal_10818[148] = 5'h10;
  assign literal_10818[149] = 5'h10;
  assign literal_10818[150] = 5'h10;
  assign literal_10818[151] = 5'h10;
  assign literal_10818[152] = 5'h10;
  assign literal_10818[153] = 5'h10;
  assign literal_10818[154] = 5'h10;
  assign literal_10818[155] = 5'h00;
  assign literal_10818[156] = 5'h00;
  assign literal_10818[157] = 5'h00;
  assign literal_10818[158] = 5'h00;
  assign literal_10818[159] = 5'h00;
  assign literal_10818[160] = 5'h00;
  assign literal_10818[161] = 5'h09;
  assign literal_10818[162] = 5'h0d;
  assign literal_10818[163] = 5'h10;
  assign literal_10818[164] = 5'h10;
  assign literal_10818[165] = 5'h10;
  assign literal_10818[166] = 5'h10;
  assign literal_10818[167] = 5'h10;
  assign literal_10818[168] = 5'h10;
  assign literal_10818[169] = 5'h10;
  assign literal_10818[170] = 5'h10;
  assign literal_10818[171] = 5'h00;
  assign literal_10818[172] = 5'h00;
  assign literal_10818[173] = 5'h00;
  assign literal_10818[174] = 5'h00;
  assign literal_10818[175] = 5'h00;
  assign literal_10818[176] = 5'h00;
  assign literal_10818[177] = 5'h09;
  assign literal_10818[178] = 5'h0d;
  assign literal_10818[179] = 5'h10;
  assign literal_10818[180] = 5'h10;
  assign literal_10818[181] = 5'h10;
  assign literal_10818[182] = 5'h10;
  assign literal_10818[183] = 5'h10;
  assign literal_10818[184] = 5'h10;
  assign literal_10818[185] = 5'h10;
  assign literal_10818[186] = 5'h10;
  assign literal_10818[187] = 5'h00;
  assign literal_10818[188] = 5'h00;
  assign literal_10818[189] = 5'h00;
  assign literal_10818[190] = 5'h00;
  assign literal_10818[191] = 5'h00;
  assign literal_10818[192] = 5'h00;
  assign literal_10818[193] = 5'h0a;
  assign literal_10818[194] = 5'h0d;
  assign literal_10818[195] = 5'h10;
  assign literal_10818[196] = 5'h10;
  assign literal_10818[197] = 5'h10;
  assign literal_10818[198] = 5'h10;
  assign literal_10818[199] = 5'h10;
  assign literal_10818[200] = 5'h10;
  assign literal_10818[201] = 5'h10;
  assign literal_10818[202] = 5'h10;
  assign literal_10818[203] = 5'h00;
  assign literal_10818[204] = 5'h00;
  assign literal_10818[205] = 5'h00;
  assign literal_10818[206] = 5'h00;
  assign literal_10818[207] = 5'h00;
  assign literal_10818[208] = 5'h00;
  assign literal_10818[209] = 5'h0a;
  assign literal_10818[210] = 5'h0e;
  assign literal_10818[211] = 5'h10;
  assign literal_10818[212] = 5'h10;
  assign literal_10818[213] = 5'h10;
  assign literal_10818[214] = 5'h10;
  assign literal_10818[215] = 5'h10;
  assign literal_10818[216] = 5'h10;
  assign literal_10818[217] = 5'h10;
  assign literal_10818[218] = 5'h10;
  assign literal_10818[219] = 5'h00;
  assign literal_10818[220] = 5'h00;
  assign literal_10818[221] = 5'h00;
  assign literal_10818[222] = 5'h00;
  assign literal_10818[223] = 5'h00;
  assign literal_10818[224] = 5'h00;
  assign literal_10818[225] = 5'h0a;
  assign literal_10818[226] = 5'h0f;
  assign literal_10818[227] = 5'h10;
  assign literal_10818[228] = 5'h10;
  assign literal_10818[229] = 5'h10;
  assign literal_10818[230] = 5'h10;
  assign literal_10818[231] = 5'h10;
  assign literal_10818[232] = 5'h10;
  assign literal_10818[233] = 5'h10;
  assign literal_10818[234] = 5'h10;
  assign literal_10818[235] = 5'h00;
  assign literal_10818[236] = 5'h00;
  assign literal_10818[237] = 5'h00;
  assign literal_10818[238] = 5'h00;
  assign literal_10818[239] = 5'h00;
  assign literal_10818[240] = 5'h09;
  assign literal_10818[241] = 5'h0b;
  assign literal_10818[242] = 5'h10;
  assign literal_10818[243] = 5'h10;
  assign literal_10818[244] = 5'h10;
  assign literal_10818[245] = 5'h10;
  assign literal_10818[246] = 5'h10;
  assign literal_10818[247] = 5'h10;
  assign literal_10818[248] = 5'h10;
  assign literal_10818[249] = 5'h10;
  assign literal_10818[250] = 5'h10;
  assign literal_10818[251] = 5'h00;
  wire [15:0] literal_10822[0:251];
  assign literal_10822[0] = 16'h0001;
  assign literal_10822[1] = 16'h0000;
  assign literal_10822[2] = 16'h0004;
  assign literal_10822[3] = 16'h000c;
  assign literal_10822[4] = 16'h001a;
  assign literal_10822[5] = 16'h0076;
  assign literal_10822[6] = 16'h00f6;
  assign literal_10822[7] = 16'h3fe0;
  assign literal_10822[8] = 16'hff96;
  assign literal_10822[9] = 16'hff97;
  assign literal_10822[10] = 16'hff98;
  assign literal_10822[11] = 16'h0000;
  assign literal_10822[12] = 16'h0000;
  assign literal_10822[13] = 16'h0000;
  assign literal_10822[14] = 16'h0000;
  assign literal_10822[15] = 16'h0000;
  assign literal_10822[16] = 16'h0000;
  assign literal_10822[17] = 16'h0005;
  assign literal_10822[18] = 16'h0038;
  assign literal_10822[19] = 16'h0078;
  assign literal_10822[20] = 16'h01f9;
  assign literal_10822[21] = 16'h07f2;
  assign literal_10822[22] = 16'h1fe8;
  assign literal_10822[23] = 16'hff93;
  assign literal_10822[24] = 16'hff99;
  assign literal_10822[25] = 16'hff9a;
  assign literal_10822[26] = 16'hff9e;
  assign literal_10822[27] = 16'h0000;
  assign literal_10822[28] = 16'h0000;
  assign literal_10822[29] = 16'h0000;
  assign literal_10822[30] = 16'h0000;
  assign literal_10822[31] = 16'h0000;
  assign literal_10822[32] = 16'h0000;
  assign literal_10822[33] = 16'h001b;
  assign literal_10822[34] = 16'h007a;
  assign literal_10822[35] = 16'h03f7;
  assign literal_10822[36] = 16'h0ff0;
  assign literal_10822[37] = 16'h1feb;
  assign literal_10822[38] = 16'hff9b;
  assign literal_10822[39] = 16'hff9f;
  assign literal_10822[40] = 16'hffa8;
  assign literal_10822[41] = 16'hffa9;
  assign literal_10822[42] = 16'hfff1;
  assign literal_10822[43] = 16'h0000;
  assign literal_10822[44] = 16'h0000;
  assign literal_10822[45] = 16'h0000;
  assign literal_10822[46] = 16'h0000;
  assign literal_10822[47] = 16'h0000;
  assign literal_10822[48] = 16'h0000;
  assign literal_10822[49] = 16'h0039;
  assign literal_10822[50] = 16'h00fa;
  assign literal_10822[51] = 16'h07f7;
  assign literal_10822[52] = 16'h0ff1;
  assign literal_10822[53] = 16'h7fc6;
  assign literal_10822[54] = 16'hff9c;
  assign literal_10822[55] = 16'hffa3;
  assign literal_10822[56] = 16'hffd7;
  assign literal_10822[57] = 16'hffe4;
  assign literal_10822[58] = 16'hfff2;
  assign literal_10822[59] = 16'h0000;
  assign literal_10822[60] = 16'h0000;
  assign literal_10822[61] = 16'h0000;
  assign literal_10822[62] = 16'h0000;
  assign literal_10822[63] = 16'h0000;
  assign literal_10822[64] = 16'h0000;
  assign literal_10822[65] = 16'h003a;
  assign literal_10822[66] = 16'h03f8;
  assign literal_10822[67] = 16'h0ff2;
  assign literal_10822[68] = 16'h7fc8;
  assign literal_10822[69] = 16'hff9d;
  assign literal_10822[70] = 16'hffbf;
  assign literal_10822[71] = 16'hffcb;
  assign literal_10822[72] = 16'hffd8;
  assign literal_10822[73] = 16'hffe5;
  assign literal_10822[74] = 16'hfff3;
  assign literal_10822[75] = 16'h0000;
  assign literal_10822[76] = 16'h0000;
  assign literal_10822[77] = 16'h0000;
  assign literal_10822[78] = 16'h0000;
  assign literal_10822[79] = 16'h0000;
  assign literal_10822[80] = 16'h0000;
  assign literal_10822[81] = 16'h0077;
  assign literal_10822[82] = 16'h07f3;
  assign literal_10822[83] = 16'h1fea;
  assign literal_10822[84] = 16'hff94;
  assign literal_10822[85] = 16'hffa2;
  assign literal_10822[86] = 16'hffc0;
  assign literal_10822[87] = 16'hffcc;
  assign literal_10822[88] = 16'hffd9;
  assign literal_10822[89] = 16'hffe6;
  assign literal_10822[90] = 16'hfff4;
  assign literal_10822[91] = 16'h0000;
  assign literal_10822[92] = 16'h0000;
  assign literal_10822[93] = 16'h0000;
  assign literal_10822[94] = 16'h0000;
  assign literal_10822[95] = 16'h0000;
  assign literal_10822[96] = 16'h0000;
  assign literal_10822[97] = 16'h0079;
  assign literal_10822[98] = 16'h07f4;
  assign literal_10822[99] = 16'h1fed;
  assign literal_10822[100] = 16'hffa0;
  assign literal_10822[101] = 16'hffb5;
  assign literal_10822[102] = 16'hffc1;
  assign literal_10822[103] = 16'hffcd;
  assign literal_10822[104] = 16'hffda;
  assign literal_10822[105] = 16'hffe7;
  assign literal_10822[106] = 16'hfff5;
  assign literal_10822[107] = 16'h0000;
  assign literal_10822[108] = 16'h0000;
  assign literal_10822[109] = 16'h0000;
  assign literal_10822[110] = 16'h0000;
  assign literal_10822[111] = 16'h0000;
  assign literal_10822[112] = 16'h0000;
  assign literal_10822[113] = 16'h00f7;
  assign literal_10822[114] = 16'h07f5;
  assign literal_10822[115] = 16'h3fe1;
  assign literal_10822[116] = 16'hffa1;
  assign literal_10822[117] = 16'hffb6;
  assign literal_10822[118] = 16'hffc2;
  assign literal_10822[119] = 16'hffce;
  assign literal_10822[120] = 16'hffdb;
  assign literal_10822[121] = 16'hffe8;
  assign literal_10822[122] = 16'hfff6;
  assign literal_10822[123] = 16'h0000;
  assign literal_10822[124] = 16'h0000;
  assign literal_10822[125] = 16'h0000;
  assign literal_10822[126] = 16'h0000;
  assign literal_10822[127] = 16'h0000;
  assign literal_10822[128] = 16'h0000;
  assign literal_10822[129] = 16'h00f8;
  assign literal_10822[130] = 16'h0ff3;
  assign literal_10822[131] = 16'hff92;
  assign literal_10822[132] = 16'hffad;
  assign literal_10822[133] = 16'hffb7;
  assign literal_10822[134] = 16'hffc3;
  assign literal_10822[135] = 16'hffcf;
  assign literal_10822[136] = 16'hffdc;
  assign literal_10822[137] = 16'hffe9;
  assign literal_10822[138] = 16'hfff7;
  assign literal_10822[139] = 16'h0000;
  assign literal_10822[140] = 16'h0000;
  assign literal_10822[141] = 16'h0000;
  assign literal_10822[142] = 16'h0000;
  assign literal_10822[143] = 16'h0000;
  assign literal_10822[144] = 16'h0000;
  assign literal_10822[145] = 16'h00f9;
  assign literal_10822[146] = 16'h1fe9;
  assign literal_10822[147] = 16'hff95;
  assign literal_10822[148] = 16'hffae;
  assign literal_10822[149] = 16'hffb8;
  assign literal_10822[150] = 16'hffc4;
  assign literal_10822[151] = 16'hffd0;
  assign literal_10822[152] = 16'hffdd;
  assign literal_10822[153] = 16'hffea;
  assign literal_10822[154] = 16'hfff8;
  assign literal_10822[155] = 16'h0000;
  assign literal_10822[156] = 16'h0000;
  assign literal_10822[157] = 16'h0000;
  assign literal_10822[158] = 16'h0000;
  assign literal_10822[159] = 16'h0000;
  assign literal_10822[160] = 16'h0000;
  assign literal_10822[161] = 16'h01f6;
  assign literal_10822[162] = 16'h1fec;
  assign literal_10822[163] = 16'hffa5;
  assign literal_10822[164] = 16'hffaf;
  assign literal_10822[165] = 16'hffb9;
  assign literal_10822[166] = 16'hffc5;
  assign literal_10822[167] = 16'hffd1;
  assign literal_10822[168] = 16'hffde;
  assign literal_10822[169] = 16'hffeb;
  assign literal_10822[170] = 16'hfff9;
  assign literal_10822[171] = 16'h0000;
  assign literal_10822[172] = 16'h0000;
  assign literal_10822[173] = 16'h0000;
  assign literal_10822[174] = 16'h0000;
  assign literal_10822[175] = 16'h0000;
  assign literal_10822[176] = 16'h0000;
  assign literal_10822[177] = 16'h01f7;
  assign literal_10822[178] = 16'h1fee;
  assign literal_10822[179] = 16'hffa6;
  assign literal_10822[180] = 16'hffb0;
  assign literal_10822[181] = 16'hffba;
  assign literal_10822[182] = 16'hffc6;
  assign literal_10822[183] = 16'hffd2;
  assign literal_10822[184] = 16'hffdf;
  assign literal_10822[185] = 16'hffec;
  assign literal_10822[186] = 16'hfffa;
  assign literal_10822[187] = 16'h0000;
  assign literal_10822[188] = 16'h0000;
  assign literal_10822[189] = 16'h0000;
  assign literal_10822[190] = 16'h0000;
  assign literal_10822[191] = 16'h0000;
  assign literal_10822[192] = 16'h0000;
  assign literal_10822[193] = 16'h03f4;
  assign literal_10822[194] = 16'h1fef;
  assign literal_10822[195] = 16'hffa7;
  assign literal_10822[196] = 16'hffb1;
  assign literal_10822[197] = 16'hffbb;
  assign literal_10822[198] = 16'hffc7;
  assign literal_10822[199] = 16'hffd3;
  assign literal_10822[200] = 16'hffe0;
  assign literal_10822[201] = 16'hffed;
  assign literal_10822[202] = 16'hfffb;
  assign literal_10822[203] = 16'h0000;
  assign literal_10822[204] = 16'h0000;
  assign literal_10822[205] = 16'h0000;
  assign literal_10822[206] = 16'h0000;
  assign literal_10822[207] = 16'h0000;
  assign literal_10822[208] = 16'h0000;
  assign literal_10822[209] = 16'h03f5;
  assign literal_10822[210] = 16'h3fe2;
  assign literal_10822[211] = 16'hffaa;
  assign literal_10822[212] = 16'hffb2;
  assign literal_10822[213] = 16'hffbc;
  assign literal_10822[214] = 16'hffc8;
  assign literal_10822[215] = 16'hffd4;
  assign literal_10822[216] = 16'hffe1;
  assign literal_10822[217] = 16'hffee;
  assign literal_10822[218] = 16'hfffc;
  assign literal_10822[219] = 16'h0000;
  assign literal_10822[220] = 16'h0000;
  assign literal_10822[221] = 16'h0000;
  assign literal_10822[222] = 16'h0000;
  assign literal_10822[223] = 16'h0000;
  assign literal_10822[224] = 16'h0000;
  assign literal_10822[225] = 16'h03f6;
  assign literal_10822[226] = 16'h7fc7;
  assign literal_10822[227] = 16'hffab;
  assign literal_10822[228] = 16'hffb3;
  assign literal_10822[229] = 16'hffbd;
  assign literal_10822[230] = 16'hffc9;
  assign literal_10822[231] = 16'hffd5;
  assign literal_10822[232] = 16'hffe2;
  assign literal_10822[233] = 16'hffef;
  assign literal_10822[234] = 16'hfffd;
  assign literal_10822[235] = 16'h0000;
  assign literal_10822[236] = 16'h0000;
  assign literal_10822[237] = 16'h0000;
  assign literal_10822[238] = 16'h0000;
  assign literal_10822[239] = 16'h0000;
  assign literal_10822[240] = 16'h01f8;
  assign literal_10822[241] = 16'h07f6;
  assign literal_10822[242] = 16'hffa4;
  assign literal_10822[243] = 16'hffac;
  assign literal_10822[244] = 16'hffb4;
  assign literal_10822[245] = 16'hffbe;
  assign literal_10822[246] = 16'hffca;
  assign literal_10822[247] = 16'hffd6;
  assign literal_10822[248] = 16'hffe3;
  assign literal_10822[249] = 16'hfff0;
  assign literal_10822[250] = 16'hfffe;
  assign literal_10822[251] = 16'h0000;
  wire [7:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[7:0];
  assign matrix_unflattened[0][1] = matrix[15:8];
  assign matrix_unflattened[0][2] = matrix[23:16];
  assign matrix_unflattened[0][3] = matrix[31:24];
  assign matrix_unflattened[0][4] = matrix[39:32];
  assign matrix_unflattened[0][5] = matrix[47:40];
  assign matrix_unflattened[0][6] = matrix[55:48];
  assign matrix_unflattened[0][7] = matrix[63:56];
  assign matrix_unflattened[1][0] = matrix[71:64];
  assign matrix_unflattened[1][1] = matrix[79:72];
  assign matrix_unflattened[1][2] = matrix[87:80];
  assign matrix_unflattened[1][3] = matrix[95:88];
  assign matrix_unflattened[1][4] = matrix[103:96];
  assign matrix_unflattened[1][5] = matrix[111:104];
  assign matrix_unflattened[1][6] = matrix[119:112];
  assign matrix_unflattened[1][7] = matrix[127:120];
  assign matrix_unflattened[2][0] = matrix[135:128];
  assign matrix_unflattened[2][1] = matrix[143:136];
  assign matrix_unflattened[2][2] = matrix[151:144];
  assign matrix_unflattened[2][3] = matrix[159:152];
  assign matrix_unflattened[2][4] = matrix[167:160];
  assign matrix_unflattened[2][5] = matrix[175:168];
  assign matrix_unflattened[2][6] = matrix[183:176];
  assign matrix_unflattened[2][7] = matrix[191:184];
  assign matrix_unflattened[3][0] = matrix[199:192];
  assign matrix_unflattened[3][1] = matrix[207:200];
  assign matrix_unflattened[3][2] = matrix[215:208];
  assign matrix_unflattened[3][3] = matrix[223:216];
  assign matrix_unflattened[3][4] = matrix[231:224];
  assign matrix_unflattened[3][5] = matrix[239:232];
  assign matrix_unflattened[3][6] = matrix[247:240];
  assign matrix_unflattened[3][7] = matrix[255:248];
  assign matrix_unflattened[4][0] = matrix[263:256];
  assign matrix_unflattened[4][1] = matrix[271:264];
  assign matrix_unflattened[4][2] = matrix[279:272];
  assign matrix_unflattened[4][3] = matrix[287:280];
  assign matrix_unflattened[4][4] = matrix[295:288];
  assign matrix_unflattened[4][5] = matrix[303:296];
  assign matrix_unflattened[4][6] = matrix[311:304];
  assign matrix_unflattened[4][7] = matrix[319:312];
  assign matrix_unflattened[5][0] = matrix[327:320];
  assign matrix_unflattened[5][1] = matrix[335:328];
  assign matrix_unflattened[5][2] = matrix[343:336];
  assign matrix_unflattened[5][3] = matrix[351:344];
  assign matrix_unflattened[5][4] = matrix[359:352];
  assign matrix_unflattened[5][5] = matrix[367:360];
  assign matrix_unflattened[5][6] = matrix[375:368];
  assign matrix_unflattened[5][7] = matrix[383:376];
  assign matrix_unflattened[6][0] = matrix[391:384];
  assign matrix_unflattened[6][1] = matrix[399:392];
  assign matrix_unflattened[6][2] = matrix[407:400];
  assign matrix_unflattened[6][3] = matrix[415:408];
  assign matrix_unflattened[6][4] = matrix[423:416];
  assign matrix_unflattened[6][5] = matrix[431:424];
  assign matrix_unflattened[6][6] = matrix[439:432];
  assign matrix_unflattened[6][7] = matrix[447:440];
  assign matrix_unflattened[7][0] = matrix[455:448];
  assign matrix_unflattened[7][1] = matrix[463:456];
  assign matrix_unflattened[7][2] = matrix[471:464];
  assign matrix_unflattened[7][3] = matrix[479:472];
  assign matrix_unflattened[7][4] = matrix[487:480];
  assign matrix_unflattened[7][5] = matrix[495:488];
  assign matrix_unflattened[7][6] = matrix[503:496];
  assign matrix_unflattened[7][7] = matrix[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_row0_comb[0:7];
  wire [7:0] p1_row1_comb[0:7];
  wire [7:0] p1_array_concat_9825_comb[0:15];
  wire [7:0] p1_row2_comb[0:7];
  wire [7:0] p1_array_concat_9828_comb[0:23];
  wire [7:0] p1_row3_comb[0:7];
  wire [2:0] p1_idx_u8__4_squeezed_comb;
  wire [7:0] p1_array_concat_9831_comb[0:31];
  wire [7:0] p1_row4_comb[0:7];
  wire [2:0] p1_idx_u8__5_squeezed_comb;
  wire [7:0] p1_array_concat_9834_comb[0:39];
  wire [7:0] p1_row5_comb[0:7];
  wire [2:0] p1_idx_u8__6_squeezed_comb;
  wire [7:0] p1_idx_u8__13_comb;
  wire [7:0] p1_array_concat_9840_comb[0:47];
  wire [7:0] p1_row6_comb[0:7];
  wire [2:0] p1_idx_u8__7_squeezed_comb;
  wire [6:0] p1_add_9843_comb;
  wire [7:0] p1_actual_index__13_comb;
  wire [7:0] p1_array_concat_9847_comb[0:55];
  wire [7:0] p1_row7_comb[0:7];
  wire [5:0] p1_add_9852_comb;
  wire [7:0] p1_flat_comb[0:63];
  wire [7:0] p1_actual_index__14_comb;
  wire [7:0] p1_idx_u8__11_comb;
  wire [7:0] p1_actual_index__12_comb;
  wire [7:0] p1_actual_index__11_comb;
  wire [7:0] p1_and_9871_comb;
  wire [7:0] p1_idx_u8__1_comb;
  wire [7:0] p1_idx_u8__3_comb;
  wire [7:0] p1_idx_u8__5_comb;
  wire [7:0] p1_idx_u8__7_comb;
  wire [7:0] p1_idx_u8__9_comb;
  wire [6:0] p1_add_9876_comb;
  wire [7:0] p1_and_9879_comb;
  wire p1_eq_9882_comb;
  wire [7:0] p1_and_9883_comb;
  wire [7:0] p1_actual_index__1_comb;
  wire [6:0] p1_add_9967_comb;
  wire [7:0] p1_actual_index__3_comb;
  wire [5:0] p1_add_9949_comb;
  wire [7:0] p1_actual_index__5_comb;
  wire [6:0] p1_add_9929_comb;
  wire [7:0] p1_actual_index__7_comb;
  wire [7:0] p1_actual_index__9_comb;
  wire [7:0] p1_idx_u8__15_comb;
  wire [7:0] p1_idx_u8__17_comb;
  wire [7:0] p1_idx_u8__19_comb;
  wire [7:0] p1_idx_u8__21_comb;
  wire [7:0] p1_idx_u8__23_comb;
  wire [7:0] p1_idx_u8__25_comb;
  wire [7:0] p1_idx_u8__27_comb;
  wire [7:0] p1_idx_u8__29_comb;
  wire [7:0] p1_idx_u8__31_comb;
  wire [7:0] p1_idx_u8__33_comb;
  wire [7:0] p1_idx_u8__35_comb;
  wire [7:0] p1_idx_u8__37_comb;
  wire [7:0] p1_idx_u8__39_comb;
  wire [7:0] p1_idx_u8__41_comb;
  wire [7:0] p1_idx_u8__43_comb;
  wire [7:0] p1_idx_u8__45_comb;
  wire [7:0] p1_idx_u8__47_comb;
  wire [7:0] p1_idx_u8__49_comb;
  wire [7:0] p1_idx_u8__51_comb;
  wire [7:0] p1_idx_u8__53_comb;
  wire [7:0] p1_idx_u8__55_comb;
  wire [7:0] p1_idx_u8__57_comb;
  wire [7:0] p1_idx_u8__59_comb;
  wire [7:0] p1_idx_u8__61_comb;
  wire p1_ne_9891_comb;
  wire [1:0] p1_idx_u8__1_squeezed_comb;
  wire p1_eq_9894_comb;
  wire [4:0] p1_add_9895_comb;
  wire [7:0] p1_actual_index__15_comb;
  wire [3:0] p1_add_10070_comb;
  wire [7:0] p1_actual_index__17_comb;
  wire [6:0] p1_add_10072_comb;
  wire [7:0] p1_actual_index__19_comb;
  wire [5:0] p1_add_10074_comb;
  wire [7:0] p1_actual_index__21_comb;
  wire [6:0] p1_add_10076_comb;
  wire [7:0] p1_actual_index__23_comb;
  wire [4:0] p1_add_10078_comb;
  wire [7:0] p1_actual_index__25_comb;
  wire [6:0] p1_add_10080_comb;
  wire [7:0] p1_actual_index__27_comb;
  wire [5:0] p1_add_10082_comb;
  wire [7:0] p1_actual_index__29_comb;
  wire [6:0] p1_add_10084_comb;
  wire [7:0] p1_actual_index__31_comb;
  wire [2:0] p1_add_10086_comb;
  wire [7:0] p1_actual_index__33_comb;
  wire [6:0] p1_add_10088_comb;
  wire [7:0] p1_actual_index__35_comb;
  wire [5:0] p1_add_10090_comb;
  wire [7:0] p1_actual_index__37_comb;
  wire [6:0] p1_add_10092_comb;
  wire [7:0] p1_actual_index__39_comb;
  wire [4:0] p1_add_10094_comb;
  wire [7:0] p1_actual_index__41_comb;
  wire [6:0] p1_add_10096_comb;
  wire [7:0] p1_actual_index__43_comb;
  wire [5:0] p1_add_10098_comb;
  wire [7:0] p1_actual_index__45_comb;
  wire [6:0] p1_add_10100_comb;
  wire [7:0] p1_actual_index__47_comb;
  wire [3:0] p1_add_10102_comb;
  wire [7:0] p1_actual_index__49_comb;
  wire [6:0] p1_add_10104_comb;
  wire [7:0] p1_actual_index__51_comb;
  wire [5:0] p1_add_10106_comb;
  wire [7:0] p1_actual_index__53_comb;
  wire [6:0] p1_add_10108_comb;
  wire [7:0] p1_actual_index__55_comb;
  wire [4:0] p1_add_10110_comb;
  wire [7:0] p1_actual_index__57_comb;
  wire [6:0] p1_add_10112_comb;
  wire [7:0] p1_actual_index__59_comb;
  wire [5:0] p1_add_10114_comb;
  wire [7:0] p1_actual_index__61_comb;
  wire [6:0] p1_add_10116_comb;
  wire [7:0] p1_actual_index__10_comb;
  wire [7:0] p1_actual_index__2_comb;
  wire [7:0] p1_actual_index__4_comb;
  wire [7:0] p1_actual_index__6_comb;
  wire [7:0] p1_and_9911_comb;
  wire [7:0] p1_actual_index__8_comb;
  wire [7:0] p1_actual_index__16_comb;
  wire [7:0] p1_actual_index__18_comb;
  wire [7:0] p1_actual_index__20_comb;
  wire [7:0] p1_actual_index__22_comb;
  wire [7:0] p1_actual_index__24_comb;
  wire [7:0] p1_actual_index__26_comb;
  wire [7:0] p1_actual_index__28_comb;
  wire [7:0] p1_actual_index__30_comb;
  wire [7:0] p1_actual_index__32_comb;
  wire [7:0] p1_actual_index__34_comb;
  wire [7:0] p1_actual_index__36_comb;
  wire [7:0] p1_actual_index__38_comb;
  wire [7:0] p1_actual_index__40_comb;
  wire [7:0] p1_actual_index__42_comb;
  wire [7:0] p1_actual_index__44_comb;
  wire [7:0] p1_actual_index__46_comb;
  wire [7:0] p1_actual_index__48_comb;
  wire [7:0] p1_actual_index__50_comb;
  wire [7:0] p1_actual_index__52_comb;
  wire [7:0] p1_actual_index__54_comb;
  wire [7:0] p1_actual_index__56_comb;
  wire [7:0] p1_actual_index__58_comb;
  wire [7:0] p1_actual_index__60_comb;
  wire [7:0] p1_actual_index__62_comb;
  wire [7:0] p1_and_9921_comb;
  wire p1_ne_9923_comb;
  wire [7:0] p1_and_10011_comb;
  wire [7:0] p1_and_10013_comb;
  wire [7:0] p1_and_10008_comb;
  wire [7:0] p1_and_10001_comb;
  wire [7:0] p1_and_9994_comb;
  wire [7:0] p1_and_9983_comb;
  wire [7:0] p1_and_9974_comb;
  wire [7:0] p1_and_9964_comb;
  wire [7:0] p1_and_9932_comb;
  wire p1_ne_9934_comb;
  wire [2:0] p1_sel_9935_comb;
  wire p1_ne_10016_comb;
  wire p1_ne_10017_comb;
  wire p1_ne_10015_comb;
  wire p1_ne_10010_comb;
  wire p1_ne_10003_comb;
  wire p1_ne_9996_comb;
  wire p1_ne_9985_comb;
  wire p1_ne_9976_comb;
  wire [7:0] p1_and_9937_comb;
  wire p1_ne_9944_comb;
  wire p1_not_10018_comb;
  wire p1_eq_9947_comb;
  wire [2:0] p1_sel_9956_comb;
  wire p1_and_10538_comb;
  wire [7:0] p1_value_comb;
  assign p1_row0_comb[0] = p0_matrix[3'h0][0];
  assign p1_row0_comb[1] = p0_matrix[3'h0][1];
  assign p1_row0_comb[2] = p0_matrix[3'h0][2];
  assign p1_row0_comb[3] = p0_matrix[3'h0][3];
  assign p1_row0_comb[4] = p0_matrix[3'h0][4];
  assign p1_row0_comb[5] = p0_matrix[3'h0][5];
  assign p1_row0_comb[6] = p0_matrix[3'h0][6];
  assign p1_row0_comb[7] = p0_matrix[3'h0][7];
  assign p1_row1_comb[0] = p0_matrix[3'h1][0];
  assign p1_row1_comb[1] = p0_matrix[3'h1][1];
  assign p1_row1_comb[2] = p0_matrix[3'h1][2];
  assign p1_row1_comb[3] = p0_matrix[3'h1][3];
  assign p1_row1_comb[4] = p0_matrix[3'h1][4];
  assign p1_row1_comb[5] = p0_matrix[3'h1][5];
  assign p1_row1_comb[6] = p0_matrix[3'h1][6];
  assign p1_row1_comb[7] = p0_matrix[3'h1][7];
  assign p1_array_concat_9825_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_9825_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_9825_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_9825_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_9825_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_9825_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_9825_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_9825_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_9825_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_9825_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_9825_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_9825_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_9825_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_9825_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_9825_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_9825_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_9828_comb[0] = p1_array_concat_9825_comb[0];
  assign p1_array_concat_9828_comb[1] = p1_array_concat_9825_comb[1];
  assign p1_array_concat_9828_comb[2] = p1_array_concat_9825_comb[2];
  assign p1_array_concat_9828_comb[3] = p1_array_concat_9825_comb[3];
  assign p1_array_concat_9828_comb[4] = p1_array_concat_9825_comb[4];
  assign p1_array_concat_9828_comb[5] = p1_array_concat_9825_comb[5];
  assign p1_array_concat_9828_comb[6] = p1_array_concat_9825_comb[6];
  assign p1_array_concat_9828_comb[7] = p1_array_concat_9825_comb[7];
  assign p1_array_concat_9828_comb[8] = p1_array_concat_9825_comb[8];
  assign p1_array_concat_9828_comb[9] = p1_array_concat_9825_comb[9];
  assign p1_array_concat_9828_comb[10] = p1_array_concat_9825_comb[10];
  assign p1_array_concat_9828_comb[11] = p1_array_concat_9825_comb[11];
  assign p1_array_concat_9828_comb[12] = p1_array_concat_9825_comb[12];
  assign p1_array_concat_9828_comb[13] = p1_array_concat_9825_comb[13];
  assign p1_array_concat_9828_comb[14] = p1_array_concat_9825_comb[14];
  assign p1_array_concat_9828_comb[15] = p1_array_concat_9825_comb[15];
  assign p1_array_concat_9828_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_9828_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_9828_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_9828_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_9828_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_9828_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_9828_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_9828_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_idx_u8__4_squeezed_comb = 3'h4;
  assign p1_array_concat_9831_comb[0] = p1_array_concat_9828_comb[0];
  assign p1_array_concat_9831_comb[1] = p1_array_concat_9828_comb[1];
  assign p1_array_concat_9831_comb[2] = p1_array_concat_9828_comb[2];
  assign p1_array_concat_9831_comb[3] = p1_array_concat_9828_comb[3];
  assign p1_array_concat_9831_comb[4] = p1_array_concat_9828_comb[4];
  assign p1_array_concat_9831_comb[5] = p1_array_concat_9828_comb[5];
  assign p1_array_concat_9831_comb[6] = p1_array_concat_9828_comb[6];
  assign p1_array_concat_9831_comb[7] = p1_array_concat_9828_comb[7];
  assign p1_array_concat_9831_comb[8] = p1_array_concat_9828_comb[8];
  assign p1_array_concat_9831_comb[9] = p1_array_concat_9828_comb[9];
  assign p1_array_concat_9831_comb[10] = p1_array_concat_9828_comb[10];
  assign p1_array_concat_9831_comb[11] = p1_array_concat_9828_comb[11];
  assign p1_array_concat_9831_comb[12] = p1_array_concat_9828_comb[12];
  assign p1_array_concat_9831_comb[13] = p1_array_concat_9828_comb[13];
  assign p1_array_concat_9831_comb[14] = p1_array_concat_9828_comb[14];
  assign p1_array_concat_9831_comb[15] = p1_array_concat_9828_comb[15];
  assign p1_array_concat_9831_comb[16] = p1_array_concat_9828_comb[16];
  assign p1_array_concat_9831_comb[17] = p1_array_concat_9828_comb[17];
  assign p1_array_concat_9831_comb[18] = p1_array_concat_9828_comb[18];
  assign p1_array_concat_9831_comb[19] = p1_array_concat_9828_comb[19];
  assign p1_array_concat_9831_comb[20] = p1_array_concat_9828_comb[20];
  assign p1_array_concat_9831_comb[21] = p1_array_concat_9828_comb[21];
  assign p1_array_concat_9831_comb[22] = p1_array_concat_9828_comb[22];
  assign p1_array_concat_9831_comb[23] = p1_array_concat_9828_comb[23];
  assign p1_array_concat_9831_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_9831_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_9831_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_9831_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_9831_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_9831_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_9831_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_9831_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[p1_idx_u8__4_squeezed_comb][0];
  assign p1_row4_comb[1] = p0_matrix[p1_idx_u8__4_squeezed_comb][1];
  assign p1_row4_comb[2] = p0_matrix[p1_idx_u8__4_squeezed_comb][2];
  assign p1_row4_comb[3] = p0_matrix[p1_idx_u8__4_squeezed_comb][3];
  assign p1_row4_comb[4] = p0_matrix[p1_idx_u8__4_squeezed_comb][4];
  assign p1_row4_comb[5] = p0_matrix[p1_idx_u8__4_squeezed_comb][5];
  assign p1_row4_comb[6] = p0_matrix[p1_idx_u8__4_squeezed_comb][6];
  assign p1_row4_comb[7] = p0_matrix[p1_idx_u8__4_squeezed_comb][7];
  assign p1_idx_u8__5_squeezed_comb = 3'h5;
  assign p1_array_concat_9834_comb[0] = p1_array_concat_9831_comb[0];
  assign p1_array_concat_9834_comb[1] = p1_array_concat_9831_comb[1];
  assign p1_array_concat_9834_comb[2] = p1_array_concat_9831_comb[2];
  assign p1_array_concat_9834_comb[3] = p1_array_concat_9831_comb[3];
  assign p1_array_concat_9834_comb[4] = p1_array_concat_9831_comb[4];
  assign p1_array_concat_9834_comb[5] = p1_array_concat_9831_comb[5];
  assign p1_array_concat_9834_comb[6] = p1_array_concat_9831_comb[6];
  assign p1_array_concat_9834_comb[7] = p1_array_concat_9831_comb[7];
  assign p1_array_concat_9834_comb[8] = p1_array_concat_9831_comb[8];
  assign p1_array_concat_9834_comb[9] = p1_array_concat_9831_comb[9];
  assign p1_array_concat_9834_comb[10] = p1_array_concat_9831_comb[10];
  assign p1_array_concat_9834_comb[11] = p1_array_concat_9831_comb[11];
  assign p1_array_concat_9834_comb[12] = p1_array_concat_9831_comb[12];
  assign p1_array_concat_9834_comb[13] = p1_array_concat_9831_comb[13];
  assign p1_array_concat_9834_comb[14] = p1_array_concat_9831_comb[14];
  assign p1_array_concat_9834_comb[15] = p1_array_concat_9831_comb[15];
  assign p1_array_concat_9834_comb[16] = p1_array_concat_9831_comb[16];
  assign p1_array_concat_9834_comb[17] = p1_array_concat_9831_comb[17];
  assign p1_array_concat_9834_comb[18] = p1_array_concat_9831_comb[18];
  assign p1_array_concat_9834_comb[19] = p1_array_concat_9831_comb[19];
  assign p1_array_concat_9834_comb[20] = p1_array_concat_9831_comb[20];
  assign p1_array_concat_9834_comb[21] = p1_array_concat_9831_comb[21];
  assign p1_array_concat_9834_comb[22] = p1_array_concat_9831_comb[22];
  assign p1_array_concat_9834_comb[23] = p1_array_concat_9831_comb[23];
  assign p1_array_concat_9834_comb[24] = p1_array_concat_9831_comb[24];
  assign p1_array_concat_9834_comb[25] = p1_array_concat_9831_comb[25];
  assign p1_array_concat_9834_comb[26] = p1_array_concat_9831_comb[26];
  assign p1_array_concat_9834_comb[27] = p1_array_concat_9831_comb[27];
  assign p1_array_concat_9834_comb[28] = p1_array_concat_9831_comb[28];
  assign p1_array_concat_9834_comb[29] = p1_array_concat_9831_comb[29];
  assign p1_array_concat_9834_comb[30] = p1_array_concat_9831_comb[30];
  assign p1_array_concat_9834_comb[31] = p1_array_concat_9831_comb[31];
  assign p1_array_concat_9834_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_9834_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_9834_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_9834_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_9834_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_9834_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_9834_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_9834_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[p1_idx_u8__5_squeezed_comb][0];
  assign p1_row5_comb[1] = p0_matrix[p1_idx_u8__5_squeezed_comb][1];
  assign p1_row5_comb[2] = p0_matrix[p1_idx_u8__5_squeezed_comb][2];
  assign p1_row5_comb[3] = p0_matrix[p1_idx_u8__5_squeezed_comb][3];
  assign p1_row5_comb[4] = p0_matrix[p1_idx_u8__5_squeezed_comb][4];
  assign p1_row5_comb[5] = p0_matrix[p1_idx_u8__5_squeezed_comb][5];
  assign p1_row5_comb[6] = p0_matrix[p1_idx_u8__5_squeezed_comb][6];
  assign p1_row5_comb[7] = p0_matrix[p1_idx_u8__5_squeezed_comb][7];
  assign p1_idx_u8__6_squeezed_comb = 3'h6;
  assign p1_idx_u8__13_comb = 8'h0d;
  assign p1_array_concat_9840_comb[0] = p1_array_concat_9834_comb[0];
  assign p1_array_concat_9840_comb[1] = p1_array_concat_9834_comb[1];
  assign p1_array_concat_9840_comb[2] = p1_array_concat_9834_comb[2];
  assign p1_array_concat_9840_comb[3] = p1_array_concat_9834_comb[3];
  assign p1_array_concat_9840_comb[4] = p1_array_concat_9834_comb[4];
  assign p1_array_concat_9840_comb[5] = p1_array_concat_9834_comb[5];
  assign p1_array_concat_9840_comb[6] = p1_array_concat_9834_comb[6];
  assign p1_array_concat_9840_comb[7] = p1_array_concat_9834_comb[7];
  assign p1_array_concat_9840_comb[8] = p1_array_concat_9834_comb[8];
  assign p1_array_concat_9840_comb[9] = p1_array_concat_9834_comb[9];
  assign p1_array_concat_9840_comb[10] = p1_array_concat_9834_comb[10];
  assign p1_array_concat_9840_comb[11] = p1_array_concat_9834_comb[11];
  assign p1_array_concat_9840_comb[12] = p1_array_concat_9834_comb[12];
  assign p1_array_concat_9840_comb[13] = p1_array_concat_9834_comb[13];
  assign p1_array_concat_9840_comb[14] = p1_array_concat_9834_comb[14];
  assign p1_array_concat_9840_comb[15] = p1_array_concat_9834_comb[15];
  assign p1_array_concat_9840_comb[16] = p1_array_concat_9834_comb[16];
  assign p1_array_concat_9840_comb[17] = p1_array_concat_9834_comb[17];
  assign p1_array_concat_9840_comb[18] = p1_array_concat_9834_comb[18];
  assign p1_array_concat_9840_comb[19] = p1_array_concat_9834_comb[19];
  assign p1_array_concat_9840_comb[20] = p1_array_concat_9834_comb[20];
  assign p1_array_concat_9840_comb[21] = p1_array_concat_9834_comb[21];
  assign p1_array_concat_9840_comb[22] = p1_array_concat_9834_comb[22];
  assign p1_array_concat_9840_comb[23] = p1_array_concat_9834_comb[23];
  assign p1_array_concat_9840_comb[24] = p1_array_concat_9834_comb[24];
  assign p1_array_concat_9840_comb[25] = p1_array_concat_9834_comb[25];
  assign p1_array_concat_9840_comb[26] = p1_array_concat_9834_comb[26];
  assign p1_array_concat_9840_comb[27] = p1_array_concat_9834_comb[27];
  assign p1_array_concat_9840_comb[28] = p1_array_concat_9834_comb[28];
  assign p1_array_concat_9840_comb[29] = p1_array_concat_9834_comb[29];
  assign p1_array_concat_9840_comb[30] = p1_array_concat_9834_comb[30];
  assign p1_array_concat_9840_comb[31] = p1_array_concat_9834_comb[31];
  assign p1_array_concat_9840_comb[32] = p1_array_concat_9834_comb[32];
  assign p1_array_concat_9840_comb[33] = p1_array_concat_9834_comb[33];
  assign p1_array_concat_9840_comb[34] = p1_array_concat_9834_comb[34];
  assign p1_array_concat_9840_comb[35] = p1_array_concat_9834_comb[35];
  assign p1_array_concat_9840_comb[36] = p1_array_concat_9834_comb[36];
  assign p1_array_concat_9840_comb[37] = p1_array_concat_9834_comb[37];
  assign p1_array_concat_9840_comb[38] = p1_array_concat_9834_comb[38];
  assign p1_array_concat_9840_comb[39] = p1_array_concat_9834_comb[39];
  assign p1_array_concat_9840_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_9840_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_9840_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_9840_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_9840_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_9840_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_9840_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_9840_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[p1_idx_u8__6_squeezed_comb][0];
  assign p1_row6_comb[1] = p0_matrix[p1_idx_u8__6_squeezed_comb][1];
  assign p1_row6_comb[2] = p0_matrix[p1_idx_u8__6_squeezed_comb][2];
  assign p1_row6_comb[3] = p0_matrix[p1_idx_u8__6_squeezed_comb][3];
  assign p1_row6_comb[4] = p0_matrix[p1_idx_u8__6_squeezed_comb][4];
  assign p1_row6_comb[5] = p0_matrix[p1_idx_u8__6_squeezed_comb][5];
  assign p1_row6_comb[6] = p0_matrix[p1_idx_u8__6_squeezed_comb][6];
  assign p1_row6_comb[7] = p0_matrix[p1_idx_u8__6_squeezed_comb][7];
  assign p1_idx_u8__7_squeezed_comb = 3'h7;
  assign p1_add_9843_comb = p0_start_pix[7:1] + 7'h07;
  assign p1_actual_index__13_comb = p0_start_pix + p1_idx_u8__13_comb;
  assign p1_array_concat_9847_comb[0] = p1_array_concat_9840_comb[0];
  assign p1_array_concat_9847_comb[1] = p1_array_concat_9840_comb[1];
  assign p1_array_concat_9847_comb[2] = p1_array_concat_9840_comb[2];
  assign p1_array_concat_9847_comb[3] = p1_array_concat_9840_comb[3];
  assign p1_array_concat_9847_comb[4] = p1_array_concat_9840_comb[4];
  assign p1_array_concat_9847_comb[5] = p1_array_concat_9840_comb[5];
  assign p1_array_concat_9847_comb[6] = p1_array_concat_9840_comb[6];
  assign p1_array_concat_9847_comb[7] = p1_array_concat_9840_comb[7];
  assign p1_array_concat_9847_comb[8] = p1_array_concat_9840_comb[8];
  assign p1_array_concat_9847_comb[9] = p1_array_concat_9840_comb[9];
  assign p1_array_concat_9847_comb[10] = p1_array_concat_9840_comb[10];
  assign p1_array_concat_9847_comb[11] = p1_array_concat_9840_comb[11];
  assign p1_array_concat_9847_comb[12] = p1_array_concat_9840_comb[12];
  assign p1_array_concat_9847_comb[13] = p1_array_concat_9840_comb[13];
  assign p1_array_concat_9847_comb[14] = p1_array_concat_9840_comb[14];
  assign p1_array_concat_9847_comb[15] = p1_array_concat_9840_comb[15];
  assign p1_array_concat_9847_comb[16] = p1_array_concat_9840_comb[16];
  assign p1_array_concat_9847_comb[17] = p1_array_concat_9840_comb[17];
  assign p1_array_concat_9847_comb[18] = p1_array_concat_9840_comb[18];
  assign p1_array_concat_9847_comb[19] = p1_array_concat_9840_comb[19];
  assign p1_array_concat_9847_comb[20] = p1_array_concat_9840_comb[20];
  assign p1_array_concat_9847_comb[21] = p1_array_concat_9840_comb[21];
  assign p1_array_concat_9847_comb[22] = p1_array_concat_9840_comb[22];
  assign p1_array_concat_9847_comb[23] = p1_array_concat_9840_comb[23];
  assign p1_array_concat_9847_comb[24] = p1_array_concat_9840_comb[24];
  assign p1_array_concat_9847_comb[25] = p1_array_concat_9840_comb[25];
  assign p1_array_concat_9847_comb[26] = p1_array_concat_9840_comb[26];
  assign p1_array_concat_9847_comb[27] = p1_array_concat_9840_comb[27];
  assign p1_array_concat_9847_comb[28] = p1_array_concat_9840_comb[28];
  assign p1_array_concat_9847_comb[29] = p1_array_concat_9840_comb[29];
  assign p1_array_concat_9847_comb[30] = p1_array_concat_9840_comb[30];
  assign p1_array_concat_9847_comb[31] = p1_array_concat_9840_comb[31];
  assign p1_array_concat_9847_comb[32] = p1_array_concat_9840_comb[32];
  assign p1_array_concat_9847_comb[33] = p1_array_concat_9840_comb[33];
  assign p1_array_concat_9847_comb[34] = p1_array_concat_9840_comb[34];
  assign p1_array_concat_9847_comb[35] = p1_array_concat_9840_comb[35];
  assign p1_array_concat_9847_comb[36] = p1_array_concat_9840_comb[36];
  assign p1_array_concat_9847_comb[37] = p1_array_concat_9840_comb[37];
  assign p1_array_concat_9847_comb[38] = p1_array_concat_9840_comb[38];
  assign p1_array_concat_9847_comb[39] = p1_array_concat_9840_comb[39];
  assign p1_array_concat_9847_comb[40] = p1_array_concat_9840_comb[40];
  assign p1_array_concat_9847_comb[41] = p1_array_concat_9840_comb[41];
  assign p1_array_concat_9847_comb[42] = p1_array_concat_9840_comb[42];
  assign p1_array_concat_9847_comb[43] = p1_array_concat_9840_comb[43];
  assign p1_array_concat_9847_comb[44] = p1_array_concat_9840_comb[44];
  assign p1_array_concat_9847_comb[45] = p1_array_concat_9840_comb[45];
  assign p1_array_concat_9847_comb[46] = p1_array_concat_9840_comb[46];
  assign p1_array_concat_9847_comb[47] = p1_array_concat_9840_comb[47];
  assign p1_array_concat_9847_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_9847_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_9847_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_9847_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_9847_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_9847_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_9847_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_9847_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[p1_idx_u8__7_squeezed_comb][0];
  assign p1_row7_comb[1] = p0_matrix[p1_idx_u8__7_squeezed_comb][1];
  assign p1_row7_comb[2] = p0_matrix[p1_idx_u8__7_squeezed_comb][2];
  assign p1_row7_comb[3] = p0_matrix[p1_idx_u8__7_squeezed_comb][3];
  assign p1_row7_comb[4] = p0_matrix[p1_idx_u8__7_squeezed_comb][4];
  assign p1_row7_comb[5] = p0_matrix[p1_idx_u8__7_squeezed_comb][5];
  assign p1_row7_comb[6] = p0_matrix[p1_idx_u8__7_squeezed_comb][6];
  assign p1_row7_comb[7] = p0_matrix[p1_idx_u8__7_squeezed_comb][7];
  assign p1_add_9852_comb = p0_start_pix[7:2] + 6'h03;
  assign p1_flat_comb[0] = p1_array_concat_9847_comb[0];
  assign p1_flat_comb[1] = p1_array_concat_9847_comb[1];
  assign p1_flat_comb[2] = p1_array_concat_9847_comb[2];
  assign p1_flat_comb[3] = p1_array_concat_9847_comb[3];
  assign p1_flat_comb[4] = p1_array_concat_9847_comb[4];
  assign p1_flat_comb[5] = p1_array_concat_9847_comb[5];
  assign p1_flat_comb[6] = p1_array_concat_9847_comb[6];
  assign p1_flat_comb[7] = p1_array_concat_9847_comb[7];
  assign p1_flat_comb[8] = p1_array_concat_9847_comb[8];
  assign p1_flat_comb[9] = p1_array_concat_9847_comb[9];
  assign p1_flat_comb[10] = p1_array_concat_9847_comb[10];
  assign p1_flat_comb[11] = p1_array_concat_9847_comb[11];
  assign p1_flat_comb[12] = p1_array_concat_9847_comb[12];
  assign p1_flat_comb[13] = p1_array_concat_9847_comb[13];
  assign p1_flat_comb[14] = p1_array_concat_9847_comb[14];
  assign p1_flat_comb[15] = p1_array_concat_9847_comb[15];
  assign p1_flat_comb[16] = p1_array_concat_9847_comb[16];
  assign p1_flat_comb[17] = p1_array_concat_9847_comb[17];
  assign p1_flat_comb[18] = p1_array_concat_9847_comb[18];
  assign p1_flat_comb[19] = p1_array_concat_9847_comb[19];
  assign p1_flat_comb[20] = p1_array_concat_9847_comb[20];
  assign p1_flat_comb[21] = p1_array_concat_9847_comb[21];
  assign p1_flat_comb[22] = p1_array_concat_9847_comb[22];
  assign p1_flat_comb[23] = p1_array_concat_9847_comb[23];
  assign p1_flat_comb[24] = p1_array_concat_9847_comb[24];
  assign p1_flat_comb[25] = p1_array_concat_9847_comb[25];
  assign p1_flat_comb[26] = p1_array_concat_9847_comb[26];
  assign p1_flat_comb[27] = p1_array_concat_9847_comb[27];
  assign p1_flat_comb[28] = p1_array_concat_9847_comb[28];
  assign p1_flat_comb[29] = p1_array_concat_9847_comb[29];
  assign p1_flat_comb[30] = p1_array_concat_9847_comb[30];
  assign p1_flat_comb[31] = p1_array_concat_9847_comb[31];
  assign p1_flat_comb[32] = p1_array_concat_9847_comb[32];
  assign p1_flat_comb[33] = p1_array_concat_9847_comb[33];
  assign p1_flat_comb[34] = p1_array_concat_9847_comb[34];
  assign p1_flat_comb[35] = p1_array_concat_9847_comb[35];
  assign p1_flat_comb[36] = p1_array_concat_9847_comb[36];
  assign p1_flat_comb[37] = p1_array_concat_9847_comb[37];
  assign p1_flat_comb[38] = p1_array_concat_9847_comb[38];
  assign p1_flat_comb[39] = p1_array_concat_9847_comb[39];
  assign p1_flat_comb[40] = p1_array_concat_9847_comb[40];
  assign p1_flat_comb[41] = p1_array_concat_9847_comb[41];
  assign p1_flat_comb[42] = p1_array_concat_9847_comb[42];
  assign p1_flat_comb[43] = p1_array_concat_9847_comb[43];
  assign p1_flat_comb[44] = p1_array_concat_9847_comb[44];
  assign p1_flat_comb[45] = p1_array_concat_9847_comb[45];
  assign p1_flat_comb[46] = p1_array_concat_9847_comb[46];
  assign p1_flat_comb[47] = p1_array_concat_9847_comb[47];
  assign p1_flat_comb[48] = p1_array_concat_9847_comb[48];
  assign p1_flat_comb[49] = p1_array_concat_9847_comb[49];
  assign p1_flat_comb[50] = p1_array_concat_9847_comb[50];
  assign p1_flat_comb[51] = p1_array_concat_9847_comb[51];
  assign p1_flat_comb[52] = p1_array_concat_9847_comb[52];
  assign p1_flat_comb[53] = p1_array_concat_9847_comb[53];
  assign p1_flat_comb[54] = p1_array_concat_9847_comb[54];
  assign p1_flat_comb[55] = p1_array_concat_9847_comb[55];
  assign p1_flat_comb[56] = p1_row7_comb[0];
  assign p1_flat_comb[57] = p1_row7_comb[1];
  assign p1_flat_comb[58] = p1_row7_comb[2];
  assign p1_flat_comb[59] = p1_row7_comb[3];
  assign p1_flat_comb[60] = p1_row7_comb[4];
  assign p1_flat_comb[61] = p1_row7_comb[5];
  assign p1_flat_comb[62] = p1_row7_comb[6];
  assign p1_flat_comb[63] = p1_row7_comb[7];
  assign p1_actual_index__14_comb = {p1_add_9843_comb, p0_start_pix[0]};
  assign p1_idx_u8__11_comb = 8'h0b;
  assign p1_actual_index__12_comb = {p1_add_9852_comb, p0_start_pix[1:0]};
  assign p1_actual_index__11_comb = p0_start_pix + p1_idx_u8__11_comb;
  assign p1_and_9871_comb = p1_flat_comb[p1_actual_index__14_comb > 8'h3f ? 6'h3f : p1_actual_index__14_comb[5:0]] & {8{~(p1_add_9843_comb[5] | p1_add_9843_comb[6])}};
  assign p1_idx_u8__1_comb = 8'h01;
  assign p1_idx_u8__3_comb = 8'h03;
  assign p1_idx_u8__5_comb = 8'h05;
  assign p1_idx_u8__7_comb = 8'h07;
  assign p1_idx_u8__9_comb = 8'h09;
  assign p1_add_9876_comb = p0_start_pix[7:1] + 7'h05;
  assign p1_and_9879_comb = p1_flat_comb[p1_actual_index__13_comb > 8'h3f ? 6'h3f : p1_actual_index__13_comb[5:0]] & {8{~(p1_actual_index__13_comb[6] | p1_actual_index__13_comb[7])}};
  assign p1_eq_9882_comb = p1_and_9871_comb == 8'h00;
  assign p1_and_9883_comb = p1_flat_comb[p1_actual_index__12_comb > 8'h3f ? 6'h3f : p1_actual_index__12_comb[5:0]] & {8{~(p1_add_9852_comb[4] | p1_add_9852_comb[5])}};
  assign p1_actual_index__1_comb = p0_start_pix + p1_idx_u8__1_comb;
  assign p1_add_9967_comb = p0_start_pix[7:1] + 7'h01;
  assign p1_actual_index__3_comb = p0_start_pix + p1_idx_u8__3_comb;
  assign p1_add_9949_comb = p0_start_pix[7:2] + 6'h01;
  assign p1_actual_index__5_comb = p0_start_pix + p1_idx_u8__5_comb;
  assign p1_add_9929_comb = p0_start_pix[7:1] + 7'h03;
  assign p1_actual_index__7_comb = p0_start_pix + p1_idx_u8__7_comb;
  assign p1_actual_index__9_comb = p0_start_pix + p1_idx_u8__9_comb;
  assign p1_idx_u8__15_comb = 8'h0f;
  assign p1_idx_u8__17_comb = 8'h11;
  assign p1_idx_u8__19_comb = 8'h13;
  assign p1_idx_u8__21_comb = 8'h15;
  assign p1_idx_u8__23_comb = 8'h17;
  assign p1_idx_u8__25_comb = 8'h19;
  assign p1_idx_u8__27_comb = 8'h1b;
  assign p1_idx_u8__29_comb = 8'h1d;
  assign p1_idx_u8__31_comb = 8'h1f;
  assign p1_idx_u8__33_comb = 8'h21;
  assign p1_idx_u8__35_comb = 8'h23;
  assign p1_idx_u8__37_comb = 8'h25;
  assign p1_idx_u8__39_comb = 8'h27;
  assign p1_idx_u8__41_comb = 8'h29;
  assign p1_idx_u8__43_comb = 8'h2b;
  assign p1_idx_u8__45_comb = 8'h2d;
  assign p1_idx_u8__47_comb = 8'h2f;
  assign p1_idx_u8__49_comb = 8'h31;
  assign p1_idx_u8__51_comb = 8'h33;
  assign p1_idx_u8__53_comb = 8'h35;
  assign p1_idx_u8__55_comb = 8'h37;
  assign p1_idx_u8__57_comb = 8'h39;
  assign p1_idx_u8__59_comb = 8'h3b;
  assign p1_idx_u8__61_comb = 8'h3d;
  assign p1_ne_9891_comb = p1_and_9879_comb != 8'h00;
  assign p1_idx_u8__1_squeezed_comb = 2'h1;
  assign p1_eq_9894_comb = p1_and_9883_comb == 8'h00;
  assign p1_add_9895_comb = p0_start_pix[7:3] + 5'h01;
  assign p1_actual_index__15_comb = p0_start_pix + p1_idx_u8__15_comb;
  assign p1_add_10070_comb = p0_start_pix[7:4] + 4'h1;
  assign p1_actual_index__17_comb = p0_start_pix + p1_idx_u8__17_comb;
  assign p1_add_10072_comb = p0_start_pix[7:1] + 7'h09;
  assign p1_actual_index__19_comb = p0_start_pix + p1_idx_u8__19_comb;
  assign p1_add_10074_comb = p0_start_pix[7:2] + 6'h05;
  assign p1_actual_index__21_comb = p0_start_pix + p1_idx_u8__21_comb;
  assign p1_add_10076_comb = p0_start_pix[7:1] + 7'h0b;
  assign p1_actual_index__23_comb = p0_start_pix + p1_idx_u8__23_comb;
  assign p1_add_10078_comb = p0_start_pix[7:3] + 5'h03;
  assign p1_actual_index__25_comb = p0_start_pix + p1_idx_u8__25_comb;
  assign p1_add_10080_comb = p0_start_pix[7:1] + 7'h0d;
  assign p1_actual_index__27_comb = p0_start_pix + p1_idx_u8__27_comb;
  assign p1_add_10082_comb = p0_start_pix[7:2] + 6'h07;
  assign p1_actual_index__29_comb = p0_start_pix + p1_idx_u8__29_comb;
  assign p1_add_10084_comb = p0_start_pix[7:1] + 7'h0f;
  assign p1_actual_index__31_comb = p0_start_pix + p1_idx_u8__31_comb;
  assign p1_add_10086_comb = p0_start_pix[7:5] + 3'h1;
  assign p1_actual_index__33_comb = p0_start_pix + p1_idx_u8__33_comb;
  assign p1_add_10088_comb = p0_start_pix[7:1] + 7'h11;
  assign p1_actual_index__35_comb = p0_start_pix + p1_idx_u8__35_comb;
  assign p1_add_10090_comb = p0_start_pix[7:2] + 6'h09;
  assign p1_actual_index__37_comb = p0_start_pix + p1_idx_u8__37_comb;
  assign p1_add_10092_comb = p0_start_pix[7:1] + 7'h13;
  assign p1_actual_index__39_comb = p0_start_pix + p1_idx_u8__39_comb;
  assign p1_add_10094_comb = p0_start_pix[7:3] + 5'h05;
  assign p1_actual_index__41_comb = p0_start_pix + p1_idx_u8__41_comb;
  assign p1_add_10096_comb = p0_start_pix[7:1] + 7'h15;
  assign p1_actual_index__43_comb = p0_start_pix + p1_idx_u8__43_comb;
  assign p1_add_10098_comb = p0_start_pix[7:2] + 6'h0b;
  assign p1_actual_index__45_comb = p0_start_pix + p1_idx_u8__45_comb;
  assign p1_add_10100_comb = p0_start_pix[7:1] + 7'h17;
  assign p1_actual_index__47_comb = p0_start_pix + p1_idx_u8__47_comb;
  assign p1_add_10102_comb = p0_start_pix[7:4] + 4'h3;
  assign p1_actual_index__49_comb = p0_start_pix + p1_idx_u8__49_comb;
  assign p1_add_10104_comb = p0_start_pix[7:1] + 7'h19;
  assign p1_actual_index__51_comb = p0_start_pix + p1_idx_u8__51_comb;
  assign p1_add_10106_comb = p0_start_pix[7:2] + 6'h0d;
  assign p1_actual_index__53_comb = p0_start_pix + p1_idx_u8__53_comb;
  assign p1_add_10108_comb = p0_start_pix[7:1] + 7'h1b;
  assign p1_actual_index__55_comb = p0_start_pix + p1_idx_u8__55_comb;
  assign p1_add_10110_comb = p0_start_pix[7:3] + 5'h07;
  assign p1_actual_index__57_comb = p0_start_pix + p1_idx_u8__57_comb;
  assign p1_add_10112_comb = p0_start_pix[7:1] + 7'h1d;
  assign p1_actual_index__59_comb = p0_start_pix + p1_idx_u8__59_comb;
  assign p1_add_10114_comb = p0_start_pix[7:2] + 6'h0f;
  assign p1_actual_index__61_comb = p0_start_pix + p1_idx_u8__61_comb;
  assign p1_add_10116_comb = p0_start_pix[7:1] + 7'h1f;
  assign p1_actual_index__10_comb = {p1_add_9876_comb, p0_start_pix[0]};
  assign p1_actual_index__2_comb = {p1_add_9967_comb, p0_start_pix[0]};
  assign p1_actual_index__4_comb = {p1_add_9949_comb, p0_start_pix[1:0]};
  assign p1_actual_index__6_comb = {p1_add_9929_comb, p0_start_pix[0]};
  assign p1_and_9911_comb = p1_flat_comb[p1_actual_index__11_comb > 8'h3f ? 6'h3f : p1_actual_index__11_comb[5:0]] & {8{~(p1_actual_index__11_comb[6] | p1_actual_index__11_comb[7])}};
  assign p1_actual_index__8_comb = {p1_add_9895_comb, p0_start_pix[2:0]};
  assign p1_actual_index__16_comb = {p1_add_10070_comb, p0_start_pix[3:0]};
  assign p1_actual_index__18_comb = {p1_add_10072_comb, p0_start_pix[0]};
  assign p1_actual_index__20_comb = {p1_add_10074_comb, p0_start_pix[1:0]};
  assign p1_actual_index__22_comb = {p1_add_10076_comb, p0_start_pix[0]};
  assign p1_actual_index__24_comb = {p1_add_10078_comb, p0_start_pix[2:0]};
  assign p1_actual_index__26_comb = {p1_add_10080_comb, p0_start_pix[0]};
  assign p1_actual_index__28_comb = {p1_add_10082_comb, p0_start_pix[1:0]};
  assign p1_actual_index__30_comb = {p1_add_10084_comb, p0_start_pix[0]};
  assign p1_actual_index__32_comb = {p1_add_10086_comb, p0_start_pix[4:0]};
  assign p1_actual_index__34_comb = {p1_add_10088_comb, p0_start_pix[0]};
  assign p1_actual_index__36_comb = {p1_add_10090_comb, p0_start_pix[1:0]};
  assign p1_actual_index__38_comb = {p1_add_10092_comb, p0_start_pix[0]};
  assign p1_actual_index__40_comb = {p1_add_10094_comb, p0_start_pix[2:0]};
  assign p1_actual_index__42_comb = {p1_add_10096_comb, p0_start_pix[0]};
  assign p1_actual_index__44_comb = {p1_add_10098_comb, p0_start_pix[1:0]};
  assign p1_actual_index__46_comb = {p1_add_10100_comb, p0_start_pix[0]};
  assign p1_actual_index__48_comb = {p1_add_10102_comb, p0_start_pix[3:0]};
  assign p1_actual_index__50_comb = {p1_add_10104_comb, p0_start_pix[0]};
  assign p1_actual_index__52_comb = {p1_add_10106_comb, p0_start_pix[1:0]};
  assign p1_actual_index__54_comb = {p1_add_10108_comb, p0_start_pix[0]};
  assign p1_actual_index__56_comb = {p1_add_10110_comb, p0_start_pix[2:0]};
  assign p1_actual_index__58_comb = {p1_add_10112_comb, p0_start_pix[0]};
  assign p1_actual_index__60_comb = {p1_add_10114_comb, p0_start_pix[1:0]};
  assign p1_actual_index__62_comb = {p1_add_10116_comb, p0_start_pix[0]};
  assign p1_and_9921_comb = p1_flat_comb[p1_actual_index__10_comb > 8'h3f ? 6'h3f : p1_actual_index__10_comb[5:0]] & {8{~(p1_add_9876_comb[5] | p1_add_9876_comb[6])}};
  assign p1_ne_9923_comb = p1_and_9911_comb != 8'h00;
  assign p1_and_10011_comb = p1_flat_comb[p0_start_pix > 8'h3f ? 6'h3f : p0_start_pix[5:0]] & {8{~(p0_start_pix[6] | p0_start_pix[7])}};
  assign p1_and_10013_comb = p1_flat_comb[p1_actual_index__1_comb > 8'h3f ? 6'h3f : p1_actual_index__1_comb[5:0]] & {8{~(p1_actual_index__1_comb[6] | p1_actual_index__1_comb[7])}};
  assign p1_and_10008_comb = p1_flat_comb[p1_actual_index__2_comb > 8'h3f ? 6'h3f : p1_actual_index__2_comb[5:0]] & {8{~(p1_add_9967_comb[5] | p1_add_9967_comb[6])}};
  assign p1_and_10001_comb = p1_flat_comb[p1_actual_index__3_comb > 8'h3f ? 6'h3f : p1_actual_index__3_comb[5:0]] & {8{~(p1_actual_index__3_comb[6] | p1_actual_index__3_comb[7])}};
  assign p1_and_9994_comb = p1_flat_comb[p1_actual_index__4_comb > 8'h3f ? 6'h3f : p1_actual_index__4_comb[5:0]] & {8{~(p1_add_9949_comb[4] | p1_add_9949_comb[5])}};
  assign p1_and_9983_comb = p1_flat_comb[p1_actual_index__5_comb > 8'h3f ? 6'h3f : p1_actual_index__5_comb[5:0]] & {8{~(p1_actual_index__5_comb[6] | p1_actual_index__5_comb[7])}};
  assign p1_and_9974_comb = p1_flat_comb[p1_actual_index__6_comb > 8'h3f ? 6'h3f : p1_actual_index__6_comb[5:0]] & {8{~(p1_add_9929_comb[5] | p1_add_9929_comb[6])}};
  assign p1_and_9964_comb = p1_flat_comb[p1_actual_index__7_comb > 8'h3f ? 6'h3f : p1_actual_index__7_comb[5:0]] & {8{~(p1_actual_index__7_comb[6] | p1_actual_index__7_comb[7])}};
  assign p1_and_9932_comb = p1_flat_comb[p1_actual_index__9_comb > 8'h3f ? 6'h3f : p1_actual_index__9_comb[5:0]] & {8{~(p1_actual_index__9_comb[6] | p1_actual_index__9_comb[7])}};
  assign p1_ne_9934_comb = p1_and_9921_comb != 8'h00;
  assign p1_sel_9935_comb = p1_ne_9923_comb ? 3'h3 : {1'h1, (p1_ne_9891_comb ? p1_idx_u8__1_squeezed_comb : {1'h1, p1_eq_9882_comb}) & {2{p1_eq_9894_comb}}};
  assign p1_ne_10016_comb = p1_and_10011_comb != 8'h00;
  assign p1_ne_10017_comb = p1_and_10013_comb != 8'h00;
  assign p1_ne_10015_comb = p1_and_10008_comb != 8'h00;
  assign p1_ne_10010_comb = p1_and_10001_comb != 8'h00;
  assign p1_ne_10003_comb = p1_and_9994_comb != 8'h00;
  assign p1_ne_9996_comb = p1_and_9983_comb != 8'h00;
  assign p1_ne_9985_comb = p1_and_9974_comb != 8'h00;
  assign p1_ne_9976_comb = p1_and_9964_comb != 8'h00;
  assign p1_and_9937_comb = p1_flat_comb[p1_actual_index__8_comb > 8'h3f ? 6'h3f : p1_actual_index__8_comb[5:0]] & {8{~(p1_add_9895_comb[3] | p1_add_9895_comb[4])}};
  assign p1_ne_9944_comb = p1_and_9932_comb != 8'h00;
  assign p1_not_10018_comb = ~p1_ne_10016_comb;
  assign p1_eq_9947_comb = p1_and_9937_comb == 8'h00;
  assign p1_sel_9956_comb = p1_ne_9944_comb ? 3'h1 : (p1_ne_9934_comb ? 3'h2 : p1_sel_9935_comb);
  assign p1_and_10538_comb = p1_not_10018_comb & ~p1_ne_10017_comb & ~p1_ne_10015_comb & ~p1_ne_10010_comb & ~p1_ne_10003_comb & ~p1_ne_9996_comb & ~p1_ne_9985_comb & ~p1_ne_9976_comb & p1_eq_9947_comb & ~p1_ne_9944_comb & ~p1_ne_9934_comb & ~p1_ne_9923_comb & p1_eq_9894_comb & ~p1_ne_9891_comb & p1_eq_9882_comb & (p1_flat_comb[p1_actual_index__15_comb > 8'h3f ? 6'h3f : p1_actual_index__15_comb[5:0]] & {8{~(p1_actual_index__15_comb[6] | p1_actual_index__15_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__16_comb > 8'h3f ? 6'h3f : p1_actual_index__16_comb[5:0]] & {8{~(p1_add_10070_comb[2] | p1_add_10070_comb[3])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__17_comb > 8'h3f ? 6'h3f : p1_actual_index__17_comb[5:0]] & {8{~(p1_actual_index__17_comb[6] | p1_actual_index__17_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__18_comb > 8'h3f ? 6'h3f : p1_actual_index__18_comb[5:0]] & {8{~(p1_add_10072_comb[5] | p1_add_10072_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__19_comb > 8'h3f ? 6'h3f : p1_actual_index__19_comb[5:0]] & {8{~(p1_actual_index__19_comb[6] | p1_actual_index__19_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__20_comb > 8'h3f ? 6'h3f : p1_actual_index__20_comb[5:0]] & {8{~(p1_add_10074_comb[4] | p1_add_10074_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__21_comb > 8'h3f ? 6'h3f : p1_actual_index__21_comb[5:0]] & {8{~(p1_actual_index__21_comb[6] | p1_actual_index__21_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__22_comb > 8'h3f ? 6'h3f : p1_actual_index__22_comb[5:0]] & {8{~(p1_add_10076_comb[5] | p1_add_10076_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__23_comb > 8'h3f ? 6'h3f : p1_actual_index__23_comb[5:0]] & {8{~(p1_actual_index__23_comb[6] | p1_actual_index__23_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__24_comb > 8'h3f ? 6'h3f : p1_actual_index__24_comb[5:0]] & {8{~(p1_add_10078_comb[3] | p1_add_10078_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__25_comb > 8'h3f ? 6'h3f : p1_actual_index__25_comb[5:0]] & {8{~(p1_actual_index__25_comb[6] | p1_actual_index__25_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__26_comb > 8'h3f ? 6'h3f : p1_actual_index__26_comb[5:0]] & {8{~(p1_add_10080_comb[5] | p1_add_10080_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__27_comb > 8'h3f ? 6'h3f : p1_actual_index__27_comb[5:0]] & {8{~(p1_actual_index__27_comb[6] | p1_actual_index__27_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__28_comb > 8'h3f ? 6'h3f : p1_actual_index__28_comb[5:0]] & {8{~(p1_add_10082_comb[4] | p1_add_10082_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__29_comb > 8'h3f ? 6'h3f : p1_actual_index__29_comb[5:0]] & {8{~(p1_actual_index__29_comb[6] | p1_actual_index__29_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__30_comb > 8'h3f ? 6'h3f : p1_actual_index__30_comb[5:0]] & {8{~(p1_add_10084_comb[5] | p1_add_10084_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__31_comb > 8'h3f ? 6'h3f : p1_actual_index__31_comb[5:0]] & {8{~(p1_actual_index__31_comb[6] | p1_actual_index__31_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__32_comb > 8'h3f ? 6'h3f : p1_actual_index__32_comb[5:0]] & {8{~(p1_add_10086_comb[1] | p1_add_10086_comb[2])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__33_comb > 8'h3f ? 6'h3f : p1_actual_index__33_comb[5:0]] & {8{~(p1_actual_index__33_comb[6] | p1_actual_index__33_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__34_comb > 8'h3f ? 6'h3f : p1_actual_index__34_comb[5:0]] & {8{~(p1_add_10088_comb[5] | p1_add_10088_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__35_comb > 8'h3f ? 6'h3f : p1_actual_index__35_comb[5:0]] & {8{~(p1_actual_index__35_comb[6] | p1_actual_index__35_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__36_comb > 8'h3f ? 6'h3f : p1_actual_index__36_comb[5:0]] & {8{~(p1_add_10090_comb[4] | p1_add_10090_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__37_comb > 8'h3f ? 6'h3f : p1_actual_index__37_comb[5:0]] & {8{~(p1_actual_index__37_comb[6] | p1_actual_index__37_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__38_comb > 8'h3f ? 6'h3f : p1_actual_index__38_comb[5:0]] & {8{~(p1_add_10092_comb[5] | p1_add_10092_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__39_comb > 8'h3f ? 6'h3f : p1_actual_index__39_comb[5:0]] & {8{~(p1_actual_index__39_comb[6] | p1_actual_index__39_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__40_comb > 8'h3f ? 6'h3f : p1_actual_index__40_comb[5:0]] & {8{~(p1_add_10094_comb[3] | p1_add_10094_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__41_comb > 8'h3f ? 6'h3f : p1_actual_index__41_comb[5:0]] & {8{~(p1_actual_index__41_comb[6] | p1_actual_index__41_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__42_comb > 8'h3f ? 6'h3f : p1_actual_index__42_comb[5:0]] & {8{~(p1_add_10096_comb[5] | p1_add_10096_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__43_comb > 8'h3f ? 6'h3f : p1_actual_index__43_comb[5:0]] & {8{~(p1_actual_index__43_comb[6] | p1_actual_index__43_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__44_comb > 8'h3f ? 6'h3f : p1_actual_index__44_comb[5:0]] & {8{~(p1_add_10098_comb[4] | p1_add_10098_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__45_comb > 8'h3f ? 6'h3f : p1_actual_index__45_comb[5:0]] & {8{~(p1_actual_index__45_comb[6] | p1_actual_index__45_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__46_comb > 8'h3f ? 6'h3f : p1_actual_index__46_comb[5:0]] & {8{~(p1_add_10100_comb[5] | p1_add_10100_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__47_comb > 8'h3f ? 6'h3f : p1_actual_index__47_comb[5:0]] & {8{~(p1_actual_index__47_comb[6] | p1_actual_index__47_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__48_comb > 8'h3f ? 6'h3f : p1_actual_index__48_comb[5:0]] & {8{~(p1_add_10102_comb[2] | p1_add_10102_comb[3])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__49_comb > 8'h3f ? 6'h3f : p1_actual_index__49_comb[5:0]] & {8{~(p1_actual_index__49_comb[6] | p1_actual_index__49_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__50_comb > 8'h3f ? 6'h3f : p1_actual_index__50_comb[5:0]] & {8{~(p1_add_10104_comb[5] | p1_add_10104_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__51_comb > 8'h3f ? 6'h3f : p1_actual_index__51_comb[5:0]] & {8{~(p1_actual_index__51_comb[6] | p1_actual_index__51_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__52_comb > 8'h3f ? 6'h3f : p1_actual_index__52_comb[5:0]] & {8{~(p1_add_10106_comb[4] | p1_add_10106_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__53_comb > 8'h3f ? 6'h3f : p1_actual_index__53_comb[5:0]] & {8{~(p1_actual_index__53_comb[6] | p1_actual_index__53_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__54_comb > 8'h3f ? 6'h3f : p1_actual_index__54_comb[5:0]] & {8{~(p1_add_10108_comb[5] | p1_add_10108_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__55_comb > 8'h3f ? 6'h3f : p1_actual_index__55_comb[5:0]] & {8{~(p1_actual_index__55_comb[6] | p1_actual_index__55_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__56_comb > 8'h3f ? 6'h3f : p1_actual_index__56_comb[5:0]] & {8{~(p1_add_10110_comb[3] | p1_add_10110_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__57_comb > 8'h3f ? 6'h3f : p1_actual_index__57_comb[5:0]] & {8{~(p1_actual_index__57_comb[6] | p1_actual_index__57_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__58_comb > 8'h3f ? 6'h3f : p1_actual_index__58_comb[5:0]] & {8{~(p1_add_10112_comb[5] | p1_add_10112_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__59_comb > 8'h3f ? 6'h3f : p1_actual_index__59_comb[5:0]] & {8{~(p1_actual_index__59_comb[6] | p1_actual_index__59_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__60_comb > 8'h3f ? 6'h3f : p1_actual_index__60_comb[5:0]] & {8{~(p1_add_10114_comb[4] | p1_add_10114_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__61_comb > 8'h3f ? 6'h3f : p1_actual_index__61_comb[5:0]] & {8{~(p1_actual_index__61_comb[6] | p1_actual_index__61_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__62_comb > 8'h3f ? 6'h3f : p1_actual_index__62_comb[5:0]] & {8{~(p1_add_10116_comb[5] | p1_add_10116_comb[6])}}) == 8'h00;
  assign p1_value_comb = p0_matrix[3'h0][3'h0];

  // Registers for pipe stage 1:
  reg p1_is_luminance;
  reg [7:0] p1_and_9871;
  reg [7:0] p1_and_9879;
  reg [7:0] p1_and_9883;
  reg [7:0] p1_and_9911;
  reg [7:0] p1_and_9921;
  reg [7:0] p1_and_9932;
  reg [7:0] p1_and_9937;
  reg p1_eq_9947;
  reg [2:0] p1_sel_9956;
  reg [7:0] p1_and_9964;
  reg [7:0] p1_and_9974;
  reg p1_ne_9976;
  reg [7:0] p1_and_9983;
  reg p1_ne_9985;
  reg [7:0] p1_and_9994;
  reg p1_ne_9996;
  reg [7:0] p1_and_10001;
  reg p1_ne_10003;
  reg [7:0] p1_and_10008;
  reg p1_ne_10010;
  reg [7:0] p1_and_10011;
  reg [7:0] p1_and_10013;
  reg p1_ne_10015;
  reg p1_ne_10016;
  reg p1_ne_10017;
  reg p1_not_10018;
  reg p1_and_10538;
  reg [7:0] p1_value;
  always @ (posedge clk) begin
    p1_is_luminance <= p0_is_luminance;
    p1_and_9871 <= p1_and_9871_comb;
    p1_and_9879 <= p1_and_9879_comb;
    p1_and_9883 <= p1_and_9883_comb;
    p1_and_9911 <= p1_and_9911_comb;
    p1_and_9921 <= p1_and_9921_comb;
    p1_and_9932 <= p1_and_9932_comb;
    p1_and_9937 <= p1_and_9937_comb;
    p1_eq_9947 <= p1_eq_9947_comb;
    p1_sel_9956 <= p1_sel_9956_comb;
    p1_and_9964 <= p1_and_9964_comb;
    p1_and_9974 <= p1_and_9974_comb;
    p1_ne_9976 <= p1_ne_9976_comb;
    p1_and_9983 <= p1_and_9983_comb;
    p1_ne_9985 <= p1_ne_9985_comb;
    p1_and_9994 <= p1_and_9994_comb;
    p1_ne_9996 <= p1_ne_9996_comb;
    p1_and_10001 <= p1_and_10001_comb;
    p1_ne_10003 <= p1_ne_10003_comb;
    p1_and_10008 <= p1_and_10008_comb;
    p1_ne_10010 <= p1_ne_10010_comb;
    p1_and_10011 <= p1_and_10011_comb;
    p1_and_10013 <= p1_and_10013_comb;
    p1_ne_10015 <= p1_ne_10015_comb;
    p1_ne_10016 <= p1_ne_10016_comb;
    p1_ne_10017 <= p1_ne_10017_comb;
    p1_not_10018 <= p1_not_10018_comb;
    p1_and_10538 <= p1_and_10538_comb;
    p1_value <= p1_value_comb;
  end

  // ===== Pipe stage 2:
  wire [3:0] p2_sel_10609_comb;
  wire [3:0] p2_sel_10613_comb;
  wire [3:0] p2_sel_10617_comb;
  wire [3:0] p2_run_comb;
  wire [7:0] p2_value__1_comb;
  wire [1:0] p2_idx_u8__1_squeezed__1_comb;
  wire [1:0] p2_idx_u8__2_squeezed_comb;
  wire p2_eq_10653_comb;
  wire [1:0] p2_idx_u8__3_squeezed_comb;
  wire p2_eq_10647_comb;
  wire [7:0] p2_flipped__1_comb;
  wire [7:0] p2_code_list__1_comb;
  wire [2:0] p2_idx_u8__4_squeezed__1_comb;
  wire [3:0] p2_add_10649_comb;
  wire p2_or_reduce_10638_comb;
  wire [2:0] p2_sel_10639_comb;
  wire p2_or_reduce_10641_comb;
  wire p2_or_reduce_10642_comb;
  wire p2_bit_slice_10646_comb;
  wire p2_not_10650_comb;
  wire [3:0] p2_run_u8__1_comb;
  wire p2_or_10654_comb;
  wire [7:0] p2_sel_10664_comb;
  wire [3:0] p2_sel_10665_comb;
  assign p2_sel_10609_comb = p1_ne_9996 ? 4'h5 : (p1_ne_9985 ? 4'h6 : (p1_ne_9976 ? 4'h7 : {1'h1, p1_sel_9956 & {3{p1_eq_9947}}}));
  assign p2_sel_10613_comb = p1_ne_10010 ? 4'h3 : (p1_ne_10003 ? 4'h4 : p2_sel_10609_comb);
  assign p2_sel_10617_comb = p1_ne_10017 ? 4'h1 : (p1_ne_10015 ? 4'h2 : p2_sel_10613_comb);
  assign p2_run_comb = p2_sel_10617_comb & {4{p1_not_10018}};
  assign p2_value__1_comb = p2_run_comb == 4'h0 ? p1_and_10011 : (p2_run_comb == 4'h1 ? p1_and_10013 : (p2_run_comb == 4'h2 ? p1_and_10008 : (p2_run_comb == 4'h3 ? p1_and_10001 : (p2_run_comb == 4'h4 ? p1_and_9994 : (p2_run_comb == 4'h5 ? p1_and_9983 : (p2_run_comb == 4'h6 ? p1_and_9974 : (p2_run_comb == 4'h7 ? p1_and_9964 : (p2_run_comb == 4'h8 ? p1_and_9937 : (p2_run_comb == 4'h9 ? p1_and_9932 : (p2_run_comb == 4'ha ? p1_and_9921 : (p2_run_comb == 4'hb ? p1_and_9911 : (p2_run_comb == 4'hc ? p1_and_9883 : (p2_run_comb == 4'hd ? p1_and_9879 : (p2_run_comb == 4'he ? p1_and_9871 : 8'h00))))))))))))));
  assign p2_idx_u8__1_squeezed__1_comb = 2'h1;
  assign p2_idx_u8__2_squeezed_comb = 2'h2;
  assign p2_eq_10653_comb = p2_run_comb == 4'hf;
  assign p2_idx_u8__3_squeezed_comb = 2'h3;
  assign p2_eq_10647_comb = p2_value__1_comb == 8'h00;
  assign p2_flipped__1_comb = 8'hff;
  assign p2_code_list__1_comb = p2_eq_10647_comb ? p2_flipped__1_comb : p2_value__1_comb;
  assign p2_idx_u8__4_squeezed__1_comb = 3'h4;
  assign p2_add_10649_comb = p2_sel_10613_comb + 4'h7;
  assign p2_or_reduce_10638_comb = |p2_value__1_comb[7:4];
  assign p2_sel_10639_comb = |p2_value__1_comb[7:3] ? p2_idx_u8__4_squeezed__1_comb : {1'h0, |p2_value__1_comb[7:2] ? p2_idx_u8__3_squeezed_comb : (|p2_value__1_comb[7:1] ? p2_idx_u8__2_squeezed_comb : p2_idx_u8__1_squeezed__1_comb)};
  assign p2_or_reduce_10641_comb = |p2_value__1_comb[7:5];
  assign p2_or_reduce_10642_comb = |p2_value__1_comb[7:6];
  assign p2_bit_slice_10646_comb = p2_value__1_comb[7];
  assign p2_not_10650_comb = ~p2_eq_10647_comb;
  assign p2_run_u8__1_comb = p2_run_comb < 4'ha ? p2_run_comb : p2_add_10649_comb;
  assign p2_or_10654_comb = p1_and_10538 | p2_eq_10653_comb;
  assign p2_sel_10664_comb = p1_and_10538 ? p1_value : p2_code_list__1_comb & {8{~p2_eq_10653_comb}};
  assign p2_sel_10665_comb = p1_and_10538 ? 4'hf : p2_sel_10617_comb & {4{~(p2_eq_10653_comb | p1_ne_10016)}};

  // Registers for pipe stage 2:
  reg p2_is_luminance;
  reg p2_or_reduce_10638;
  reg [2:0] p2_sel_10639;
  reg p2_or_reduce_10641;
  reg p2_or_reduce_10642;
  reg p2_bit_slice_10646;
  reg p2_not_10650;
  reg [3:0] p2_run_u8__1;
  reg p2_or_10654;
  reg [7:0] p2_sel_10664;
  reg [3:0] p2_sel_10665;
  always @ (posedge clk) begin
    p2_is_luminance <= p1_is_luminance;
    p2_or_reduce_10638 <= p2_or_reduce_10638_comb;
    p2_sel_10639 <= p2_sel_10639_comb;
    p2_or_reduce_10641 <= p2_or_reduce_10641_comb;
    p2_or_reduce_10642 <= p2_or_reduce_10642_comb;
    p2_bit_slice_10646 <= p2_bit_slice_10646_comb;
    p2_not_10650 <= p2_not_10650_comb;
    p2_run_u8__1 <= p2_run_u8__1_comb;
    p2_or_10654 <= p2_or_10654_comb;
    p2_sel_10664 <= p2_sel_10664_comb;
    p2_sel_10665 <= p2_sel_10665_comb;
  end

  // ===== Pipe stage 3:
  wire [2:0] p3_idx_u8__5_squeezed__1_comb;
  wire [2:0] p3_idx_u8__6_squeezed__1_comb;
  wire [2:0] p3_idx_u8__7_squeezed__1_comb;
  wire [3:0] p3_idx_u8__8_squeezed_comb;
  wire [7:0] p3_concat_10700_comb;
  wire [7:0] p3_size__1_comb;
  wire [7:0] p3_idx_u8__48_comb;
  wire [7:0] p3_run_size_str_u8__1_comb;
  wire [7:0] p3_idx_u8__8_comb;
  wire [7:0] p3_idx_u8__56_comb;
  wire [7:0] p3_idx_u8__54_comb;
  wire [7:0] p3_idx_u8__6_comb;
  wire [7:0] p3_idx_u8__52_comb;
  wire [7:0] p3_idx_u8__4_comb;
  wire [7:0] p3_idx_u8__50_comb;
  wire [7:0] p3_idx_u8__2_comb;
  wire p3_eq_10734_comb;
  wire p3_eq_10735_comb;
  wire p3_eq_10736_comb;
  wire p3_eq_10737_comb;
  wire p3_eq_10738_comb;
  wire p3_eq_10739_comb;
  wire p3_eq_10740_comb;
  wire p3_eq_10741_comb;
  wire p3_eq_10742_comb;
  wire p3_eq_10743_comb;
  wire p3_eq_10744_comb;
  wire p3_eq_10745_comb;
  wire p3_eq_10746_comb;
  wire p3_eq_10747_comb;
  wire p3_eq_10748_comb;
  wire p3_eq_10749_comb;
  wire p3_eq_10750_comb;
  wire p3_eq_10751_comb;
  wire p3_eq_10752_comb;
  wire p3_eq_10753_comb;
  wire p3_eq_10754_comb;
  wire p3_eq_10755_comb;
  wire p3_eq_10756_comb;
  wire p3_eq_10757_comb;
  wire p3_eq_10758_comb;
  wire p3_eq_10759_comb;
  wire p3_eq_10760_comb;
  wire p3_eq_10761_comb;
  wire p3_or_10762_comb;
  wire [2:0] p3_concat_10767_comb;
  wire [1:0] p3_idx_u8__1_squeezed__2_comb;
  wire [1:0] p3_idx_u8__3_squeezed__1_comb;
  wire [8:0] p3_concat_10776_comb;
  wire [2:0] p3_idx_u8__6_squeezed__2_comb;
  wire [2:0] p3_idx_u8__4_squeezed__2_comb;
  wire [2:0] p3_idx_u8__5_squeezed__2_comb;
  wire [2:0] p3_idx_u8__6_squeezed__3_comb;
  wire [2:0] p3_idx_u8__7_squeezed__2_comb;
  wire [1:0] p3_one_hot_sel_10859_comb;
  wire [27:0] p3_concat_10788_comb;
  wire [4:0] p3_huffman_length_squeezed_comb;
  wire [4:0] p3_idx_u8__2_squeezed__1_comb;
  wire [15:0] p3_huffman_code_full_comb;
  wire [28:0] p3_one_hot_10842_comb;
  wire [9:0] p3_one_hot_10848_comb;
  wire [3:0] p3_one_hot_10854_comb;
  wire [35:0] p3_tuple_10838_comb;
  assign p3_idx_u8__5_squeezed__1_comb = 3'h5;
  assign p3_idx_u8__6_squeezed__1_comb = 3'h6;
  assign p3_idx_u8__7_squeezed__1_comb = 3'h7;
  assign p3_idx_u8__8_squeezed_comb = 4'h8;
  assign p3_concat_10700_comb = {4'h0, p2_bit_slice_10646 ? p3_idx_u8__8_squeezed_comb : {1'h0, p2_or_reduce_10642 ? p3_idx_u8__7_squeezed__1_comb : (p2_or_reduce_10641 ? p3_idx_u8__6_squeezed__1_comb : (p2_or_reduce_10638 ? p3_idx_u8__5_squeezed__1_comb : p2_sel_10639))}};
  assign p3_size__1_comb = p3_concat_10700_comb & {8{p2_not_10650}};
  assign p3_idx_u8__48_comb = 8'h30;
  assign p3_run_size_str_u8__1_comb = {p2_run_u8__1, 4'h0} | p3_size__1_comb | p3_idx_u8__48_comb;
  assign p3_idx_u8__8_comb = 8'h37;
  assign p3_idx_u8__56_comb = 8'h38;
  assign p3_idx_u8__54_comb = 8'h36;
  assign p3_idx_u8__6_comb = 8'h35;
  assign p3_idx_u8__52_comb = 8'h34;
  assign p3_idx_u8__4_comb = 8'h33;
  assign p3_idx_u8__50_comb = 8'h32;
  assign p3_idx_u8__2_comb = 8'h31;
  assign p3_eq_10734_comb = p3_run_size_str_u8__1_comb == 8'h72;
  assign p3_eq_10735_comb = p3_run_size_str_u8__1_comb == 8'hf0;
  assign p3_eq_10736_comb = p3_run_size_str_u8__1_comb == 8'hb7;
  assign p3_eq_10737_comb = p3_run_size_str_u8__1_comb == 8'h77;
  assign p3_eq_10738_comb = p3_run_size_str_u8__1_comb == p3_idx_u8__8_comb;
  assign p3_eq_10739_comb = p3_run_size_str_u8__1_comb == 8'hf6;
  assign p3_eq_10740_comb = p3_run_size_str_u8__1_comb == 8'hb6;
  assign p3_eq_10741_comb = p3_run_size_str_u8__1_comb == 8'h76;
  assign p3_eq_10742_comb = p3_run_size_str_u8__1_comb == 8'hf5;
  assign p3_eq_10743_comb = p3_run_size_str_u8__1_comb == 8'hf4;
  assign p3_eq_10744_comb = p3_run_size_str_u8__1_comb == 8'hf3;
  assign p3_eq_10745_comb = p3_run_size_str_u8__1_comb == 8'hf2;
  assign p3_eq_10746_comb = p3_run_size_str_u8__1_comb == 8'hb5;
  assign p3_eq_10747_comb = p3_run_size_str_u8__1_comb == 8'h75;
  assign p3_eq_10748_comb = p3_run_size_str_u8__1_comb == p3_idx_u8__56_comb;
  assign p3_eq_10749_comb = p3_run_size_str_u8__1_comb == 8'h74;
  assign p3_eq_10750_comb = p3_run_size_str_u8__1_comb == p3_idx_u8__54_comb;
  assign p3_eq_10751_comb = p3_run_size_str_u8__1_comb == 8'hb3;
  assign p3_eq_10752_comb = p3_run_size_str_u8__1_comb == p3_idx_u8__6_comb;
  assign p3_eq_10753_comb = p3_run_size_str_u8__1_comb == 8'h73;
  assign p3_eq_10754_comb = p3_run_size_str_u8__1_comb == 8'hb2;
  assign p3_eq_10755_comb = p3_run_size_str_u8__1_comb == p3_idx_u8__52_comb;
  assign p3_eq_10756_comb = p3_run_size_str_u8__1_comb == 8'hf1;
  assign p3_eq_10757_comb = p3_run_size_str_u8__1_comb == p3_idx_u8__4_comb;
  assign p3_eq_10758_comb = p3_run_size_str_u8__1_comb == 8'hb1;
  assign p3_eq_10759_comb = p3_run_size_str_u8__1_comb == p3_idx_u8__50_comb;
  assign p3_eq_10760_comb = p3_run_size_str_u8__1_comb == 8'h71;
  assign p3_eq_10761_comb = p3_run_size_str_u8__1_comb == p3_idx_u8__2_comb;
  assign p3_or_10762_comb = p3_eq_10734_comb | p3_eq_10735_comb;
  assign p3_concat_10767_comb = {p3_eq_10736_comb | p3_eq_10737_comb | p3_eq_10738_comb | p3_eq_10739_comb | p3_eq_10740_comb | p3_eq_10741_comb | p3_eq_10742_comb | p3_eq_10743_comb | p3_eq_10744_comb | p3_eq_10745_comb | p3_eq_10746_comb | p3_eq_10747_comb | p3_eq_10748_comb, p3_eq_10749_comb | p3_eq_10750_comb | p3_eq_10751_comb | p3_eq_10752_comb | p3_eq_10753_comb | p3_eq_10754_comb | p3_eq_10755_comb, p3_eq_10756_comb | p3_eq_10734_comb | p3_eq_10735_comb | p3_eq_10757_comb | p3_eq_10758_comb | p3_eq_10759_comb | p3_eq_10760_comb | p3_eq_10761_comb};
  assign p3_idx_u8__1_squeezed__2_comb = 2'h1;
  assign p3_idx_u8__3_squeezed__1_comb = 2'h3;
  assign p3_concat_10776_comb = {p3_eq_10754_comb, p3_eq_10755_comb, p3_eq_10756_comb, p3_or_10762_comb, p3_eq_10757_comb, p3_eq_10758_comb, p3_eq_10759_comb, p3_eq_10760_comb, p3_eq_10761_comb};
  assign p3_idx_u8__6_squeezed__2_comb = 3'h6;
  assign p3_idx_u8__4_squeezed__2_comb = 3'h4;
  assign p3_idx_u8__5_squeezed__2_comb = 3'h5;
  assign p3_idx_u8__6_squeezed__3_comb = 3'h6;
  assign p3_idx_u8__7_squeezed__2_comb = 3'h7;
  assign p3_one_hot_sel_10859_comb = 2'h0 & {2{p3_concat_10767_comb[0]}} | p3_idx_u8__1_squeezed__2_comb & {2{p3_concat_10767_comb[1]}} | p3_idx_u8__3_squeezed__1_comb & {2{p3_concat_10767_comb[2]}};
  assign p3_concat_10788_comb = {p3_eq_10736_comb, p3_eq_10737_comb, p3_eq_10738_comb, p3_eq_10739_comb, p3_eq_10740_comb, p3_eq_10741_comb, p3_eq_10742_comb, p3_eq_10743_comb, p3_eq_10744_comb, p3_eq_10745_comb, p3_eq_10746_comb, p3_eq_10747_comb, p3_eq_10748_comb, p3_eq_10749_comb, p3_eq_10750_comb, p3_eq_10751_comb, p3_eq_10752_comb, p3_eq_10753_comb, p3_eq_10754_comb, p3_eq_10755_comb, p3_eq_10756_comb, p3_eq_10734_comb, p3_eq_10735_comb, p3_eq_10757_comb, p3_eq_10758_comb, p3_eq_10759_comb, p3_eq_10760_comb, p3_eq_10761_comb};
  assign p3_huffman_length_squeezed_comb = p2_is_luminance ? {(p3_eq_10736_comb | p3_eq_10737_comb | p3_eq_10738_comb | p3_eq_10739_comb | p3_eq_10740_comb | p3_eq_10741_comb | p3_eq_10742_comb | p3_eq_10743_comb | p3_eq_10744_comb | p3_eq_10745_comb | p3_eq_10746_comb | p3_eq_10747_comb | p3_eq_10748_comb | p3_eq_10749_comb | p3_eq_10750_comb | p3_eq_10751_comb | p3_eq_10752_comb | p3_eq_10753_comb) & ~(p3_eq_10754_comb | p3_eq_10755_comb | p3_eq_10756_comb | p3_or_10762_comb | p3_eq_10757_comb | p3_eq_10758_comb | p3_eq_10759_comb | p3_eq_10760_comb | p3_eq_10761_comb), (p3_eq_10754_comb | p3_eq_10755_comb | p3_eq_10756_comb | p3_or_10762_comb | p3_eq_10757_comb | p3_eq_10758_comb | p3_eq_10759_comb | p3_eq_10760_comb) & ~p3_eq_10761_comb, p3_idx_u8__6_squeezed__2_comb & {3{p3_concat_10776_comb[0]}} | 3'h0 & {3{p3_concat_10776_comb[1]}} | 3'h1 & {3{p3_concat_10776_comb[2]}} | 3'h2 & {3{p3_concat_10776_comb[3]}} | 3'h3 & {3{p3_concat_10776_comb[4]}} | p3_idx_u8__4_squeezed__2_comb & {3{p3_concat_10776_comb[5]}} | p3_idx_u8__5_squeezed__2_comb & {3{p3_concat_10776_comb[6]}} | p3_idx_u8__6_squeezed__3_comb & {3{p3_concat_10776_comb[7]}} | p3_idx_u8__7_squeezed__2_comb & {3{p3_concat_10776_comb[8]}}} : literal_10818[p3_run_size_str_u8__1_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8__1_comb];
  assign p3_idx_u8__2_squeezed__1_comb = 5'h02;
  assign p3_huffman_code_full_comb = p2_is_luminance ? {{{1{p3_one_hot_sel_10859_comb[1]}}, p3_one_hot_sel_10859_comb}, 13'h003a & {13{p3_concat_10788_comb[0]}} | 13'h00f9 & {13{p3_concat_10788_comb[1]}} | 13'h01f6 & {13{p3_concat_10788_comb[2]}} | 13'h03f5 & {13{p3_concat_10788_comb[3]}} | 13'h07f7 & {13{p3_concat_10788_comb[4]}} | 13'h0ff3 & {13{p3_concat_10788_comb[5]}} | 13'h0ff5 & {13{p3_concat_10788_comb[6]}} | 13'h1fed & {13{p3_concat_10788_comb[7]}} | 13'h1fe0 & {13{p3_concat_10788_comb[8]}} | 13'h1fe4 & {13{p3_concat_10788_comb[9]}} | 13'h1fe6 & {13{p3_concat_10788_comb[10]}} | 13'h1fe8 & {13{p3_concat_10788_comb[11]}} | 13'h1fed & {13{p3_concat_10788_comb[12]}} | 13'h1fee & {13{p3_concat_10788_comb[13]}} | 13'h1ff2 & {13{p3_concat_10788_comb[14]}} | 13'h1fd6 & {13{p3_concat_10788_comb[15]}} | 13'h1fd4 & {13{p3_concat_10788_comb[16]}} | 13'h1fd8 & {13{p3_concat_10788_comb[17]}} | 13'h1fdb & {13{p3_concat_10788_comb[18]}} | 13'h1fdd & {13{p3_concat_10788_comb[19]}} | 13'h1fe1 & {13{p3_concat_10788_comb[20]}} | 13'h1fea & {13{p3_concat_10788_comb[21]}} | 13'h1fec & {13{p3_concat_10788_comb[22]}} | 13'h1ff0 & {13{p3_concat_10788_comb[23]}} | 13'h1ff4 & {13{p3_concat_10788_comb[24]}} | 13'h1ff5 & {13{p3_concat_10788_comb[25]}} | 13'h1ff9 & {13{p3_concat_10788_comb[26]}} | 13'h1ffd & {13{p3_concat_10788_comb[27]}}} : literal_10822[p3_run_size_str_u8__1_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8__1_comb];
  assign p3_one_hot_10842_comb = {p3_concat_10788_comb[27:0] == 28'h000_0000, p3_concat_10788_comb[27] && p3_concat_10788_comb[26:0] == 27'h000_0000, p3_concat_10788_comb[26] && p3_concat_10788_comb[25:0] == 26'h000_0000, p3_concat_10788_comb[25] && p3_concat_10788_comb[24:0] == 25'h000_0000, p3_concat_10788_comb[24] && p3_concat_10788_comb[23:0] == 24'h00_0000, p3_concat_10788_comb[23] && p3_concat_10788_comb[22:0] == 23'h00_0000, p3_concat_10788_comb[22] && p3_concat_10788_comb[21:0] == 22'h00_0000, p3_concat_10788_comb[21] && p3_concat_10788_comb[20:0] == 21'h00_0000, p3_concat_10788_comb[20] && p3_concat_10788_comb[19:0] == 20'h0_0000, p3_concat_10788_comb[19] && p3_concat_10788_comb[18:0] == 19'h0_0000, p3_concat_10788_comb[18] && p3_concat_10788_comb[17:0] == 18'h0_0000, p3_concat_10788_comb[17] && p3_concat_10788_comb[16:0] == 17'h0_0000, p3_concat_10788_comb[16] && p3_concat_10788_comb[15:0] == 16'h0000, p3_concat_10788_comb[15] && p3_concat_10788_comb[14:0] == 15'h0000, p3_concat_10788_comb[14] && p3_concat_10788_comb[13:0] == 14'h0000, p3_concat_10788_comb[13] && p3_concat_10788_comb[12:0] == 13'h0000, p3_concat_10788_comb[12] && p3_concat_10788_comb[11:0] == 12'h000, p3_concat_10788_comb[11] && p3_concat_10788_comb[10:0] == 11'h000, p3_concat_10788_comb[10] && p3_concat_10788_comb[9:0] == 10'h000, p3_concat_10788_comb[9] && p3_concat_10788_comb[8:0] == 9'h000, p3_concat_10788_comb[8] && p3_concat_10788_comb[7:0] == 8'h00, p3_concat_10788_comb[7] && p3_concat_10788_comb[6:0] == 7'h00, p3_concat_10788_comb[6] && p3_concat_10788_comb[5:0] == 6'h00, p3_concat_10788_comb[5] && p3_concat_10788_comb[4:0] == 5'h00, p3_concat_10788_comb[4] && p3_concat_10788_comb[3:0] == 4'h0, p3_concat_10788_comb[3] && p3_concat_10788_comb[2:0] == 3'h0, p3_concat_10788_comb[2] && p3_concat_10788_comb[1:0] == 2'h0, p3_concat_10788_comb[1] && !p3_concat_10788_comb[0], p3_concat_10788_comb[0]};
  assign p3_one_hot_10848_comb = {p3_concat_10776_comb[8:0] == 9'h000, p3_concat_10776_comb[8] && p3_concat_10776_comb[7:0] == 8'h00, p3_concat_10776_comb[7] && p3_concat_10776_comb[6:0] == 7'h00, p3_concat_10776_comb[6] && p3_concat_10776_comb[5:0] == 6'h00, p3_concat_10776_comb[5] && p3_concat_10776_comb[4:0] == 5'h00, p3_concat_10776_comb[4] && p3_concat_10776_comb[3:0] == 4'h0, p3_concat_10776_comb[3] && p3_concat_10776_comb[2:0] == 3'h0, p3_concat_10776_comb[2] && p3_concat_10776_comb[1:0] == 2'h0, p3_concat_10776_comb[1] && !p3_concat_10776_comb[0], p3_concat_10776_comb[0]};
  assign p3_one_hot_10854_comb = {p3_concat_10767_comb[2:0] == 3'h0, p3_concat_10767_comb[2] && p3_concat_10767_comb[1:0] == 2'h0, p3_concat_10767_comb[1] && !p3_concat_10767_comb[0], p3_concat_10767_comb[0]};
  assign p3_tuple_10838_comb = {p3_huffman_code_full_comb & {16{~p2_or_10654}}, {3'h0, p2_or_10654 ? p3_idx_u8__2_squeezed__1_comb : p3_huffman_length_squeezed_comb}, p2_sel_10664, p2_sel_10665};

  // Registers for pipe stage 3:
  reg [35:0] p3_tuple_10838;
  always @ (posedge clk) begin
    p3_tuple_10838 <= p3_tuple_10838_comb;
  end
  assign out = p3_tuple_10838;
endmodule
