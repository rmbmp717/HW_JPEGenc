module Huffman_enc_controller(
  input  wire               clock,
  input  wire               reset_n,
  input  wire               Huffman_start,
  input  wire  [511:0]      zigzag_pix_in,
  output reg   [511:0]      dc_matrix,
  output reg   [511:0]      ac_matrix,
  output reg   [7:0]        start_pix,
  // from enc module
  input  wire  [23:0]       dc_out,
  input  wire  [15:0]       ac_out,
  input  wire  [7:0]        length,
  input  wire  [7:0]        code,
  input  wire  [3:0]        run,
  // final output 
  output reg                jpeg_out_enable,
  output reg   [23:0]       jpeg_dc_out,
  output reg   [15:0]       jpeg_out,
  output reg   [3:0]        jpeg_data_length,
  output reg   [7:0]        code_out
);

  // 状態レジスタ: 初回はDCを出力、その後はACを出力
  reg [3:0] state;  // 0: DC, 1: AC
  always @(posedge clock or negedge reset_n) begin
    if (!reset_n) begin
      state <= 0;
      dc_matrix <= 0;
      ac_matrix <= 0;
      start_pix <= 0;
      jpeg_out_enable <= 0;
      jpeg_dc_out <= 0;
      jpeg_out <= 0;
      jpeg_data_length <= 0;
      code_out <= 0;
    end else begin
      case(state)
        0: begin
          dc_matrix <= 0;
          jpeg_out_enable <= 0;
          if(Huffman_start) begin
            state <= 1;
          end
        end
        // DC enc Start
        1: begin
          jpeg_out_enable <= 0;
          dc_matrix <= zigzag_pix_in;
          state <= 2;
        end
        2: begin
          state <= 3;
          start_pix <= 1;
          jpeg_dc_out <= dc_out;
        end
        // AC enc Start
        3: begin
          if(start_pix >= 63) begin
            state <= 0;
          end else begin
            jpeg_out_enable <= 0;
            ac_matrix <= zigzag_pix_in;
            state <= 4;
          end
        end
        4: begin
          state <= 5;
        end
        5: begin
          state <= 6;
        end
        6: begin
          state <= 7;
        end
        7: begin
          state <= 8;
        end
        8: begin
          jpeg_out_enable <= 1;
          start_pix <= start_pix + run + 1;
          jpeg_out <= ac_out;
          jpeg_data_length <= length;
          state <= 3;
          code_out <= code; 
        end
      endcase
    end
  end

  //assign jpeg_out = 0;
  //assign jpeg_data_bits = 0;

endmodule
