module Quantize(
  input wire clk,
  input wire [639:0] dct_coeffs,
  input wire [7:0] matrix_row,
  input wire is_luminance,
  input wire quantize_off,
  output wire [79:0] out
);
  function automatic [31:0] sdiv_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    begin
      sdiv_32b = rhs == 32'h0000_0000 ? (lhs[31] ? 32'h8000_0000 : 32'h7fff_ffff) : (lhs == 32'h8000_0000 && rhs == 32'hffff_ffff ? 32'h8000_0000 : $unsigned($signed(lhs) / $signed(rhs)));
    end
  endfunction
  wire [15:0] CHROMINANCE_QUANT_TBL[0:7][0:7];
  assign CHROMINANCE_QUANT_TBL[0][0] = 16'h0022;
  assign CHROMINANCE_QUANT_TBL[0][1] = 16'h0024;
  assign CHROMINANCE_QUANT_TBL[0][2] = 16'h0030;
  assign CHROMINANCE_QUANT_TBL[0][3] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[0][4] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[0][5] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[0][6] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[0][7] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[1][0] = 16'h0024;
  assign CHROMINANCE_QUANT_TBL[1][1] = 16'h002a;
  assign CHROMINANCE_QUANT_TBL[1][2] = 16'h0034;
  assign CHROMINANCE_QUANT_TBL[1][3] = 16'h0084;
  assign CHROMINANCE_QUANT_TBL[1][4] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[1][5] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[1][6] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[1][7] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[2][0] = 16'h0030;
  assign CHROMINANCE_QUANT_TBL[2][1] = 16'h0034;
  assign CHROMINANCE_QUANT_TBL[2][2] = 16'h0070;
  assign CHROMINANCE_QUANT_TBL[2][3] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[2][4] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[2][5] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[2][6] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[2][7] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[3][0] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[3][1] = 16'h0084;
  assign CHROMINANCE_QUANT_TBL[3][2] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[3][3] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[3][4] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[3][5] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[3][6] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[3][7] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[4][0] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[4][1] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[4][2] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[4][3] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[4][4] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[4][5] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[4][6] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[4][7] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[5][0] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[5][1] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[5][2] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[5][3] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[5][4] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[5][5] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[5][6] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[5][7] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[6][0] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[6][1] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[6][2] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[6][3] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[6][4] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[6][5] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[6][6] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[6][7] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[7][0] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[7][1] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[7][2] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[7][3] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[7][4] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[7][5] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[7][6] = 16'h00c6;
  assign CHROMINANCE_QUANT_TBL[7][7] = 16'h00c6;
  wire [15:0] LUMINANCE_QUANT_TBL[0:7][0:7];
  assign LUMINANCE_QUANT_TBL[0][0] = 16'h0020;
  assign LUMINANCE_QUANT_TBL[0][1] = 16'h0016;
  assign LUMINANCE_QUANT_TBL[0][2] = 16'h0014;
  assign LUMINANCE_QUANT_TBL[0][3] = 16'h0020;
  assign LUMINANCE_QUANT_TBL[0][4] = 16'h0030;
  assign LUMINANCE_QUANT_TBL[0][5] = 16'h0050;
  assign LUMINANCE_QUANT_TBL[0][6] = 16'h0066;
  assign LUMINANCE_QUANT_TBL[0][7] = 16'h007a;
  assign LUMINANCE_QUANT_TBL[1][0] = 16'h0018;
  assign LUMINANCE_QUANT_TBL[1][1] = 16'h0018;
  assign LUMINANCE_QUANT_TBL[1][2] = 16'h001c;
  assign LUMINANCE_QUANT_TBL[1][3] = 16'h0026;
  assign LUMINANCE_QUANT_TBL[1][4] = 16'h0034;
  assign LUMINANCE_QUANT_TBL[1][5] = 16'h0074;
  assign LUMINANCE_QUANT_TBL[1][6] = 16'h0078;
  assign LUMINANCE_QUANT_TBL[1][7] = 16'h006e;
  assign LUMINANCE_QUANT_TBL[2][0] = 16'h001c;
  assign LUMINANCE_QUANT_TBL[2][1] = 16'h001a;
  assign LUMINANCE_QUANT_TBL[2][2] = 16'h0020;
  assign LUMINANCE_QUANT_TBL[2][3] = 16'h0030;
  assign LUMINANCE_QUANT_TBL[2][4] = 16'h0050;
  assign LUMINANCE_QUANT_TBL[2][5] = 16'h0072;
  assign LUMINANCE_QUANT_TBL[2][6] = 16'h008a;
  assign LUMINANCE_QUANT_TBL[2][7] = 16'h0070;
  assign LUMINANCE_QUANT_TBL[3][0] = 16'h001c;
  assign LUMINANCE_QUANT_TBL[3][1] = 16'h0022;
  assign LUMINANCE_QUANT_TBL[3][2] = 16'h002c;
  assign LUMINANCE_QUANT_TBL[3][3] = 16'h003a;
  assign LUMINANCE_QUANT_TBL[3][4] = 16'h0066;
  assign LUMINANCE_QUANT_TBL[3][5] = 16'h00ae;
  assign LUMINANCE_QUANT_TBL[3][6] = 16'h00a0;
  assign LUMINANCE_QUANT_TBL[3][7] = 16'h007c;
  assign LUMINANCE_QUANT_TBL[4][0] = 16'h0024;
  assign LUMINANCE_QUANT_TBL[4][1] = 16'h002c;
  assign LUMINANCE_QUANT_TBL[4][2] = 16'h004a;
  assign LUMINANCE_QUANT_TBL[4][3] = 16'h0070;
  assign LUMINANCE_QUANT_TBL[4][4] = 16'h0088;
  assign LUMINANCE_QUANT_TBL[4][5] = 16'h00da;
  assign LUMINANCE_QUANT_TBL[4][6] = 16'h00ce;
  assign LUMINANCE_QUANT_TBL[4][7] = 16'h009a;
  assign LUMINANCE_QUANT_TBL[5][0] = 16'h0030;
  assign LUMINANCE_QUANT_TBL[5][1] = 16'h0046;
  assign LUMINANCE_QUANT_TBL[5][2] = 16'h006e;
  assign LUMINANCE_QUANT_TBL[5][3] = 16'h0080;
  assign LUMINANCE_QUANT_TBL[5][4] = 16'h00a2;
  assign LUMINANCE_QUANT_TBL[5][5] = 16'h00d0;
  assign LUMINANCE_QUANT_TBL[5][6] = 16'h00e2;
  assign LUMINANCE_QUANT_TBL[5][7] = 16'h00b8;
  assign LUMINANCE_QUANT_TBL[6][0] = 16'h0062;
  assign LUMINANCE_QUANT_TBL[6][1] = 16'h0080;
  assign LUMINANCE_QUANT_TBL[6][2] = 16'h009c;
  assign LUMINANCE_QUANT_TBL[6][3] = 16'h00ae;
  assign LUMINANCE_QUANT_TBL[6][4] = 16'h00ce;
  assign LUMINANCE_QUANT_TBL[6][5] = 16'h00f2;
  assign LUMINANCE_QUANT_TBL[6][6] = 16'h00f0;
  assign LUMINANCE_QUANT_TBL[6][7] = 16'h00ca;
  assign LUMINANCE_QUANT_TBL[7][0] = 16'h0090;
  assign LUMINANCE_QUANT_TBL[7][1] = 16'h00b8;
  assign LUMINANCE_QUANT_TBL[7][2] = 16'h00be;
  assign LUMINANCE_QUANT_TBL[7][3] = 16'h00c4;
  assign LUMINANCE_QUANT_TBL[7][4] = 16'h00e0;
  assign LUMINANCE_QUANT_TBL[7][5] = 16'h00c8;
  assign LUMINANCE_QUANT_TBL[7][6] = 16'h00ce;
  assign LUMINANCE_QUANT_TBL[7][7] = 16'h00c6;
  wire [9:0] dct_coeffs_unflattened[0:7][0:7];
  assign dct_coeffs_unflattened[0][0] = dct_coeffs[9:0];
  assign dct_coeffs_unflattened[0][1] = dct_coeffs[19:10];
  assign dct_coeffs_unflattened[0][2] = dct_coeffs[29:20];
  assign dct_coeffs_unflattened[0][3] = dct_coeffs[39:30];
  assign dct_coeffs_unflattened[0][4] = dct_coeffs[49:40];
  assign dct_coeffs_unflattened[0][5] = dct_coeffs[59:50];
  assign dct_coeffs_unflattened[0][6] = dct_coeffs[69:60];
  assign dct_coeffs_unflattened[0][7] = dct_coeffs[79:70];
  assign dct_coeffs_unflattened[1][0] = dct_coeffs[89:80];
  assign dct_coeffs_unflattened[1][1] = dct_coeffs[99:90];
  assign dct_coeffs_unflattened[1][2] = dct_coeffs[109:100];
  assign dct_coeffs_unflattened[1][3] = dct_coeffs[119:110];
  assign dct_coeffs_unflattened[1][4] = dct_coeffs[129:120];
  assign dct_coeffs_unflattened[1][5] = dct_coeffs[139:130];
  assign dct_coeffs_unflattened[1][6] = dct_coeffs[149:140];
  assign dct_coeffs_unflattened[1][7] = dct_coeffs[159:150];
  assign dct_coeffs_unflattened[2][0] = dct_coeffs[169:160];
  assign dct_coeffs_unflattened[2][1] = dct_coeffs[179:170];
  assign dct_coeffs_unflattened[2][2] = dct_coeffs[189:180];
  assign dct_coeffs_unflattened[2][3] = dct_coeffs[199:190];
  assign dct_coeffs_unflattened[2][4] = dct_coeffs[209:200];
  assign dct_coeffs_unflattened[2][5] = dct_coeffs[219:210];
  assign dct_coeffs_unflattened[2][6] = dct_coeffs[229:220];
  assign dct_coeffs_unflattened[2][7] = dct_coeffs[239:230];
  assign dct_coeffs_unflattened[3][0] = dct_coeffs[249:240];
  assign dct_coeffs_unflattened[3][1] = dct_coeffs[259:250];
  assign dct_coeffs_unflattened[3][2] = dct_coeffs[269:260];
  assign dct_coeffs_unflattened[3][3] = dct_coeffs[279:270];
  assign dct_coeffs_unflattened[3][4] = dct_coeffs[289:280];
  assign dct_coeffs_unflattened[3][5] = dct_coeffs[299:290];
  assign dct_coeffs_unflattened[3][6] = dct_coeffs[309:300];
  assign dct_coeffs_unflattened[3][7] = dct_coeffs[319:310];
  assign dct_coeffs_unflattened[4][0] = dct_coeffs[329:320];
  assign dct_coeffs_unflattened[4][1] = dct_coeffs[339:330];
  assign dct_coeffs_unflattened[4][2] = dct_coeffs[349:340];
  assign dct_coeffs_unflattened[4][3] = dct_coeffs[359:350];
  assign dct_coeffs_unflattened[4][4] = dct_coeffs[369:360];
  assign dct_coeffs_unflattened[4][5] = dct_coeffs[379:370];
  assign dct_coeffs_unflattened[4][6] = dct_coeffs[389:380];
  assign dct_coeffs_unflattened[4][7] = dct_coeffs[399:390];
  assign dct_coeffs_unflattened[5][0] = dct_coeffs[409:400];
  assign dct_coeffs_unflattened[5][1] = dct_coeffs[419:410];
  assign dct_coeffs_unflattened[5][2] = dct_coeffs[429:420];
  assign dct_coeffs_unflattened[5][3] = dct_coeffs[439:430];
  assign dct_coeffs_unflattened[5][4] = dct_coeffs[449:440];
  assign dct_coeffs_unflattened[5][5] = dct_coeffs[459:450];
  assign dct_coeffs_unflattened[5][6] = dct_coeffs[469:460];
  assign dct_coeffs_unflattened[5][7] = dct_coeffs[479:470];
  assign dct_coeffs_unflattened[6][0] = dct_coeffs[489:480];
  assign dct_coeffs_unflattened[6][1] = dct_coeffs[499:490];
  assign dct_coeffs_unflattened[6][2] = dct_coeffs[509:500];
  assign dct_coeffs_unflattened[6][3] = dct_coeffs[519:510];
  assign dct_coeffs_unflattened[6][4] = dct_coeffs[529:520];
  assign dct_coeffs_unflattened[6][5] = dct_coeffs[539:530];
  assign dct_coeffs_unflattened[6][6] = dct_coeffs[549:540];
  assign dct_coeffs_unflattened[6][7] = dct_coeffs[559:550];
  assign dct_coeffs_unflattened[7][0] = dct_coeffs[569:560];
  assign dct_coeffs_unflattened[7][1] = dct_coeffs[579:570];
  assign dct_coeffs_unflattened[7][2] = dct_coeffs[589:580];
  assign dct_coeffs_unflattened[7][3] = dct_coeffs[599:590];
  assign dct_coeffs_unflattened[7][4] = dct_coeffs[609:600];
  assign dct_coeffs_unflattened[7][5] = dct_coeffs[619:610];
  assign dct_coeffs_unflattened[7][6] = dct_coeffs[629:620];
  assign dct_coeffs_unflattened[7][7] = dct_coeffs[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_dct_coeffs[0:7][0:7];
  reg [7:0] p0_matrix_row;
  reg p0_is_luminance;
  reg p0_quantize_off;
  always @ (posedge clk) begin
    p0_dct_coeffs[0][0] <= dct_coeffs_unflattened[0][0];
    p0_dct_coeffs[0][1] <= dct_coeffs_unflattened[0][1];
    p0_dct_coeffs[0][2] <= dct_coeffs_unflattened[0][2];
    p0_dct_coeffs[0][3] <= dct_coeffs_unflattened[0][3];
    p0_dct_coeffs[0][4] <= dct_coeffs_unflattened[0][4];
    p0_dct_coeffs[0][5] <= dct_coeffs_unflattened[0][5];
    p0_dct_coeffs[0][6] <= dct_coeffs_unflattened[0][6];
    p0_dct_coeffs[0][7] <= dct_coeffs_unflattened[0][7];
    p0_dct_coeffs[1][0] <= dct_coeffs_unflattened[1][0];
    p0_dct_coeffs[1][1] <= dct_coeffs_unflattened[1][1];
    p0_dct_coeffs[1][2] <= dct_coeffs_unflattened[1][2];
    p0_dct_coeffs[1][3] <= dct_coeffs_unflattened[1][3];
    p0_dct_coeffs[1][4] <= dct_coeffs_unflattened[1][4];
    p0_dct_coeffs[1][5] <= dct_coeffs_unflattened[1][5];
    p0_dct_coeffs[1][6] <= dct_coeffs_unflattened[1][6];
    p0_dct_coeffs[1][7] <= dct_coeffs_unflattened[1][7];
    p0_dct_coeffs[2][0] <= dct_coeffs_unflattened[2][0];
    p0_dct_coeffs[2][1] <= dct_coeffs_unflattened[2][1];
    p0_dct_coeffs[2][2] <= dct_coeffs_unflattened[2][2];
    p0_dct_coeffs[2][3] <= dct_coeffs_unflattened[2][3];
    p0_dct_coeffs[2][4] <= dct_coeffs_unflattened[2][4];
    p0_dct_coeffs[2][5] <= dct_coeffs_unflattened[2][5];
    p0_dct_coeffs[2][6] <= dct_coeffs_unflattened[2][6];
    p0_dct_coeffs[2][7] <= dct_coeffs_unflattened[2][7];
    p0_dct_coeffs[3][0] <= dct_coeffs_unflattened[3][0];
    p0_dct_coeffs[3][1] <= dct_coeffs_unflattened[3][1];
    p0_dct_coeffs[3][2] <= dct_coeffs_unflattened[3][2];
    p0_dct_coeffs[3][3] <= dct_coeffs_unflattened[3][3];
    p0_dct_coeffs[3][4] <= dct_coeffs_unflattened[3][4];
    p0_dct_coeffs[3][5] <= dct_coeffs_unflattened[3][5];
    p0_dct_coeffs[3][6] <= dct_coeffs_unflattened[3][6];
    p0_dct_coeffs[3][7] <= dct_coeffs_unflattened[3][7];
    p0_dct_coeffs[4][0] <= dct_coeffs_unflattened[4][0];
    p0_dct_coeffs[4][1] <= dct_coeffs_unflattened[4][1];
    p0_dct_coeffs[4][2] <= dct_coeffs_unflattened[4][2];
    p0_dct_coeffs[4][3] <= dct_coeffs_unflattened[4][3];
    p0_dct_coeffs[4][4] <= dct_coeffs_unflattened[4][4];
    p0_dct_coeffs[4][5] <= dct_coeffs_unflattened[4][5];
    p0_dct_coeffs[4][6] <= dct_coeffs_unflattened[4][6];
    p0_dct_coeffs[4][7] <= dct_coeffs_unflattened[4][7];
    p0_dct_coeffs[5][0] <= dct_coeffs_unflattened[5][0];
    p0_dct_coeffs[5][1] <= dct_coeffs_unflattened[5][1];
    p0_dct_coeffs[5][2] <= dct_coeffs_unflattened[5][2];
    p0_dct_coeffs[5][3] <= dct_coeffs_unflattened[5][3];
    p0_dct_coeffs[5][4] <= dct_coeffs_unflattened[5][4];
    p0_dct_coeffs[5][5] <= dct_coeffs_unflattened[5][5];
    p0_dct_coeffs[5][6] <= dct_coeffs_unflattened[5][6];
    p0_dct_coeffs[5][7] <= dct_coeffs_unflattened[5][7];
    p0_dct_coeffs[6][0] <= dct_coeffs_unflattened[6][0];
    p0_dct_coeffs[6][1] <= dct_coeffs_unflattened[6][1];
    p0_dct_coeffs[6][2] <= dct_coeffs_unflattened[6][2];
    p0_dct_coeffs[6][3] <= dct_coeffs_unflattened[6][3];
    p0_dct_coeffs[6][4] <= dct_coeffs_unflattened[6][4];
    p0_dct_coeffs[6][5] <= dct_coeffs_unflattened[6][5];
    p0_dct_coeffs[6][6] <= dct_coeffs_unflattened[6][6];
    p0_dct_coeffs[6][7] <= dct_coeffs_unflattened[6][7];
    p0_dct_coeffs[7][0] <= dct_coeffs_unflattened[7][0];
    p0_dct_coeffs[7][1] <= dct_coeffs_unflattened[7][1];
    p0_dct_coeffs[7][2] <= dct_coeffs_unflattened[7][2];
    p0_dct_coeffs[7][3] <= dct_coeffs_unflattened[7][3];
    p0_dct_coeffs[7][4] <= dct_coeffs_unflattened[7][4];
    p0_dct_coeffs[7][5] <= dct_coeffs_unflattened[7][5];
    p0_dct_coeffs[7][6] <= dct_coeffs_unflattened[7][6];
    p0_dct_coeffs[7][7] <= dct_coeffs_unflattened[7][7];
    p0_matrix_row <= matrix_row;
    p0_is_luminance <= is_luminance;
    p0_quantize_off <= quantize_off;
  end

  // ===== Pipe stage 1:
  wire [9:0] p1_array_index_831_comb;
  wire [6:0] p1_q_value_squeezed_comb;
  wire p1_q_value_squeezed_const_lsb_bits_comb;
  wire [9:0] p1_array_index_835_comb;
  wire [6:0] p1_q_value__1_squeezed_comb;
  wire p1_q_value_squeezed_const_lsb_bits__1_comb;
  wire [9:0] p1_array_index_839_comb;
  wire [6:0] p1_q_value__2_squeezed_comb;
  wire p1_q_value_squeezed_const_lsb_bits__2_comb;
  wire [9:0] p1_array_index_843_comb;
  wire [6:0] p1_q_value__3_squeezed_comb;
  wire p1_q_value_squeezed_const_lsb_bits__3_comb;
  wire [9:0] p1_array_index_847_comb;
  wire [6:0] p1_q_value__4_squeezed_comb;
  wire p1_q_value_squeezed_const_lsb_bits__4_comb;
  wire [9:0] p1_array_index_851_comb;
  wire [6:0] p1_q_value__5_squeezed_comb;
  wire p1_q_value_squeezed_const_lsb_bits__5_comb;
  wire [9:0] p1_array_index_855_comb;
  wire [6:0] p1_q_value__6_squeezed_comb;
  wire p1_q_value_squeezed_const_lsb_bits__6_comb;
  wire [9:0] p1_array_index_859_comb;
  wire [6:0] p1_q_value__7_squeezed_comb;
  wire p1_q_value_squeezed_const_lsb_bits__7_comb;
  wire [31:0] p1_sdiv_879_comb;
  wire [31:0] p1_sdiv_880_comb;
  wire [31:0] p1_sdiv_881_comb;
  wire [31:0] p1_sdiv_882_comb;
  wire [31:0] p1_sdiv_883_comb;
  wire [31:0] p1_sdiv_884_comb;
  wire [31:0] p1_sdiv_885_comb;
  wire [31:0] p1_sdiv_886_comb;
  wire [9:0] p1_divided_squeezed_comb;
  wire [9:0] p1_divided__1_squeezed_comb;
  wire [9:0] p1_divided__2_squeezed_comb;
  wire [9:0] p1_divided__3_squeezed_comb;
  wire [9:0] p1_divided__4_squeezed_comb;
  wire [9:0] p1_divided__5_squeezed_comb;
  wire [9:0] p1_divided__6_squeezed_comb;
  wire [9:0] p1_divided__7_squeezed_comb;
  wire [9:0] p1_clipped_comb;
  wire [9:0] p1_clipped__1_comb;
  wire [9:0] p1_clipped__2_comb;
  wire [9:0] p1_clipped__3_comb;
  wire [9:0] p1_clipped__4_comb;
  wire [9:0] p1_clipped__5_comb;
  wire [9:0] p1_clipped__6_comb;
  wire [9:0] p1_clipped__7_comb;
  wire [9:0] p1_array_967_comb[0:7];
  assign p1_array_index_831_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h0];
  assign p1_q_value_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h0][7:1] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h0][7:1];
  assign p1_q_value_squeezed_const_lsb_bits_comb = 1'h0;
  assign p1_array_index_835_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h1];
  assign p1_q_value__1_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h1][7:1] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h1][7:1];
  assign p1_q_value_squeezed_const_lsb_bits__1_comb = 1'h0;
  assign p1_array_index_839_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h2];
  assign p1_q_value__2_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h2][7:1] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h2][7:1];
  assign p1_q_value_squeezed_const_lsb_bits__2_comb = 1'h0;
  assign p1_array_index_843_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h3];
  assign p1_q_value__3_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h3][7:1] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h3][7:1];
  assign p1_q_value_squeezed_const_lsb_bits__3_comb = 1'h0;
  assign p1_array_index_847_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h4];
  assign p1_q_value__4_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h4][7:1] : 7'h63;
  assign p1_q_value_squeezed_const_lsb_bits__4_comb = 1'h0;
  assign p1_array_index_851_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h5];
  assign p1_q_value__5_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h5][7:1] : 7'h63;
  assign p1_q_value_squeezed_const_lsb_bits__5_comb = 1'h0;
  assign p1_array_index_855_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h6];
  assign p1_q_value__6_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h6][7:1] : 7'h63;
  assign p1_q_value_squeezed_const_lsb_bits__6_comb = 1'h0;
  assign p1_array_index_859_comb = p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h7];
  assign p1_q_value__7_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h7][7:1] : 7'h63;
  assign p1_q_value_squeezed_const_lsb_bits__7_comb = 1'h0;
  assign p1_sdiv_879_comb = sdiv_32b({{22{p1_array_index_831_comb[9]}}, p1_array_index_831_comb}, {24'h00_0000, p1_q_value_squeezed_comb, p1_q_value_squeezed_const_lsb_bits_comb});
  assign p1_sdiv_880_comb = sdiv_32b({{22{p1_array_index_835_comb[9]}}, p1_array_index_835_comb}, {24'h00_0000, p1_q_value__1_squeezed_comb, p1_q_value_squeezed_const_lsb_bits__1_comb});
  assign p1_sdiv_881_comb = sdiv_32b({{22{p1_array_index_839_comb[9]}}, p1_array_index_839_comb}, {24'h00_0000, p1_q_value__2_squeezed_comb, p1_q_value_squeezed_const_lsb_bits__2_comb});
  assign p1_sdiv_882_comb = sdiv_32b({{22{p1_array_index_843_comb[9]}}, p1_array_index_843_comb}, {24'h00_0000, p1_q_value__3_squeezed_comb, p1_q_value_squeezed_const_lsb_bits__3_comb});
  assign p1_sdiv_883_comb = sdiv_32b({{22{p1_array_index_847_comb[9]}}, p1_array_index_847_comb}, {24'h00_0000, p1_q_value__4_squeezed_comb, p1_q_value_squeezed_const_lsb_bits__4_comb});
  assign p1_sdiv_884_comb = sdiv_32b({{22{p1_array_index_851_comb[9]}}, p1_array_index_851_comb}, {24'h00_0000, p1_q_value__5_squeezed_comb, p1_q_value_squeezed_const_lsb_bits__5_comb});
  assign p1_sdiv_885_comb = sdiv_32b({{22{p1_array_index_855_comb[9]}}, p1_array_index_855_comb}, {24'h00_0000, p1_q_value__6_squeezed_comb, p1_q_value_squeezed_const_lsb_bits__6_comb});
  assign p1_sdiv_886_comb = sdiv_32b({{22{p1_array_index_859_comb[9]}}, p1_array_index_859_comb}, {24'h00_0000, p1_q_value__7_squeezed_comb, p1_q_value_squeezed_const_lsb_bits__7_comb});
  assign p1_divided_squeezed_comb = p0_quantize_off ? p1_array_index_831_comb : p1_sdiv_879_comb[9:0];
  assign p1_divided__1_squeezed_comb = p0_quantize_off ? p1_array_index_835_comb : p1_sdiv_880_comb[9:0];
  assign p1_divided__2_squeezed_comb = p0_quantize_off ? p1_array_index_839_comb : p1_sdiv_881_comb[9:0];
  assign p1_divided__3_squeezed_comb = p0_quantize_off ? p1_array_index_843_comb : p1_sdiv_882_comb[9:0];
  assign p1_divided__4_squeezed_comb = p0_quantize_off ? p1_array_index_847_comb : p1_sdiv_883_comb[9:0];
  assign p1_divided__5_squeezed_comb = p0_quantize_off ? p1_array_index_851_comb : p1_sdiv_884_comb[9:0];
  assign p1_divided__6_squeezed_comb = p0_quantize_off ? p1_array_index_855_comb : p1_sdiv_885_comb[9:0];
  assign p1_divided__7_squeezed_comb = p0_quantize_off ? p1_array_index_859_comb : p1_sdiv_886_comb[9:0];
  assign p1_clipped_comb = $signed(p1_divided_squeezed_comb) > $signed(10'h0ff) ? 10'h0ff : p1_divided_squeezed_comb & {10{$signed(p1_divided_squeezed_comb) >= $signed(10'h301)}};
  assign p1_clipped__1_comb = $signed(p1_divided__1_squeezed_comb) > $signed(10'h0ff) ? 10'h0ff : p1_divided__1_squeezed_comb & {10{$signed(p1_divided__1_squeezed_comb) >= $signed(10'h301)}};
  assign p1_clipped__2_comb = $signed(p1_divided__2_squeezed_comb) > $signed(10'h0ff) ? 10'h0ff : p1_divided__2_squeezed_comb & {10{$signed(p1_divided__2_squeezed_comb) >= $signed(10'h301)}};
  assign p1_clipped__3_comb = $signed(p1_divided__3_squeezed_comb) > $signed(10'h0ff) ? 10'h0ff : p1_divided__3_squeezed_comb & {10{$signed(p1_divided__3_squeezed_comb) >= $signed(10'h301)}};
  assign p1_clipped__4_comb = $signed(p1_divided__4_squeezed_comb) > $signed(10'h0ff) ? 10'h0ff : p1_divided__4_squeezed_comb & {10{$signed(p1_divided__4_squeezed_comb) >= $signed(10'h301)}};
  assign p1_clipped__5_comb = $signed(p1_divided__5_squeezed_comb) > $signed(10'h0ff) ? 10'h0ff : p1_divided__5_squeezed_comb & {10{$signed(p1_divided__5_squeezed_comb) >= $signed(10'h301)}};
  assign p1_clipped__6_comb = $signed(p1_divided__6_squeezed_comb) > $signed(10'h0ff) ? 10'h0ff : p1_divided__6_squeezed_comb & {10{$signed(p1_divided__6_squeezed_comb) >= $signed(10'h301)}};
  assign p1_clipped__7_comb = $signed(p1_divided__7_squeezed_comb) > $signed(10'h0ff) ? 10'h0ff : p1_divided__7_squeezed_comb & {10{$signed(p1_divided__7_squeezed_comb) >= $signed(10'h301)}};
  assign p1_array_967_comb[0] = p1_clipped_comb;
  assign p1_array_967_comb[1] = p1_clipped__1_comb;
  assign p1_array_967_comb[2] = p1_clipped__2_comb;
  assign p1_array_967_comb[3] = p1_clipped__3_comb;
  assign p1_array_967_comb[4] = p1_clipped__4_comb;
  assign p1_array_967_comb[5] = p1_clipped__5_comb;
  assign p1_array_967_comb[6] = p1_clipped__6_comb;
  assign p1_array_967_comb[7] = p1_clipped__7_comb;

  // Registers for pipe stage 1:
  reg [9:0] p1_array_967[0:7];
  always @ (posedge clk) begin
    p1_array_967[0] <= p1_array_967_comb[0];
    p1_array_967[1] <= p1_array_967_comb[1];
    p1_array_967[2] <= p1_array_967_comb[2];
    p1_array_967[3] <= p1_array_967_comb[3];
    p1_array_967[4] <= p1_array_967_comb[4];
    p1_array_967[5] <= p1_array_967_comb[5];
    p1_array_967[6] <= p1_array_967_comb[6];
    p1_array_967[7] <= p1_array_967_comb[7];
  end
  assign out = {p1_array_967[7], p1_array_967[6], p1_array_967[5], p1_array_967[4], p1_array_967[3], p1_array_967[2], p1_array_967[1], p1_array_967[0]};
endmodule
