module Huffman_ACenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [57:0] out
);
  wire [4:0] literal_10861[0:251];
  assign literal_10861[0] = 5'h02;
  assign literal_10861[1] = 5'h02;
  assign literal_10861[2] = 5'h03;
  assign literal_10861[3] = 5'h04;
  assign literal_10861[4] = 5'h05;
  assign literal_10861[5] = 5'h07;
  assign literal_10861[6] = 5'h08;
  assign literal_10861[7] = 5'h0e;
  assign literal_10861[8] = 5'h10;
  assign literal_10861[9] = 5'h10;
  assign literal_10861[10] = 5'h10;
  assign literal_10861[11] = 5'h00;
  assign literal_10861[12] = 5'h00;
  assign literal_10861[13] = 5'h00;
  assign literal_10861[14] = 5'h00;
  assign literal_10861[15] = 5'h00;
  assign literal_10861[16] = 5'h00;
  assign literal_10861[17] = 5'h03;
  assign literal_10861[18] = 5'h06;
  assign literal_10861[19] = 5'h07;
  assign literal_10861[20] = 5'h09;
  assign literal_10861[21] = 5'h0b;
  assign literal_10861[22] = 5'h0d;
  assign literal_10861[23] = 5'h10;
  assign literal_10861[24] = 5'h10;
  assign literal_10861[25] = 5'h10;
  assign literal_10861[26] = 5'h10;
  assign literal_10861[27] = 5'h00;
  assign literal_10861[28] = 5'h00;
  assign literal_10861[29] = 5'h00;
  assign literal_10861[30] = 5'h00;
  assign literal_10861[31] = 5'h00;
  assign literal_10861[32] = 5'h00;
  assign literal_10861[33] = 5'h05;
  assign literal_10861[34] = 5'h07;
  assign literal_10861[35] = 5'h0a;
  assign literal_10861[36] = 5'h0c;
  assign literal_10861[37] = 5'h0d;
  assign literal_10861[38] = 5'h10;
  assign literal_10861[39] = 5'h10;
  assign literal_10861[40] = 5'h10;
  assign literal_10861[41] = 5'h10;
  assign literal_10861[42] = 5'h10;
  assign literal_10861[43] = 5'h00;
  assign literal_10861[44] = 5'h00;
  assign literal_10861[45] = 5'h00;
  assign literal_10861[46] = 5'h00;
  assign literal_10861[47] = 5'h00;
  assign literal_10861[48] = 5'h00;
  assign literal_10861[49] = 5'h06;
  assign literal_10861[50] = 5'h08;
  assign literal_10861[51] = 5'h0b;
  assign literal_10861[52] = 5'h0c;
  assign literal_10861[53] = 5'h0f;
  assign literal_10861[54] = 5'h10;
  assign literal_10861[55] = 5'h10;
  assign literal_10861[56] = 5'h10;
  assign literal_10861[57] = 5'h10;
  assign literal_10861[58] = 5'h10;
  assign literal_10861[59] = 5'h00;
  assign literal_10861[60] = 5'h00;
  assign literal_10861[61] = 5'h00;
  assign literal_10861[62] = 5'h00;
  assign literal_10861[63] = 5'h00;
  assign literal_10861[64] = 5'h00;
  assign literal_10861[65] = 5'h06;
  assign literal_10861[66] = 5'h0a;
  assign literal_10861[67] = 5'h0c;
  assign literal_10861[68] = 5'h0f;
  assign literal_10861[69] = 5'h10;
  assign literal_10861[70] = 5'h10;
  assign literal_10861[71] = 5'h10;
  assign literal_10861[72] = 5'h10;
  assign literal_10861[73] = 5'h10;
  assign literal_10861[74] = 5'h10;
  assign literal_10861[75] = 5'h00;
  assign literal_10861[76] = 5'h00;
  assign literal_10861[77] = 5'h00;
  assign literal_10861[78] = 5'h00;
  assign literal_10861[79] = 5'h00;
  assign literal_10861[80] = 5'h00;
  assign literal_10861[81] = 5'h07;
  assign literal_10861[82] = 5'h0b;
  assign literal_10861[83] = 5'h0d;
  assign literal_10861[84] = 5'h10;
  assign literal_10861[85] = 5'h10;
  assign literal_10861[86] = 5'h10;
  assign literal_10861[87] = 5'h10;
  assign literal_10861[88] = 5'h10;
  assign literal_10861[89] = 5'h10;
  assign literal_10861[90] = 5'h10;
  assign literal_10861[91] = 5'h00;
  assign literal_10861[92] = 5'h00;
  assign literal_10861[93] = 5'h00;
  assign literal_10861[94] = 5'h00;
  assign literal_10861[95] = 5'h00;
  assign literal_10861[96] = 5'h00;
  assign literal_10861[97] = 5'h07;
  assign literal_10861[98] = 5'h0b;
  assign literal_10861[99] = 5'h0d;
  assign literal_10861[100] = 5'h10;
  assign literal_10861[101] = 5'h10;
  assign literal_10861[102] = 5'h10;
  assign literal_10861[103] = 5'h10;
  assign literal_10861[104] = 5'h10;
  assign literal_10861[105] = 5'h10;
  assign literal_10861[106] = 5'h10;
  assign literal_10861[107] = 5'h00;
  assign literal_10861[108] = 5'h00;
  assign literal_10861[109] = 5'h00;
  assign literal_10861[110] = 5'h00;
  assign literal_10861[111] = 5'h00;
  assign literal_10861[112] = 5'h00;
  assign literal_10861[113] = 5'h08;
  assign literal_10861[114] = 5'h0b;
  assign literal_10861[115] = 5'h0e;
  assign literal_10861[116] = 5'h10;
  assign literal_10861[117] = 5'h10;
  assign literal_10861[118] = 5'h10;
  assign literal_10861[119] = 5'h10;
  assign literal_10861[120] = 5'h10;
  assign literal_10861[121] = 5'h10;
  assign literal_10861[122] = 5'h10;
  assign literal_10861[123] = 5'h00;
  assign literal_10861[124] = 5'h00;
  assign literal_10861[125] = 5'h00;
  assign literal_10861[126] = 5'h00;
  assign literal_10861[127] = 5'h00;
  assign literal_10861[128] = 5'h00;
  assign literal_10861[129] = 5'h08;
  assign literal_10861[130] = 5'h0c;
  assign literal_10861[131] = 5'h10;
  assign literal_10861[132] = 5'h10;
  assign literal_10861[133] = 5'h10;
  assign literal_10861[134] = 5'h10;
  assign literal_10861[135] = 5'h10;
  assign literal_10861[136] = 5'h10;
  assign literal_10861[137] = 5'h10;
  assign literal_10861[138] = 5'h10;
  assign literal_10861[139] = 5'h00;
  assign literal_10861[140] = 5'h00;
  assign literal_10861[141] = 5'h00;
  assign literal_10861[142] = 5'h00;
  assign literal_10861[143] = 5'h00;
  assign literal_10861[144] = 5'h00;
  assign literal_10861[145] = 5'h08;
  assign literal_10861[146] = 5'h0d;
  assign literal_10861[147] = 5'h10;
  assign literal_10861[148] = 5'h10;
  assign literal_10861[149] = 5'h10;
  assign literal_10861[150] = 5'h10;
  assign literal_10861[151] = 5'h10;
  assign literal_10861[152] = 5'h10;
  assign literal_10861[153] = 5'h10;
  assign literal_10861[154] = 5'h10;
  assign literal_10861[155] = 5'h00;
  assign literal_10861[156] = 5'h00;
  assign literal_10861[157] = 5'h00;
  assign literal_10861[158] = 5'h00;
  assign literal_10861[159] = 5'h00;
  assign literal_10861[160] = 5'h00;
  assign literal_10861[161] = 5'h09;
  assign literal_10861[162] = 5'h0d;
  assign literal_10861[163] = 5'h10;
  assign literal_10861[164] = 5'h10;
  assign literal_10861[165] = 5'h10;
  assign literal_10861[166] = 5'h10;
  assign literal_10861[167] = 5'h10;
  assign literal_10861[168] = 5'h10;
  assign literal_10861[169] = 5'h10;
  assign literal_10861[170] = 5'h10;
  assign literal_10861[171] = 5'h00;
  assign literal_10861[172] = 5'h00;
  assign literal_10861[173] = 5'h00;
  assign literal_10861[174] = 5'h00;
  assign literal_10861[175] = 5'h00;
  assign literal_10861[176] = 5'h00;
  assign literal_10861[177] = 5'h09;
  assign literal_10861[178] = 5'h0d;
  assign literal_10861[179] = 5'h10;
  assign literal_10861[180] = 5'h10;
  assign literal_10861[181] = 5'h10;
  assign literal_10861[182] = 5'h10;
  assign literal_10861[183] = 5'h10;
  assign literal_10861[184] = 5'h10;
  assign literal_10861[185] = 5'h10;
  assign literal_10861[186] = 5'h10;
  assign literal_10861[187] = 5'h00;
  assign literal_10861[188] = 5'h00;
  assign literal_10861[189] = 5'h00;
  assign literal_10861[190] = 5'h00;
  assign literal_10861[191] = 5'h00;
  assign literal_10861[192] = 5'h00;
  assign literal_10861[193] = 5'h0a;
  assign literal_10861[194] = 5'h0d;
  assign literal_10861[195] = 5'h10;
  assign literal_10861[196] = 5'h10;
  assign literal_10861[197] = 5'h10;
  assign literal_10861[198] = 5'h10;
  assign literal_10861[199] = 5'h10;
  assign literal_10861[200] = 5'h10;
  assign literal_10861[201] = 5'h10;
  assign literal_10861[202] = 5'h10;
  assign literal_10861[203] = 5'h00;
  assign literal_10861[204] = 5'h00;
  assign literal_10861[205] = 5'h00;
  assign literal_10861[206] = 5'h00;
  assign literal_10861[207] = 5'h00;
  assign literal_10861[208] = 5'h00;
  assign literal_10861[209] = 5'h0a;
  assign literal_10861[210] = 5'h0e;
  assign literal_10861[211] = 5'h10;
  assign literal_10861[212] = 5'h10;
  assign literal_10861[213] = 5'h10;
  assign literal_10861[214] = 5'h10;
  assign literal_10861[215] = 5'h10;
  assign literal_10861[216] = 5'h10;
  assign literal_10861[217] = 5'h10;
  assign literal_10861[218] = 5'h10;
  assign literal_10861[219] = 5'h00;
  assign literal_10861[220] = 5'h00;
  assign literal_10861[221] = 5'h00;
  assign literal_10861[222] = 5'h00;
  assign literal_10861[223] = 5'h00;
  assign literal_10861[224] = 5'h00;
  assign literal_10861[225] = 5'h0a;
  assign literal_10861[226] = 5'h0f;
  assign literal_10861[227] = 5'h10;
  assign literal_10861[228] = 5'h10;
  assign literal_10861[229] = 5'h10;
  assign literal_10861[230] = 5'h10;
  assign literal_10861[231] = 5'h10;
  assign literal_10861[232] = 5'h10;
  assign literal_10861[233] = 5'h10;
  assign literal_10861[234] = 5'h10;
  assign literal_10861[235] = 5'h00;
  assign literal_10861[236] = 5'h00;
  assign literal_10861[237] = 5'h00;
  assign literal_10861[238] = 5'h00;
  assign literal_10861[239] = 5'h00;
  assign literal_10861[240] = 5'h09;
  assign literal_10861[241] = 5'h0b;
  assign literal_10861[242] = 5'h10;
  assign literal_10861[243] = 5'h10;
  assign literal_10861[244] = 5'h10;
  assign literal_10861[245] = 5'h10;
  assign literal_10861[246] = 5'h10;
  assign literal_10861[247] = 5'h10;
  assign literal_10861[248] = 5'h10;
  assign literal_10861[249] = 5'h10;
  assign literal_10861[250] = 5'h10;
  assign literal_10861[251] = 5'h00;
  wire [4:0] literal_10863[0:251];
  assign literal_10863[0] = 5'h04;
  assign literal_10863[1] = 5'h02;
  assign literal_10863[2] = 5'h02;
  assign literal_10863[3] = 5'h03;
  assign literal_10863[4] = 5'h04;
  assign literal_10863[5] = 5'h05;
  assign literal_10863[6] = 5'h07;
  assign literal_10863[7] = 5'h09;
  assign literal_10863[8] = 5'h10;
  assign literal_10863[9] = 5'h10;
  assign literal_10863[10] = 5'h10;
  assign literal_10863[11] = 5'h00;
  assign literal_10863[12] = 5'h00;
  assign literal_10863[13] = 5'h00;
  assign literal_10863[14] = 5'h00;
  assign literal_10863[15] = 5'h00;
  assign literal_10863[16] = 5'h00;
  assign literal_10863[17] = 5'h04;
  assign literal_10863[18] = 5'h05;
  assign literal_10863[19] = 5'h07;
  assign literal_10863[20] = 5'h09;
  assign literal_10863[21] = 5'h0a;
  assign literal_10863[22] = 5'h0b;
  assign literal_10863[23] = 5'h10;
  assign literal_10863[24] = 5'h10;
  assign literal_10863[25] = 5'h10;
  assign literal_10863[26] = 5'h10;
  assign literal_10863[27] = 5'h00;
  assign literal_10863[28] = 5'h00;
  assign literal_10863[29] = 5'h00;
  assign literal_10863[30] = 5'h00;
  assign literal_10863[31] = 5'h00;
  assign literal_10863[32] = 5'h00;
  assign literal_10863[33] = 5'h05;
  assign literal_10863[34] = 5'h08;
  assign literal_10863[35] = 5'h0a;
  assign literal_10863[36] = 5'h0c;
  assign literal_10863[37] = 5'h0e;
  assign literal_10863[38] = 5'h10;
  assign literal_10863[39] = 5'h10;
  assign literal_10863[40] = 5'h10;
  assign literal_10863[41] = 5'h10;
  assign literal_10863[42] = 5'h10;
  assign literal_10863[43] = 5'h00;
  assign literal_10863[44] = 5'h00;
  assign literal_10863[45] = 5'h00;
  assign literal_10863[46] = 5'h00;
  assign literal_10863[47] = 5'h00;
  assign literal_10863[48] = 5'h00;
  assign literal_10863[49] = 5'h06;
  assign literal_10863[50] = 5'h09;
  assign literal_10863[51] = 5'h0b;
  assign literal_10863[52] = 5'h0e;
  assign literal_10863[53] = 5'h10;
  assign literal_10863[54] = 5'h10;
  assign literal_10863[55] = 5'h10;
  assign literal_10863[56] = 5'h10;
  assign literal_10863[57] = 5'h10;
  assign literal_10863[58] = 5'h10;
  assign literal_10863[59] = 5'h00;
  assign literal_10863[60] = 5'h00;
  assign literal_10863[61] = 5'h00;
  assign literal_10863[62] = 5'h00;
  assign literal_10863[63] = 5'h00;
  assign literal_10863[64] = 5'h00;
  assign literal_10863[65] = 5'h06;
  assign literal_10863[66] = 5'h0a;
  assign literal_10863[67] = 5'h0e;
  assign literal_10863[68] = 5'h10;
  assign literal_10863[69] = 5'h10;
  assign literal_10863[70] = 5'h10;
  assign literal_10863[71] = 5'h10;
  assign literal_10863[72] = 5'h10;
  assign literal_10863[73] = 5'h10;
  assign literal_10863[74] = 5'h10;
  assign literal_10863[75] = 5'h00;
  assign literal_10863[76] = 5'h00;
  assign literal_10863[77] = 5'h00;
  assign literal_10863[78] = 5'h00;
  assign literal_10863[79] = 5'h00;
  assign literal_10863[80] = 5'h00;
  assign literal_10863[81] = 5'h07;
  assign literal_10863[82] = 5'h0a;
  assign literal_10863[83] = 5'h0e;
  assign literal_10863[84] = 5'h10;
  assign literal_10863[85] = 5'h10;
  assign literal_10863[86] = 5'h10;
  assign literal_10863[87] = 5'h10;
  assign literal_10863[88] = 5'h10;
  assign literal_10863[89] = 5'h10;
  assign literal_10863[90] = 5'h10;
  assign literal_10863[91] = 5'h00;
  assign literal_10863[92] = 5'h00;
  assign literal_10863[93] = 5'h00;
  assign literal_10863[94] = 5'h00;
  assign literal_10863[95] = 5'h00;
  assign literal_10863[96] = 5'h00;
  assign literal_10863[97] = 5'h07;
  assign literal_10863[98] = 5'h0c;
  assign literal_10863[99] = 5'h0f;
  assign literal_10863[100] = 5'h10;
  assign literal_10863[101] = 5'h10;
  assign literal_10863[102] = 5'h10;
  assign literal_10863[103] = 5'h10;
  assign literal_10863[104] = 5'h10;
  assign literal_10863[105] = 5'h10;
  assign literal_10863[106] = 5'h10;
  assign literal_10863[107] = 5'h00;
  assign literal_10863[108] = 5'h00;
  assign literal_10863[109] = 5'h00;
  assign literal_10863[110] = 5'h00;
  assign literal_10863[111] = 5'h00;
  assign literal_10863[112] = 5'h00;
  assign literal_10863[113] = 5'h08;
  assign literal_10863[114] = 5'h0c;
  assign literal_10863[115] = 5'h10;
  assign literal_10863[116] = 5'h10;
  assign literal_10863[117] = 5'h10;
  assign literal_10863[118] = 5'h10;
  assign literal_10863[119] = 5'h10;
  assign literal_10863[120] = 5'h10;
  assign literal_10863[121] = 5'h10;
  assign literal_10863[122] = 5'h10;
  assign literal_10863[123] = 5'h00;
  assign literal_10863[124] = 5'h00;
  assign literal_10863[125] = 5'h00;
  assign literal_10863[126] = 5'h00;
  assign literal_10863[127] = 5'h00;
  assign literal_10863[128] = 5'h00;
  assign literal_10863[129] = 5'h09;
  assign literal_10863[130] = 5'h0d;
  assign literal_10863[131] = 5'h10;
  assign literal_10863[132] = 5'h10;
  assign literal_10863[133] = 5'h10;
  assign literal_10863[134] = 5'h10;
  assign literal_10863[135] = 5'h10;
  assign literal_10863[136] = 5'h10;
  assign literal_10863[137] = 5'h10;
  assign literal_10863[138] = 5'h10;
  assign literal_10863[139] = 5'h00;
  assign literal_10863[140] = 5'h00;
  assign literal_10863[141] = 5'h00;
  assign literal_10863[142] = 5'h00;
  assign literal_10863[143] = 5'h00;
  assign literal_10863[144] = 5'h00;
  assign literal_10863[145] = 5'h09;
  assign literal_10863[146] = 5'h0e;
  assign literal_10863[147] = 5'h10;
  assign literal_10863[148] = 5'h10;
  assign literal_10863[149] = 5'h10;
  assign literal_10863[150] = 5'h10;
  assign literal_10863[151] = 5'h10;
  assign literal_10863[152] = 5'h10;
  assign literal_10863[153] = 5'h10;
  assign literal_10863[154] = 5'h10;
  assign literal_10863[155] = 5'h00;
  assign literal_10863[156] = 5'h00;
  assign literal_10863[157] = 5'h00;
  assign literal_10863[158] = 5'h00;
  assign literal_10863[159] = 5'h00;
  assign literal_10863[160] = 5'h00;
  assign literal_10863[161] = 5'h09;
  assign literal_10863[162] = 5'h0e;
  assign literal_10863[163] = 5'h10;
  assign literal_10863[164] = 5'h10;
  assign literal_10863[165] = 5'h10;
  assign literal_10863[166] = 5'h10;
  assign literal_10863[167] = 5'h10;
  assign literal_10863[168] = 5'h10;
  assign literal_10863[169] = 5'h10;
  assign literal_10863[170] = 5'h10;
  assign literal_10863[171] = 5'h00;
  assign literal_10863[172] = 5'h00;
  assign literal_10863[173] = 5'h00;
  assign literal_10863[174] = 5'h00;
  assign literal_10863[175] = 5'h00;
  assign literal_10863[176] = 5'h00;
  assign literal_10863[177] = 5'h0a;
  assign literal_10863[178] = 5'h0f;
  assign literal_10863[179] = 5'h10;
  assign literal_10863[180] = 5'h10;
  assign literal_10863[181] = 5'h10;
  assign literal_10863[182] = 5'h10;
  assign literal_10863[183] = 5'h10;
  assign literal_10863[184] = 5'h10;
  assign literal_10863[185] = 5'h10;
  assign literal_10863[186] = 5'h10;
  assign literal_10863[187] = 5'h00;
  assign literal_10863[188] = 5'h00;
  assign literal_10863[189] = 5'h00;
  assign literal_10863[190] = 5'h00;
  assign literal_10863[191] = 5'h00;
  assign literal_10863[192] = 5'h00;
  assign literal_10863[193] = 5'h0a;
  assign literal_10863[194] = 5'h10;
  assign literal_10863[195] = 5'h10;
  assign literal_10863[196] = 5'h10;
  assign literal_10863[197] = 5'h10;
  assign literal_10863[198] = 5'h10;
  assign literal_10863[199] = 5'h10;
  assign literal_10863[200] = 5'h10;
  assign literal_10863[201] = 5'h10;
  assign literal_10863[202] = 5'h10;
  assign literal_10863[203] = 5'h00;
  assign literal_10863[204] = 5'h00;
  assign literal_10863[205] = 5'h00;
  assign literal_10863[206] = 5'h00;
  assign literal_10863[207] = 5'h00;
  assign literal_10863[208] = 5'h00;
  assign literal_10863[209] = 5'h0a;
  assign literal_10863[210] = 5'h10;
  assign literal_10863[211] = 5'h10;
  assign literal_10863[212] = 5'h10;
  assign literal_10863[213] = 5'h10;
  assign literal_10863[214] = 5'h10;
  assign literal_10863[215] = 5'h10;
  assign literal_10863[216] = 5'h10;
  assign literal_10863[217] = 5'h10;
  assign literal_10863[218] = 5'h10;
  assign literal_10863[219] = 5'h00;
  assign literal_10863[220] = 5'h00;
  assign literal_10863[221] = 5'h00;
  assign literal_10863[222] = 5'h00;
  assign literal_10863[223] = 5'h00;
  assign literal_10863[224] = 5'h00;
  assign literal_10863[225] = 5'h0b;
  assign literal_10863[226] = 5'h10;
  assign literal_10863[227] = 5'h10;
  assign literal_10863[228] = 5'h10;
  assign literal_10863[229] = 5'h10;
  assign literal_10863[230] = 5'h10;
  assign literal_10863[231] = 5'h10;
  assign literal_10863[232] = 5'h10;
  assign literal_10863[233] = 5'h10;
  assign literal_10863[234] = 5'h10;
  assign literal_10863[235] = 5'h00;
  assign literal_10863[236] = 5'h00;
  assign literal_10863[237] = 5'h00;
  assign literal_10863[238] = 5'h00;
  assign literal_10863[239] = 5'h00;
  assign literal_10863[240] = 5'h0c;
  assign literal_10863[241] = 5'h0d;
  assign literal_10863[242] = 5'h10;
  assign literal_10863[243] = 5'h10;
  assign literal_10863[244] = 5'h10;
  assign literal_10863[245] = 5'h10;
  assign literal_10863[246] = 5'h10;
  assign literal_10863[247] = 5'h10;
  assign literal_10863[248] = 5'h10;
  assign literal_10863[249] = 5'h10;
  assign literal_10863[250] = 5'h10;
  assign literal_10863[251] = 5'h00;
  wire [15:0] literal_10869[0:251];
  assign literal_10869[0] = 16'h0001;
  assign literal_10869[1] = 16'h0000;
  assign literal_10869[2] = 16'h0004;
  assign literal_10869[3] = 16'h000c;
  assign literal_10869[4] = 16'h001a;
  assign literal_10869[5] = 16'h0076;
  assign literal_10869[6] = 16'h00f6;
  assign literal_10869[7] = 16'h3fe0;
  assign literal_10869[8] = 16'hff96;
  assign literal_10869[9] = 16'hff97;
  assign literal_10869[10] = 16'hff98;
  assign literal_10869[11] = 16'h0000;
  assign literal_10869[12] = 16'h0000;
  assign literal_10869[13] = 16'h0000;
  assign literal_10869[14] = 16'h0000;
  assign literal_10869[15] = 16'h0000;
  assign literal_10869[16] = 16'h0000;
  assign literal_10869[17] = 16'h0005;
  assign literal_10869[18] = 16'h0038;
  assign literal_10869[19] = 16'h0078;
  assign literal_10869[20] = 16'h01f9;
  assign literal_10869[21] = 16'h07f2;
  assign literal_10869[22] = 16'h1fe8;
  assign literal_10869[23] = 16'hff93;
  assign literal_10869[24] = 16'hff99;
  assign literal_10869[25] = 16'hff9a;
  assign literal_10869[26] = 16'hff9e;
  assign literal_10869[27] = 16'h0000;
  assign literal_10869[28] = 16'h0000;
  assign literal_10869[29] = 16'h0000;
  assign literal_10869[30] = 16'h0000;
  assign literal_10869[31] = 16'h0000;
  assign literal_10869[32] = 16'h0000;
  assign literal_10869[33] = 16'h001b;
  assign literal_10869[34] = 16'h007a;
  assign literal_10869[35] = 16'h03f7;
  assign literal_10869[36] = 16'h0ff0;
  assign literal_10869[37] = 16'h1feb;
  assign literal_10869[38] = 16'hff9b;
  assign literal_10869[39] = 16'hff9f;
  assign literal_10869[40] = 16'hffa8;
  assign literal_10869[41] = 16'hffa9;
  assign literal_10869[42] = 16'hfff1;
  assign literal_10869[43] = 16'h0000;
  assign literal_10869[44] = 16'h0000;
  assign literal_10869[45] = 16'h0000;
  assign literal_10869[46] = 16'h0000;
  assign literal_10869[47] = 16'h0000;
  assign literal_10869[48] = 16'h0000;
  assign literal_10869[49] = 16'h0039;
  assign literal_10869[50] = 16'h00fa;
  assign literal_10869[51] = 16'h07f7;
  assign literal_10869[52] = 16'h0ff1;
  assign literal_10869[53] = 16'h7fc6;
  assign literal_10869[54] = 16'hff9c;
  assign literal_10869[55] = 16'hffa3;
  assign literal_10869[56] = 16'hffd7;
  assign literal_10869[57] = 16'hffe4;
  assign literal_10869[58] = 16'hfff2;
  assign literal_10869[59] = 16'h0000;
  assign literal_10869[60] = 16'h0000;
  assign literal_10869[61] = 16'h0000;
  assign literal_10869[62] = 16'h0000;
  assign literal_10869[63] = 16'h0000;
  assign literal_10869[64] = 16'h0000;
  assign literal_10869[65] = 16'h003a;
  assign literal_10869[66] = 16'h03f8;
  assign literal_10869[67] = 16'h0ff2;
  assign literal_10869[68] = 16'h7fc8;
  assign literal_10869[69] = 16'hff9d;
  assign literal_10869[70] = 16'hffbf;
  assign literal_10869[71] = 16'hffcb;
  assign literal_10869[72] = 16'hffd8;
  assign literal_10869[73] = 16'hffe5;
  assign literal_10869[74] = 16'hfff3;
  assign literal_10869[75] = 16'h0000;
  assign literal_10869[76] = 16'h0000;
  assign literal_10869[77] = 16'h0000;
  assign literal_10869[78] = 16'h0000;
  assign literal_10869[79] = 16'h0000;
  assign literal_10869[80] = 16'h0000;
  assign literal_10869[81] = 16'h0077;
  assign literal_10869[82] = 16'h07f3;
  assign literal_10869[83] = 16'h1fea;
  assign literal_10869[84] = 16'hff94;
  assign literal_10869[85] = 16'hffa2;
  assign literal_10869[86] = 16'hffc0;
  assign literal_10869[87] = 16'hffcc;
  assign literal_10869[88] = 16'hffd9;
  assign literal_10869[89] = 16'hffe6;
  assign literal_10869[90] = 16'hfff4;
  assign literal_10869[91] = 16'h0000;
  assign literal_10869[92] = 16'h0000;
  assign literal_10869[93] = 16'h0000;
  assign literal_10869[94] = 16'h0000;
  assign literal_10869[95] = 16'h0000;
  assign literal_10869[96] = 16'h0000;
  assign literal_10869[97] = 16'h0079;
  assign literal_10869[98] = 16'h07f4;
  assign literal_10869[99] = 16'h1fed;
  assign literal_10869[100] = 16'hffa0;
  assign literal_10869[101] = 16'hffb5;
  assign literal_10869[102] = 16'hffc1;
  assign literal_10869[103] = 16'hffcd;
  assign literal_10869[104] = 16'hffda;
  assign literal_10869[105] = 16'hffe7;
  assign literal_10869[106] = 16'hfff5;
  assign literal_10869[107] = 16'h0000;
  assign literal_10869[108] = 16'h0000;
  assign literal_10869[109] = 16'h0000;
  assign literal_10869[110] = 16'h0000;
  assign literal_10869[111] = 16'h0000;
  assign literal_10869[112] = 16'h0000;
  assign literal_10869[113] = 16'h00f7;
  assign literal_10869[114] = 16'h07f5;
  assign literal_10869[115] = 16'h3fe1;
  assign literal_10869[116] = 16'hffa1;
  assign literal_10869[117] = 16'hffb6;
  assign literal_10869[118] = 16'hffc2;
  assign literal_10869[119] = 16'hffce;
  assign literal_10869[120] = 16'hffdb;
  assign literal_10869[121] = 16'hffe8;
  assign literal_10869[122] = 16'hfff6;
  assign literal_10869[123] = 16'h0000;
  assign literal_10869[124] = 16'h0000;
  assign literal_10869[125] = 16'h0000;
  assign literal_10869[126] = 16'h0000;
  assign literal_10869[127] = 16'h0000;
  assign literal_10869[128] = 16'h0000;
  assign literal_10869[129] = 16'h00f8;
  assign literal_10869[130] = 16'h0ff3;
  assign literal_10869[131] = 16'hff92;
  assign literal_10869[132] = 16'hffad;
  assign literal_10869[133] = 16'hffb7;
  assign literal_10869[134] = 16'hffc3;
  assign literal_10869[135] = 16'hffcf;
  assign literal_10869[136] = 16'hffdc;
  assign literal_10869[137] = 16'hffe9;
  assign literal_10869[138] = 16'hfff7;
  assign literal_10869[139] = 16'h0000;
  assign literal_10869[140] = 16'h0000;
  assign literal_10869[141] = 16'h0000;
  assign literal_10869[142] = 16'h0000;
  assign literal_10869[143] = 16'h0000;
  assign literal_10869[144] = 16'h0000;
  assign literal_10869[145] = 16'h00f9;
  assign literal_10869[146] = 16'h1fe9;
  assign literal_10869[147] = 16'hff95;
  assign literal_10869[148] = 16'hffae;
  assign literal_10869[149] = 16'hffb8;
  assign literal_10869[150] = 16'hffc4;
  assign literal_10869[151] = 16'hffd0;
  assign literal_10869[152] = 16'hffdd;
  assign literal_10869[153] = 16'hffea;
  assign literal_10869[154] = 16'hfff8;
  assign literal_10869[155] = 16'h0000;
  assign literal_10869[156] = 16'h0000;
  assign literal_10869[157] = 16'h0000;
  assign literal_10869[158] = 16'h0000;
  assign literal_10869[159] = 16'h0000;
  assign literal_10869[160] = 16'h0000;
  assign literal_10869[161] = 16'h01f6;
  assign literal_10869[162] = 16'h1fec;
  assign literal_10869[163] = 16'hffa5;
  assign literal_10869[164] = 16'hffaf;
  assign literal_10869[165] = 16'hffb9;
  assign literal_10869[166] = 16'hffc5;
  assign literal_10869[167] = 16'hffd1;
  assign literal_10869[168] = 16'hffde;
  assign literal_10869[169] = 16'hffeb;
  assign literal_10869[170] = 16'hfff9;
  assign literal_10869[171] = 16'h0000;
  assign literal_10869[172] = 16'h0000;
  assign literal_10869[173] = 16'h0000;
  assign literal_10869[174] = 16'h0000;
  assign literal_10869[175] = 16'h0000;
  assign literal_10869[176] = 16'h0000;
  assign literal_10869[177] = 16'h01f7;
  assign literal_10869[178] = 16'h1fee;
  assign literal_10869[179] = 16'hffa6;
  assign literal_10869[180] = 16'hffb0;
  assign literal_10869[181] = 16'hffba;
  assign literal_10869[182] = 16'hffc6;
  assign literal_10869[183] = 16'hffd2;
  assign literal_10869[184] = 16'hffdf;
  assign literal_10869[185] = 16'hffec;
  assign literal_10869[186] = 16'hfffa;
  assign literal_10869[187] = 16'h0000;
  assign literal_10869[188] = 16'h0000;
  assign literal_10869[189] = 16'h0000;
  assign literal_10869[190] = 16'h0000;
  assign literal_10869[191] = 16'h0000;
  assign literal_10869[192] = 16'h0000;
  assign literal_10869[193] = 16'h03f4;
  assign literal_10869[194] = 16'h1fef;
  assign literal_10869[195] = 16'hffa7;
  assign literal_10869[196] = 16'hffb1;
  assign literal_10869[197] = 16'hffbb;
  assign literal_10869[198] = 16'hffc7;
  assign literal_10869[199] = 16'hffd3;
  assign literal_10869[200] = 16'hffe0;
  assign literal_10869[201] = 16'hffed;
  assign literal_10869[202] = 16'hfffb;
  assign literal_10869[203] = 16'h0000;
  assign literal_10869[204] = 16'h0000;
  assign literal_10869[205] = 16'h0000;
  assign literal_10869[206] = 16'h0000;
  assign literal_10869[207] = 16'h0000;
  assign literal_10869[208] = 16'h0000;
  assign literal_10869[209] = 16'h03f5;
  assign literal_10869[210] = 16'h3fe2;
  assign literal_10869[211] = 16'hffaa;
  assign literal_10869[212] = 16'hffb2;
  assign literal_10869[213] = 16'hffbc;
  assign literal_10869[214] = 16'hffc8;
  assign literal_10869[215] = 16'hffd4;
  assign literal_10869[216] = 16'hffe1;
  assign literal_10869[217] = 16'hffee;
  assign literal_10869[218] = 16'hfffc;
  assign literal_10869[219] = 16'h0000;
  assign literal_10869[220] = 16'h0000;
  assign literal_10869[221] = 16'h0000;
  assign literal_10869[222] = 16'h0000;
  assign literal_10869[223] = 16'h0000;
  assign literal_10869[224] = 16'h0000;
  assign literal_10869[225] = 16'h03f6;
  assign literal_10869[226] = 16'h7fc7;
  assign literal_10869[227] = 16'hffab;
  assign literal_10869[228] = 16'hffb3;
  assign literal_10869[229] = 16'hffbd;
  assign literal_10869[230] = 16'hffc9;
  assign literal_10869[231] = 16'hffd5;
  assign literal_10869[232] = 16'hffe2;
  assign literal_10869[233] = 16'hffef;
  assign literal_10869[234] = 16'hfffd;
  assign literal_10869[235] = 16'h0000;
  assign literal_10869[236] = 16'h0000;
  assign literal_10869[237] = 16'h0000;
  assign literal_10869[238] = 16'h0000;
  assign literal_10869[239] = 16'h0000;
  assign literal_10869[240] = 16'h01f8;
  assign literal_10869[241] = 16'h07f6;
  assign literal_10869[242] = 16'hffa4;
  assign literal_10869[243] = 16'hffac;
  assign literal_10869[244] = 16'hffb4;
  assign literal_10869[245] = 16'hffbe;
  assign literal_10869[246] = 16'hffca;
  assign literal_10869[247] = 16'hffd6;
  assign literal_10869[248] = 16'hffe3;
  assign literal_10869[249] = 16'hfff0;
  assign literal_10869[250] = 16'hfffe;
  assign literal_10869[251] = 16'h0000;
  wire [15:0] literal_10870[0:251];
  assign literal_10870[0] = 16'h000c;
  assign literal_10870[1] = 16'h0000;
  assign literal_10870[2] = 16'h0001;
  assign literal_10870[3] = 16'h0004;
  assign literal_10870[4] = 16'h000b;
  assign literal_10870[5] = 16'h001a;
  assign literal_10870[6] = 16'h0079;
  assign literal_10870[7] = 16'h01f9;
  assign literal_10870[8] = 16'hff9c;
  assign literal_10870[9] = 16'hff9f;
  assign literal_10870[10] = 16'hffa0;
  assign literal_10870[11] = 16'h0000;
  assign literal_10870[12] = 16'h0000;
  assign literal_10870[13] = 16'h0000;
  assign literal_10870[14] = 16'h0000;
  assign literal_10870[15] = 16'h0000;
  assign literal_10870[16] = 16'h0000;
  assign literal_10870[17] = 16'h000a;
  assign literal_10870[18] = 16'h001c;
  assign literal_10870[19] = 16'h007a;
  assign literal_10870[20] = 16'h01f5;
  assign literal_10870[21] = 16'h03f4;
  assign literal_10870[22] = 16'h07f8;
  assign literal_10870[23] = 16'hff95;
  assign literal_10870[24] = 16'hffa1;
  assign literal_10870[25] = 16'hffa2;
  assign literal_10870[26] = 16'hffad;
  assign literal_10870[27] = 16'h0000;
  assign literal_10870[28] = 16'h0000;
  assign literal_10870[29] = 16'h0000;
  assign literal_10870[30] = 16'h0000;
  assign literal_10870[31] = 16'h0000;
  assign literal_10870[32] = 16'h0000;
  assign literal_10870[33] = 16'h001b;
  assign literal_10870[34] = 16'h00f8;
  assign literal_10870[35] = 16'h03f7;
  assign literal_10870[36] = 16'h0ff4;
  assign literal_10870[37] = 16'h3fdc;
  assign literal_10870[38] = 16'hff9d;
  assign literal_10870[39] = 16'hff90;
  assign literal_10870[40] = 16'hffac;
  assign literal_10870[41] = 16'hffe3;
  assign literal_10870[42] = 16'hfff1;
  assign literal_10870[43] = 16'h0000;
  assign literal_10870[44] = 16'h0000;
  assign literal_10870[45] = 16'h0000;
  assign literal_10870[46] = 16'h0000;
  assign literal_10870[47] = 16'h0000;
  assign literal_10870[48] = 16'h0000;
  assign literal_10870[49] = 16'h003a;
  assign literal_10870[50] = 16'h01f6;
  assign literal_10870[51] = 16'h07f7;
  assign literal_10870[52] = 16'h3fde;
  assign literal_10870[53] = 16'hff8e;
  assign literal_10870[54] = 16'hff94;
  assign literal_10870[55] = 16'hffc9;
  assign literal_10870[56] = 16'hffd6;
  assign literal_10870[57] = 16'hffe4;
  assign literal_10870[58] = 16'hfff2;
  assign literal_10870[59] = 16'h0000;
  assign literal_10870[60] = 16'h0000;
  assign literal_10870[61] = 16'h0000;
  assign literal_10870[62] = 16'h0000;
  assign literal_10870[63] = 16'h0000;
  assign literal_10870[64] = 16'h0000;
  assign literal_10870[65] = 16'h003b;
  assign literal_10870[66] = 16'h03f6;
  assign literal_10870[67] = 16'h3fdd;
  assign literal_10870[68] = 16'hff8f;
  assign literal_10870[69] = 16'hffa5;
  assign literal_10870[70] = 16'hffa6;
  assign literal_10870[71] = 16'hffca;
  assign literal_10870[72] = 16'hffd7;
  assign literal_10870[73] = 16'hffe5;
  assign literal_10870[74] = 16'hfff3;
  assign literal_10870[75] = 16'h0000;
  assign literal_10870[76] = 16'h0000;
  assign literal_10870[77] = 16'h0000;
  assign literal_10870[78] = 16'h0000;
  assign literal_10870[79] = 16'h0000;
  assign literal_10870[80] = 16'h0000;
  assign literal_10870[81] = 16'h0078;
  assign literal_10870[82] = 16'h03f9;
  assign literal_10870[83] = 16'h3fdf;
  assign literal_10870[84] = 16'hff96;
  assign literal_10870[85] = 16'hffab;
  assign literal_10870[86] = 16'hffa9;
  assign literal_10870[87] = 16'hffcb;
  assign literal_10870[88] = 16'hffd8;
  assign literal_10870[89] = 16'hffe6;
  assign literal_10870[90] = 16'hfff4;
  assign literal_10870[91] = 16'h0000;
  assign literal_10870[92] = 16'h0000;
  assign literal_10870[93] = 16'h0000;
  assign literal_10870[94] = 16'h0000;
  assign literal_10870[95] = 16'h0000;
  assign literal_10870[96] = 16'h0000;
  assign literal_10870[97] = 16'h007b;
  assign literal_10870[98] = 16'h0ff2;
  assign literal_10870[99] = 16'h7fc5;
  assign literal_10870[100] = 16'hff97;
  assign literal_10870[101] = 16'hffb5;
  assign literal_10870[102] = 16'hffbf;
  assign literal_10870[103] = 16'hffcc;
  assign literal_10870[104] = 16'hffd9;
  assign literal_10870[105] = 16'hffe7;
  assign literal_10870[106] = 16'hfff5;
  assign literal_10870[107] = 16'h0000;
  assign literal_10870[108] = 16'h0000;
  assign literal_10870[109] = 16'h0000;
  assign literal_10870[110] = 16'h0000;
  assign literal_10870[111] = 16'h0000;
  assign literal_10870[112] = 16'h0000;
  assign literal_10870[113] = 16'h00f9;
  assign literal_10870[114] = 16'h0ff5;
  assign literal_10870[115] = 16'hff8c;
  assign literal_10870[116] = 16'hff98;
  assign literal_10870[117] = 16'hffb6;
  assign literal_10870[118] = 16'hffc0;
  assign literal_10870[119] = 16'hffcd;
  assign literal_10870[120] = 16'hffda;
  assign literal_10870[121] = 16'hffe8;
  assign literal_10870[122] = 16'hfff6;
  assign literal_10870[123] = 16'h0000;
  assign literal_10870[124] = 16'h0000;
  assign literal_10870[125] = 16'h0000;
  assign literal_10870[126] = 16'h0000;
  assign literal_10870[127] = 16'h0000;
  assign literal_10870[128] = 16'h0000;
  assign literal_10870[129] = 16'h01f4;
  assign literal_10870[130] = 16'h1fec;
  assign literal_10870[131] = 16'hff9e;
  assign literal_10870[132] = 16'hffa3;
  assign literal_10870[133] = 16'hffb7;
  assign literal_10870[134] = 16'hffc1;
  assign literal_10870[135] = 16'hffce;
  assign literal_10870[136] = 16'hffdb;
  assign literal_10870[137] = 16'hffe9;
  assign literal_10870[138] = 16'hfff7;
  assign literal_10870[139] = 16'h0000;
  assign literal_10870[140] = 16'h0000;
  assign literal_10870[141] = 16'h0000;
  assign literal_10870[142] = 16'h0000;
  assign literal_10870[143] = 16'h0000;
  assign literal_10870[144] = 16'h0000;
  assign literal_10870[145] = 16'h01f7;
  assign literal_10870[146] = 16'h3fe0;
  assign literal_10870[147] = 16'hff91;
  assign literal_10870[148] = 16'hffa4;
  assign literal_10870[149] = 16'hffb8;
  assign literal_10870[150] = 16'hffc2;
  assign literal_10870[151] = 16'hffcf;
  assign literal_10870[152] = 16'hffdc;
  assign literal_10870[153] = 16'hffea;
  assign literal_10870[154] = 16'hfff8;
  assign literal_10870[155] = 16'h0000;
  assign literal_10870[156] = 16'h0000;
  assign literal_10870[157] = 16'h0000;
  assign literal_10870[158] = 16'h0000;
  assign literal_10870[159] = 16'h0000;
  assign literal_10870[160] = 16'h0000;
  assign literal_10870[161] = 16'h01f8;
  assign literal_10870[162] = 16'h3fe1;
  assign literal_10870[163] = 16'hff92;
  assign literal_10870[164] = 16'hffa7;
  assign literal_10870[165] = 16'hffb9;
  assign literal_10870[166] = 16'hffc3;
  assign literal_10870[167] = 16'hffd0;
  assign literal_10870[168] = 16'hffdd;
  assign literal_10870[169] = 16'hffeb;
  assign literal_10870[170] = 16'hfff9;
  assign literal_10870[171] = 16'h0000;
  assign literal_10870[172] = 16'h0000;
  assign literal_10870[173] = 16'h0000;
  assign literal_10870[174] = 16'h0000;
  assign literal_10870[175] = 16'h0000;
  assign literal_10870[176] = 16'h0000;
  assign literal_10870[177] = 16'h03f5;
  assign literal_10870[178] = 16'h7fc4;
  assign literal_10870[179] = 16'hff93;
  assign literal_10870[180] = 16'hffa8;
  assign literal_10870[181] = 16'hffba;
  assign literal_10870[182] = 16'hffc4;
  assign literal_10870[183] = 16'hffd1;
  assign literal_10870[184] = 16'hffde;
  assign literal_10870[185] = 16'hffec;
  assign literal_10870[186] = 16'hfffa;
  assign literal_10870[187] = 16'h0000;
  assign literal_10870[188] = 16'h0000;
  assign literal_10870[189] = 16'h0000;
  assign literal_10870[190] = 16'h0000;
  assign literal_10870[191] = 16'h0000;
  assign literal_10870[192] = 16'h0000;
  assign literal_10870[193] = 16'h03f8;
  assign literal_10870[194] = 16'hff8d;
  assign literal_10870[195] = 16'hff99;
  assign literal_10870[196] = 16'hffb1;
  assign literal_10870[197] = 16'hffbb;
  assign literal_10870[198] = 16'hffc5;
  assign literal_10870[199] = 16'hffd2;
  assign literal_10870[200] = 16'hffdf;
  assign literal_10870[201] = 16'hffed;
  assign literal_10870[202] = 16'hfffb;
  assign literal_10870[203] = 16'h0000;
  assign literal_10870[204] = 16'h0000;
  assign literal_10870[205] = 16'h0000;
  assign literal_10870[206] = 16'h0000;
  assign literal_10870[207] = 16'h0000;
  assign literal_10870[208] = 16'h0000;
  assign literal_10870[209] = 16'h03fa;
  assign literal_10870[210] = 16'hff9a;
  assign literal_10870[211] = 16'hffaa;
  assign literal_10870[212] = 16'hffb2;
  assign literal_10870[213] = 16'hffbc;
  assign literal_10870[214] = 16'hffc6;
  assign literal_10870[215] = 16'hffd3;
  assign literal_10870[216] = 16'hffe0;
  assign literal_10870[217] = 16'hffee;
  assign literal_10870[218] = 16'hfffc;
  assign literal_10870[219] = 16'h0000;
  assign literal_10870[220] = 16'h0000;
  assign literal_10870[221] = 16'h0000;
  assign literal_10870[222] = 16'h0000;
  assign literal_10870[223] = 16'h0000;
  assign literal_10870[224] = 16'h0000;
  assign literal_10870[225] = 16'h07f6;
  assign literal_10870[226] = 16'hff9b;
  assign literal_10870[227] = 16'hffaf;
  assign literal_10870[228] = 16'hffb3;
  assign literal_10870[229] = 16'hffbd;
  assign literal_10870[230] = 16'hffc7;
  assign literal_10870[231] = 16'hffd4;
  assign literal_10870[232] = 16'hffe1;
  assign literal_10870[233] = 16'hffef;
  assign literal_10870[234] = 16'hfffd;
  assign literal_10870[235] = 16'h0000;
  assign literal_10870[236] = 16'h0000;
  assign literal_10870[237] = 16'h0000;
  assign literal_10870[238] = 16'h0000;
  assign literal_10870[239] = 16'h0000;
  assign literal_10870[240] = 16'h0ff3;
  assign literal_10870[241] = 16'h1fed;
  assign literal_10870[242] = 16'hffae;
  assign literal_10870[243] = 16'hffb0;
  assign literal_10870[244] = 16'hffb4;
  assign literal_10870[245] = 16'hffbe;
  assign literal_10870[246] = 16'hffc8;
  assign literal_10870[247] = 16'hffd5;
  assign literal_10870[248] = 16'hffe2;
  assign literal_10870[249] = 16'hfff0;
  assign literal_10870[250] = 16'hfffe;
  assign literal_10870[251] = 16'h0000;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [4:0] p1_concat_9933_comb;
  wire [7:0] p1_concat_9940_comb;
  wire [6:0] p1_concat_10141_comb;
  wire [5:0] p1_concat_10203_comb;
  wire [7:0] p1_flipped__2_comb;
  wire [4:0] p1_add_9938_comb;
  wire [8:0] p1_concat_9942_comb;
  wire [7:0] p1_add_10073_comb;
  wire [6:0] p1_add_10152_comb;
  wire [7:0] p1_add_10185_comb;
  wire [5:0] p1_add_10226_comb;
  wire [7:0] p1_add_10267_comb;
  wire [6:0] p1_add_10307_comb;
  wire [7:0] p1_add_10347_comb;
  wire [8:0] p1_concat_9944_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed_comb;
  wire [2:0] p1_huff_length_squeezed_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__1_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__2_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__3_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__4_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__5_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__6_comb;
  wire [2:0] p1_huff_length_squeezed__1_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__7_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__8_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__9_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__10_comb;
  wire [2:0] p1_huff_length_squeezed__3_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__11_comb;
  wire [2:0] p1_huff_length_squeezed__4_comb;
  wire [2:0] p1_huff_length_squeezed__5_comb;
  wire [2:0] p1_huff_length_squeezed__6_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__12_comb;
  wire [2:0] p1_huff_length_squeezed__7_comb;
  wire [2:0] p1_huff_length_squeezed__8_comb;
  wire [2:0] p1_huff_length_squeezed__9_comb;
  wire [2:0] p1_huff_length_squeezed__10_comb;
  wire [2:0] p1_huff_length_squeezed__11_comb;
  wire [2:0] p1_huff_length_squeezed__12_comb;
  wire [2:0] p1_huff_length_squeezed__13_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__13_comb;
  wire [2:0] p1_huff_length_squeezed__14_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__14_comb;
  wire [2:0] p1_huff_length_squeezed__15_comb;
  wire [2:0] p1_huff_code__1_squeezed_squeezed__15_comb;
  wire [2:0] p1_huff_length_squeezed__16_comb;
  wire [8:0] p1_add_10075_comb;
  wire [8:0] p1_concat_10144_comb;
  wire [4:0] p1_add_10151_comb;
  wire [8:0] p1_add_10154_comb;
  wire [8:0] p1_add_10163_comb;
  wire [8:0] p1_concat_10167_comb;
  wire [7:0] p1_add_10177_comb;
  wire [8:0] p1_add_10186_comb;
  wire [8:0] p1_add_10196_comb;
  wire [8:0] p1_concat_10206_comb;
  wire [6:0] p1_add_10217_comb;
  wire [8:0] p1_add_10228_comb;
  wire [8:0] p1_add_10238_comb;
  wire [8:0] p1_concat_10248_comb;
  wire [7:0] p1_add_10258_comb;
  wire [8:0] p1_add_10268_comb;
  wire [8:0] p1_add_10278_comb;
  wire [8:0] p1_concat_10288_comb;
  wire [5:0] p1_add_10298_comb;
  wire [8:0] p1_add_10308_comb;
  wire [8:0] p1_add_10318_comb;
  wire [8:0] p1_concat_10328_comb;
  wire [7:0] p1_add_10338_comb;
  wire [8:0] p1_add_10348_comb;
  wire [8:0] p1_add_10359_comb;
  wire [8:0] p1_concat_10367_comb;
  wire [8:0] p1_add_10375_comb;
  wire [6:0] p1_add_10378_comb;
  wire [8:0] p1_add_10397_comb;
  wire [7:0] p1_add_10415_comb;
  wire [8:0] p1_add_10438_comb;
  wire [9:0] p1_array_index_10077_comb;
  wire [9:0] p1_array_index_10078_comb;
  wire [9:0] p1_array_index_10079_comb;
  wire [9:0] p1_array_index_10080_comb;
  wire [9:0] p1_array_index_10081_comb;
  wire [9:0] p1_array_index_10082_comb;
  wire [9:0] p1_array_index_10083_comb;
  wire [9:0] p1_array_index_10084_comb;
  wire [9:0] p1_array_index_10085_comb;
  wire [9:0] p1_array_index_10086_comb;
  wire [9:0] p1_array_index_10087_comb;
  wire [9:0] p1_array_index_10088_comb;
  wire [9:0] p1_array_index_10089_comb;
  wire [9:0] p1_array_index_10090_comb;
  wire [9:0] p1_array_index_10091_comb;
  wire [9:0] p1_array_index_10092_comb;
  wire [9:0] p1_array_index_10093_comb;
  wire [9:0] p1_array_index_10094_comb;
  wire [9:0] p1_array_index_10095_comb;
  wire [9:0] p1_array_index_10096_comb;
  wire [9:0] p1_array_index_10097_comb;
  wire [9:0] p1_array_index_10098_comb;
  wire [9:0] p1_array_index_10099_comb;
  wire [9:0] p1_array_index_10100_comb;
  wire [9:0] p1_array_index_10101_comb;
  wire [9:0] p1_array_index_10102_comb;
  wire [9:0] p1_array_index_10103_comb;
  wire [9:0] p1_array_index_10104_comb;
  wire [9:0] p1_array_index_10105_comb;
  wire [9:0] p1_array_index_10106_comb;
  wire [9:0] p1_array_index_10107_comb;
  wire [9:0] p1_array_index_10108_comb;
  wire [9:0] p1_array_index_10109_comb;
  wire [9:0] p1_array_index_10110_comb;
  wire [9:0] p1_array_index_10111_comb;
  wire [9:0] p1_array_index_10112_comb;
  wire [9:0] p1_array_index_10113_comb;
  wire [9:0] p1_array_index_10114_comb;
  wire [9:0] p1_array_index_10115_comb;
  wire [9:0] p1_array_index_10116_comb;
  wire [9:0] p1_array_index_10117_comb;
  wire [9:0] p1_array_index_10118_comb;
  wire [9:0] p1_array_index_10119_comb;
  wire [9:0] p1_array_index_10120_comb;
  wire [9:0] p1_array_index_10121_comb;
  wire [9:0] p1_array_index_10122_comb;
  wire [9:0] p1_array_index_10123_comb;
  wire [9:0] p1_array_index_10124_comb;
  wire [9:0] p1_array_index_10125_comb;
  wire [9:0] p1_array_index_10126_comb;
  wire [9:0] p1_array_index_10127_comb;
  wire [9:0] p1_array_index_10128_comb;
  wire [9:0] p1_array_index_10129_comb;
  wire [9:0] p1_array_index_10130_comb;
  wire [9:0] p1_array_index_10131_comb;
  wire [9:0] p1_array_index_10132_comb;
  wire [9:0] p1_array_index_10133_comb;
  wire [9:0] p1_array_index_10134_comb;
  wire [9:0] p1_array_index_10135_comb;
  wire [9:0] p1_array_index_10136_comb;
  wire [9:0] p1_array_index_10137_comb;
  wire [9:0] p1_array_index_10138_comb;
  wire [9:0] p1_array_index_10139_comb;
  wire [7:0] p1_huff_length_comb;
  wire [7:0] p1_huff_length__1_comb;
  wire p1_or_10174_comb;
  wire p1_or_10193_comb;
  wire p1_or_10213_comb;
  wire [9:0] p1_value__1_comb;
  wire p1_or_10225_comb;
  wire p1_or_10235_comb;
  wire p1_or_10245_comb;
  wire p1_or_10255_comb;
  wire p1_or_10266_comb;
  wire p1_or_10275_comb;
  wire p1_or_10285_comb;
  wire p1_or_10295_comb;
  wire p1_or_10306_comb;
  wire p1_or_10315_comb;
  wire p1_or_10325_comb;
  wire p1_or_10335_comb;
  wire p1_or_10346_comb;
  wire p1_or_10355_comb;
  wire p1_or_10366_comb;
  wire p1_or_10374_comb;
  wire p1_or_10386_comb;
  wire p1_or_10393_comb;
  wire p1_or_10404_comb;
  wire p1_or_10410_comb;
  wire p1_or_10423_comb;
  wire p1_or_10427_comb;
  wire p1_or_10436_comb;
  wire p1_or_10439_comb;
  wire p1_nor_10440_comb;
  wire p1_or_10447_comb;
  wire p1_or_10451_comb;
  wire p1_or_10455_comb;
  wire p1_nor_10458_comb;
  wire p1_and_10585_comb;
  assign p1_concat_9933_comb = {1'h0, p0_start_pix[7:4]};
  assign p1_concat_9940_comb = {1'h0, p0_start_pix[7:1]};
  assign p1_concat_10141_comb = {1'h0, p0_start_pix[7:2]};
  assign p1_concat_10203_comb = {1'h0, p0_start_pix[7:3]};
  assign p1_flipped__2_comb = 8'hff;
  assign p1_add_9938_comb = p1_concat_9933_comb + 5'h1f;
  assign p1_concat_9942_comb = {1'h0, p0_start_pix};
  assign p1_add_10073_comb = p1_concat_9940_comb + 8'hf9;
  assign p1_add_10152_comb = p1_concat_10141_comb + 7'h7d;
  assign p1_add_10185_comb = p1_concat_9940_comb + 8'hfb;
  assign p1_add_10226_comb = p1_concat_10203_comb + 6'h3f;
  assign p1_add_10267_comb = p1_concat_9940_comb + 8'hfd;
  assign p1_add_10307_comb = p1_concat_10141_comb + 7'h7f;
  assign p1_add_10347_comb = p1_concat_9940_comb + p1_flipped__2_comb;
  assign p1_concat_9944_comb = {p1_add_9938_comb, p0_start_pix[3:0]};
  assign p1_huff_code__1_squeezed_squeezed_comb = 3'h1;
  assign p1_huff_length_squeezed_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__1_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__2_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__3_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__4_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__5_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__6_comb = 3'h1;
  assign p1_huff_length_squeezed__1_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__7_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__8_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__9_comb = 3'h1;
  assign p1_huff_code__1_squeezed_squeezed__10_comb = 3'h1;
  assign p1_huff_length_squeezed__3_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__11_comb = 3'h1;
  assign p1_huff_length_squeezed__4_comb = 3'h4;
  assign p1_huff_length_squeezed__5_comb = 3'h4;
  assign p1_huff_length_squeezed__6_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__12_comb = 3'h1;
  assign p1_huff_length_squeezed__7_comb = 3'h4;
  assign p1_huff_length_squeezed__8_comb = 3'h4;
  assign p1_huff_length_squeezed__9_comb = 3'h4;
  assign p1_huff_length_squeezed__10_comb = 3'h4;
  assign p1_huff_length_squeezed__11_comb = 3'h4;
  assign p1_huff_length_squeezed__12_comb = 3'h4;
  assign p1_huff_length_squeezed__13_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__13_comb = 3'h1;
  assign p1_huff_length_squeezed__14_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__14_comb = 3'h1;
  assign p1_huff_length_squeezed__15_comb = 3'h4;
  assign p1_huff_code__1_squeezed_squeezed__15_comb = 3'h1;
  assign p1_huff_length_squeezed__16_comb = 3'h4;
  assign p1_add_10075_comb = p1_concat_9942_comb + 9'h1f1;
  assign p1_concat_10144_comb = {p1_add_10073_comb, p0_start_pix[0]};
  assign p1_add_10151_comb = p1_concat_9933_comb + 5'h01;
  assign p1_add_10154_comb = p1_concat_9942_comb + 9'h1f3;
  assign p1_add_10163_comb = p1_concat_9942_comb + 9'h00f;
  assign p1_concat_10167_comb = {p1_add_10152_comb, p0_start_pix[1:0]};
  assign p1_add_10177_comb = p1_concat_9940_comb + 8'h07;
  assign p1_add_10186_comb = p1_concat_9942_comb + 9'h1f5;
  assign p1_add_10196_comb = p1_concat_9942_comb + 9'h00d;
  assign p1_concat_10206_comb = {p1_add_10185_comb, p0_start_pix[0]};
  assign p1_add_10217_comb = p1_concat_10141_comb + 7'h03;
  assign p1_add_10228_comb = p1_concat_9942_comb + 9'h1f7;
  assign p1_add_10238_comb = p1_concat_9942_comb + 9'h00b;
  assign p1_concat_10248_comb = {p1_add_10226_comb, p0_start_pix[2:0]};
  assign p1_add_10258_comb = p1_concat_9940_comb + 8'h05;
  assign p1_add_10268_comb = p1_concat_9942_comb + 9'h1f9;
  assign p1_add_10278_comb = p1_concat_9942_comb + 9'h009;
  assign p1_concat_10288_comb = {p1_add_10267_comb, p0_start_pix[0]};
  assign p1_add_10298_comb = p1_concat_10203_comb + 6'h01;
  assign p1_add_10308_comb = p1_concat_9942_comb + 9'h1fb;
  assign p1_add_10318_comb = p1_concat_9942_comb + 9'h007;
  assign p1_concat_10328_comb = {p1_add_10307_comb, p0_start_pix[1:0]};
  assign p1_add_10338_comb = p1_concat_9940_comb + 8'h03;
  assign p1_add_10348_comb = p1_concat_9942_comb + 9'h1fd;
  assign p1_add_10359_comb = p1_concat_9942_comb + 9'h005;
  assign p1_concat_10367_comb = {p1_add_10347_comb, p0_start_pix[0]};
  assign p1_add_10375_comb = p1_concat_9942_comb + 9'h1ff;
  assign p1_add_10378_comb = p1_concat_10141_comb + 7'h01;
  assign p1_add_10397_comb = p1_concat_9942_comb + 9'h003;
  assign p1_add_10415_comb = p1_concat_9940_comb + 8'h01;
  assign p1_add_10438_comb = p1_concat_9942_comb + 9'h001;
  assign p1_array_index_10077_comb = p0_matrix[3'h0][3'h0];
  assign p1_array_index_10078_comb = p0_matrix[3'h0][p1_huff_code__1_squeezed_squeezed_comb];
  assign p1_array_index_10079_comb = p0_matrix[3'h0][3'h2];
  assign p1_array_index_10080_comb = p0_matrix[3'h0][3'h3];
  assign p1_array_index_10081_comb = p0_matrix[3'h0][p1_huff_length_squeezed_comb];
  assign p1_array_index_10082_comb = p0_matrix[3'h0][3'h5];
  assign p1_array_index_10083_comb = p0_matrix[3'h0][3'h6];
  assign p1_array_index_10084_comb = p0_matrix[3'h0][3'h7];
  assign p1_array_index_10085_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__1_comb][3'h0];
  assign p1_array_index_10086_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__2_comb][p1_huff_code__1_squeezed_squeezed__3_comb];
  assign p1_array_index_10087_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__4_comb][3'h2];
  assign p1_array_index_10088_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__5_comb][3'h3];
  assign p1_array_index_10089_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__6_comb][p1_huff_length_squeezed__1_comb];
  assign p1_array_index_10090_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__7_comb][3'h5];
  assign p1_array_index_10091_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__8_comb][3'h6];
  assign p1_array_index_10092_comb = p0_matrix[p1_huff_code__1_squeezed_squeezed__9_comb][3'h7];
  assign p1_array_index_10093_comb = p0_matrix[3'h2][3'h0];
  assign p1_array_index_10094_comb = p0_matrix[3'h2][p1_huff_code__1_squeezed_squeezed__10_comb];
  assign p1_array_index_10095_comb = p0_matrix[3'h2][3'h2];
  assign p1_array_index_10096_comb = p0_matrix[3'h2][3'h3];
  assign p1_array_index_10097_comb = p0_matrix[3'h2][p1_huff_length_squeezed__3_comb];
  assign p1_array_index_10098_comb = p0_matrix[3'h2][3'h5];
  assign p1_array_index_10099_comb = p0_matrix[3'h2][3'h6];
  assign p1_array_index_10100_comb = p0_matrix[3'h2][3'h7];
  assign p1_array_index_10101_comb = p0_matrix[3'h3][3'h0];
  assign p1_array_index_10102_comb = p0_matrix[3'h3][p1_huff_code__1_squeezed_squeezed__11_comb];
  assign p1_array_index_10103_comb = p0_matrix[3'h3][3'h2];
  assign p1_array_index_10104_comb = p0_matrix[3'h3][3'h3];
  assign p1_array_index_10105_comb = p0_matrix[3'h3][p1_huff_length_squeezed__4_comb];
  assign p1_array_index_10106_comb = p0_matrix[3'h3][3'h5];
  assign p1_array_index_10107_comb = p0_matrix[3'h3][3'h6];
  assign p1_array_index_10108_comb = p0_matrix[3'h3][3'h7];
  assign p1_array_index_10109_comb = p0_matrix[p1_huff_length_squeezed__5_comb][3'h0];
  assign p1_array_index_10110_comb = p0_matrix[p1_huff_length_squeezed__6_comb][p1_huff_code__1_squeezed_squeezed__12_comb];
  assign p1_array_index_10111_comb = p0_matrix[p1_huff_length_squeezed__7_comb][3'h2];
  assign p1_array_index_10112_comb = p0_matrix[p1_huff_length_squeezed__8_comb][3'h3];
  assign p1_array_index_10113_comb = p0_matrix[p1_huff_length_squeezed__9_comb][p1_huff_length_squeezed__10_comb];
  assign p1_array_index_10114_comb = p0_matrix[p1_huff_length_squeezed__11_comb][3'h5];
  assign p1_array_index_10115_comb = p0_matrix[p1_huff_length_squeezed__12_comb][3'h6];
  assign p1_array_index_10116_comb = p0_matrix[p1_huff_length_squeezed__13_comb][3'h7];
  assign p1_array_index_10117_comb = p0_matrix[3'h5][3'h0];
  assign p1_array_index_10118_comb = p0_matrix[3'h5][p1_huff_code__1_squeezed_squeezed__13_comb];
  assign p1_array_index_10119_comb = p0_matrix[3'h5][3'h2];
  assign p1_array_index_10120_comb = p0_matrix[3'h5][3'h3];
  assign p1_array_index_10121_comb = p0_matrix[3'h5][p1_huff_length_squeezed__14_comb];
  assign p1_array_index_10122_comb = p0_matrix[3'h5][3'h5];
  assign p1_array_index_10123_comb = p0_matrix[3'h5][3'h6];
  assign p1_array_index_10124_comb = p0_matrix[3'h5][3'h7];
  assign p1_array_index_10125_comb = p0_matrix[3'h6][3'h0];
  assign p1_array_index_10126_comb = p0_matrix[3'h6][p1_huff_code__1_squeezed_squeezed__14_comb];
  assign p1_array_index_10127_comb = p0_matrix[3'h6][3'h2];
  assign p1_array_index_10128_comb = p0_matrix[3'h6][3'h3];
  assign p1_array_index_10129_comb = p0_matrix[3'h6][p1_huff_length_squeezed__15_comb];
  assign p1_array_index_10130_comb = p0_matrix[3'h6][3'h5];
  assign p1_array_index_10131_comb = p0_matrix[3'h6][3'h6];
  assign p1_array_index_10132_comb = p0_matrix[3'h6][3'h7];
  assign p1_array_index_10133_comb = p0_matrix[3'h7][3'h0];
  assign p1_array_index_10134_comb = p0_matrix[3'h7][p1_huff_code__1_squeezed_squeezed__15_comb];
  assign p1_array_index_10135_comb = p0_matrix[3'h7][3'h2];
  assign p1_array_index_10136_comb = p0_matrix[3'h7][3'h3];
  assign p1_array_index_10137_comb = p0_matrix[3'h7][p1_huff_length_squeezed__16_comb];
  assign p1_array_index_10138_comb = p0_matrix[3'h7][3'h5];
  assign p1_array_index_10139_comb = p0_matrix[3'h7][3'h6];
  assign p1_huff_length_comb = 8'h04;
  assign p1_huff_length__1_comb = 8'h02;
  assign p1_or_10174_comb = p0_start_pix == 8'h0f | ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_concat_9944_comb[8]}}, p1_concat_9944_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10193_comb = p0_start_pix == 8'h0e | ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_add_10075_comb[8]}}, p1_add_10075_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10213_comb = p0_start_pix == 8'h0d | ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_concat_10144_comb[8]}}, p1_concat_10144_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_value__1_comb = p0_start_pix == 8'h00 ? p1_array_index_10077_comb : (p0_start_pix == 8'h01 ? p1_array_index_10078_comb : (p0_start_pix == 8'h02 ? p1_array_index_10079_comb : (p0_start_pix == 8'h03 ? p1_array_index_10080_comb : (p0_start_pix == 8'h04 ? p1_array_index_10081_comb : (p0_start_pix == 8'h05 ? p1_array_index_10082_comb : (p0_start_pix == 8'h06 ? p1_array_index_10083_comb : (p0_start_pix == 8'h07 ? p1_array_index_10084_comb : (p0_start_pix == 8'h08 ? p1_array_index_10085_comb : (p0_start_pix == 8'h09 ? p1_array_index_10086_comb : (p0_start_pix == 8'h0a ? p1_array_index_10087_comb : (p0_start_pix == 8'h0b ? p1_array_index_10088_comb : (p0_start_pix == 8'h0c ? p1_array_index_10089_comb : (p0_start_pix == 8'h0d ? p1_array_index_10090_comb : (p0_start_pix == 8'h0e ? p1_array_index_10091_comb : (p0_start_pix == 8'h0f ? p1_array_index_10092_comb : (p0_start_pix == 8'h10 ? p1_array_index_10093_comb : (p0_start_pix == 8'h11 ? p1_array_index_10094_comb : (p0_start_pix == 8'h12 ? p1_array_index_10095_comb : (p0_start_pix == 8'h13 ? p1_array_index_10096_comb : (p0_start_pix == 8'h14 ? p1_array_index_10097_comb : (p0_start_pix == 8'h15 ? p1_array_index_10098_comb : (p0_start_pix == 8'h16 ? p1_array_index_10099_comb : (p0_start_pix == 8'h17 ? p1_array_index_10100_comb : (p0_start_pix == 8'h18 ? p1_array_index_10101_comb : (p0_start_pix == 8'h19 ? p1_array_index_10102_comb : (p0_start_pix == 8'h1a ? p1_array_index_10103_comb : (p0_start_pix == 8'h1b ? p1_array_index_10104_comb : (p0_start_pix == 8'h1c ? p1_array_index_10105_comb : (p0_start_pix == 8'h1d ? p1_array_index_10106_comb : (p0_start_pix == 8'h1e ? p1_array_index_10107_comb : (p0_start_pix == 8'h1f ? p1_array_index_10108_comb : (p0_start_pix == 8'h20 ? p1_array_index_10109_comb : (p0_start_pix == 8'h21 ? p1_array_index_10110_comb : (p0_start_pix == 8'h22 ? p1_array_index_10111_comb : (p0_start_pix == 8'h23 ? p1_array_index_10112_comb : (p0_start_pix == 8'h24 ? p1_array_index_10113_comb : (p0_start_pix == 8'h25 ? p1_array_index_10114_comb : (p0_start_pix == 8'h26 ? p1_array_index_10115_comb : (p0_start_pix == 8'h27 ? p1_array_index_10116_comb : (p0_start_pix == 8'h28 ? p1_array_index_10117_comb : (p0_start_pix == 8'h29 ? p1_array_index_10118_comb : (p0_start_pix == 8'h2a ? p1_array_index_10119_comb : (p0_start_pix == 8'h2b ? p1_array_index_10120_comb : (p0_start_pix == 8'h2c ? p1_array_index_10121_comb : (p0_start_pix == 8'h2d ? p1_array_index_10122_comb : (p0_start_pix == 8'h2e ? p1_array_index_10123_comb : (p0_start_pix == 8'h2f ? p1_array_index_10124_comb : (p0_start_pix == 8'h30 ? p1_array_index_10125_comb : (p0_start_pix == 8'h31 ? p1_array_index_10126_comb : (p0_start_pix == 8'h32 ? p1_array_index_10127_comb : (p0_start_pix == 8'h33 ? p1_array_index_10128_comb : (p0_start_pix == 8'h34 ? p1_array_index_10129_comb : (p0_start_pix == 8'h35 ? p1_array_index_10130_comb : (p0_start_pix == 8'h36 ? p1_array_index_10131_comb : (p0_start_pix == 8'h37 ? p1_array_index_10132_comb : (p0_start_pix == 8'h38 ? p1_array_index_10133_comb : (p0_start_pix == 8'h39 ? p1_array_index_10134_comb : (p0_start_pix == 8'h3a ? p1_array_index_10135_comb : (p0_start_pix == 8'h3b ? p1_array_index_10136_comb : (p0_start_pix == 8'h3c ? p1_array_index_10137_comb : (p0_start_pix == 8'h3d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign p1_or_10225_comb = {p1_add_10151_comb, p0_start_pix[3:0]} > 9'h03e | ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10151_comb, p0_start_pix[3:0]} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10235_comb = p0_start_pix == 8'h0c | ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_add_10154_comb[8]}}, p1_add_10154_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10245_comb = p1_add_10163_comb > 9'h03e | ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10163_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10255_comb = p0_start_pix == 8'h0b | ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_concat_10167_comb[8]}}, p1_concat_10167_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10266_comb = {p1_add_10177_comb, p0_start_pix[0]} > 9'h03e | ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10177_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10275_comb = p0_start_pix == 8'h0a | ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_add_10186_comb[8]}}, p1_add_10186_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10285_comb = p1_add_10196_comb > 9'h03e | ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10196_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10295_comb = p0_start_pix == 8'h09 | ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_concat_10206_comb[8]}}, p1_concat_10206_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10306_comb = {p1_add_10217_comb, p0_start_pix[1:0]} > 9'h03e | ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10217_comb, p0_start_pix[1:0]} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10315_comb = p0_start_pix == 8'h08 | ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_add_10228_comb[8]}}, p1_add_10228_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10325_comb = p1_add_10238_comb > 9'h03e | ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10238_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10335_comb = p0_start_pix == 8'h07 | ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_concat_10248_comb[8]}}, p1_concat_10248_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10346_comb = {p1_add_10258_comb, p0_start_pix[0]} > 9'h03e | ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10258_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10355_comb = p0_start_pix == 8'h06 | ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_add_10268_comb[8]}}, p1_add_10268_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10366_comb = p1_add_10278_comb > 9'h03e | ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10278_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10374_comb = p0_start_pix == 8'h05 | ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_concat_10288_comb[8]}}, p1_concat_10288_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10386_comb = {p1_add_10298_comb, p0_start_pix[2:0]} > 9'h03e | ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10298_comb, p0_start_pix[2:0]} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10393_comb = p0_start_pix == p1_huff_length_comb | ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_add_10308_comb[8]}}, p1_add_10308_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10404_comb = p1_add_10318_comb > 9'h03e | ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10318_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10410_comb = p0_start_pix == 8'h03 | ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_concat_10328_comb[8]}}, p1_concat_10328_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10423_comb = {p1_add_10338_comb, p0_start_pix[0]} > 9'h03e | ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10338_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10427_comb = p0_start_pix == p1_huff_length__1_comb | ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_add_10348_comb[8]}}, p1_add_10348_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10436_comb = p1_add_10359_comb > 9'h03e | ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10359_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10439_comb = p0_start_pix == 8'h01 | ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_concat_10367_comb[8]}}, p1_concat_10367_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_nor_10440_comb = ~(p0_start_pix == 8'h00 | ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({{23{p1_add_10375_comb[8]}}, p1_add_10375_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000);
  assign p1_or_10447_comb = {p1_add_10378_comb, p0_start_pix[1:0]} > 9'h03e | ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10378_comb, p0_start_pix[1:0]} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10451_comb = p1_add_10397_comb > 9'h03e | ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10397_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_or_10455_comb = {p1_add_10415_comb, p0_start_pix[0]} > 9'h03e | ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10415_comb, p0_start_pix[0]} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000;
  assign p1_nor_10458_comb = ~(p1_add_10438_comb > 9'h03e | ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0000 ? p1_array_index_10077_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0001 ? p1_array_index_10078_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0002 ? p1_array_index_10079_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0003 ? p1_array_index_10080_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0004 ? p1_array_index_10081_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0005 ? p1_array_index_10082_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0006 ? p1_array_index_10083_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0007 ? p1_array_index_10084_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0008 ? p1_array_index_10085_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0009 ? p1_array_index_10086_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_000a ? p1_array_index_10087_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_000b ? p1_array_index_10088_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_000c ? p1_array_index_10089_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_000d ? p1_array_index_10090_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_000e ? p1_array_index_10091_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_000f ? p1_array_index_10092_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0010 ? p1_array_index_10093_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0011 ? p1_array_index_10094_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0012 ? p1_array_index_10095_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0013 ? p1_array_index_10096_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0014 ? p1_array_index_10097_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0015 ? p1_array_index_10098_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0016 ? p1_array_index_10099_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0017 ? p1_array_index_10100_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0018 ? p1_array_index_10101_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0019 ? p1_array_index_10102_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_001a ? p1_array_index_10103_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_001b ? p1_array_index_10104_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_001c ? p1_array_index_10105_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_001d ? p1_array_index_10106_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_001e ? p1_array_index_10107_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_001f ? p1_array_index_10108_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0020 ? p1_array_index_10109_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0021 ? p1_array_index_10110_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0022 ? p1_array_index_10111_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0023 ? p1_array_index_10112_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0024 ? p1_array_index_10113_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0025 ? p1_array_index_10114_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0026 ? p1_array_index_10115_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0027 ? p1_array_index_10116_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0028 ? p1_array_index_10117_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0029 ? p1_array_index_10118_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_002a ? p1_array_index_10119_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_002b ? p1_array_index_10120_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_002c ? p1_array_index_10121_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_002d ? p1_array_index_10122_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_002e ? p1_array_index_10123_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_002f ? p1_array_index_10124_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0030 ? p1_array_index_10125_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0031 ? p1_array_index_10126_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0032 ? p1_array_index_10127_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0033 ? p1_array_index_10128_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0034 ? p1_array_index_10129_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0035 ? p1_array_index_10130_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0036 ? p1_array_index_10131_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0037 ? p1_array_index_10132_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0038 ? p1_array_index_10133_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_0039 ? p1_array_index_10134_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_003a ? p1_array_index_10135_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_003b ? p1_array_index_10136_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_003c ? p1_array_index_10137_comb : ({23'h00_0000, p1_add_10438_comb} == 32'h0000_003d ? p1_array_index_10138_comb : p1_array_index_10139_comb)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) != 10'h000);
  assign p1_and_10585_comb = p1_array_index_10077_comb == 10'h000 & p1_array_index_10078_comb == 10'h000 & p1_array_index_10079_comb == 10'h000 & p1_array_index_10080_comb == 10'h000 & p1_array_index_10081_comb == 10'h000 & p1_array_index_10082_comb == 10'h000 & p1_array_index_10083_comb == 10'h000 & p1_array_index_10084_comb == 10'h000 & p1_array_index_10085_comb == 10'h000 & p1_array_index_10086_comb == 10'h000 & p1_array_index_10087_comb == 10'h000 & p1_array_index_10088_comb == 10'h000 & p1_array_index_10089_comb == 10'h000 & p1_array_index_10090_comb == 10'h000 & p1_array_index_10091_comb == 10'h000 & p1_array_index_10092_comb == 10'h000 & p1_array_index_10093_comb == 10'h000 & p1_array_index_10094_comb == 10'h000 & p1_array_index_10095_comb == 10'h000 & p1_array_index_10096_comb == 10'h000 & p1_array_index_10097_comb == 10'h000 & p1_array_index_10098_comb == 10'h000 & p1_array_index_10099_comb == 10'h000 & p1_array_index_10100_comb == 10'h000 & p1_array_index_10101_comb == 10'h000 & p1_array_index_10102_comb == 10'h000 & p1_array_index_10103_comb == 10'h000 & p1_array_index_10104_comb == 10'h000 & p1_array_index_10105_comb == 10'h000 & p1_array_index_10106_comb == 10'h000 & p1_array_index_10107_comb == 10'h000 & p1_array_index_10108_comb == 10'h000 & p1_array_index_10109_comb == 10'h000 & p1_array_index_10110_comb == 10'h000 & p1_array_index_10111_comb == 10'h000 & p1_array_index_10112_comb == 10'h000 & p1_array_index_10113_comb == 10'h000 & p1_array_index_10114_comb == 10'h000 & p1_array_index_10115_comb == 10'h000 & p1_array_index_10116_comb == 10'h000 & p1_array_index_10117_comb == 10'h000 & p1_array_index_10118_comb == 10'h000 & p1_array_index_10119_comb == 10'h000 & p1_array_index_10120_comb == 10'h000 & p1_array_index_10121_comb == 10'h000 & p1_array_index_10122_comb == 10'h000 & p1_array_index_10123_comb == 10'h000 & p1_array_index_10124_comb == 10'h000 & p1_array_index_10125_comb == 10'h000 & p1_array_index_10126_comb == 10'h000 & p1_array_index_10127_comb == 10'h000 & p1_array_index_10128_comb == 10'h000 & p1_array_index_10129_comb == 10'h000 & p1_array_index_10130_comb == 10'h000 & p1_array_index_10131_comb == 10'h000 & p1_array_index_10132_comb == 10'h000 & p1_array_index_10133_comb == 10'h000 & p1_array_index_10134_comb == 10'h000 & p1_array_index_10135_comb == 10'h000 & p1_array_index_10136_comb == 10'h000 & p1_array_index_10137_comb == 10'h000 & p1_array_index_10138_comb == 10'h000 & p1_array_index_10139_comb == 10'h000;

  // Registers for pipe stage 1:
  reg p1_is_luminance;
  reg p1_or_10174;
  reg p1_or_10193;
  reg p1_or_10213;
  reg [9:0] p1_value__1;
  reg p1_or_10225;
  reg p1_or_10235;
  reg p1_or_10245;
  reg p1_or_10255;
  reg p1_or_10266;
  reg p1_or_10275;
  reg p1_or_10285;
  reg p1_or_10295;
  reg p1_or_10306;
  reg p1_or_10315;
  reg p1_or_10325;
  reg p1_or_10335;
  reg p1_or_10346;
  reg p1_or_10355;
  reg p1_or_10366;
  reg p1_or_10374;
  reg p1_or_10386;
  reg p1_or_10393;
  reg p1_or_10404;
  reg p1_or_10410;
  reg p1_or_10423;
  reg p1_or_10427;
  reg p1_or_10436;
  reg p1_or_10439;
  reg p1_nor_10440;
  reg p1_or_10447;
  reg p1_or_10451;
  reg p1_or_10455;
  reg p1_nor_10458;
  reg p1_and_10585;
  always @ (posedge clk) begin
    p1_is_luminance <= p0_is_luminance;
    p1_or_10174 <= p1_or_10174_comb;
    p1_or_10193 <= p1_or_10193_comb;
    p1_or_10213 <= p1_or_10213_comb;
    p1_value__1 <= p1_value__1_comb;
    p1_or_10225 <= p1_or_10225_comb;
    p1_or_10235 <= p1_or_10235_comb;
    p1_or_10245 <= p1_or_10245_comb;
    p1_or_10255 <= p1_or_10255_comb;
    p1_or_10266 <= p1_or_10266_comb;
    p1_or_10275 <= p1_or_10275_comb;
    p1_or_10285 <= p1_or_10285_comb;
    p1_or_10295 <= p1_or_10295_comb;
    p1_or_10306 <= p1_or_10306_comb;
    p1_or_10315 <= p1_or_10315_comb;
    p1_or_10325 <= p1_or_10325_comb;
    p1_or_10335 <= p1_or_10335_comb;
    p1_or_10346 <= p1_or_10346_comb;
    p1_or_10355 <= p1_or_10355_comb;
    p1_or_10366 <= p1_or_10366_comb;
    p1_or_10374 <= p1_or_10374_comb;
    p1_or_10386 <= p1_or_10386_comb;
    p1_or_10393 <= p1_or_10393_comb;
    p1_or_10404 <= p1_or_10404_comb;
    p1_or_10410 <= p1_or_10410_comb;
    p1_or_10423 <= p1_or_10423_comb;
    p1_or_10427 <= p1_or_10427_comb;
    p1_or_10436 <= p1_or_10436_comb;
    p1_or_10439 <= p1_or_10439_comb;
    p1_nor_10440 <= p1_nor_10440_comb;
    p1_or_10447 <= p1_or_10447_comb;
    p1_or_10451 <= p1_or_10451_comb;
    p1_or_10455 <= p1_or_10455_comb;
    p1_nor_10458 <= p1_nor_10458_comb;
    p1_and_10585 <= p1_and_10585_comb;
  end

  // ===== Pipe stage 2:
  wire [7:0] p2_bin_value__2_comb;
  wire [7:0] p2_bin_value__3_comb;
  wire [7:0] p2_value_abs_comb;
  wire [4:0] p2_sel_10675_comb;
  wire [4:0] p2_sel_10691_comb;
  wire [1:0] p2_huff_length__1_squeezed__1_comb;
  wire [1:0] p2_huff_length__1_squeezed_comb;
  wire [7:0] p2_flipped__1_comb;
  wire [7:0] p2_flipped_comb;
  wire [4:0] p2_sel_10693_comb;
  wire [1:0] p2_sel_10700_comb;
  wire p2_or_reduce_10704_comb;
  wire [4:0] p2_sel_10705_comb;
  wire p2_or_reduce_10707_comb;
  wire p2_or_reduce_10709_comb;
  wire p2_or_reduce_10710_comb;
  wire p2_bit_slice_10711_comb;
  wire p2_ne_10713_comb;
  wire [7:0] p2_Code_list_comb;
  wire [7:0] p2_code_list_comb;
  assign p2_bin_value__2_comb = p1_value__1[7:0];
  assign p2_bin_value__3_comb = -p2_bin_value__2_comb;
  assign p2_value_abs_comb = p1_value__1[9] ? p2_bin_value__3_comb : p2_bin_value__2_comb;
  assign p2_sel_10675_comb = p1_or_10255 ? 5'h0b : (p1_or_10235 ? 5'h0c : (p1_or_10213 ? 5'h0d : (p1_or_10193 ? 5'h0e : (p1_or_10174 ? 5'h0f : 5'h10))));
  assign p2_sel_10691_comb = p1_or_10306 ? 5'h0b : (p1_or_10285 ? 5'h0c : (p1_or_10266 ? 5'h0d : (p1_or_10245 ? 5'h0e : (p1_or_10225 ? 5'h0f : 5'h10))));
  assign p2_huff_length__1_squeezed__1_comb = 2'h1;
  assign p2_huff_length__1_squeezed_comb = 2'h2;
  assign p2_flipped__1_comb = ~p2_bin_value__3_comb;
  assign p2_flipped_comb = 8'hff;
  assign p2_sel_10693_comb = p1_or_10315 ? 5'h08 : (p1_or_10295 ? 5'h09 : (p1_or_10275 ? 5'h0a : p2_sel_10675_comb));
  assign p2_sel_10700_comb = |p2_value_abs_comb[7:2] ? 2'h3 : (|p2_value_abs_comb[7:1] ? p2_huff_length__1_squeezed_comb : p2_huff_length__1_squeezed__1_comb);
  assign p2_or_reduce_10704_comb = |p2_value_abs_comb[7:3];
  assign p2_sel_10705_comb = p1_or_10366 ? 5'h08 : (p1_or_10346 ? 5'h09 : (p1_or_10325 ? 5'h0a : p2_sel_10691_comb));
  assign p2_or_reduce_10707_comb = |p2_value_abs_comb[7:4];
  assign p2_or_reduce_10709_comb = |p2_value_abs_comb[7:5];
  assign p2_or_reduce_10710_comb = |p2_value_abs_comb[7:6];
  assign p2_bit_slice_10711_comb = p2_value_abs_comb[7];
  assign p2_ne_10713_comb = p2_value_abs_comb != 8'h00;
  assign p2_Code_list_comb = $signed(p1_value__1) <= $signed(10'h000) ? p2_flipped__1_comb : p2_bin_value__2_comb;
  assign p2_code_list_comb = p1_value__1 == 10'h000 ? p2_flipped_comb : p2_bin_value__2_comb;

  // Registers for pipe stage 2:
  reg p2_is_luminance;
  reg [9:0] p2_value__1;
  reg p2_or_10335;
  reg [4:0] p2_sel_10693;
  reg p2_or_10355;
  reg [1:0] p2_sel_10700;
  reg p2_or_10374;
  reg p2_or_reduce_10704;
  reg p2_or_10386;
  reg [4:0] p2_sel_10705;
  reg p2_or_10393;
  reg p2_or_reduce_10707;
  reg p2_or_10404;
  reg p2_or_10410;
  reg p2_or_reduce_10709;
  reg p2_or_10423;
  reg p2_or_10427;
  reg p2_or_reduce_10710;
  reg p2_or_10436;
  reg p2_or_10439;
  reg p2_nor_10440;
  reg p2_or_10447;
  reg p2_bit_slice_10711;
  reg p2_or_10451;
  reg p2_ne_10713;
  reg p2_or_10455;
  reg p2_nor_10458;
  reg p2_and_10585;
  reg [7:0] p2_Code_list;
  reg [7:0] p2_code_list;
  always @ (posedge clk) begin
    p2_is_luminance <= p1_is_luminance;
    p2_value__1 <= p1_value__1;
    p2_or_10335 <= p1_or_10335;
    p2_sel_10693 <= p2_sel_10693_comb;
    p2_or_10355 <= p1_or_10355;
    p2_sel_10700 <= p2_sel_10700_comb;
    p2_or_10374 <= p1_or_10374;
    p2_or_reduce_10704 <= p2_or_reduce_10704_comb;
    p2_or_10386 <= p1_or_10386;
    p2_sel_10705 <= p2_sel_10705_comb;
    p2_or_10393 <= p1_or_10393;
    p2_or_reduce_10707 <= p2_or_reduce_10707_comb;
    p2_or_10404 <= p1_or_10404;
    p2_or_10410 <= p1_or_10410;
    p2_or_reduce_10709 <= p2_or_reduce_10709_comb;
    p2_or_10423 <= p1_or_10423;
    p2_or_10427 <= p1_or_10427;
    p2_or_reduce_10710 <= p2_or_reduce_10710_comb;
    p2_or_10436 <= p1_or_10436;
    p2_or_10439 <= p1_or_10439;
    p2_nor_10440 <= p1_nor_10440;
    p2_or_10447 <= p1_or_10447;
    p2_bit_slice_10711 <= p2_bit_slice_10711_comb;
    p2_or_10451 <= p1_or_10451;
    p2_ne_10713 <= p2_ne_10713_comb;
    p2_or_10455 <= p1_or_10455;
    p2_nor_10458 <= p1_nor_10458;
    p2_and_10585 <= p1_and_10585;
    p2_Code_list <= p2_Code_list_comb;
    p2_code_list <= p2_code_list_comb;
  end

  // ===== Pipe stage 3:
  wire [2:0] p3_huff_length_squeezed__17_comb;
  wire [4:0] p3_sel_10803_comb;
  wire [2:0] p3_sel_10812_comb;
  wire [4:0] p3_sel_10819_comb;
  wire [4:0] p3_run__1_comb;
  wire [3:0] p3_sel_10822_comb;
  wire [4:0] p3_sel_10825_comb;
  assign p3_huff_length_squeezed__17_comb = 3'h4;
  assign p3_sel_10803_comb = p2_or_10410 ? 5'h03 : (p2_or_10393 ? 5'h04 : (p2_or_10374 ? 5'h05 : (p2_or_10355 ? 5'h06 : (p2_or_10335 ? 5'h07 : p2_sel_10693))));
  assign p3_sel_10812_comb = p2_or_reduce_10710 ? 3'h7 : (p2_or_reduce_10709 ? 3'h6 : (p2_or_reduce_10707 ? 3'h5 : (p2_or_reduce_10704 ? p3_huff_length_squeezed__17_comb : {1'h0, p2_sel_10700})));
  assign p3_sel_10819_comb = p2_or_10447 ? 5'h03 : (p2_or_10436 ? 5'h04 : (p2_or_10423 ? 5'h05 : (p2_or_10404 ? 5'h06 : (p2_or_10386 ? 5'h07 : p2_sel_10705))));
  assign p3_run__1_comb = (p2_or_10439 ? 5'h01 : (p2_or_10427 ? 5'h02 : p3_sel_10803_comb)) & {5{p2_nor_10440}};
  assign p3_sel_10822_comb = p2_bit_slice_10711 ? 4'h8 : {1'h0, p3_sel_10812_comb};
  assign p3_sel_10825_comb = p2_or_10455 ? 5'h01 : (p2_or_10451 ? 5'h02 : p3_sel_10819_comb);

  // Registers for pipe stage 3:
  reg p3_is_luminance;
  reg [9:0] p3_value__1;
  reg [4:0] p3_run__1;
  reg [3:0] p3_sel_10822;
  reg p3_ne_10713;
  reg [4:0] p3_sel_10825;
  reg p3_nor_10458;
  reg p3_and_10585;
  reg [7:0] p3_Code_list;
  reg [7:0] p3_code_list;
  always @ (posedge clk) begin
    p3_is_luminance <= p2_is_luminance;
    p3_value__1 <= p2_value__1;
    p3_run__1 <= p3_run__1_comb;
    p3_sel_10822 <= p3_sel_10822_comb;
    p3_ne_10713 <= p2_ne_10713;
    p3_sel_10825 <= p3_sel_10825_comb;
    p3_nor_10458 <= p2_nor_10458;
    p3_and_10585 <= p2_and_10585;
    p3_Code_list <= p2_Code_list;
    p3_code_list <= p2_code_list;
  end

  // ===== Pipe stage 4:
  wire [3:0] p4_next_pix_squeezed_const_msb_bits__1_comb;
  wire [3:0] p4_next_pix_squeezed_const_msb_bits_comb;
  wire p4_eq_10853_comb;
  wire [7:0] p4_Code_size_comb;
  wire [2:0] p4_huff_code__1_squeezed_squeezed__16_comb;
  wire [2:0] p4_huff_length_squeezed__18_comb;
  wire [7:0] p4_run_size_str_u8_comb;
  wire [1:0] p4_huff_length__1_squeezed__2_comb;
  wire [1:0] p4_huff_length__1_squeezed__3_comb;
  wire [7:0] p4_sign_ext_10868_comb;
  wire [2:0] p4_sel_10871_comb;
  wire [3:0] p4_Code_size_squeezed_comb;
  wire [3:0] p4_huff_length_squeezed__2_comb;
  wire [5:0] p4_add_10879_comb;
  wire p4_or_10885_comb;
  wire [4:0] p4_Huffman_length_squeezed_comb;
  wire [3:0] p4_next_pix_squeezed_const_msb_bits__2_comb;
  wire [3:0] p4_next_pix_squeezed_comb;
  wire [5:0] p4_now_pix_data__1_comb;
  wire [15:0] p4_Huffman_code_full_comb;
  wire [7:0] p4_code_list__1_comb;
  wire [7:0] p4_next_pix_comb;
  wire [57:0] p4_tuple_10907_comb;
  assign p4_next_pix_squeezed_const_msb_bits__1_comb = 4'h0;
  assign p4_next_pix_squeezed_const_msb_bits_comb = 4'h0;
  assign p4_eq_10853_comb = p3_run__1 == 5'h10;
  assign p4_Code_size_comb = {p4_next_pix_squeezed_const_msb_bits__1_comb, p3_sel_10822} & {8{p3_ne_10713}};
  assign p4_huff_code__1_squeezed_squeezed__16_comb = 3'h1;
  assign p4_huff_length_squeezed__18_comb = 3'h4;
  assign p4_run_size_str_u8_comb = {p3_run__1[3:0], p4_next_pix_squeezed_const_msb_bits_comb} | p4_Code_size_comb;
  assign p4_huff_length__1_squeezed__2_comb = 2'h1;
  assign p4_huff_length__1_squeezed__3_comb = 2'h2;
  assign p4_sign_ext_10868_comb = {8{~p4_eq_10853_comb}};
  assign p4_sel_10871_comb = p3_is_luminance ? p4_huff_length_squeezed__18_comb : p4_huff_code__1_squeezed_squeezed__16_comb;
  assign p4_Code_size_squeezed_comb = p4_Code_size_comb[3:0];
  assign p4_huff_length_squeezed__2_comb = 4'h4;
  assign p4_add_10879_comb = ({1'h0, p3_sel_10825} & {6{p3_nor_10458}}) + 6'h01;
  assign p4_or_10885_comb = p3_and_10585 | p4_eq_10853_comb;
  assign p4_Huffman_length_squeezed_comb = p3_is_luminance ? literal_10863[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_10861[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_next_pix_squeezed_const_msb_bits__2_comb = 4'h0;
  assign p4_next_pix_squeezed_comb = p4_eq_10853_comb ? p4_huff_length_squeezed__2_comb : p4_Code_size_squeezed_comb;
  assign p4_now_pix_data__1_comb = p4_add_10879_comb & p4_sign_ext_10868_comb[5:0];
  assign p4_Huffman_code_full_comb = p3_is_luminance ? literal_10870[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_10869[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_code_list__1_comb = p3_Code_list & p4_sign_ext_10868_comb;
  assign p4_next_pix_comb = {p4_next_pix_squeezed_const_msb_bits__2_comb, p4_next_pix_squeezed_comb};
  assign p4_tuple_10907_comb = {p4_or_10885_comb ? {12'h000, {{1{p4_sel_10871_comb[2]}}, p4_sel_10871_comb}} : p4_Huffman_code_full_comb, {3'h0, p4_or_10885_comb ? {2'h0, p3_is_luminance ? p4_huff_length__1_squeezed__3_comb : p4_huff_length__1_squeezed__2_comb, 1'h0} : p4_Huffman_length_squeezed_comb}, p3_and_10585 ? p3_code_list : p4_code_list__1_comb, p4_next_pix_comb & {8{~p3_and_10585}}, {2'h0, p3_and_10585 ? 6'h3f : p4_now_pix_data__1_comb}, p3_value__1};

  // Registers for pipe stage 4:
  reg [57:0] p4_tuple_10907;
  always @ (posedge clk) begin
    p4_tuple_10907 <= p4_tuple_10907_comb;
  end
  assign out = p4_tuple_10907;
endmodule
