module Huffman_ACenc(
  input wire clk,
  input wire [511:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [35:0] out
);
  wire [4:0] literal_9180[0:251];
  assign literal_9180[0] = 5'h02;
  assign literal_9180[1] = 5'h02;
  assign literal_9180[2] = 5'h03;
  assign literal_9180[3] = 5'h04;
  assign literal_9180[4] = 5'h05;
  assign literal_9180[5] = 5'h07;
  assign literal_9180[6] = 5'h08;
  assign literal_9180[7] = 5'h0e;
  assign literal_9180[8] = 5'h10;
  assign literal_9180[9] = 5'h10;
  assign literal_9180[10] = 5'h10;
  assign literal_9180[11] = 5'h00;
  assign literal_9180[12] = 5'h00;
  assign literal_9180[13] = 5'h00;
  assign literal_9180[14] = 5'h00;
  assign literal_9180[15] = 5'h00;
  assign literal_9180[16] = 5'h00;
  assign literal_9180[17] = 5'h03;
  assign literal_9180[18] = 5'h06;
  assign literal_9180[19] = 5'h07;
  assign literal_9180[20] = 5'h09;
  assign literal_9180[21] = 5'h0b;
  assign literal_9180[22] = 5'h0d;
  assign literal_9180[23] = 5'h10;
  assign literal_9180[24] = 5'h10;
  assign literal_9180[25] = 5'h10;
  assign literal_9180[26] = 5'h10;
  assign literal_9180[27] = 5'h00;
  assign literal_9180[28] = 5'h00;
  assign literal_9180[29] = 5'h00;
  assign literal_9180[30] = 5'h00;
  assign literal_9180[31] = 5'h00;
  assign literal_9180[32] = 5'h00;
  assign literal_9180[33] = 5'h05;
  assign literal_9180[34] = 5'h07;
  assign literal_9180[35] = 5'h0a;
  assign literal_9180[36] = 5'h0c;
  assign literal_9180[37] = 5'h0d;
  assign literal_9180[38] = 5'h10;
  assign literal_9180[39] = 5'h10;
  assign literal_9180[40] = 5'h10;
  assign literal_9180[41] = 5'h10;
  assign literal_9180[42] = 5'h10;
  assign literal_9180[43] = 5'h00;
  assign literal_9180[44] = 5'h00;
  assign literal_9180[45] = 5'h00;
  assign literal_9180[46] = 5'h00;
  assign literal_9180[47] = 5'h00;
  assign literal_9180[48] = 5'h00;
  assign literal_9180[49] = 5'h06;
  assign literal_9180[50] = 5'h08;
  assign literal_9180[51] = 5'h0b;
  assign literal_9180[52] = 5'h0c;
  assign literal_9180[53] = 5'h0f;
  assign literal_9180[54] = 5'h10;
  assign literal_9180[55] = 5'h10;
  assign literal_9180[56] = 5'h10;
  assign literal_9180[57] = 5'h10;
  assign literal_9180[58] = 5'h10;
  assign literal_9180[59] = 5'h00;
  assign literal_9180[60] = 5'h00;
  assign literal_9180[61] = 5'h00;
  assign literal_9180[62] = 5'h00;
  assign literal_9180[63] = 5'h00;
  assign literal_9180[64] = 5'h00;
  assign literal_9180[65] = 5'h06;
  assign literal_9180[66] = 5'h0a;
  assign literal_9180[67] = 5'h0c;
  assign literal_9180[68] = 5'h0f;
  assign literal_9180[69] = 5'h10;
  assign literal_9180[70] = 5'h10;
  assign literal_9180[71] = 5'h10;
  assign literal_9180[72] = 5'h10;
  assign literal_9180[73] = 5'h10;
  assign literal_9180[74] = 5'h10;
  assign literal_9180[75] = 5'h00;
  assign literal_9180[76] = 5'h00;
  assign literal_9180[77] = 5'h00;
  assign literal_9180[78] = 5'h00;
  assign literal_9180[79] = 5'h00;
  assign literal_9180[80] = 5'h00;
  assign literal_9180[81] = 5'h07;
  assign literal_9180[82] = 5'h0b;
  assign literal_9180[83] = 5'h0d;
  assign literal_9180[84] = 5'h10;
  assign literal_9180[85] = 5'h10;
  assign literal_9180[86] = 5'h10;
  assign literal_9180[87] = 5'h10;
  assign literal_9180[88] = 5'h10;
  assign literal_9180[89] = 5'h10;
  assign literal_9180[90] = 5'h10;
  assign literal_9180[91] = 5'h00;
  assign literal_9180[92] = 5'h00;
  assign literal_9180[93] = 5'h00;
  assign literal_9180[94] = 5'h00;
  assign literal_9180[95] = 5'h00;
  assign literal_9180[96] = 5'h00;
  assign literal_9180[97] = 5'h07;
  assign literal_9180[98] = 5'h0b;
  assign literal_9180[99] = 5'h0d;
  assign literal_9180[100] = 5'h10;
  assign literal_9180[101] = 5'h10;
  assign literal_9180[102] = 5'h10;
  assign literal_9180[103] = 5'h10;
  assign literal_9180[104] = 5'h10;
  assign literal_9180[105] = 5'h10;
  assign literal_9180[106] = 5'h10;
  assign literal_9180[107] = 5'h00;
  assign literal_9180[108] = 5'h00;
  assign literal_9180[109] = 5'h00;
  assign literal_9180[110] = 5'h00;
  assign literal_9180[111] = 5'h00;
  assign literal_9180[112] = 5'h00;
  assign literal_9180[113] = 5'h08;
  assign literal_9180[114] = 5'h0b;
  assign literal_9180[115] = 5'h0e;
  assign literal_9180[116] = 5'h10;
  assign literal_9180[117] = 5'h10;
  assign literal_9180[118] = 5'h10;
  assign literal_9180[119] = 5'h10;
  assign literal_9180[120] = 5'h10;
  assign literal_9180[121] = 5'h10;
  assign literal_9180[122] = 5'h10;
  assign literal_9180[123] = 5'h00;
  assign literal_9180[124] = 5'h00;
  assign literal_9180[125] = 5'h00;
  assign literal_9180[126] = 5'h00;
  assign literal_9180[127] = 5'h00;
  assign literal_9180[128] = 5'h00;
  assign literal_9180[129] = 5'h08;
  assign literal_9180[130] = 5'h0c;
  assign literal_9180[131] = 5'h10;
  assign literal_9180[132] = 5'h10;
  assign literal_9180[133] = 5'h10;
  assign literal_9180[134] = 5'h10;
  assign literal_9180[135] = 5'h10;
  assign literal_9180[136] = 5'h10;
  assign literal_9180[137] = 5'h10;
  assign literal_9180[138] = 5'h10;
  assign literal_9180[139] = 5'h00;
  assign literal_9180[140] = 5'h00;
  assign literal_9180[141] = 5'h00;
  assign literal_9180[142] = 5'h00;
  assign literal_9180[143] = 5'h00;
  assign literal_9180[144] = 5'h00;
  assign literal_9180[145] = 5'h08;
  assign literal_9180[146] = 5'h0d;
  assign literal_9180[147] = 5'h10;
  assign literal_9180[148] = 5'h10;
  assign literal_9180[149] = 5'h10;
  assign literal_9180[150] = 5'h10;
  assign literal_9180[151] = 5'h10;
  assign literal_9180[152] = 5'h10;
  assign literal_9180[153] = 5'h10;
  assign literal_9180[154] = 5'h10;
  assign literal_9180[155] = 5'h00;
  assign literal_9180[156] = 5'h00;
  assign literal_9180[157] = 5'h00;
  assign literal_9180[158] = 5'h00;
  assign literal_9180[159] = 5'h00;
  assign literal_9180[160] = 5'h00;
  assign literal_9180[161] = 5'h09;
  assign literal_9180[162] = 5'h0d;
  assign literal_9180[163] = 5'h10;
  assign literal_9180[164] = 5'h10;
  assign literal_9180[165] = 5'h10;
  assign literal_9180[166] = 5'h10;
  assign literal_9180[167] = 5'h10;
  assign literal_9180[168] = 5'h10;
  assign literal_9180[169] = 5'h10;
  assign literal_9180[170] = 5'h10;
  assign literal_9180[171] = 5'h00;
  assign literal_9180[172] = 5'h00;
  assign literal_9180[173] = 5'h00;
  assign literal_9180[174] = 5'h00;
  assign literal_9180[175] = 5'h00;
  assign literal_9180[176] = 5'h00;
  assign literal_9180[177] = 5'h09;
  assign literal_9180[178] = 5'h0d;
  assign literal_9180[179] = 5'h10;
  assign literal_9180[180] = 5'h10;
  assign literal_9180[181] = 5'h10;
  assign literal_9180[182] = 5'h10;
  assign literal_9180[183] = 5'h10;
  assign literal_9180[184] = 5'h10;
  assign literal_9180[185] = 5'h10;
  assign literal_9180[186] = 5'h10;
  assign literal_9180[187] = 5'h00;
  assign literal_9180[188] = 5'h00;
  assign literal_9180[189] = 5'h00;
  assign literal_9180[190] = 5'h00;
  assign literal_9180[191] = 5'h00;
  assign literal_9180[192] = 5'h00;
  assign literal_9180[193] = 5'h0a;
  assign literal_9180[194] = 5'h0d;
  assign literal_9180[195] = 5'h10;
  assign literal_9180[196] = 5'h10;
  assign literal_9180[197] = 5'h10;
  assign literal_9180[198] = 5'h10;
  assign literal_9180[199] = 5'h10;
  assign literal_9180[200] = 5'h10;
  assign literal_9180[201] = 5'h10;
  assign literal_9180[202] = 5'h10;
  assign literal_9180[203] = 5'h00;
  assign literal_9180[204] = 5'h00;
  assign literal_9180[205] = 5'h00;
  assign literal_9180[206] = 5'h00;
  assign literal_9180[207] = 5'h00;
  assign literal_9180[208] = 5'h00;
  assign literal_9180[209] = 5'h0a;
  assign literal_9180[210] = 5'h0e;
  assign literal_9180[211] = 5'h10;
  assign literal_9180[212] = 5'h10;
  assign literal_9180[213] = 5'h10;
  assign literal_9180[214] = 5'h10;
  assign literal_9180[215] = 5'h10;
  assign literal_9180[216] = 5'h10;
  assign literal_9180[217] = 5'h10;
  assign literal_9180[218] = 5'h10;
  assign literal_9180[219] = 5'h00;
  assign literal_9180[220] = 5'h00;
  assign literal_9180[221] = 5'h00;
  assign literal_9180[222] = 5'h00;
  assign literal_9180[223] = 5'h00;
  assign literal_9180[224] = 5'h00;
  assign literal_9180[225] = 5'h0a;
  assign literal_9180[226] = 5'h0f;
  assign literal_9180[227] = 5'h10;
  assign literal_9180[228] = 5'h10;
  assign literal_9180[229] = 5'h10;
  assign literal_9180[230] = 5'h10;
  assign literal_9180[231] = 5'h10;
  assign literal_9180[232] = 5'h10;
  assign literal_9180[233] = 5'h10;
  assign literal_9180[234] = 5'h10;
  assign literal_9180[235] = 5'h00;
  assign literal_9180[236] = 5'h00;
  assign literal_9180[237] = 5'h00;
  assign literal_9180[238] = 5'h00;
  assign literal_9180[239] = 5'h00;
  assign literal_9180[240] = 5'h09;
  assign literal_9180[241] = 5'h0b;
  assign literal_9180[242] = 5'h10;
  assign literal_9180[243] = 5'h10;
  assign literal_9180[244] = 5'h10;
  assign literal_9180[245] = 5'h10;
  assign literal_9180[246] = 5'h10;
  assign literal_9180[247] = 5'h10;
  assign literal_9180[248] = 5'h10;
  assign literal_9180[249] = 5'h10;
  assign literal_9180[250] = 5'h10;
  assign literal_9180[251] = 5'h00;
  wire [4:0] literal_9182[0:251];
  assign literal_9182[0] = 5'h04;
  assign literal_9182[1] = 5'h02;
  assign literal_9182[2] = 5'h02;
  assign literal_9182[3] = 5'h03;
  assign literal_9182[4] = 5'h04;
  assign literal_9182[5] = 5'h05;
  assign literal_9182[6] = 5'h07;
  assign literal_9182[7] = 5'h09;
  assign literal_9182[8] = 5'h10;
  assign literal_9182[9] = 5'h10;
  assign literal_9182[10] = 5'h10;
  assign literal_9182[11] = 5'h00;
  assign literal_9182[12] = 5'h00;
  assign literal_9182[13] = 5'h00;
  assign literal_9182[14] = 5'h00;
  assign literal_9182[15] = 5'h00;
  assign literal_9182[16] = 5'h00;
  assign literal_9182[17] = 5'h04;
  assign literal_9182[18] = 5'h05;
  assign literal_9182[19] = 5'h07;
  assign literal_9182[20] = 5'h09;
  assign literal_9182[21] = 5'h0a;
  assign literal_9182[22] = 5'h0b;
  assign literal_9182[23] = 5'h10;
  assign literal_9182[24] = 5'h10;
  assign literal_9182[25] = 5'h10;
  assign literal_9182[26] = 5'h10;
  assign literal_9182[27] = 5'h00;
  assign literal_9182[28] = 5'h00;
  assign literal_9182[29] = 5'h00;
  assign literal_9182[30] = 5'h00;
  assign literal_9182[31] = 5'h00;
  assign literal_9182[32] = 5'h00;
  assign literal_9182[33] = 5'h05;
  assign literal_9182[34] = 5'h08;
  assign literal_9182[35] = 5'h0a;
  assign literal_9182[36] = 5'h0c;
  assign literal_9182[37] = 5'h0e;
  assign literal_9182[38] = 5'h10;
  assign literal_9182[39] = 5'h10;
  assign literal_9182[40] = 5'h10;
  assign literal_9182[41] = 5'h10;
  assign literal_9182[42] = 5'h10;
  assign literal_9182[43] = 5'h00;
  assign literal_9182[44] = 5'h00;
  assign literal_9182[45] = 5'h00;
  assign literal_9182[46] = 5'h00;
  assign literal_9182[47] = 5'h00;
  assign literal_9182[48] = 5'h00;
  assign literal_9182[49] = 5'h06;
  assign literal_9182[50] = 5'h09;
  assign literal_9182[51] = 5'h0b;
  assign literal_9182[52] = 5'h0e;
  assign literal_9182[53] = 5'h10;
  assign literal_9182[54] = 5'h10;
  assign literal_9182[55] = 5'h10;
  assign literal_9182[56] = 5'h10;
  assign literal_9182[57] = 5'h10;
  assign literal_9182[58] = 5'h10;
  assign literal_9182[59] = 5'h00;
  assign literal_9182[60] = 5'h00;
  assign literal_9182[61] = 5'h00;
  assign literal_9182[62] = 5'h00;
  assign literal_9182[63] = 5'h00;
  assign literal_9182[64] = 5'h00;
  assign literal_9182[65] = 5'h06;
  assign literal_9182[66] = 5'h0a;
  assign literal_9182[67] = 5'h0e;
  assign literal_9182[68] = 5'h10;
  assign literal_9182[69] = 5'h10;
  assign literal_9182[70] = 5'h10;
  assign literal_9182[71] = 5'h10;
  assign literal_9182[72] = 5'h10;
  assign literal_9182[73] = 5'h10;
  assign literal_9182[74] = 5'h10;
  assign literal_9182[75] = 5'h00;
  assign literal_9182[76] = 5'h00;
  assign literal_9182[77] = 5'h00;
  assign literal_9182[78] = 5'h00;
  assign literal_9182[79] = 5'h00;
  assign literal_9182[80] = 5'h00;
  assign literal_9182[81] = 5'h07;
  assign literal_9182[82] = 5'h0a;
  assign literal_9182[83] = 5'h0e;
  assign literal_9182[84] = 5'h10;
  assign literal_9182[85] = 5'h10;
  assign literal_9182[86] = 5'h10;
  assign literal_9182[87] = 5'h10;
  assign literal_9182[88] = 5'h10;
  assign literal_9182[89] = 5'h10;
  assign literal_9182[90] = 5'h10;
  assign literal_9182[91] = 5'h00;
  assign literal_9182[92] = 5'h00;
  assign literal_9182[93] = 5'h00;
  assign literal_9182[94] = 5'h00;
  assign literal_9182[95] = 5'h00;
  assign literal_9182[96] = 5'h00;
  assign literal_9182[97] = 5'h07;
  assign literal_9182[98] = 5'h0c;
  assign literal_9182[99] = 5'h0f;
  assign literal_9182[100] = 5'h10;
  assign literal_9182[101] = 5'h10;
  assign literal_9182[102] = 5'h10;
  assign literal_9182[103] = 5'h10;
  assign literal_9182[104] = 5'h10;
  assign literal_9182[105] = 5'h10;
  assign literal_9182[106] = 5'h10;
  assign literal_9182[107] = 5'h00;
  assign literal_9182[108] = 5'h00;
  assign literal_9182[109] = 5'h00;
  assign literal_9182[110] = 5'h00;
  assign literal_9182[111] = 5'h00;
  assign literal_9182[112] = 5'h00;
  assign literal_9182[113] = 5'h08;
  assign literal_9182[114] = 5'h0c;
  assign literal_9182[115] = 5'h10;
  assign literal_9182[116] = 5'h10;
  assign literal_9182[117] = 5'h10;
  assign literal_9182[118] = 5'h10;
  assign literal_9182[119] = 5'h10;
  assign literal_9182[120] = 5'h10;
  assign literal_9182[121] = 5'h10;
  assign literal_9182[122] = 5'h10;
  assign literal_9182[123] = 5'h00;
  assign literal_9182[124] = 5'h00;
  assign literal_9182[125] = 5'h00;
  assign literal_9182[126] = 5'h00;
  assign literal_9182[127] = 5'h00;
  assign literal_9182[128] = 5'h00;
  assign literal_9182[129] = 5'h09;
  assign literal_9182[130] = 5'h0d;
  assign literal_9182[131] = 5'h10;
  assign literal_9182[132] = 5'h10;
  assign literal_9182[133] = 5'h10;
  assign literal_9182[134] = 5'h10;
  assign literal_9182[135] = 5'h10;
  assign literal_9182[136] = 5'h10;
  assign literal_9182[137] = 5'h10;
  assign literal_9182[138] = 5'h10;
  assign literal_9182[139] = 5'h00;
  assign literal_9182[140] = 5'h00;
  assign literal_9182[141] = 5'h00;
  assign literal_9182[142] = 5'h00;
  assign literal_9182[143] = 5'h00;
  assign literal_9182[144] = 5'h00;
  assign literal_9182[145] = 5'h09;
  assign literal_9182[146] = 5'h0e;
  assign literal_9182[147] = 5'h10;
  assign literal_9182[148] = 5'h10;
  assign literal_9182[149] = 5'h10;
  assign literal_9182[150] = 5'h10;
  assign literal_9182[151] = 5'h10;
  assign literal_9182[152] = 5'h10;
  assign literal_9182[153] = 5'h10;
  assign literal_9182[154] = 5'h10;
  assign literal_9182[155] = 5'h00;
  assign literal_9182[156] = 5'h00;
  assign literal_9182[157] = 5'h00;
  assign literal_9182[158] = 5'h00;
  assign literal_9182[159] = 5'h00;
  assign literal_9182[160] = 5'h00;
  assign literal_9182[161] = 5'h09;
  assign literal_9182[162] = 5'h0e;
  assign literal_9182[163] = 5'h10;
  assign literal_9182[164] = 5'h10;
  assign literal_9182[165] = 5'h10;
  assign literal_9182[166] = 5'h10;
  assign literal_9182[167] = 5'h10;
  assign literal_9182[168] = 5'h10;
  assign literal_9182[169] = 5'h10;
  assign literal_9182[170] = 5'h10;
  assign literal_9182[171] = 5'h00;
  assign literal_9182[172] = 5'h00;
  assign literal_9182[173] = 5'h00;
  assign literal_9182[174] = 5'h00;
  assign literal_9182[175] = 5'h00;
  assign literal_9182[176] = 5'h00;
  assign literal_9182[177] = 5'h0a;
  assign literal_9182[178] = 5'h0f;
  assign literal_9182[179] = 5'h10;
  assign literal_9182[180] = 5'h10;
  assign literal_9182[181] = 5'h10;
  assign literal_9182[182] = 5'h10;
  assign literal_9182[183] = 5'h10;
  assign literal_9182[184] = 5'h10;
  assign literal_9182[185] = 5'h10;
  assign literal_9182[186] = 5'h10;
  assign literal_9182[187] = 5'h00;
  assign literal_9182[188] = 5'h00;
  assign literal_9182[189] = 5'h00;
  assign literal_9182[190] = 5'h00;
  assign literal_9182[191] = 5'h00;
  assign literal_9182[192] = 5'h00;
  assign literal_9182[193] = 5'h0a;
  assign literal_9182[194] = 5'h10;
  assign literal_9182[195] = 5'h10;
  assign literal_9182[196] = 5'h10;
  assign literal_9182[197] = 5'h10;
  assign literal_9182[198] = 5'h10;
  assign literal_9182[199] = 5'h10;
  assign literal_9182[200] = 5'h10;
  assign literal_9182[201] = 5'h10;
  assign literal_9182[202] = 5'h10;
  assign literal_9182[203] = 5'h00;
  assign literal_9182[204] = 5'h00;
  assign literal_9182[205] = 5'h00;
  assign literal_9182[206] = 5'h00;
  assign literal_9182[207] = 5'h00;
  assign literal_9182[208] = 5'h00;
  assign literal_9182[209] = 5'h0a;
  assign literal_9182[210] = 5'h10;
  assign literal_9182[211] = 5'h10;
  assign literal_9182[212] = 5'h10;
  assign literal_9182[213] = 5'h10;
  assign literal_9182[214] = 5'h10;
  assign literal_9182[215] = 5'h10;
  assign literal_9182[216] = 5'h10;
  assign literal_9182[217] = 5'h10;
  assign literal_9182[218] = 5'h10;
  assign literal_9182[219] = 5'h00;
  assign literal_9182[220] = 5'h00;
  assign literal_9182[221] = 5'h00;
  assign literal_9182[222] = 5'h00;
  assign literal_9182[223] = 5'h00;
  assign literal_9182[224] = 5'h00;
  assign literal_9182[225] = 5'h0b;
  assign literal_9182[226] = 5'h10;
  assign literal_9182[227] = 5'h10;
  assign literal_9182[228] = 5'h10;
  assign literal_9182[229] = 5'h10;
  assign literal_9182[230] = 5'h10;
  assign literal_9182[231] = 5'h10;
  assign literal_9182[232] = 5'h10;
  assign literal_9182[233] = 5'h10;
  assign literal_9182[234] = 5'h10;
  assign literal_9182[235] = 5'h00;
  assign literal_9182[236] = 5'h00;
  assign literal_9182[237] = 5'h00;
  assign literal_9182[238] = 5'h00;
  assign literal_9182[239] = 5'h00;
  assign literal_9182[240] = 5'h0c;
  assign literal_9182[241] = 5'h0d;
  assign literal_9182[242] = 5'h10;
  assign literal_9182[243] = 5'h10;
  assign literal_9182[244] = 5'h10;
  assign literal_9182[245] = 5'h10;
  assign literal_9182[246] = 5'h10;
  assign literal_9182[247] = 5'h10;
  assign literal_9182[248] = 5'h10;
  assign literal_9182[249] = 5'h10;
  assign literal_9182[250] = 5'h10;
  assign literal_9182[251] = 5'h00;
  wire [15:0] literal_9183[0:251];
  assign literal_9183[0] = 16'h0001;
  assign literal_9183[1] = 16'h0000;
  assign literal_9183[2] = 16'h0004;
  assign literal_9183[3] = 16'h000c;
  assign literal_9183[4] = 16'h001a;
  assign literal_9183[5] = 16'h0076;
  assign literal_9183[6] = 16'h00f6;
  assign literal_9183[7] = 16'h3fe0;
  assign literal_9183[8] = 16'hff96;
  assign literal_9183[9] = 16'hff97;
  assign literal_9183[10] = 16'hff98;
  assign literal_9183[11] = 16'h0000;
  assign literal_9183[12] = 16'h0000;
  assign literal_9183[13] = 16'h0000;
  assign literal_9183[14] = 16'h0000;
  assign literal_9183[15] = 16'h0000;
  assign literal_9183[16] = 16'h0000;
  assign literal_9183[17] = 16'h0005;
  assign literal_9183[18] = 16'h0038;
  assign literal_9183[19] = 16'h0078;
  assign literal_9183[20] = 16'h01f9;
  assign literal_9183[21] = 16'h07f2;
  assign literal_9183[22] = 16'h1fe8;
  assign literal_9183[23] = 16'hff93;
  assign literal_9183[24] = 16'hff99;
  assign literal_9183[25] = 16'hff9a;
  assign literal_9183[26] = 16'hff9e;
  assign literal_9183[27] = 16'h0000;
  assign literal_9183[28] = 16'h0000;
  assign literal_9183[29] = 16'h0000;
  assign literal_9183[30] = 16'h0000;
  assign literal_9183[31] = 16'h0000;
  assign literal_9183[32] = 16'h0000;
  assign literal_9183[33] = 16'h001b;
  assign literal_9183[34] = 16'h007a;
  assign literal_9183[35] = 16'h03f7;
  assign literal_9183[36] = 16'h0ff0;
  assign literal_9183[37] = 16'h1feb;
  assign literal_9183[38] = 16'hff9b;
  assign literal_9183[39] = 16'hff9f;
  assign literal_9183[40] = 16'hffa8;
  assign literal_9183[41] = 16'hffa9;
  assign literal_9183[42] = 16'hfff1;
  assign literal_9183[43] = 16'h0000;
  assign literal_9183[44] = 16'h0000;
  assign literal_9183[45] = 16'h0000;
  assign literal_9183[46] = 16'h0000;
  assign literal_9183[47] = 16'h0000;
  assign literal_9183[48] = 16'h0000;
  assign literal_9183[49] = 16'h0039;
  assign literal_9183[50] = 16'h00fa;
  assign literal_9183[51] = 16'h07f7;
  assign literal_9183[52] = 16'h0ff1;
  assign literal_9183[53] = 16'h7fc6;
  assign literal_9183[54] = 16'hff9c;
  assign literal_9183[55] = 16'hffa3;
  assign literal_9183[56] = 16'hffd7;
  assign literal_9183[57] = 16'hffe4;
  assign literal_9183[58] = 16'hfff2;
  assign literal_9183[59] = 16'h0000;
  assign literal_9183[60] = 16'h0000;
  assign literal_9183[61] = 16'h0000;
  assign literal_9183[62] = 16'h0000;
  assign literal_9183[63] = 16'h0000;
  assign literal_9183[64] = 16'h0000;
  assign literal_9183[65] = 16'h003a;
  assign literal_9183[66] = 16'h03f8;
  assign literal_9183[67] = 16'h0ff2;
  assign literal_9183[68] = 16'h7fc8;
  assign literal_9183[69] = 16'hff9d;
  assign literal_9183[70] = 16'hffbf;
  assign literal_9183[71] = 16'hffcb;
  assign literal_9183[72] = 16'hffd8;
  assign literal_9183[73] = 16'hffe5;
  assign literal_9183[74] = 16'hfff3;
  assign literal_9183[75] = 16'h0000;
  assign literal_9183[76] = 16'h0000;
  assign literal_9183[77] = 16'h0000;
  assign literal_9183[78] = 16'h0000;
  assign literal_9183[79] = 16'h0000;
  assign literal_9183[80] = 16'h0000;
  assign literal_9183[81] = 16'h0077;
  assign literal_9183[82] = 16'h07f3;
  assign literal_9183[83] = 16'h1fea;
  assign literal_9183[84] = 16'hff94;
  assign literal_9183[85] = 16'hffa2;
  assign literal_9183[86] = 16'hffc0;
  assign literal_9183[87] = 16'hffcc;
  assign literal_9183[88] = 16'hffd9;
  assign literal_9183[89] = 16'hffe6;
  assign literal_9183[90] = 16'hfff4;
  assign literal_9183[91] = 16'h0000;
  assign literal_9183[92] = 16'h0000;
  assign literal_9183[93] = 16'h0000;
  assign literal_9183[94] = 16'h0000;
  assign literal_9183[95] = 16'h0000;
  assign literal_9183[96] = 16'h0000;
  assign literal_9183[97] = 16'h0079;
  assign literal_9183[98] = 16'h07f4;
  assign literal_9183[99] = 16'h1fed;
  assign literal_9183[100] = 16'hffa0;
  assign literal_9183[101] = 16'hffb5;
  assign literal_9183[102] = 16'hffc1;
  assign literal_9183[103] = 16'hffcd;
  assign literal_9183[104] = 16'hffda;
  assign literal_9183[105] = 16'hffe7;
  assign literal_9183[106] = 16'hfff5;
  assign literal_9183[107] = 16'h0000;
  assign literal_9183[108] = 16'h0000;
  assign literal_9183[109] = 16'h0000;
  assign literal_9183[110] = 16'h0000;
  assign literal_9183[111] = 16'h0000;
  assign literal_9183[112] = 16'h0000;
  assign literal_9183[113] = 16'h00f7;
  assign literal_9183[114] = 16'h07f5;
  assign literal_9183[115] = 16'h3fe1;
  assign literal_9183[116] = 16'hffa1;
  assign literal_9183[117] = 16'hffb6;
  assign literal_9183[118] = 16'hffc2;
  assign literal_9183[119] = 16'hffce;
  assign literal_9183[120] = 16'hffdb;
  assign literal_9183[121] = 16'hffe8;
  assign literal_9183[122] = 16'hfff6;
  assign literal_9183[123] = 16'h0000;
  assign literal_9183[124] = 16'h0000;
  assign literal_9183[125] = 16'h0000;
  assign literal_9183[126] = 16'h0000;
  assign literal_9183[127] = 16'h0000;
  assign literal_9183[128] = 16'h0000;
  assign literal_9183[129] = 16'h00f8;
  assign literal_9183[130] = 16'h0ff3;
  assign literal_9183[131] = 16'hff92;
  assign literal_9183[132] = 16'hffad;
  assign literal_9183[133] = 16'hffb7;
  assign literal_9183[134] = 16'hffc3;
  assign literal_9183[135] = 16'hffcf;
  assign literal_9183[136] = 16'hffdc;
  assign literal_9183[137] = 16'hffe9;
  assign literal_9183[138] = 16'hfff7;
  assign literal_9183[139] = 16'h0000;
  assign literal_9183[140] = 16'h0000;
  assign literal_9183[141] = 16'h0000;
  assign literal_9183[142] = 16'h0000;
  assign literal_9183[143] = 16'h0000;
  assign literal_9183[144] = 16'h0000;
  assign literal_9183[145] = 16'h00f9;
  assign literal_9183[146] = 16'h1fe9;
  assign literal_9183[147] = 16'hff95;
  assign literal_9183[148] = 16'hffae;
  assign literal_9183[149] = 16'hffb8;
  assign literal_9183[150] = 16'hffc4;
  assign literal_9183[151] = 16'hffd0;
  assign literal_9183[152] = 16'hffdd;
  assign literal_9183[153] = 16'hffea;
  assign literal_9183[154] = 16'hfff8;
  assign literal_9183[155] = 16'h0000;
  assign literal_9183[156] = 16'h0000;
  assign literal_9183[157] = 16'h0000;
  assign literal_9183[158] = 16'h0000;
  assign literal_9183[159] = 16'h0000;
  assign literal_9183[160] = 16'h0000;
  assign literal_9183[161] = 16'h01f6;
  assign literal_9183[162] = 16'h1fec;
  assign literal_9183[163] = 16'hffa5;
  assign literal_9183[164] = 16'hffaf;
  assign literal_9183[165] = 16'hffb9;
  assign literal_9183[166] = 16'hffc5;
  assign literal_9183[167] = 16'hffd1;
  assign literal_9183[168] = 16'hffde;
  assign literal_9183[169] = 16'hffeb;
  assign literal_9183[170] = 16'hfff9;
  assign literal_9183[171] = 16'h0000;
  assign literal_9183[172] = 16'h0000;
  assign literal_9183[173] = 16'h0000;
  assign literal_9183[174] = 16'h0000;
  assign literal_9183[175] = 16'h0000;
  assign literal_9183[176] = 16'h0000;
  assign literal_9183[177] = 16'h01f7;
  assign literal_9183[178] = 16'h1fee;
  assign literal_9183[179] = 16'hffa6;
  assign literal_9183[180] = 16'hffb0;
  assign literal_9183[181] = 16'hffba;
  assign literal_9183[182] = 16'hffc6;
  assign literal_9183[183] = 16'hffd2;
  assign literal_9183[184] = 16'hffdf;
  assign literal_9183[185] = 16'hffec;
  assign literal_9183[186] = 16'hfffa;
  assign literal_9183[187] = 16'h0000;
  assign literal_9183[188] = 16'h0000;
  assign literal_9183[189] = 16'h0000;
  assign literal_9183[190] = 16'h0000;
  assign literal_9183[191] = 16'h0000;
  assign literal_9183[192] = 16'h0000;
  assign literal_9183[193] = 16'h03f4;
  assign literal_9183[194] = 16'h1fef;
  assign literal_9183[195] = 16'hffa7;
  assign literal_9183[196] = 16'hffb1;
  assign literal_9183[197] = 16'hffbb;
  assign literal_9183[198] = 16'hffc7;
  assign literal_9183[199] = 16'hffd3;
  assign literal_9183[200] = 16'hffe0;
  assign literal_9183[201] = 16'hffed;
  assign literal_9183[202] = 16'hfffb;
  assign literal_9183[203] = 16'h0000;
  assign literal_9183[204] = 16'h0000;
  assign literal_9183[205] = 16'h0000;
  assign literal_9183[206] = 16'h0000;
  assign literal_9183[207] = 16'h0000;
  assign literal_9183[208] = 16'h0000;
  assign literal_9183[209] = 16'h03f5;
  assign literal_9183[210] = 16'h3fe2;
  assign literal_9183[211] = 16'hffaa;
  assign literal_9183[212] = 16'hffb2;
  assign literal_9183[213] = 16'hffbc;
  assign literal_9183[214] = 16'hffc8;
  assign literal_9183[215] = 16'hffd4;
  assign literal_9183[216] = 16'hffe1;
  assign literal_9183[217] = 16'hffee;
  assign literal_9183[218] = 16'hfffc;
  assign literal_9183[219] = 16'h0000;
  assign literal_9183[220] = 16'h0000;
  assign literal_9183[221] = 16'h0000;
  assign literal_9183[222] = 16'h0000;
  assign literal_9183[223] = 16'h0000;
  assign literal_9183[224] = 16'h0000;
  assign literal_9183[225] = 16'h03f6;
  assign literal_9183[226] = 16'h7fc7;
  assign literal_9183[227] = 16'hffab;
  assign literal_9183[228] = 16'hffb3;
  assign literal_9183[229] = 16'hffbd;
  assign literal_9183[230] = 16'hffc9;
  assign literal_9183[231] = 16'hffd5;
  assign literal_9183[232] = 16'hffe2;
  assign literal_9183[233] = 16'hffef;
  assign literal_9183[234] = 16'hfffd;
  assign literal_9183[235] = 16'h0000;
  assign literal_9183[236] = 16'h0000;
  assign literal_9183[237] = 16'h0000;
  assign literal_9183[238] = 16'h0000;
  assign literal_9183[239] = 16'h0000;
  assign literal_9183[240] = 16'h01f8;
  assign literal_9183[241] = 16'h07f6;
  assign literal_9183[242] = 16'hffa4;
  assign literal_9183[243] = 16'hffac;
  assign literal_9183[244] = 16'hffb4;
  assign literal_9183[245] = 16'hffbe;
  assign literal_9183[246] = 16'hffca;
  assign literal_9183[247] = 16'hffd6;
  assign literal_9183[248] = 16'hffe3;
  assign literal_9183[249] = 16'hfff0;
  assign literal_9183[250] = 16'hfffe;
  assign literal_9183[251] = 16'h0000;
  wire [15:0] literal_9184[0:251];
  assign literal_9184[0] = 16'h000c;
  assign literal_9184[1] = 16'h0000;
  assign literal_9184[2] = 16'h0001;
  assign literal_9184[3] = 16'h0004;
  assign literal_9184[4] = 16'h000b;
  assign literal_9184[5] = 16'h001a;
  assign literal_9184[6] = 16'h0079;
  assign literal_9184[7] = 16'h01f9;
  assign literal_9184[8] = 16'hff9c;
  assign literal_9184[9] = 16'hff9f;
  assign literal_9184[10] = 16'hffa0;
  assign literal_9184[11] = 16'h0000;
  assign literal_9184[12] = 16'h0000;
  assign literal_9184[13] = 16'h0000;
  assign literal_9184[14] = 16'h0000;
  assign literal_9184[15] = 16'h0000;
  assign literal_9184[16] = 16'h0000;
  assign literal_9184[17] = 16'h000a;
  assign literal_9184[18] = 16'h001c;
  assign literal_9184[19] = 16'h007a;
  assign literal_9184[20] = 16'h01f5;
  assign literal_9184[21] = 16'h03f4;
  assign literal_9184[22] = 16'h07f8;
  assign literal_9184[23] = 16'hff95;
  assign literal_9184[24] = 16'hffa1;
  assign literal_9184[25] = 16'hffa2;
  assign literal_9184[26] = 16'hffad;
  assign literal_9184[27] = 16'h0000;
  assign literal_9184[28] = 16'h0000;
  assign literal_9184[29] = 16'h0000;
  assign literal_9184[30] = 16'h0000;
  assign literal_9184[31] = 16'h0000;
  assign literal_9184[32] = 16'h0000;
  assign literal_9184[33] = 16'h001b;
  assign literal_9184[34] = 16'h00f8;
  assign literal_9184[35] = 16'h03f7;
  assign literal_9184[36] = 16'h0ff4;
  assign literal_9184[37] = 16'h3fdc;
  assign literal_9184[38] = 16'hff9d;
  assign literal_9184[39] = 16'hff90;
  assign literal_9184[40] = 16'hffac;
  assign literal_9184[41] = 16'hffe3;
  assign literal_9184[42] = 16'hfff1;
  assign literal_9184[43] = 16'h0000;
  assign literal_9184[44] = 16'h0000;
  assign literal_9184[45] = 16'h0000;
  assign literal_9184[46] = 16'h0000;
  assign literal_9184[47] = 16'h0000;
  assign literal_9184[48] = 16'h0000;
  assign literal_9184[49] = 16'h003a;
  assign literal_9184[50] = 16'h01f6;
  assign literal_9184[51] = 16'h07f7;
  assign literal_9184[52] = 16'h3fde;
  assign literal_9184[53] = 16'hff8e;
  assign literal_9184[54] = 16'hff94;
  assign literal_9184[55] = 16'hffc9;
  assign literal_9184[56] = 16'hffd6;
  assign literal_9184[57] = 16'hffe4;
  assign literal_9184[58] = 16'hfff2;
  assign literal_9184[59] = 16'h0000;
  assign literal_9184[60] = 16'h0000;
  assign literal_9184[61] = 16'h0000;
  assign literal_9184[62] = 16'h0000;
  assign literal_9184[63] = 16'h0000;
  assign literal_9184[64] = 16'h0000;
  assign literal_9184[65] = 16'h003b;
  assign literal_9184[66] = 16'h03f6;
  assign literal_9184[67] = 16'h3fdd;
  assign literal_9184[68] = 16'hff8f;
  assign literal_9184[69] = 16'hffa5;
  assign literal_9184[70] = 16'hffa6;
  assign literal_9184[71] = 16'hffca;
  assign literal_9184[72] = 16'hffd7;
  assign literal_9184[73] = 16'hffe5;
  assign literal_9184[74] = 16'hfff3;
  assign literal_9184[75] = 16'h0000;
  assign literal_9184[76] = 16'h0000;
  assign literal_9184[77] = 16'h0000;
  assign literal_9184[78] = 16'h0000;
  assign literal_9184[79] = 16'h0000;
  assign literal_9184[80] = 16'h0000;
  assign literal_9184[81] = 16'h0078;
  assign literal_9184[82] = 16'h03f9;
  assign literal_9184[83] = 16'h3fdf;
  assign literal_9184[84] = 16'hff96;
  assign literal_9184[85] = 16'hffab;
  assign literal_9184[86] = 16'hffa9;
  assign literal_9184[87] = 16'hffcb;
  assign literal_9184[88] = 16'hffd8;
  assign literal_9184[89] = 16'hffe6;
  assign literal_9184[90] = 16'hfff4;
  assign literal_9184[91] = 16'h0000;
  assign literal_9184[92] = 16'h0000;
  assign literal_9184[93] = 16'h0000;
  assign literal_9184[94] = 16'h0000;
  assign literal_9184[95] = 16'h0000;
  assign literal_9184[96] = 16'h0000;
  assign literal_9184[97] = 16'h007b;
  assign literal_9184[98] = 16'h0ff2;
  assign literal_9184[99] = 16'h7fc5;
  assign literal_9184[100] = 16'hff97;
  assign literal_9184[101] = 16'hffb5;
  assign literal_9184[102] = 16'hffbf;
  assign literal_9184[103] = 16'hffcc;
  assign literal_9184[104] = 16'hffd9;
  assign literal_9184[105] = 16'hffe7;
  assign literal_9184[106] = 16'hfff5;
  assign literal_9184[107] = 16'h0000;
  assign literal_9184[108] = 16'h0000;
  assign literal_9184[109] = 16'h0000;
  assign literal_9184[110] = 16'h0000;
  assign literal_9184[111] = 16'h0000;
  assign literal_9184[112] = 16'h0000;
  assign literal_9184[113] = 16'h00f9;
  assign literal_9184[114] = 16'h0ff5;
  assign literal_9184[115] = 16'hff8c;
  assign literal_9184[116] = 16'hff98;
  assign literal_9184[117] = 16'hffb6;
  assign literal_9184[118] = 16'hffc0;
  assign literal_9184[119] = 16'hffcd;
  assign literal_9184[120] = 16'hffda;
  assign literal_9184[121] = 16'hffe8;
  assign literal_9184[122] = 16'hfff6;
  assign literal_9184[123] = 16'h0000;
  assign literal_9184[124] = 16'h0000;
  assign literal_9184[125] = 16'h0000;
  assign literal_9184[126] = 16'h0000;
  assign literal_9184[127] = 16'h0000;
  assign literal_9184[128] = 16'h0000;
  assign literal_9184[129] = 16'h01f4;
  assign literal_9184[130] = 16'h1fec;
  assign literal_9184[131] = 16'hff9e;
  assign literal_9184[132] = 16'hffa3;
  assign literal_9184[133] = 16'hffb7;
  assign literal_9184[134] = 16'hffc1;
  assign literal_9184[135] = 16'hffce;
  assign literal_9184[136] = 16'hffdb;
  assign literal_9184[137] = 16'hffe9;
  assign literal_9184[138] = 16'hfff7;
  assign literal_9184[139] = 16'h0000;
  assign literal_9184[140] = 16'h0000;
  assign literal_9184[141] = 16'h0000;
  assign literal_9184[142] = 16'h0000;
  assign literal_9184[143] = 16'h0000;
  assign literal_9184[144] = 16'h0000;
  assign literal_9184[145] = 16'h01f7;
  assign literal_9184[146] = 16'h3fe0;
  assign literal_9184[147] = 16'hff91;
  assign literal_9184[148] = 16'hffa4;
  assign literal_9184[149] = 16'hffb8;
  assign literal_9184[150] = 16'hffc2;
  assign literal_9184[151] = 16'hffcf;
  assign literal_9184[152] = 16'hffdc;
  assign literal_9184[153] = 16'hffea;
  assign literal_9184[154] = 16'hfff8;
  assign literal_9184[155] = 16'h0000;
  assign literal_9184[156] = 16'h0000;
  assign literal_9184[157] = 16'h0000;
  assign literal_9184[158] = 16'h0000;
  assign literal_9184[159] = 16'h0000;
  assign literal_9184[160] = 16'h0000;
  assign literal_9184[161] = 16'h01f8;
  assign literal_9184[162] = 16'h3fe1;
  assign literal_9184[163] = 16'hff92;
  assign literal_9184[164] = 16'hffa7;
  assign literal_9184[165] = 16'hffb9;
  assign literal_9184[166] = 16'hffc3;
  assign literal_9184[167] = 16'hffd0;
  assign literal_9184[168] = 16'hffdd;
  assign literal_9184[169] = 16'hffeb;
  assign literal_9184[170] = 16'hfff9;
  assign literal_9184[171] = 16'h0000;
  assign literal_9184[172] = 16'h0000;
  assign literal_9184[173] = 16'h0000;
  assign literal_9184[174] = 16'h0000;
  assign literal_9184[175] = 16'h0000;
  assign literal_9184[176] = 16'h0000;
  assign literal_9184[177] = 16'h03f5;
  assign literal_9184[178] = 16'h7fc4;
  assign literal_9184[179] = 16'hff93;
  assign literal_9184[180] = 16'hffa8;
  assign literal_9184[181] = 16'hffba;
  assign literal_9184[182] = 16'hffc4;
  assign literal_9184[183] = 16'hffd1;
  assign literal_9184[184] = 16'hffde;
  assign literal_9184[185] = 16'hffec;
  assign literal_9184[186] = 16'hfffa;
  assign literal_9184[187] = 16'h0000;
  assign literal_9184[188] = 16'h0000;
  assign literal_9184[189] = 16'h0000;
  assign literal_9184[190] = 16'h0000;
  assign literal_9184[191] = 16'h0000;
  assign literal_9184[192] = 16'h0000;
  assign literal_9184[193] = 16'h03f8;
  assign literal_9184[194] = 16'hff8d;
  assign literal_9184[195] = 16'hff99;
  assign literal_9184[196] = 16'hffb1;
  assign literal_9184[197] = 16'hffbb;
  assign literal_9184[198] = 16'hffc5;
  assign literal_9184[199] = 16'hffd2;
  assign literal_9184[200] = 16'hffdf;
  assign literal_9184[201] = 16'hffed;
  assign literal_9184[202] = 16'hfffb;
  assign literal_9184[203] = 16'h0000;
  assign literal_9184[204] = 16'h0000;
  assign literal_9184[205] = 16'h0000;
  assign literal_9184[206] = 16'h0000;
  assign literal_9184[207] = 16'h0000;
  assign literal_9184[208] = 16'h0000;
  assign literal_9184[209] = 16'h03fa;
  assign literal_9184[210] = 16'hff9a;
  assign literal_9184[211] = 16'hffaa;
  assign literal_9184[212] = 16'hffb2;
  assign literal_9184[213] = 16'hffbc;
  assign literal_9184[214] = 16'hffc6;
  assign literal_9184[215] = 16'hffd3;
  assign literal_9184[216] = 16'hffe0;
  assign literal_9184[217] = 16'hffee;
  assign literal_9184[218] = 16'hfffc;
  assign literal_9184[219] = 16'h0000;
  assign literal_9184[220] = 16'h0000;
  assign literal_9184[221] = 16'h0000;
  assign literal_9184[222] = 16'h0000;
  assign literal_9184[223] = 16'h0000;
  assign literal_9184[224] = 16'h0000;
  assign literal_9184[225] = 16'h07f6;
  assign literal_9184[226] = 16'hff9b;
  assign literal_9184[227] = 16'hffaf;
  assign literal_9184[228] = 16'hffb3;
  assign literal_9184[229] = 16'hffbd;
  assign literal_9184[230] = 16'hffc7;
  assign literal_9184[231] = 16'hffd4;
  assign literal_9184[232] = 16'hffe1;
  assign literal_9184[233] = 16'hffef;
  assign literal_9184[234] = 16'hfffd;
  assign literal_9184[235] = 16'h0000;
  assign literal_9184[236] = 16'h0000;
  assign literal_9184[237] = 16'h0000;
  assign literal_9184[238] = 16'h0000;
  assign literal_9184[239] = 16'h0000;
  assign literal_9184[240] = 16'h0ff3;
  assign literal_9184[241] = 16'h1fed;
  assign literal_9184[242] = 16'hffae;
  assign literal_9184[243] = 16'hffb0;
  assign literal_9184[244] = 16'hffb4;
  assign literal_9184[245] = 16'hffbe;
  assign literal_9184[246] = 16'hffc8;
  assign literal_9184[247] = 16'hffd5;
  assign literal_9184[248] = 16'hffe2;
  assign literal_9184[249] = 16'hfff0;
  assign literal_9184[250] = 16'hfffe;
  assign literal_9184[251] = 16'h0000;
  wire [7:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[7:0];
  assign matrix_unflattened[0][1] = matrix[15:8];
  assign matrix_unflattened[0][2] = matrix[23:16];
  assign matrix_unflattened[0][3] = matrix[31:24];
  assign matrix_unflattened[0][4] = matrix[39:32];
  assign matrix_unflattened[0][5] = matrix[47:40];
  assign matrix_unflattened[0][6] = matrix[55:48];
  assign matrix_unflattened[0][7] = matrix[63:56];
  assign matrix_unflattened[1][0] = matrix[71:64];
  assign matrix_unflattened[1][1] = matrix[79:72];
  assign matrix_unflattened[1][2] = matrix[87:80];
  assign matrix_unflattened[1][3] = matrix[95:88];
  assign matrix_unflattened[1][4] = matrix[103:96];
  assign matrix_unflattened[1][5] = matrix[111:104];
  assign matrix_unflattened[1][6] = matrix[119:112];
  assign matrix_unflattened[1][7] = matrix[127:120];
  assign matrix_unflattened[2][0] = matrix[135:128];
  assign matrix_unflattened[2][1] = matrix[143:136];
  assign matrix_unflattened[2][2] = matrix[151:144];
  assign matrix_unflattened[2][3] = matrix[159:152];
  assign matrix_unflattened[2][4] = matrix[167:160];
  assign matrix_unflattened[2][5] = matrix[175:168];
  assign matrix_unflattened[2][6] = matrix[183:176];
  assign matrix_unflattened[2][7] = matrix[191:184];
  assign matrix_unflattened[3][0] = matrix[199:192];
  assign matrix_unflattened[3][1] = matrix[207:200];
  assign matrix_unflattened[3][2] = matrix[215:208];
  assign matrix_unflattened[3][3] = matrix[223:216];
  assign matrix_unflattened[3][4] = matrix[231:224];
  assign matrix_unflattened[3][5] = matrix[239:232];
  assign matrix_unflattened[3][6] = matrix[247:240];
  assign matrix_unflattened[3][7] = matrix[255:248];
  assign matrix_unflattened[4][0] = matrix[263:256];
  assign matrix_unflattened[4][1] = matrix[271:264];
  assign matrix_unflattened[4][2] = matrix[279:272];
  assign matrix_unflattened[4][3] = matrix[287:280];
  assign matrix_unflattened[4][4] = matrix[295:288];
  assign matrix_unflattened[4][5] = matrix[303:296];
  assign matrix_unflattened[4][6] = matrix[311:304];
  assign matrix_unflattened[4][7] = matrix[319:312];
  assign matrix_unflattened[5][0] = matrix[327:320];
  assign matrix_unflattened[5][1] = matrix[335:328];
  assign matrix_unflattened[5][2] = matrix[343:336];
  assign matrix_unflattened[5][3] = matrix[351:344];
  assign matrix_unflattened[5][4] = matrix[359:352];
  assign matrix_unflattened[5][5] = matrix[367:360];
  assign matrix_unflattened[5][6] = matrix[375:368];
  assign matrix_unflattened[5][7] = matrix[383:376];
  assign matrix_unflattened[6][0] = matrix[391:384];
  assign matrix_unflattened[6][1] = matrix[399:392];
  assign matrix_unflattened[6][2] = matrix[407:400];
  assign matrix_unflattened[6][3] = matrix[415:408];
  assign matrix_unflattened[6][4] = matrix[423:416];
  assign matrix_unflattened[6][5] = matrix[431:424];
  assign matrix_unflattened[6][6] = matrix[439:432];
  assign matrix_unflattened[6][7] = matrix[447:440];
  assign matrix_unflattened[7][0] = matrix[455:448];
  assign matrix_unflattened[7][1] = matrix[463:456];
  assign matrix_unflattened[7][2] = matrix[471:464];
  assign matrix_unflattened[7][3] = matrix[479:472];
  assign matrix_unflattened[7][4] = matrix[487:480];
  assign matrix_unflattened[7][5] = matrix[495:488];
  assign matrix_unflattened[7][6] = matrix[503:496];
  assign matrix_unflattened[7][7] = matrix[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_row0_comb[0:7];
  wire [7:0] p1_row1_comb[0:7];
  wire [7:0] p1_array_concat_8180_comb[0:15];
  wire [7:0] p1_row2_comb[0:7];
  wire [7:0] p1_array_concat_8183_comb[0:23];
  wire [7:0] p1_row3_comb[0:7];
  wire [2:0] p1_idx_u8__4_squeezed_comb;
  wire [7:0] p1_array_concat_8186_comb[0:31];
  wire [7:0] p1_row4_comb[0:7];
  wire [2:0] p1_idx_u8__5_squeezed_comb;
  wire [7:0] p1_array_concat_8189_comb[0:39];
  wire [7:0] p1_row5_comb[0:7];
  wire [2:0] p1_idx_u8__6_squeezed_comb;
  wire [7:0] p1_idx_u8__13_comb;
  wire [7:0] p1_array_concat_8195_comb[0:47];
  wire [7:0] p1_row6_comb[0:7];
  wire [2:0] p1_idx_u8__7_squeezed_comb;
  wire [6:0] p1_add_8198_comb;
  wire [7:0] p1_idx_u8__15_comb;
  wire [7:0] p1_idx_u8__17_comb;
  wire [7:0] p1_idx_u8__19_comb;
  wire [7:0] p1_idx_u8__21_comb;
  wire [7:0] p1_idx_u8__23_comb;
  wire [7:0] p1_idx_u8__25_comb;
  wire [7:0] p1_idx_u8__27_comb;
  wire [7:0] p1_idx_u8__29_comb;
  wire [7:0] p1_idx_u8__31_comb;
  wire [7:0] p1_idx_u8__33_comb;
  wire [7:0] p1_idx_u8__35_comb;
  wire [7:0] p1_idx_u8__37_comb;
  wire [7:0] p1_idx_u8__39_comb;
  wire [7:0] p1_idx_u8__41_comb;
  wire [7:0] p1_idx_u8__43_comb;
  wire [7:0] p1_idx_u8__45_comb;
  wire [7:0] p1_idx_u8__47_comb;
  wire [7:0] p1_idx_u8__49_comb;
  wire [7:0] p1_idx_u8__51_comb;
  wire [7:0] p1_idx_u8__53_comb;
  wire [7:0] p1_idx_u8__55_comb;
  wire [7:0] p1_idx_u8__57_comb;
  wire [7:0] p1_idx_u8__59_comb;
  wire [7:0] p1_idx_u8__61_comb;
  wire [7:0] p1_actual_index__13_comb;
  wire [7:0] p1_array_concat_8202_comb[0:55];
  wire [7:0] p1_row7_comb[0:7];
  wire [5:0] p1_add_8207_comb;
  wire [7:0] p1_idx_u8__11_comb;
  wire [7:0] p1_idx_u8__9_comb;
  wire [7:0] p1_idx_u8__7_comb;
  wire [7:0] p1_idx_u8__5_comb;
  wire [7:0] p1_idx_u8__3_comb;
  wire [7:0] p1_idx_u8__1_comb;
  wire [7:0] p1_actual_index__15_comb;
  wire [3:0] p1_add_8388_comb;
  wire [7:0] p1_actual_index__17_comb;
  wire [6:0] p1_add_8390_comb;
  wire [7:0] p1_actual_index__19_comb;
  wire [5:0] p1_add_8392_comb;
  wire [7:0] p1_actual_index__21_comb;
  wire [6:0] p1_add_8394_comb;
  wire [7:0] p1_actual_index__23_comb;
  wire [4:0] p1_add_8396_comb;
  wire [7:0] p1_actual_index__25_comb;
  wire [6:0] p1_add_8398_comb;
  wire [7:0] p1_actual_index__27_comb;
  wire [5:0] p1_add_8400_comb;
  wire [7:0] p1_actual_index__29_comb;
  wire [6:0] p1_add_8402_comb;
  wire [7:0] p1_actual_index__31_comb;
  wire [2:0] p1_add_8404_comb;
  wire [7:0] p1_actual_index__33_comb;
  wire [6:0] p1_add_8406_comb;
  wire [7:0] p1_actual_index__35_comb;
  wire [5:0] p1_add_8408_comb;
  wire [7:0] p1_actual_index__37_comb;
  wire [6:0] p1_add_8410_comb;
  wire [7:0] p1_actual_index__39_comb;
  wire [4:0] p1_add_8412_comb;
  wire [7:0] p1_actual_index__41_comb;
  wire [6:0] p1_add_8414_comb;
  wire [7:0] p1_actual_index__43_comb;
  wire [5:0] p1_add_8416_comb;
  wire [7:0] p1_actual_index__45_comb;
  wire [6:0] p1_add_8418_comb;
  wire [7:0] p1_actual_index__47_comb;
  wire [3:0] p1_add_8420_comb;
  wire [7:0] p1_actual_index__49_comb;
  wire [6:0] p1_add_8422_comb;
  wire [7:0] p1_actual_index__51_comb;
  wire [5:0] p1_add_8424_comb;
  wire [7:0] p1_actual_index__53_comb;
  wire [6:0] p1_add_8426_comb;
  wire [7:0] p1_actual_index__55_comb;
  wire [4:0] p1_add_8428_comb;
  wire [7:0] p1_actual_index__57_comb;
  wire [6:0] p1_add_8430_comb;
  wire [7:0] p1_actual_index__59_comb;
  wire [5:0] p1_add_8432_comb;
  wire [7:0] p1_actual_index__61_comb;
  wire [6:0] p1_add_8434_comb;
  wire [7:0] p1_flat_comb[0:63];
  wire [7:0] p1_actual_index__14_comb;
  wire [7:0] p1_actual_index__11_comb;
  wire [6:0] p1_add_8231_comb;
  wire [7:0] p1_actual_index__9_comb;
  wire [4:0] p1_add_8249_comb;
  wire [7:0] p1_actual_index__7_comb;
  wire [6:0] p1_add_8274_comb;
  wire [7:0] p1_actual_index__5_comb;
  wire [5:0] p1_add_8285_comb;
  wire [7:0] p1_actual_index__3_comb;
  wire [6:0] p1_add_8301_comb;
  wire [7:0] p1_actual_index__1_comb;
  wire [7:0] p1_actual_index__12_comb;
  wire [7:0] p1_actual_index__16_comb;
  wire [7:0] p1_actual_index__18_comb;
  wire [7:0] p1_actual_index__20_comb;
  wire [7:0] p1_actual_index__22_comb;
  wire [7:0] p1_actual_index__24_comb;
  wire [7:0] p1_actual_index__26_comb;
  wire [7:0] p1_actual_index__28_comb;
  wire [7:0] p1_actual_index__30_comb;
  wire [7:0] p1_actual_index__32_comb;
  wire [7:0] p1_actual_index__34_comb;
  wire [7:0] p1_actual_index__36_comb;
  wire [7:0] p1_actual_index__38_comb;
  wire [7:0] p1_actual_index__40_comb;
  wire [7:0] p1_actual_index__42_comb;
  wire [7:0] p1_actual_index__44_comb;
  wire [7:0] p1_actual_index__46_comb;
  wire [7:0] p1_actual_index__48_comb;
  wire [7:0] p1_actual_index__50_comb;
  wire [7:0] p1_actual_index__52_comb;
  wire [7:0] p1_actual_index__54_comb;
  wire [7:0] p1_actual_index__56_comb;
  wire [7:0] p1_actual_index__58_comb;
  wire [7:0] p1_actual_index__60_comb;
  wire [7:0] p1_actual_index__62_comb;
  wire [7:0] p1_and_8226_comb;
  wire [7:0] p1_actual_index__10_comb;
  wire [7:0] p1_actual_index__8_comb;
  wire [7:0] p1_actual_index__6_comb;
  wire [7:0] p1_actual_index__4_comb;
  wire [7:0] p1_actual_index__2_comb;
  wire [7:0] p1_and_8234_comb;
  wire p1_eq_8237_comb;
  wire [7:0] p1_and_8238_comb;
  wire p1_ne_8246_comb;
  wire [1:0] p1_concat_8247_comb;
  wire p1_eq_8248_comb;
  wire [7:0] p1_and_8263_comb;
  wire [7:0] p1_and_8270_comb;
  wire [7:0] p1_and_8277_comb;
  wire [7:0] p1_and_8278_comb;
  wire [7:0] p1_and_8299_comb;
  wire [7:0] p1_and_8308_comb;
  wire [7:0] p1_and_8315_comb;
  wire [7:0] p1_and_8324_comb;
  wire [7:0] p1_and_8329_comb;
  wire [7:0] p1_and_8334_comb;
  wire [7:0] p1_and_8335_comb;
  wire [7:0] p1_and_8336_comb;
  wire p1_eq_8797_comb;
  wire p1_eq_8798_comb;
  wire p1_eq_8799_comb;
  wire p1_eq_8800_comb;
  wire p1_eq_8801_comb;
  wire p1_eq_8802_comb;
  wire p1_eq_8803_comb;
  wire p1_eq_8804_comb;
  wire p1_eq_8805_comb;
  wire p1_eq_8806_comb;
  wire p1_eq_8807_comb;
  wire p1_eq_8808_comb;
  wire p1_eq_8809_comb;
  wire p1_eq_8810_comb;
  wire p1_eq_8811_comb;
  wire p1_eq_8812_comb;
  wire p1_eq_8813_comb;
  wire p1_eq_8814_comb;
  wire p1_eq_8815_comb;
  wire p1_eq_8816_comb;
  wire p1_eq_8817_comb;
  wire p1_eq_8818_comb;
  wire p1_eq_8819_comb;
  wire p1_eq_8820_comb;
  wire p1_eq_8821_comb;
  wire p1_eq_8822_comb;
  wire p1_eq_8823_comb;
  wire p1_eq_8824_comb;
  wire p1_eq_8825_comb;
  wire p1_eq_8826_comb;
  wire p1_eq_8827_comb;
  wire p1_eq_8828_comb;
  wire p1_eq_8829_comb;
  wire p1_eq_8830_comb;
  wire p1_eq_8831_comb;
  wire p1_eq_8832_comb;
  wire p1_eq_8833_comb;
  wire p1_eq_8834_comb;
  wire p1_eq_8835_comb;
  wire p1_eq_8836_comb;
  wire p1_eq_8837_comb;
  wire p1_eq_8838_comb;
  wire p1_eq_8839_comb;
  wire p1_eq_8840_comb;
  wire p1_eq_8841_comb;
  wire p1_eq_8842_comb;
  wire p1_eq_8843_comb;
  wire p1_eq_8844_comb;
  wire [7:0] p1_value_comb;
  assign p1_row0_comb[0] = p0_matrix[3'h0][0];
  assign p1_row0_comb[1] = p0_matrix[3'h0][1];
  assign p1_row0_comb[2] = p0_matrix[3'h0][2];
  assign p1_row0_comb[3] = p0_matrix[3'h0][3];
  assign p1_row0_comb[4] = p0_matrix[3'h0][4];
  assign p1_row0_comb[5] = p0_matrix[3'h0][5];
  assign p1_row0_comb[6] = p0_matrix[3'h0][6];
  assign p1_row0_comb[7] = p0_matrix[3'h0][7];
  assign p1_row1_comb[0] = p0_matrix[3'h1][0];
  assign p1_row1_comb[1] = p0_matrix[3'h1][1];
  assign p1_row1_comb[2] = p0_matrix[3'h1][2];
  assign p1_row1_comb[3] = p0_matrix[3'h1][3];
  assign p1_row1_comb[4] = p0_matrix[3'h1][4];
  assign p1_row1_comb[5] = p0_matrix[3'h1][5];
  assign p1_row1_comb[6] = p0_matrix[3'h1][6];
  assign p1_row1_comb[7] = p0_matrix[3'h1][7];
  assign p1_array_concat_8180_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_8180_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_8180_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_8180_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_8180_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_8180_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_8180_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_8180_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_8180_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_8180_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_8180_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_8180_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_8180_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_8180_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_8180_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_8180_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_8183_comb[0] = p1_array_concat_8180_comb[0];
  assign p1_array_concat_8183_comb[1] = p1_array_concat_8180_comb[1];
  assign p1_array_concat_8183_comb[2] = p1_array_concat_8180_comb[2];
  assign p1_array_concat_8183_comb[3] = p1_array_concat_8180_comb[3];
  assign p1_array_concat_8183_comb[4] = p1_array_concat_8180_comb[4];
  assign p1_array_concat_8183_comb[5] = p1_array_concat_8180_comb[5];
  assign p1_array_concat_8183_comb[6] = p1_array_concat_8180_comb[6];
  assign p1_array_concat_8183_comb[7] = p1_array_concat_8180_comb[7];
  assign p1_array_concat_8183_comb[8] = p1_array_concat_8180_comb[8];
  assign p1_array_concat_8183_comb[9] = p1_array_concat_8180_comb[9];
  assign p1_array_concat_8183_comb[10] = p1_array_concat_8180_comb[10];
  assign p1_array_concat_8183_comb[11] = p1_array_concat_8180_comb[11];
  assign p1_array_concat_8183_comb[12] = p1_array_concat_8180_comb[12];
  assign p1_array_concat_8183_comb[13] = p1_array_concat_8180_comb[13];
  assign p1_array_concat_8183_comb[14] = p1_array_concat_8180_comb[14];
  assign p1_array_concat_8183_comb[15] = p1_array_concat_8180_comb[15];
  assign p1_array_concat_8183_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_8183_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_8183_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_8183_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_8183_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_8183_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_8183_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_8183_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_idx_u8__4_squeezed_comb = 3'h4;
  assign p1_array_concat_8186_comb[0] = p1_array_concat_8183_comb[0];
  assign p1_array_concat_8186_comb[1] = p1_array_concat_8183_comb[1];
  assign p1_array_concat_8186_comb[2] = p1_array_concat_8183_comb[2];
  assign p1_array_concat_8186_comb[3] = p1_array_concat_8183_comb[3];
  assign p1_array_concat_8186_comb[4] = p1_array_concat_8183_comb[4];
  assign p1_array_concat_8186_comb[5] = p1_array_concat_8183_comb[5];
  assign p1_array_concat_8186_comb[6] = p1_array_concat_8183_comb[6];
  assign p1_array_concat_8186_comb[7] = p1_array_concat_8183_comb[7];
  assign p1_array_concat_8186_comb[8] = p1_array_concat_8183_comb[8];
  assign p1_array_concat_8186_comb[9] = p1_array_concat_8183_comb[9];
  assign p1_array_concat_8186_comb[10] = p1_array_concat_8183_comb[10];
  assign p1_array_concat_8186_comb[11] = p1_array_concat_8183_comb[11];
  assign p1_array_concat_8186_comb[12] = p1_array_concat_8183_comb[12];
  assign p1_array_concat_8186_comb[13] = p1_array_concat_8183_comb[13];
  assign p1_array_concat_8186_comb[14] = p1_array_concat_8183_comb[14];
  assign p1_array_concat_8186_comb[15] = p1_array_concat_8183_comb[15];
  assign p1_array_concat_8186_comb[16] = p1_array_concat_8183_comb[16];
  assign p1_array_concat_8186_comb[17] = p1_array_concat_8183_comb[17];
  assign p1_array_concat_8186_comb[18] = p1_array_concat_8183_comb[18];
  assign p1_array_concat_8186_comb[19] = p1_array_concat_8183_comb[19];
  assign p1_array_concat_8186_comb[20] = p1_array_concat_8183_comb[20];
  assign p1_array_concat_8186_comb[21] = p1_array_concat_8183_comb[21];
  assign p1_array_concat_8186_comb[22] = p1_array_concat_8183_comb[22];
  assign p1_array_concat_8186_comb[23] = p1_array_concat_8183_comb[23];
  assign p1_array_concat_8186_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_8186_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_8186_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_8186_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_8186_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_8186_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_8186_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_8186_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[p1_idx_u8__4_squeezed_comb][0];
  assign p1_row4_comb[1] = p0_matrix[p1_idx_u8__4_squeezed_comb][1];
  assign p1_row4_comb[2] = p0_matrix[p1_idx_u8__4_squeezed_comb][2];
  assign p1_row4_comb[3] = p0_matrix[p1_idx_u8__4_squeezed_comb][3];
  assign p1_row4_comb[4] = p0_matrix[p1_idx_u8__4_squeezed_comb][4];
  assign p1_row4_comb[5] = p0_matrix[p1_idx_u8__4_squeezed_comb][5];
  assign p1_row4_comb[6] = p0_matrix[p1_idx_u8__4_squeezed_comb][6];
  assign p1_row4_comb[7] = p0_matrix[p1_idx_u8__4_squeezed_comb][7];
  assign p1_idx_u8__5_squeezed_comb = 3'h5;
  assign p1_array_concat_8189_comb[0] = p1_array_concat_8186_comb[0];
  assign p1_array_concat_8189_comb[1] = p1_array_concat_8186_comb[1];
  assign p1_array_concat_8189_comb[2] = p1_array_concat_8186_comb[2];
  assign p1_array_concat_8189_comb[3] = p1_array_concat_8186_comb[3];
  assign p1_array_concat_8189_comb[4] = p1_array_concat_8186_comb[4];
  assign p1_array_concat_8189_comb[5] = p1_array_concat_8186_comb[5];
  assign p1_array_concat_8189_comb[6] = p1_array_concat_8186_comb[6];
  assign p1_array_concat_8189_comb[7] = p1_array_concat_8186_comb[7];
  assign p1_array_concat_8189_comb[8] = p1_array_concat_8186_comb[8];
  assign p1_array_concat_8189_comb[9] = p1_array_concat_8186_comb[9];
  assign p1_array_concat_8189_comb[10] = p1_array_concat_8186_comb[10];
  assign p1_array_concat_8189_comb[11] = p1_array_concat_8186_comb[11];
  assign p1_array_concat_8189_comb[12] = p1_array_concat_8186_comb[12];
  assign p1_array_concat_8189_comb[13] = p1_array_concat_8186_comb[13];
  assign p1_array_concat_8189_comb[14] = p1_array_concat_8186_comb[14];
  assign p1_array_concat_8189_comb[15] = p1_array_concat_8186_comb[15];
  assign p1_array_concat_8189_comb[16] = p1_array_concat_8186_comb[16];
  assign p1_array_concat_8189_comb[17] = p1_array_concat_8186_comb[17];
  assign p1_array_concat_8189_comb[18] = p1_array_concat_8186_comb[18];
  assign p1_array_concat_8189_comb[19] = p1_array_concat_8186_comb[19];
  assign p1_array_concat_8189_comb[20] = p1_array_concat_8186_comb[20];
  assign p1_array_concat_8189_comb[21] = p1_array_concat_8186_comb[21];
  assign p1_array_concat_8189_comb[22] = p1_array_concat_8186_comb[22];
  assign p1_array_concat_8189_comb[23] = p1_array_concat_8186_comb[23];
  assign p1_array_concat_8189_comb[24] = p1_array_concat_8186_comb[24];
  assign p1_array_concat_8189_comb[25] = p1_array_concat_8186_comb[25];
  assign p1_array_concat_8189_comb[26] = p1_array_concat_8186_comb[26];
  assign p1_array_concat_8189_comb[27] = p1_array_concat_8186_comb[27];
  assign p1_array_concat_8189_comb[28] = p1_array_concat_8186_comb[28];
  assign p1_array_concat_8189_comb[29] = p1_array_concat_8186_comb[29];
  assign p1_array_concat_8189_comb[30] = p1_array_concat_8186_comb[30];
  assign p1_array_concat_8189_comb[31] = p1_array_concat_8186_comb[31];
  assign p1_array_concat_8189_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_8189_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_8189_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_8189_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_8189_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_8189_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_8189_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_8189_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[p1_idx_u8__5_squeezed_comb][0];
  assign p1_row5_comb[1] = p0_matrix[p1_idx_u8__5_squeezed_comb][1];
  assign p1_row5_comb[2] = p0_matrix[p1_idx_u8__5_squeezed_comb][2];
  assign p1_row5_comb[3] = p0_matrix[p1_idx_u8__5_squeezed_comb][3];
  assign p1_row5_comb[4] = p0_matrix[p1_idx_u8__5_squeezed_comb][4];
  assign p1_row5_comb[5] = p0_matrix[p1_idx_u8__5_squeezed_comb][5];
  assign p1_row5_comb[6] = p0_matrix[p1_idx_u8__5_squeezed_comb][6];
  assign p1_row5_comb[7] = p0_matrix[p1_idx_u8__5_squeezed_comb][7];
  assign p1_idx_u8__6_squeezed_comb = 3'h6;
  assign p1_idx_u8__13_comb = 8'h0d;
  assign p1_array_concat_8195_comb[0] = p1_array_concat_8189_comb[0];
  assign p1_array_concat_8195_comb[1] = p1_array_concat_8189_comb[1];
  assign p1_array_concat_8195_comb[2] = p1_array_concat_8189_comb[2];
  assign p1_array_concat_8195_comb[3] = p1_array_concat_8189_comb[3];
  assign p1_array_concat_8195_comb[4] = p1_array_concat_8189_comb[4];
  assign p1_array_concat_8195_comb[5] = p1_array_concat_8189_comb[5];
  assign p1_array_concat_8195_comb[6] = p1_array_concat_8189_comb[6];
  assign p1_array_concat_8195_comb[7] = p1_array_concat_8189_comb[7];
  assign p1_array_concat_8195_comb[8] = p1_array_concat_8189_comb[8];
  assign p1_array_concat_8195_comb[9] = p1_array_concat_8189_comb[9];
  assign p1_array_concat_8195_comb[10] = p1_array_concat_8189_comb[10];
  assign p1_array_concat_8195_comb[11] = p1_array_concat_8189_comb[11];
  assign p1_array_concat_8195_comb[12] = p1_array_concat_8189_comb[12];
  assign p1_array_concat_8195_comb[13] = p1_array_concat_8189_comb[13];
  assign p1_array_concat_8195_comb[14] = p1_array_concat_8189_comb[14];
  assign p1_array_concat_8195_comb[15] = p1_array_concat_8189_comb[15];
  assign p1_array_concat_8195_comb[16] = p1_array_concat_8189_comb[16];
  assign p1_array_concat_8195_comb[17] = p1_array_concat_8189_comb[17];
  assign p1_array_concat_8195_comb[18] = p1_array_concat_8189_comb[18];
  assign p1_array_concat_8195_comb[19] = p1_array_concat_8189_comb[19];
  assign p1_array_concat_8195_comb[20] = p1_array_concat_8189_comb[20];
  assign p1_array_concat_8195_comb[21] = p1_array_concat_8189_comb[21];
  assign p1_array_concat_8195_comb[22] = p1_array_concat_8189_comb[22];
  assign p1_array_concat_8195_comb[23] = p1_array_concat_8189_comb[23];
  assign p1_array_concat_8195_comb[24] = p1_array_concat_8189_comb[24];
  assign p1_array_concat_8195_comb[25] = p1_array_concat_8189_comb[25];
  assign p1_array_concat_8195_comb[26] = p1_array_concat_8189_comb[26];
  assign p1_array_concat_8195_comb[27] = p1_array_concat_8189_comb[27];
  assign p1_array_concat_8195_comb[28] = p1_array_concat_8189_comb[28];
  assign p1_array_concat_8195_comb[29] = p1_array_concat_8189_comb[29];
  assign p1_array_concat_8195_comb[30] = p1_array_concat_8189_comb[30];
  assign p1_array_concat_8195_comb[31] = p1_array_concat_8189_comb[31];
  assign p1_array_concat_8195_comb[32] = p1_array_concat_8189_comb[32];
  assign p1_array_concat_8195_comb[33] = p1_array_concat_8189_comb[33];
  assign p1_array_concat_8195_comb[34] = p1_array_concat_8189_comb[34];
  assign p1_array_concat_8195_comb[35] = p1_array_concat_8189_comb[35];
  assign p1_array_concat_8195_comb[36] = p1_array_concat_8189_comb[36];
  assign p1_array_concat_8195_comb[37] = p1_array_concat_8189_comb[37];
  assign p1_array_concat_8195_comb[38] = p1_array_concat_8189_comb[38];
  assign p1_array_concat_8195_comb[39] = p1_array_concat_8189_comb[39];
  assign p1_array_concat_8195_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_8195_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_8195_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_8195_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_8195_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_8195_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_8195_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_8195_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[p1_idx_u8__6_squeezed_comb][0];
  assign p1_row6_comb[1] = p0_matrix[p1_idx_u8__6_squeezed_comb][1];
  assign p1_row6_comb[2] = p0_matrix[p1_idx_u8__6_squeezed_comb][2];
  assign p1_row6_comb[3] = p0_matrix[p1_idx_u8__6_squeezed_comb][3];
  assign p1_row6_comb[4] = p0_matrix[p1_idx_u8__6_squeezed_comb][4];
  assign p1_row6_comb[5] = p0_matrix[p1_idx_u8__6_squeezed_comb][5];
  assign p1_row6_comb[6] = p0_matrix[p1_idx_u8__6_squeezed_comb][6];
  assign p1_row6_comb[7] = p0_matrix[p1_idx_u8__6_squeezed_comb][7];
  assign p1_idx_u8__7_squeezed_comb = 3'h7;
  assign p1_add_8198_comb = p0_start_pix[7:1] + 7'h07;
  assign p1_idx_u8__15_comb = 8'h0f;
  assign p1_idx_u8__17_comb = 8'h11;
  assign p1_idx_u8__19_comb = 8'h13;
  assign p1_idx_u8__21_comb = 8'h15;
  assign p1_idx_u8__23_comb = 8'h17;
  assign p1_idx_u8__25_comb = 8'h19;
  assign p1_idx_u8__27_comb = 8'h1b;
  assign p1_idx_u8__29_comb = 8'h1d;
  assign p1_idx_u8__31_comb = 8'h1f;
  assign p1_idx_u8__33_comb = 8'h21;
  assign p1_idx_u8__35_comb = 8'h23;
  assign p1_idx_u8__37_comb = 8'h25;
  assign p1_idx_u8__39_comb = 8'h27;
  assign p1_idx_u8__41_comb = 8'h29;
  assign p1_idx_u8__43_comb = 8'h2b;
  assign p1_idx_u8__45_comb = 8'h2d;
  assign p1_idx_u8__47_comb = 8'h2f;
  assign p1_idx_u8__49_comb = 8'h31;
  assign p1_idx_u8__51_comb = 8'h33;
  assign p1_idx_u8__53_comb = 8'h35;
  assign p1_idx_u8__55_comb = 8'h37;
  assign p1_idx_u8__57_comb = 8'h39;
  assign p1_idx_u8__59_comb = 8'h3b;
  assign p1_idx_u8__61_comb = 8'h3d;
  assign p1_actual_index__13_comb = p0_start_pix + p1_idx_u8__13_comb;
  assign p1_array_concat_8202_comb[0] = p1_array_concat_8195_comb[0];
  assign p1_array_concat_8202_comb[1] = p1_array_concat_8195_comb[1];
  assign p1_array_concat_8202_comb[2] = p1_array_concat_8195_comb[2];
  assign p1_array_concat_8202_comb[3] = p1_array_concat_8195_comb[3];
  assign p1_array_concat_8202_comb[4] = p1_array_concat_8195_comb[4];
  assign p1_array_concat_8202_comb[5] = p1_array_concat_8195_comb[5];
  assign p1_array_concat_8202_comb[6] = p1_array_concat_8195_comb[6];
  assign p1_array_concat_8202_comb[7] = p1_array_concat_8195_comb[7];
  assign p1_array_concat_8202_comb[8] = p1_array_concat_8195_comb[8];
  assign p1_array_concat_8202_comb[9] = p1_array_concat_8195_comb[9];
  assign p1_array_concat_8202_comb[10] = p1_array_concat_8195_comb[10];
  assign p1_array_concat_8202_comb[11] = p1_array_concat_8195_comb[11];
  assign p1_array_concat_8202_comb[12] = p1_array_concat_8195_comb[12];
  assign p1_array_concat_8202_comb[13] = p1_array_concat_8195_comb[13];
  assign p1_array_concat_8202_comb[14] = p1_array_concat_8195_comb[14];
  assign p1_array_concat_8202_comb[15] = p1_array_concat_8195_comb[15];
  assign p1_array_concat_8202_comb[16] = p1_array_concat_8195_comb[16];
  assign p1_array_concat_8202_comb[17] = p1_array_concat_8195_comb[17];
  assign p1_array_concat_8202_comb[18] = p1_array_concat_8195_comb[18];
  assign p1_array_concat_8202_comb[19] = p1_array_concat_8195_comb[19];
  assign p1_array_concat_8202_comb[20] = p1_array_concat_8195_comb[20];
  assign p1_array_concat_8202_comb[21] = p1_array_concat_8195_comb[21];
  assign p1_array_concat_8202_comb[22] = p1_array_concat_8195_comb[22];
  assign p1_array_concat_8202_comb[23] = p1_array_concat_8195_comb[23];
  assign p1_array_concat_8202_comb[24] = p1_array_concat_8195_comb[24];
  assign p1_array_concat_8202_comb[25] = p1_array_concat_8195_comb[25];
  assign p1_array_concat_8202_comb[26] = p1_array_concat_8195_comb[26];
  assign p1_array_concat_8202_comb[27] = p1_array_concat_8195_comb[27];
  assign p1_array_concat_8202_comb[28] = p1_array_concat_8195_comb[28];
  assign p1_array_concat_8202_comb[29] = p1_array_concat_8195_comb[29];
  assign p1_array_concat_8202_comb[30] = p1_array_concat_8195_comb[30];
  assign p1_array_concat_8202_comb[31] = p1_array_concat_8195_comb[31];
  assign p1_array_concat_8202_comb[32] = p1_array_concat_8195_comb[32];
  assign p1_array_concat_8202_comb[33] = p1_array_concat_8195_comb[33];
  assign p1_array_concat_8202_comb[34] = p1_array_concat_8195_comb[34];
  assign p1_array_concat_8202_comb[35] = p1_array_concat_8195_comb[35];
  assign p1_array_concat_8202_comb[36] = p1_array_concat_8195_comb[36];
  assign p1_array_concat_8202_comb[37] = p1_array_concat_8195_comb[37];
  assign p1_array_concat_8202_comb[38] = p1_array_concat_8195_comb[38];
  assign p1_array_concat_8202_comb[39] = p1_array_concat_8195_comb[39];
  assign p1_array_concat_8202_comb[40] = p1_array_concat_8195_comb[40];
  assign p1_array_concat_8202_comb[41] = p1_array_concat_8195_comb[41];
  assign p1_array_concat_8202_comb[42] = p1_array_concat_8195_comb[42];
  assign p1_array_concat_8202_comb[43] = p1_array_concat_8195_comb[43];
  assign p1_array_concat_8202_comb[44] = p1_array_concat_8195_comb[44];
  assign p1_array_concat_8202_comb[45] = p1_array_concat_8195_comb[45];
  assign p1_array_concat_8202_comb[46] = p1_array_concat_8195_comb[46];
  assign p1_array_concat_8202_comb[47] = p1_array_concat_8195_comb[47];
  assign p1_array_concat_8202_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_8202_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_8202_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_8202_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_8202_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_8202_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_8202_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_8202_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[p1_idx_u8__7_squeezed_comb][0];
  assign p1_row7_comb[1] = p0_matrix[p1_idx_u8__7_squeezed_comb][1];
  assign p1_row7_comb[2] = p0_matrix[p1_idx_u8__7_squeezed_comb][2];
  assign p1_row7_comb[3] = p0_matrix[p1_idx_u8__7_squeezed_comb][3];
  assign p1_row7_comb[4] = p0_matrix[p1_idx_u8__7_squeezed_comb][4];
  assign p1_row7_comb[5] = p0_matrix[p1_idx_u8__7_squeezed_comb][5];
  assign p1_row7_comb[6] = p0_matrix[p1_idx_u8__7_squeezed_comb][6];
  assign p1_row7_comb[7] = p0_matrix[p1_idx_u8__7_squeezed_comb][7];
  assign p1_add_8207_comb = p0_start_pix[7:2] + 6'h03;
  assign p1_idx_u8__11_comb = 8'h0b;
  assign p1_idx_u8__9_comb = 8'h09;
  assign p1_idx_u8__7_comb = 8'h07;
  assign p1_idx_u8__5_comb = 8'h05;
  assign p1_idx_u8__3_comb = 8'h03;
  assign p1_idx_u8__1_comb = 8'h01;
  assign p1_actual_index__15_comb = p0_start_pix + p1_idx_u8__15_comb;
  assign p1_add_8388_comb = p0_start_pix[7:4] + 4'h1;
  assign p1_actual_index__17_comb = p0_start_pix + p1_idx_u8__17_comb;
  assign p1_add_8390_comb = p0_start_pix[7:1] + 7'h09;
  assign p1_actual_index__19_comb = p0_start_pix + p1_idx_u8__19_comb;
  assign p1_add_8392_comb = p0_start_pix[7:2] + 6'h05;
  assign p1_actual_index__21_comb = p0_start_pix + p1_idx_u8__21_comb;
  assign p1_add_8394_comb = p0_start_pix[7:1] + 7'h0b;
  assign p1_actual_index__23_comb = p0_start_pix + p1_idx_u8__23_comb;
  assign p1_add_8396_comb = p0_start_pix[7:3] + 5'h03;
  assign p1_actual_index__25_comb = p0_start_pix + p1_idx_u8__25_comb;
  assign p1_add_8398_comb = p0_start_pix[7:1] + 7'h0d;
  assign p1_actual_index__27_comb = p0_start_pix + p1_idx_u8__27_comb;
  assign p1_add_8400_comb = p0_start_pix[7:2] + 6'h07;
  assign p1_actual_index__29_comb = p0_start_pix + p1_idx_u8__29_comb;
  assign p1_add_8402_comb = p0_start_pix[7:1] + 7'h0f;
  assign p1_actual_index__31_comb = p0_start_pix + p1_idx_u8__31_comb;
  assign p1_add_8404_comb = p0_start_pix[7:5] + 3'h1;
  assign p1_actual_index__33_comb = p0_start_pix + p1_idx_u8__33_comb;
  assign p1_add_8406_comb = p0_start_pix[7:1] + 7'h11;
  assign p1_actual_index__35_comb = p0_start_pix + p1_idx_u8__35_comb;
  assign p1_add_8408_comb = p0_start_pix[7:2] + 6'h09;
  assign p1_actual_index__37_comb = p0_start_pix + p1_idx_u8__37_comb;
  assign p1_add_8410_comb = p0_start_pix[7:1] + 7'h13;
  assign p1_actual_index__39_comb = p0_start_pix + p1_idx_u8__39_comb;
  assign p1_add_8412_comb = p0_start_pix[7:3] + 5'h05;
  assign p1_actual_index__41_comb = p0_start_pix + p1_idx_u8__41_comb;
  assign p1_add_8414_comb = p0_start_pix[7:1] + 7'h15;
  assign p1_actual_index__43_comb = p0_start_pix + p1_idx_u8__43_comb;
  assign p1_add_8416_comb = p0_start_pix[7:2] + 6'h0b;
  assign p1_actual_index__45_comb = p0_start_pix + p1_idx_u8__45_comb;
  assign p1_add_8418_comb = p0_start_pix[7:1] + 7'h17;
  assign p1_actual_index__47_comb = p0_start_pix + p1_idx_u8__47_comb;
  assign p1_add_8420_comb = p0_start_pix[7:4] + 4'h3;
  assign p1_actual_index__49_comb = p0_start_pix + p1_idx_u8__49_comb;
  assign p1_add_8422_comb = p0_start_pix[7:1] + 7'h19;
  assign p1_actual_index__51_comb = p0_start_pix + p1_idx_u8__51_comb;
  assign p1_add_8424_comb = p0_start_pix[7:2] + 6'h0d;
  assign p1_actual_index__53_comb = p0_start_pix + p1_idx_u8__53_comb;
  assign p1_add_8426_comb = p0_start_pix[7:1] + 7'h1b;
  assign p1_actual_index__55_comb = p0_start_pix + p1_idx_u8__55_comb;
  assign p1_add_8428_comb = p0_start_pix[7:3] + 5'h07;
  assign p1_actual_index__57_comb = p0_start_pix + p1_idx_u8__57_comb;
  assign p1_add_8430_comb = p0_start_pix[7:1] + 7'h1d;
  assign p1_actual_index__59_comb = p0_start_pix + p1_idx_u8__59_comb;
  assign p1_add_8432_comb = p0_start_pix[7:2] + 6'h0f;
  assign p1_actual_index__61_comb = p0_start_pix + p1_idx_u8__61_comb;
  assign p1_add_8434_comb = p0_start_pix[7:1] + 7'h1f;
  assign p1_flat_comb[0] = p1_array_concat_8202_comb[0];
  assign p1_flat_comb[1] = p1_array_concat_8202_comb[1];
  assign p1_flat_comb[2] = p1_array_concat_8202_comb[2];
  assign p1_flat_comb[3] = p1_array_concat_8202_comb[3];
  assign p1_flat_comb[4] = p1_array_concat_8202_comb[4];
  assign p1_flat_comb[5] = p1_array_concat_8202_comb[5];
  assign p1_flat_comb[6] = p1_array_concat_8202_comb[6];
  assign p1_flat_comb[7] = p1_array_concat_8202_comb[7];
  assign p1_flat_comb[8] = p1_array_concat_8202_comb[8];
  assign p1_flat_comb[9] = p1_array_concat_8202_comb[9];
  assign p1_flat_comb[10] = p1_array_concat_8202_comb[10];
  assign p1_flat_comb[11] = p1_array_concat_8202_comb[11];
  assign p1_flat_comb[12] = p1_array_concat_8202_comb[12];
  assign p1_flat_comb[13] = p1_array_concat_8202_comb[13];
  assign p1_flat_comb[14] = p1_array_concat_8202_comb[14];
  assign p1_flat_comb[15] = p1_array_concat_8202_comb[15];
  assign p1_flat_comb[16] = p1_array_concat_8202_comb[16];
  assign p1_flat_comb[17] = p1_array_concat_8202_comb[17];
  assign p1_flat_comb[18] = p1_array_concat_8202_comb[18];
  assign p1_flat_comb[19] = p1_array_concat_8202_comb[19];
  assign p1_flat_comb[20] = p1_array_concat_8202_comb[20];
  assign p1_flat_comb[21] = p1_array_concat_8202_comb[21];
  assign p1_flat_comb[22] = p1_array_concat_8202_comb[22];
  assign p1_flat_comb[23] = p1_array_concat_8202_comb[23];
  assign p1_flat_comb[24] = p1_array_concat_8202_comb[24];
  assign p1_flat_comb[25] = p1_array_concat_8202_comb[25];
  assign p1_flat_comb[26] = p1_array_concat_8202_comb[26];
  assign p1_flat_comb[27] = p1_array_concat_8202_comb[27];
  assign p1_flat_comb[28] = p1_array_concat_8202_comb[28];
  assign p1_flat_comb[29] = p1_array_concat_8202_comb[29];
  assign p1_flat_comb[30] = p1_array_concat_8202_comb[30];
  assign p1_flat_comb[31] = p1_array_concat_8202_comb[31];
  assign p1_flat_comb[32] = p1_array_concat_8202_comb[32];
  assign p1_flat_comb[33] = p1_array_concat_8202_comb[33];
  assign p1_flat_comb[34] = p1_array_concat_8202_comb[34];
  assign p1_flat_comb[35] = p1_array_concat_8202_comb[35];
  assign p1_flat_comb[36] = p1_array_concat_8202_comb[36];
  assign p1_flat_comb[37] = p1_array_concat_8202_comb[37];
  assign p1_flat_comb[38] = p1_array_concat_8202_comb[38];
  assign p1_flat_comb[39] = p1_array_concat_8202_comb[39];
  assign p1_flat_comb[40] = p1_array_concat_8202_comb[40];
  assign p1_flat_comb[41] = p1_array_concat_8202_comb[41];
  assign p1_flat_comb[42] = p1_array_concat_8202_comb[42];
  assign p1_flat_comb[43] = p1_array_concat_8202_comb[43];
  assign p1_flat_comb[44] = p1_array_concat_8202_comb[44];
  assign p1_flat_comb[45] = p1_array_concat_8202_comb[45];
  assign p1_flat_comb[46] = p1_array_concat_8202_comb[46];
  assign p1_flat_comb[47] = p1_array_concat_8202_comb[47];
  assign p1_flat_comb[48] = p1_array_concat_8202_comb[48];
  assign p1_flat_comb[49] = p1_array_concat_8202_comb[49];
  assign p1_flat_comb[50] = p1_array_concat_8202_comb[50];
  assign p1_flat_comb[51] = p1_array_concat_8202_comb[51];
  assign p1_flat_comb[52] = p1_array_concat_8202_comb[52];
  assign p1_flat_comb[53] = p1_array_concat_8202_comb[53];
  assign p1_flat_comb[54] = p1_array_concat_8202_comb[54];
  assign p1_flat_comb[55] = p1_array_concat_8202_comb[55];
  assign p1_flat_comb[56] = p1_row7_comb[0];
  assign p1_flat_comb[57] = p1_row7_comb[1];
  assign p1_flat_comb[58] = p1_row7_comb[2];
  assign p1_flat_comb[59] = p1_row7_comb[3];
  assign p1_flat_comb[60] = p1_row7_comb[4];
  assign p1_flat_comb[61] = p1_row7_comb[5];
  assign p1_flat_comb[62] = p1_row7_comb[6];
  assign p1_flat_comb[63] = p1_row7_comb[7];
  assign p1_actual_index__14_comb = {p1_add_8198_comb, p0_start_pix[0]};
  assign p1_actual_index__11_comb = p0_start_pix + p1_idx_u8__11_comb;
  assign p1_add_8231_comb = p0_start_pix[7:1] + 7'h05;
  assign p1_actual_index__9_comb = p0_start_pix + p1_idx_u8__9_comb;
  assign p1_add_8249_comb = p0_start_pix[7:3] + 5'h01;
  assign p1_actual_index__7_comb = p0_start_pix + p1_idx_u8__7_comb;
  assign p1_add_8274_comb = p0_start_pix[7:1] + 7'h03;
  assign p1_actual_index__5_comb = p0_start_pix + p1_idx_u8__5_comb;
  assign p1_add_8285_comb = p0_start_pix[7:2] + 6'h01;
  assign p1_actual_index__3_comb = p0_start_pix + p1_idx_u8__3_comb;
  assign p1_add_8301_comb = p0_start_pix[7:1] + 7'h01;
  assign p1_actual_index__1_comb = p0_start_pix + p1_idx_u8__1_comb;
  assign p1_actual_index__12_comb = {p1_add_8207_comb, p0_start_pix[1:0]};
  assign p1_actual_index__16_comb = {p1_add_8388_comb, p0_start_pix[3:0]};
  assign p1_actual_index__18_comb = {p1_add_8390_comb, p0_start_pix[0]};
  assign p1_actual_index__20_comb = {p1_add_8392_comb, p0_start_pix[1:0]};
  assign p1_actual_index__22_comb = {p1_add_8394_comb, p0_start_pix[0]};
  assign p1_actual_index__24_comb = {p1_add_8396_comb, p0_start_pix[2:0]};
  assign p1_actual_index__26_comb = {p1_add_8398_comb, p0_start_pix[0]};
  assign p1_actual_index__28_comb = {p1_add_8400_comb, p0_start_pix[1:0]};
  assign p1_actual_index__30_comb = {p1_add_8402_comb, p0_start_pix[0]};
  assign p1_actual_index__32_comb = {p1_add_8404_comb, p0_start_pix[4:0]};
  assign p1_actual_index__34_comb = {p1_add_8406_comb, p0_start_pix[0]};
  assign p1_actual_index__36_comb = {p1_add_8408_comb, p0_start_pix[1:0]};
  assign p1_actual_index__38_comb = {p1_add_8410_comb, p0_start_pix[0]};
  assign p1_actual_index__40_comb = {p1_add_8412_comb, p0_start_pix[2:0]};
  assign p1_actual_index__42_comb = {p1_add_8414_comb, p0_start_pix[0]};
  assign p1_actual_index__44_comb = {p1_add_8416_comb, p0_start_pix[1:0]};
  assign p1_actual_index__46_comb = {p1_add_8418_comb, p0_start_pix[0]};
  assign p1_actual_index__48_comb = {p1_add_8420_comb, p0_start_pix[3:0]};
  assign p1_actual_index__50_comb = {p1_add_8422_comb, p0_start_pix[0]};
  assign p1_actual_index__52_comb = {p1_add_8424_comb, p0_start_pix[1:0]};
  assign p1_actual_index__54_comb = {p1_add_8426_comb, p0_start_pix[0]};
  assign p1_actual_index__56_comb = {p1_add_8428_comb, p0_start_pix[2:0]};
  assign p1_actual_index__58_comb = {p1_add_8430_comb, p0_start_pix[0]};
  assign p1_actual_index__60_comb = {p1_add_8432_comb, p0_start_pix[1:0]};
  assign p1_actual_index__62_comb = {p1_add_8434_comb, p0_start_pix[0]};
  assign p1_and_8226_comb = p1_flat_comb[p1_actual_index__14_comb > 8'h3f ? 6'h3f : p1_actual_index__14_comb[5:0]] & {8{~(p1_add_8198_comb[5] | p1_add_8198_comb[6])}};
  assign p1_actual_index__10_comb = {p1_add_8231_comb, p0_start_pix[0]};
  assign p1_actual_index__8_comb = {p1_add_8249_comb, p0_start_pix[2:0]};
  assign p1_actual_index__6_comb = {p1_add_8274_comb, p0_start_pix[0]};
  assign p1_actual_index__4_comb = {p1_add_8285_comb, p0_start_pix[1:0]};
  assign p1_actual_index__2_comb = {p1_add_8301_comb, p0_start_pix[0]};
  assign p1_and_8234_comb = p1_flat_comb[p1_actual_index__13_comb > 8'h3f ? 6'h3f : p1_actual_index__13_comb[5:0]] & {8{~(p1_actual_index__13_comb[6] | p1_actual_index__13_comb[7])}};
  assign p1_eq_8237_comb = p1_and_8226_comb == 8'h00;
  assign p1_and_8238_comb = p1_flat_comb[p1_actual_index__12_comb > 8'h3f ? 6'h3f : p1_actual_index__12_comb[5:0]] & {8{~(p1_add_8207_comb[4] | p1_add_8207_comb[5])}};
  assign p1_ne_8246_comb = p1_and_8234_comb != 8'h00;
  assign p1_concat_8247_comb = {1'h1, p1_eq_8237_comb};
  assign p1_eq_8248_comb = p1_and_8238_comb == 8'h00;
  assign p1_and_8263_comb = p1_flat_comb[p1_actual_index__11_comb > 8'h3f ? 6'h3f : p1_actual_index__11_comb[5:0]] & {8{~(p1_actual_index__11_comb[6] | p1_actual_index__11_comb[7])}};
  assign p1_and_8270_comb = p1_flat_comb[p1_actual_index__10_comb > 8'h3f ? 6'h3f : p1_actual_index__10_comb[5:0]] & {8{~(p1_add_8231_comb[5] | p1_add_8231_comb[6])}};
  assign p1_and_8277_comb = p1_flat_comb[p1_actual_index__9_comb > 8'h3f ? 6'h3f : p1_actual_index__9_comb[5:0]] & {8{~(p1_actual_index__9_comb[6] | p1_actual_index__9_comb[7])}};
  assign p1_and_8278_comb = p1_flat_comb[p1_actual_index__8_comb > 8'h3f ? 6'h3f : p1_actual_index__8_comb[5:0]] & {8{~(p1_add_8249_comb[3] | p1_add_8249_comb[4])}};
  assign p1_and_8299_comb = p1_flat_comb[p1_actual_index__7_comb > 8'h3f ? 6'h3f : p1_actual_index__7_comb[5:0]] & {8{~(p1_actual_index__7_comb[6] | p1_actual_index__7_comb[7])}};
  assign p1_and_8308_comb = p1_flat_comb[p1_actual_index__6_comb > 8'h3f ? 6'h3f : p1_actual_index__6_comb[5:0]] & {8{~(p1_add_8274_comb[5] | p1_add_8274_comb[6])}};
  assign p1_and_8315_comb = p1_flat_comb[p1_actual_index__5_comb > 8'h3f ? 6'h3f : p1_actual_index__5_comb[5:0]] & {8{~(p1_actual_index__5_comb[6] | p1_actual_index__5_comb[7])}};
  assign p1_and_8324_comb = p1_flat_comb[p1_actual_index__4_comb > 8'h3f ? 6'h3f : p1_actual_index__4_comb[5:0]] & {8{~(p1_add_8285_comb[4] | p1_add_8285_comb[5])}};
  assign p1_and_8329_comb = p1_flat_comb[p1_actual_index__3_comb > 8'h3f ? 6'h3f : p1_actual_index__3_comb[5:0]] & {8{~(p1_actual_index__3_comb[6] | p1_actual_index__3_comb[7])}};
  assign p1_and_8334_comb = p1_flat_comb[p1_actual_index__2_comb > 8'h3f ? 6'h3f : p1_actual_index__2_comb[5:0]] & {8{~(p1_add_8301_comb[5] | p1_add_8301_comb[6])}};
  assign p1_and_8335_comb = p1_flat_comb[p0_start_pix > 8'h3f ? 6'h3f : p0_start_pix[5:0]] & {8{~(p0_start_pix[6] | p0_start_pix[7])}};
  assign p1_and_8336_comb = p1_flat_comb[p1_actual_index__1_comb > 8'h3f ? 6'h3f : p1_actual_index__1_comb[5:0]] & {8{~(p1_actual_index__1_comb[6] | p1_actual_index__1_comb[7])}};
  assign p1_eq_8797_comb = (p1_flat_comb[p1_actual_index__15_comb > 8'h3f ? 6'h3f : p1_actual_index__15_comb[5:0]] & {8{~(p1_actual_index__15_comb[6] | p1_actual_index__15_comb[7])}}) == 8'h00;
  assign p1_eq_8798_comb = (p1_flat_comb[p1_actual_index__16_comb > 8'h3f ? 6'h3f : p1_actual_index__16_comb[5:0]] & {8{~(p1_add_8388_comb[2] | p1_add_8388_comb[3])}}) == 8'h00;
  assign p1_eq_8799_comb = (p1_flat_comb[p1_actual_index__17_comb > 8'h3f ? 6'h3f : p1_actual_index__17_comb[5:0]] & {8{~(p1_actual_index__17_comb[6] | p1_actual_index__17_comb[7])}}) == 8'h00;
  assign p1_eq_8800_comb = (p1_flat_comb[p1_actual_index__18_comb > 8'h3f ? 6'h3f : p1_actual_index__18_comb[5:0]] & {8{~(p1_add_8390_comb[5] | p1_add_8390_comb[6])}}) == 8'h00;
  assign p1_eq_8801_comb = (p1_flat_comb[p1_actual_index__19_comb > 8'h3f ? 6'h3f : p1_actual_index__19_comb[5:0]] & {8{~(p1_actual_index__19_comb[6] | p1_actual_index__19_comb[7])}}) == 8'h00;
  assign p1_eq_8802_comb = (p1_flat_comb[p1_actual_index__20_comb > 8'h3f ? 6'h3f : p1_actual_index__20_comb[5:0]] & {8{~(p1_add_8392_comb[4] | p1_add_8392_comb[5])}}) == 8'h00;
  assign p1_eq_8803_comb = (p1_flat_comb[p1_actual_index__21_comb > 8'h3f ? 6'h3f : p1_actual_index__21_comb[5:0]] & {8{~(p1_actual_index__21_comb[6] | p1_actual_index__21_comb[7])}}) == 8'h00;
  assign p1_eq_8804_comb = (p1_flat_comb[p1_actual_index__22_comb > 8'h3f ? 6'h3f : p1_actual_index__22_comb[5:0]] & {8{~(p1_add_8394_comb[5] | p1_add_8394_comb[6])}}) == 8'h00;
  assign p1_eq_8805_comb = (p1_flat_comb[p1_actual_index__23_comb > 8'h3f ? 6'h3f : p1_actual_index__23_comb[5:0]] & {8{~(p1_actual_index__23_comb[6] | p1_actual_index__23_comb[7])}}) == 8'h00;
  assign p1_eq_8806_comb = (p1_flat_comb[p1_actual_index__24_comb > 8'h3f ? 6'h3f : p1_actual_index__24_comb[5:0]] & {8{~(p1_add_8396_comb[3] | p1_add_8396_comb[4])}}) == 8'h00;
  assign p1_eq_8807_comb = (p1_flat_comb[p1_actual_index__25_comb > 8'h3f ? 6'h3f : p1_actual_index__25_comb[5:0]] & {8{~(p1_actual_index__25_comb[6] | p1_actual_index__25_comb[7])}}) == 8'h00;
  assign p1_eq_8808_comb = (p1_flat_comb[p1_actual_index__26_comb > 8'h3f ? 6'h3f : p1_actual_index__26_comb[5:0]] & {8{~(p1_add_8398_comb[5] | p1_add_8398_comb[6])}}) == 8'h00;
  assign p1_eq_8809_comb = (p1_flat_comb[p1_actual_index__27_comb > 8'h3f ? 6'h3f : p1_actual_index__27_comb[5:0]] & {8{~(p1_actual_index__27_comb[6] | p1_actual_index__27_comb[7])}}) == 8'h00;
  assign p1_eq_8810_comb = (p1_flat_comb[p1_actual_index__28_comb > 8'h3f ? 6'h3f : p1_actual_index__28_comb[5:0]] & {8{~(p1_add_8400_comb[4] | p1_add_8400_comb[5])}}) == 8'h00;
  assign p1_eq_8811_comb = (p1_flat_comb[p1_actual_index__29_comb > 8'h3f ? 6'h3f : p1_actual_index__29_comb[5:0]] & {8{~(p1_actual_index__29_comb[6] | p1_actual_index__29_comb[7])}}) == 8'h00;
  assign p1_eq_8812_comb = (p1_flat_comb[p1_actual_index__30_comb > 8'h3f ? 6'h3f : p1_actual_index__30_comb[5:0]] & {8{~(p1_add_8402_comb[5] | p1_add_8402_comb[6])}}) == 8'h00;
  assign p1_eq_8813_comb = (p1_flat_comb[p1_actual_index__31_comb > 8'h3f ? 6'h3f : p1_actual_index__31_comb[5:0]] & {8{~(p1_actual_index__31_comb[6] | p1_actual_index__31_comb[7])}}) == 8'h00;
  assign p1_eq_8814_comb = (p1_flat_comb[p1_actual_index__32_comb > 8'h3f ? 6'h3f : p1_actual_index__32_comb[5:0]] & {8{~(p1_add_8404_comb[1] | p1_add_8404_comb[2])}}) == 8'h00;
  assign p1_eq_8815_comb = (p1_flat_comb[p1_actual_index__33_comb > 8'h3f ? 6'h3f : p1_actual_index__33_comb[5:0]] & {8{~(p1_actual_index__33_comb[6] | p1_actual_index__33_comb[7])}}) == 8'h00;
  assign p1_eq_8816_comb = (p1_flat_comb[p1_actual_index__34_comb > 8'h3f ? 6'h3f : p1_actual_index__34_comb[5:0]] & {8{~(p1_add_8406_comb[5] | p1_add_8406_comb[6])}}) == 8'h00;
  assign p1_eq_8817_comb = (p1_flat_comb[p1_actual_index__35_comb > 8'h3f ? 6'h3f : p1_actual_index__35_comb[5:0]] & {8{~(p1_actual_index__35_comb[6] | p1_actual_index__35_comb[7])}}) == 8'h00;
  assign p1_eq_8818_comb = (p1_flat_comb[p1_actual_index__36_comb > 8'h3f ? 6'h3f : p1_actual_index__36_comb[5:0]] & {8{~(p1_add_8408_comb[4] | p1_add_8408_comb[5])}}) == 8'h00;
  assign p1_eq_8819_comb = (p1_flat_comb[p1_actual_index__37_comb > 8'h3f ? 6'h3f : p1_actual_index__37_comb[5:0]] & {8{~(p1_actual_index__37_comb[6] | p1_actual_index__37_comb[7])}}) == 8'h00;
  assign p1_eq_8820_comb = (p1_flat_comb[p1_actual_index__38_comb > 8'h3f ? 6'h3f : p1_actual_index__38_comb[5:0]] & {8{~(p1_add_8410_comb[5] | p1_add_8410_comb[6])}}) == 8'h00;
  assign p1_eq_8821_comb = (p1_flat_comb[p1_actual_index__39_comb > 8'h3f ? 6'h3f : p1_actual_index__39_comb[5:0]] & {8{~(p1_actual_index__39_comb[6] | p1_actual_index__39_comb[7])}}) == 8'h00;
  assign p1_eq_8822_comb = (p1_flat_comb[p1_actual_index__40_comb > 8'h3f ? 6'h3f : p1_actual_index__40_comb[5:0]] & {8{~(p1_add_8412_comb[3] | p1_add_8412_comb[4])}}) == 8'h00;
  assign p1_eq_8823_comb = (p1_flat_comb[p1_actual_index__41_comb > 8'h3f ? 6'h3f : p1_actual_index__41_comb[5:0]] & {8{~(p1_actual_index__41_comb[6] | p1_actual_index__41_comb[7])}}) == 8'h00;
  assign p1_eq_8824_comb = (p1_flat_comb[p1_actual_index__42_comb > 8'h3f ? 6'h3f : p1_actual_index__42_comb[5:0]] & {8{~(p1_add_8414_comb[5] | p1_add_8414_comb[6])}}) == 8'h00;
  assign p1_eq_8825_comb = (p1_flat_comb[p1_actual_index__43_comb > 8'h3f ? 6'h3f : p1_actual_index__43_comb[5:0]] & {8{~(p1_actual_index__43_comb[6] | p1_actual_index__43_comb[7])}}) == 8'h00;
  assign p1_eq_8826_comb = (p1_flat_comb[p1_actual_index__44_comb > 8'h3f ? 6'h3f : p1_actual_index__44_comb[5:0]] & {8{~(p1_add_8416_comb[4] | p1_add_8416_comb[5])}}) == 8'h00;
  assign p1_eq_8827_comb = (p1_flat_comb[p1_actual_index__45_comb > 8'h3f ? 6'h3f : p1_actual_index__45_comb[5:0]] & {8{~(p1_actual_index__45_comb[6] | p1_actual_index__45_comb[7])}}) == 8'h00;
  assign p1_eq_8828_comb = (p1_flat_comb[p1_actual_index__46_comb > 8'h3f ? 6'h3f : p1_actual_index__46_comb[5:0]] & {8{~(p1_add_8418_comb[5] | p1_add_8418_comb[6])}}) == 8'h00;
  assign p1_eq_8829_comb = (p1_flat_comb[p1_actual_index__47_comb > 8'h3f ? 6'h3f : p1_actual_index__47_comb[5:0]] & {8{~(p1_actual_index__47_comb[6] | p1_actual_index__47_comb[7])}}) == 8'h00;
  assign p1_eq_8830_comb = (p1_flat_comb[p1_actual_index__48_comb > 8'h3f ? 6'h3f : p1_actual_index__48_comb[5:0]] & {8{~(p1_add_8420_comb[2] | p1_add_8420_comb[3])}}) == 8'h00;
  assign p1_eq_8831_comb = (p1_flat_comb[p1_actual_index__49_comb > 8'h3f ? 6'h3f : p1_actual_index__49_comb[5:0]] & {8{~(p1_actual_index__49_comb[6] | p1_actual_index__49_comb[7])}}) == 8'h00;
  assign p1_eq_8832_comb = (p1_flat_comb[p1_actual_index__50_comb > 8'h3f ? 6'h3f : p1_actual_index__50_comb[5:0]] & {8{~(p1_add_8422_comb[5] | p1_add_8422_comb[6])}}) == 8'h00;
  assign p1_eq_8833_comb = (p1_flat_comb[p1_actual_index__51_comb > 8'h3f ? 6'h3f : p1_actual_index__51_comb[5:0]] & {8{~(p1_actual_index__51_comb[6] | p1_actual_index__51_comb[7])}}) == 8'h00;
  assign p1_eq_8834_comb = (p1_flat_comb[p1_actual_index__52_comb > 8'h3f ? 6'h3f : p1_actual_index__52_comb[5:0]] & {8{~(p1_add_8424_comb[4] | p1_add_8424_comb[5])}}) == 8'h00;
  assign p1_eq_8835_comb = (p1_flat_comb[p1_actual_index__53_comb > 8'h3f ? 6'h3f : p1_actual_index__53_comb[5:0]] & {8{~(p1_actual_index__53_comb[6] | p1_actual_index__53_comb[7])}}) == 8'h00;
  assign p1_eq_8836_comb = (p1_flat_comb[p1_actual_index__54_comb > 8'h3f ? 6'h3f : p1_actual_index__54_comb[5:0]] & {8{~(p1_add_8426_comb[5] | p1_add_8426_comb[6])}}) == 8'h00;
  assign p1_eq_8837_comb = (p1_flat_comb[p1_actual_index__55_comb > 8'h3f ? 6'h3f : p1_actual_index__55_comb[5:0]] & {8{~(p1_actual_index__55_comb[6] | p1_actual_index__55_comb[7])}}) == 8'h00;
  assign p1_eq_8838_comb = (p1_flat_comb[p1_actual_index__56_comb > 8'h3f ? 6'h3f : p1_actual_index__56_comb[5:0]] & {8{~(p1_add_8428_comb[3] | p1_add_8428_comb[4])}}) == 8'h00;
  assign p1_eq_8839_comb = (p1_flat_comb[p1_actual_index__57_comb > 8'h3f ? 6'h3f : p1_actual_index__57_comb[5:0]] & {8{~(p1_actual_index__57_comb[6] | p1_actual_index__57_comb[7])}}) == 8'h00;
  assign p1_eq_8840_comb = (p1_flat_comb[p1_actual_index__58_comb > 8'h3f ? 6'h3f : p1_actual_index__58_comb[5:0]] & {8{~(p1_add_8430_comb[5] | p1_add_8430_comb[6])}}) == 8'h00;
  assign p1_eq_8841_comb = (p1_flat_comb[p1_actual_index__59_comb > 8'h3f ? 6'h3f : p1_actual_index__59_comb[5:0]] & {8{~(p1_actual_index__59_comb[6] | p1_actual_index__59_comb[7])}}) == 8'h00;
  assign p1_eq_8842_comb = (p1_flat_comb[p1_actual_index__60_comb > 8'h3f ? 6'h3f : p1_actual_index__60_comb[5:0]] & {8{~(p1_add_8432_comb[4] | p1_add_8432_comb[5])}}) == 8'h00;
  assign p1_eq_8843_comb = (p1_flat_comb[p1_actual_index__61_comb > 8'h3f ? 6'h3f : p1_actual_index__61_comb[5:0]] & {8{~(p1_actual_index__61_comb[6] | p1_actual_index__61_comb[7])}}) == 8'h00;
  assign p1_eq_8844_comb = (p1_flat_comb[p1_actual_index__62_comb > 8'h3f ? 6'h3f : p1_actual_index__62_comb[5:0]] & {8{~(p1_add_8434_comb[5] | p1_add_8434_comb[6])}}) == 8'h00;
  assign p1_value_comb = p0_matrix[3'h0][3'h0];

  // Registers for pipe stage 1:
  reg p1_is_luminance;
  reg [7:0] p1_and_8226;
  reg [7:0] p1_and_8234;
  reg p1_eq_8237;
  reg [7:0] p1_and_8238;
  reg p1_ne_8246;
  reg [1:0] p1_concat_8247;
  reg p1_eq_8248;
  reg [7:0] p1_and_8263;
  reg [7:0] p1_and_8270;
  reg [7:0] p1_and_8277;
  reg [7:0] p1_and_8278;
  reg [7:0] p1_and_8299;
  reg [7:0] p1_and_8308;
  reg [7:0] p1_and_8315;
  reg [7:0] p1_and_8324;
  reg [7:0] p1_and_8329;
  reg [7:0] p1_and_8334;
  reg [7:0] p1_and_8335;
  reg [7:0] p1_and_8336;
  reg p1_eq_8797;
  reg p1_eq_8798;
  reg p1_eq_8799;
  reg p1_eq_8800;
  reg p1_eq_8801;
  reg p1_eq_8802;
  reg p1_eq_8803;
  reg p1_eq_8804;
  reg p1_eq_8805;
  reg p1_eq_8806;
  reg p1_eq_8807;
  reg p1_eq_8808;
  reg p1_eq_8809;
  reg p1_eq_8810;
  reg p1_eq_8811;
  reg p1_eq_8812;
  reg p1_eq_8813;
  reg p1_eq_8814;
  reg p1_eq_8815;
  reg p1_eq_8816;
  reg p1_eq_8817;
  reg p1_eq_8818;
  reg p1_eq_8819;
  reg p1_eq_8820;
  reg p1_eq_8821;
  reg p1_eq_8822;
  reg p1_eq_8823;
  reg p1_eq_8824;
  reg p1_eq_8825;
  reg p1_eq_8826;
  reg p1_eq_8827;
  reg p1_eq_8828;
  reg p1_eq_8829;
  reg p1_eq_8830;
  reg p1_eq_8831;
  reg p1_eq_8832;
  reg p1_eq_8833;
  reg p1_eq_8834;
  reg p1_eq_8835;
  reg p1_eq_8836;
  reg p1_eq_8837;
  reg p1_eq_8838;
  reg p1_eq_8839;
  reg p1_eq_8840;
  reg p1_eq_8841;
  reg p1_eq_8842;
  reg p1_eq_8843;
  reg p1_eq_8844;
  reg [7:0] p1_value;
  always @ (posedge clk) begin
    p1_is_luminance <= p0_is_luminance;
    p1_and_8226 <= p1_and_8226_comb;
    p1_and_8234 <= p1_and_8234_comb;
    p1_eq_8237 <= p1_eq_8237_comb;
    p1_and_8238 <= p1_and_8238_comb;
    p1_ne_8246 <= p1_ne_8246_comb;
    p1_concat_8247 <= p1_concat_8247_comb;
    p1_eq_8248 <= p1_eq_8248_comb;
    p1_and_8263 <= p1_and_8263_comb;
    p1_and_8270 <= p1_and_8270_comb;
    p1_and_8277 <= p1_and_8277_comb;
    p1_and_8278 <= p1_and_8278_comb;
    p1_and_8299 <= p1_and_8299_comb;
    p1_and_8308 <= p1_and_8308_comb;
    p1_and_8315 <= p1_and_8315_comb;
    p1_and_8324 <= p1_and_8324_comb;
    p1_and_8329 <= p1_and_8329_comb;
    p1_and_8334 <= p1_and_8334_comb;
    p1_and_8335 <= p1_and_8335_comb;
    p1_and_8336 <= p1_and_8336_comb;
    p1_eq_8797 <= p1_eq_8797_comb;
    p1_eq_8798 <= p1_eq_8798_comb;
    p1_eq_8799 <= p1_eq_8799_comb;
    p1_eq_8800 <= p1_eq_8800_comb;
    p1_eq_8801 <= p1_eq_8801_comb;
    p1_eq_8802 <= p1_eq_8802_comb;
    p1_eq_8803 <= p1_eq_8803_comb;
    p1_eq_8804 <= p1_eq_8804_comb;
    p1_eq_8805 <= p1_eq_8805_comb;
    p1_eq_8806 <= p1_eq_8806_comb;
    p1_eq_8807 <= p1_eq_8807_comb;
    p1_eq_8808 <= p1_eq_8808_comb;
    p1_eq_8809 <= p1_eq_8809_comb;
    p1_eq_8810 <= p1_eq_8810_comb;
    p1_eq_8811 <= p1_eq_8811_comb;
    p1_eq_8812 <= p1_eq_8812_comb;
    p1_eq_8813 <= p1_eq_8813_comb;
    p1_eq_8814 <= p1_eq_8814_comb;
    p1_eq_8815 <= p1_eq_8815_comb;
    p1_eq_8816 <= p1_eq_8816_comb;
    p1_eq_8817 <= p1_eq_8817_comb;
    p1_eq_8818 <= p1_eq_8818_comb;
    p1_eq_8819 <= p1_eq_8819_comb;
    p1_eq_8820 <= p1_eq_8820_comb;
    p1_eq_8821 <= p1_eq_8821_comb;
    p1_eq_8822 <= p1_eq_8822_comb;
    p1_eq_8823 <= p1_eq_8823_comb;
    p1_eq_8824 <= p1_eq_8824_comb;
    p1_eq_8825 <= p1_eq_8825_comb;
    p1_eq_8826 <= p1_eq_8826_comb;
    p1_eq_8827 <= p1_eq_8827_comb;
    p1_eq_8828 <= p1_eq_8828_comb;
    p1_eq_8829 <= p1_eq_8829_comb;
    p1_eq_8830 <= p1_eq_8830_comb;
    p1_eq_8831 <= p1_eq_8831_comb;
    p1_eq_8832 <= p1_eq_8832_comb;
    p1_eq_8833 <= p1_eq_8833_comb;
    p1_eq_8834 <= p1_eq_8834_comb;
    p1_eq_8835 <= p1_eq_8835_comb;
    p1_eq_8836 <= p1_eq_8836_comb;
    p1_eq_8837 <= p1_eq_8837_comb;
    p1_eq_8838 <= p1_eq_8838_comb;
    p1_eq_8839 <= p1_eq_8839_comb;
    p1_eq_8840 <= p1_eq_8840_comb;
    p1_eq_8841 <= p1_eq_8841_comb;
    p1_eq_8842 <= p1_eq_8842_comb;
    p1_eq_8843 <= p1_eq_8843_comb;
    p1_eq_8844 <= p1_eq_8844_comb;
    p1_value <= p1_value_comb;
  end

  // ===== Pipe stage 2:
  wire [1:0] p2_idx_u8__1_squeezed_comb;
  wire p2_ne_8993_comb;
  wire p2_ne_8997_comb;
  wire p2_ne_9001_comb;
  wire p2_eq_9004_comb;
  wire [2:0] p2_sel_9005_comb;
  wire p2_ne_9011_comb;
  wire p2_ne_9015_comb;
  wire p2_ne_9019_comb;
  wire p2_ne_9032_comb;
  wire p2_ne_9033_comb;
  wire p2_ne_9031_comb;
  wire p2_ne_9027_comb;
  wire p2_ne_9023_comb;
  wire [3:0] p2_sel_9024_comb;
  wire p2_not_9034_comb;
  wire [3:0] p2_sel_9028_comb;
  wire p2_and_9046_comb;
  assign p2_idx_u8__1_squeezed_comb = 2'h1;
  assign p2_ne_8993_comb = p1_and_8263 != 8'h00;
  assign p2_ne_8997_comb = p1_and_8270 != 8'h00;
  assign p2_ne_9001_comb = p1_and_8277 != 8'h00;
  assign p2_eq_9004_comb = p1_and_8278 == 8'h00;
  assign p2_sel_9005_comb = p2_ne_9001_comb ? 3'h1 : (p2_ne_8997_comb ? 3'h2 : (p2_ne_8993_comb ? 3'h3 : {1'h1, (p1_ne_8246 ? p2_idx_u8__1_squeezed_comb : p1_concat_8247) & {2{p1_eq_8248}}}));
  assign p2_ne_9011_comb = p1_and_8299 != 8'h00;
  assign p2_ne_9015_comb = p1_and_8308 != 8'h00;
  assign p2_ne_9019_comb = p1_and_8315 != 8'h00;
  assign p2_ne_9032_comb = p1_and_8335 != 8'h00;
  assign p2_ne_9033_comb = p1_and_8336 != 8'h00;
  assign p2_ne_9031_comb = p1_and_8334 != 8'h00;
  assign p2_ne_9027_comb = p1_and_8329 != 8'h00;
  assign p2_ne_9023_comb = p1_and_8324 != 8'h00;
  assign p2_sel_9024_comb = p2_ne_9019_comb ? 4'h5 : (p2_ne_9015_comb ? 4'h6 : (p2_ne_9011_comb ? 4'h7 : {1'h1, p2_sel_9005_comb & {3{p2_eq_9004_comb}}}));
  assign p2_not_9034_comb = ~p2_ne_9032_comb;
  assign p2_sel_9028_comb = p2_ne_9023_comb ? 4'h4 : p2_sel_9024_comb;
  assign p2_and_9046_comb = p2_not_9034_comb & ~p2_ne_9033_comb & ~p2_ne_9031_comb & ~p2_ne_9027_comb & ~p2_ne_9023_comb & ~p2_ne_9019_comb & ~p2_ne_9015_comb & ~p2_ne_9011_comb & p2_eq_9004_comb & ~p2_ne_9001_comb & ~p2_ne_8997_comb & ~p2_ne_8993_comb & p1_eq_8248 & ~p1_ne_8246 & p1_eq_8237 & p1_eq_8797 & p1_eq_8798 & p1_eq_8799 & p1_eq_8800 & p1_eq_8801 & p1_eq_8802 & p1_eq_8803 & p1_eq_8804 & p1_eq_8805 & p1_eq_8806 & p1_eq_8807 & p1_eq_8808 & p1_eq_8809 & p1_eq_8810 & p1_eq_8811 & p1_eq_8812 & p1_eq_8813 & p1_eq_8814 & p1_eq_8815 & p1_eq_8816 & p1_eq_8817 & p1_eq_8818 & p1_eq_8819 & p1_eq_8820 & p1_eq_8821 & p1_eq_8822 & p1_eq_8823 & p1_eq_8824 & p1_eq_8825 & p1_eq_8826 & p1_eq_8827 & p1_eq_8828 & p1_eq_8829 & p1_eq_8830 & p1_eq_8831 & p1_eq_8832 & p1_eq_8833 & p1_eq_8834 & p1_eq_8835 & p1_eq_8836 & p1_eq_8837 & p1_eq_8838 & p1_eq_8839 & p1_eq_8840 & p1_eq_8841 & p1_eq_8842 & p1_eq_8843 & p1_eq_8844;

  // Registers for pipe stage 2:
  reg p2_is_luminance;
  reg [7:0] p2_and_8226;
  reg [7:0] p2_and_8234;
  reg [7:0] p2_and_8238;
  reg [7:0] p2_and_8263;
  reg [7:0] p2_and_8270;
  reg [7:0] p2_and_8277;
  reg [7:0] p2_and_8278;
  reg [7:0] p2_and_8299;
  reg [7:0] p2_and_8308;
  reg [7:0] p2_and_8315;
  reg [7:0] p2_and_8324;
  reg [7:0] p2_and_8329;
  reg [7:0] p2_and_8334;
  reg p2_ne_9027;
  reg [3:0] p2_sel_9028;
  reg [7:0] p2_and_8335;
  reg [7:0] p2_and_8336;
  reg p2_ne_9031;
  reg p2_ne_9032;
  reg p2_ne_9033;
  reg p2_not_9034;
  reg p2_and_9046;
  reg [7:0] p2_value;
  always @ (posedge clk) begin
    p2_is_luminance <= p1_is_luminance;
    p2_and_8226 <= p1_and_8226;
    p2_and_8234 <= p1_and_8234;
    p2_and_8238 <= p1_and_8238;
    p2_and_8263 <= p1_and_8263;
    p2_and_8270 <= p1_and_8270;
    p2_and_8277 <= p1_and_8277;
    p2_and_8278 <= p1_and_8278;
    p2_and_8299 <= p1_and_8299;
    p2_and_8308 <= p1_and_8308;
    p2_and_8315 <= p1_and_8315;
    p2_and_8324 <= p1_and_8324;
    p2_and_8329 <= p1_and_8329;
    p2_and_8334 <= p1_and_8334;
    p2_ne_9027 <= p2_ne_9027_comb;
    p2_sel_9028 <= p2_sel_9028_comb;
    p2_and_8335 <= p1_and_8335;
    p2_and_8336 <= p1_and_8336;
    p2_ne_9031 <= p2_ne_9031_comb;
    p2_ne_9032 <= p2_ne_9032_comb;
    p2_ne_9033 <= p2_ne_9033_comb;
    p2_not_9034 <= p2_not_9034_comb;
    p2_and_9046 <= p2_and_9046_comb;
    p2_value <= p1_value;
  end

  // ===== Pipe stage 3:
  wire [3:0] p3_sel_9100_comb;
  wire [3:0] p3_run_comb;
  wire [7:0] p3_value__1_comb;
  wire [1:0] p3_idx_u8__1_squeezed__1_comb;
  wire [1:0] p3_idx_u8__2_squeezed_comb;
  wire [1:0] p3_idx_u8__3_squeezed_comb;
  wire p3_eq_9133_comb;
  wire p3_eq_9130_comb;
  wire [7:0] p3_flipped__1_comb;
  wire [2:0] p3_idx_u8__4_squeezed__1_comb;
  wire [7:0] p3_code_list__1_comb;
  wire [2:0] p3_sel_9122_comb;
  wire [2:0] p3_idx_u8__5_squeezed__1_comb;
  wire p3_or_reduce_9125_comb;
  wire [2:0] p3_sel_9126_comb;
  wire p3_or_reduce_9127_comb;
  wire p3_bit_slice_9129_comb;
  wire p3_not_9131_comb;
  wire p3_or_9134_comb;
  wire [7:0] p3_sel_9144_comb;
  wire [3:0] p3_sel_9145_comb;
  assign p3_sel_9100_comb = p2_ne_9033 ? 4'h1 : (p2_ne_9031 ? 4'h2 : (p2_ne_9027 ? 4'h3 : p2_sel_9028));
  assign p3_run_comb = p3_sel_9100_comb & {4{p2_not_9034}};
  assign p3_value__1_comb = p3_run_comb == 4'h0 ? p2_and_8335 : (p3_run_comb == 4'h1 ? p2_and_8336 : (p3_run_comb == 4'h2 ? p2_and_8334 : (p3_run_comb == 4'h3 ? p2_and_8329 : (p3_run_comb == 4'h4 ? p2_and_8324 : (p3_run_comb == 4'h5 ? p2_and_8315 : (p3_run_comb == 4'h6 ? p2_and_8308 : (p3_run_comb == 4'h7 ? p2_and_8299 : (p3_run_comb == 4'h8 ? p2_and_8278 : (p3_run_comb == 4'h9 ? p2_and_8277 : (p3_run_comb == 4'ha ? p2_and_8270 : (p3_run_comb == 4'hb ? p2_and_8263 : (p3_run_comb == 4'hc ? p2_and_8238 : (p3_run_comb == 4'hd ? p2_and_8234 : (p3_run_comb == 4'he ? p2_and_8226 : 8'h00))))))))))))));
  assign p3_idx_u8__1_squeezed__1_comb = 2'h1;
  assign p3_idx_u8__2_squeezed_comb = 2'h2;
  assign p3_idx_u8__3_squeezed_comb = 2'h3;
  assign p3_eq_9133_comb = p3_run_comb == 4'hf;
  assign p3_eq_9130_comb = p3_value__1_comb == 8'h00;
  assign p3_flipped__1_comb = 8'hff;
  assign p3_idx_u8__4_squeezed__1_comb = 3'h4;
  assign p3_code_list__1_comb = p3_eq_9130_comb ? p3_flipped__1_comb : p3_value__1_comb;
  assign p3_sel_9122_comb = |p3_value__1_comb[7:3] ? p3_idx_u8__4_squeezed__1_comb : {1'h0, |p3_value__1_comb[7:2] ? p3_idx_u8__3_squeezed_comb : (|p3_value__1_comb[7:1] ? p3_idx_u8__2_squeezed_comb : p3_idx_u8__1_squeezed__1_comb)};
  assign p3_idx_u8__5_squeezed__1_comb = 3'h5;
  assign p3_or_reduce_9125_comb = |p3_value__1_comb[7:5];
  assign p3_sel_9126_comb = |p3_value__1_comb[7:4] ? p3_idx_u8__5_squeezed__1_comb : p3_sel_9122_comb;
  assign p3_or_reduce_9127_comb = |p3_value__1_comb[7:6];
  assign p3_bit_slice_9129_comb = p3_value__1_comb[7];
  assign p3_not_9131_comb = ~p3_eq_9130_comb;
  assign p3_or_9134_comb = p2_and_9046 | p3_eq_9133_comb;
  assign p3_sel_9144_comb = p2_and_9046 ? p2_value : p3_code_list__1_comb & {8{~p3_eq_9133_comb}};
  assign p3_sel_9145_comb = p2_and_9046 ? 4'hf : p3_sel_9100_comb & {4{~(p3_eq_9133_comb | p2_ne_9032)}};

  // Registers for pipe stage 3:
  reg p3_is_luminance;
  reg [3:0] p3_run;
  reg p3_or_reduce_9125;
  reg [2:0] p3_sel_9126;
  reg p3_or_reduce_9127;
  reg p3_bit_slice_9129;
  reg p3_not_9131;
  reg p3_or_9134;
  reg [7:0] p3_sel_9144;
  reg [3:0] p3_sel_9145;
  always @ (posedge clk) begin
    p3_is_luminance <= p2_is_luminance;
    p3_run <= p3_run_comb;
    p3_or_reduce_9125 <= p3_or_reduce_9125_comb;
    p3_sel_9126 <= p3_sel_9126_comb;
    p3_or_reduce_9127 <= p3_or_reduce_9127_comb;
    p3_bit_slice_9129 <= p3_bit_slice_9129_comb;
    p3_not_9131 <= p3_not_9131_comb;
    p3_or_9134 <= p3_or_9134_comb;
    p3_sel_9144 <= p3_sel_9144_comb;
    p3_sel_9145 <= p3_sel_9145_comb;
  end

  // ===== Pipe stage 4:
  wire [2:0] p4_idx_u8__6_squeezed__1_comb;
  wire [2:0] p4_idx_u8__7_squeezed__1_comb;
  wire [3:0] p4_idx_u8__8_squeezed_comb;
  wire [7:0] p4_size__1_comb;
  wire [7:0] p4_run_size_str_u8_comb;
  wire [4:0] p4_huffman_length_squeezed_comb;
  wire [4:0] p4_idx_u8__2_squeezed__1_comb;
  wire [15:0] p4_huffman_code_full_comb;
  wire [35:0] p4_tuple_9198_comb;
  assign p4_idx_u8__6_squeezed__1_comb = 3'h6;
  assign p4_idx_u8__7_squeezed__1_comb = 3'h7;
  assign p4_idx_u8__8_squeezed_comb = 4'h8;
  assign p4_size__1_comb = {4'h0, p3_bit_slice_9129 ? p4_idx_u8__8_squeezed_comb : {1'h0, p3_or_reduce_9127 ? p4_idx_u8__7_squeezed__1_comb : (p3_or_reduce_9125 ? p4_idx_u8__6_squeezed__1_comb : p3_sel_9126)}} & {8{p3_not_9131}};
  assign p4_run_size_str_u8_comb = {p3_run, 4'h0} | p4_size__1_comb;
  assign p4_huffman_length_squeezed_comb = p3_is_luminance ? literal_9182[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_9180[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_idx_u8__2_squeezed__1_comb = 5'h02;
  assign p4_huffman_code_full_comb = p3_is_luminance ? literal_9184[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_9183[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_tuple_9198_comb = {p4_huffman_code_full_comb & {16{~p3_or_9134}}, {3'h0, p3_or_9134 ? p4_idx_u8__2_squeezed__1_comb : p4_huffman_length_squeezed_comb}, p3_sel_9144, p3_sel_9145};

  // Registers for pipe stage 4:
  reg [35:0] p4_tuple_9198;
  always @ (posedge clk) begin
    p4_tuple_9198 <= p4_tuple_9198_comb;
  end
  assign out = p4_tuple_9198;
endmodule
