module Huffman_ACenc(
  input wire clk,
  input wire [511:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [35:0] out
);
  wire [4:0] literal_9174[0:251];
  assign literal_9174[0] = 5'h02;
  assign literal_9174[1] = 5'h02;
  assign literal_9174[2] = 5'h03;
  assign literal_9174[3] = 5'h04;
  assign literal_9174[4] = 5'h05;
  assign literal_9174[5] = 5'h07;
  assign literal_9174[6] = 5'h08;
  assign literal_9174[7] = 5'h0e;
  assign literal_9174[8] = 5'h10;
  assign literal_9174[9] = 5'h10;
  assign literal_9174[10] = 5'h10;
  assign literal_9174[11] = 5'h00;
  assign literal_9174[12] = 5'h00;
  assign literal_9174[13] = 5'h00;
  assign literal_9174[14] = 5'h00;
  assign literal_9174[15] = 5'h00;
  assign literal_9174[16] = 5'h00;
  assign literal_9174[17] = 5'h03;
  assign literal_9174[18] = 5'h06;
  assign literal_9174[19] = 5'h07;
  assign literal_9174[20] = 5'h09;
  assign literal_9174[21] = 5'h0b;
  assign literal_9174[22] = 5'h0d;
  assign literal_9174[23] = 5'h10;
  assign literal_9174[24] = 5'h10;
  assign literal_9174[25] = 5'h10;
  assign literal_9174[26] = 5'h10;
  assign literal_9174[27] = 5'h00;
  assign literal_9174[28] = 5'h00;
  assign literal_9174[29] = 5'h00;
  assign literal_9174[30] = 5'h00;
  assign literal_9174[31] = 5'h00;
  assign literal_9174[32] = 5'h00;
  assign literal_9174[33] = 5'h05;
  assign literal_9174[34] = 5'h07;
  assign literal_9174[35] = 5'h0a;
  assign literal_9174[36] = 5'h0c;
  assign literal_9174[37] = 5'h0d;
  assign literal_9174[38] = 5'h10;
  assign literal_9174[39] = 5'h10;
  assign literal_9174[40] = 5'h10;
  assign literal_9174[41] = 5'h10;
  assign literal_9174[42] = 5'h10;
  assign literal_9174[43] = 5'h00;
  assign literal_9174[44] = 5'h00;
  assign literal_9174[45] = 5'h00;
  assign literal_9174[46] = 5'h00;
  assign literal_9174[47] = 5'h00;
  assign literal_9174[48] = 5'h00;
  assign literal_9174[49] = 5'h06;
  assign literal_9174[50] = 5'h08;
  assign literal_9174[51] = 5'h0b;
  assign literal_9174[52] = 5'h0c;
  assign literal_9174[53] = 5'h0f;
  assign literal_9174[54] = 5'h10;
  assign literal_9174[55] = 5'h10;
  assign literal_9174[56] = 5'h10;
  assign literal_9174[57] = 5'h10;
  assign literal_9174[58] = 5'h10;
  assign literal_9174[59] = 5'h00;
  assign literal_9174[60] = 5'h00;
  assign literal_9174[61] = 5'h00;
  assign literal_9174[62] = 5'h00;
  assign literal_9174[63] = 5'h00;
  assign literal_9174[64] = 5'h00;
  assign literal_9174[65] = 5'h06;
  assign literal_9174[66] = 5'h0a;
  assign literal_9174[67] = 5'h0c;
  assign literal_9174[68] = 5'h0f;
  assign literal_9174[69] = 5'h10;
  assign literal_9174[70] = 5'h10;
  assign literal_9174[71] = 5'h10;
  assign literal_9174[72] = 5'h10;
  assign literal_9174[73] = 5'h10;
  assign literal_9174[74] = 5'h10;
  assign literal_9174[75] = 5'h00;
  assign literal_9174[76] = 5'h00;
  assign literal_9174[77] = 5'h00;
  assign literal_9174[78] = 5'h00;
  assign literal_9174[79] = 5'h00;
  assign literal_9174[80] = 5'h00;
  assign literal_9174[81] = 5'h07;
  assign literal_9174[82] = 5'h0b;
  assign literal_9174[83] = 5'h0d;
  assign literal_9174[84] = 5'h10;
  assign literal_9174[85] = 5'h10;
  assign literal_9174[86] = 5'h10;
  assign literal_9174[87] = 5'h10;
  assign literal_9174[88] = 5'h10;
  assign literal_9174[89] = 5'h10;
  assign literal_9174[90] = 5'h10;
  assign literal_9174[91] = 5'h00;
  assign literal_9174[92] = 5'h00;
  assign literal_9174[93] = 5'h00;
  assign literal_9174[94] = 5'h00;
  assign literal_9174[95] = 5'h00;
  assign literal_9174[96] = 5'h00;
  assign literal_9174[97] = 5'h07;
  assign literal_9174[98] = 5'h0b;
  assign literal_9174[99] = 5'h0d;
  assign literal_9174[100] = 5'h10;
  assign literal_9174[101] = 5'h10;
  assign literal_9174[102] = 5'h10;
  assign literal_9174[103] = 5'h10;
  assign literal_9174[104] = 5'h10;
  assign literal_9174[105] = 5'h10;
  assign literal_9174[106] = 5'h10;
  assign literal_9174[107] = 5'h00;
  assign literal_9174[108] = 5'h00;
  assign literal_9174[109] = 5'h00;
  assign literal_9174[110] = 5'h00;
  assign literal_9174[111] = 5'h00;
  assign literal_9174[112] = 5'h00;
  assign literal_9174[113] = 5'h08;
  assign literal_9174[114] = 5'h0b;
  assign literal_9174[115] = 5'h0e;
  assign literal_9174[116] = 5'h10;
  assign literal_9174[117] = 5'h10;
  assign literal_9174[118] = 5'h10;
  assign literal_9174[119] = 5'h10;
  assign literal_9174[120] = 5'h10;
  assign literal_9174[121] = 5'h10;
  assign literal_9174[122] = 5'h10;
  assign literal_9174[123] = 5'h00;
  assign literal_9174[124] = 5'h00;
  assign literal_9174[125] = 5'h00;
  assign literal_9174[126] = 5'h00;
  assign literal_9174[127] = 5'h00;
  assign literal_9174[128] = 5'h00;
  assign literal_9174[129] = 5'h08;
  assign literal_9174[130] = 5'h0c;
  assign literal_9174[131] = 5'h10;
  assign literal_9174[132] = 5'h10;
  assign literal_9174[133] = 5'h10;
  assign literal_9174[134] = 5'h10;
  assign literal_9174[135] = 5'h10;
  assign literal_9174[136] = 5'h10;
  assign literal_9174[137] = 5'h10;
  assign literal_9174[138] = 5'h10;
  assign literal_9174[139] = 5'h00;
  assign literal_9174[140] = 5'h00;
  assign literal_9174[141] = 5'h00;
  assign literal_9174[142] = 5'h00;
  assign literal_9174[143] = 5'h00;
  assign literal_9174[144] = 5'h00;
  assign literal_9174[145] = 5'h08;
  assign literal_9174[146] = 5'h0d;
  assign literal_9174[147] = 5'h10;
  assign literal_9174[148] = 5'h10;
  assign literal_9174[149] = 5'h10;
  assign literal_9174[150] = 5'h10;
  assign literal_9174[151] = 5'h10;
  assign literal_9174[152] = 5'h10;
  assign literal_9174[153] = 5'h10;
  assign literal_9174[154] = 5'h10;
  assign literal_9174[155] = 5'h00;
  assign literal_9174[156] = 5'h00;
  assign literal_9174[157] = 5'h00;
  assign literal_9174[158] = 5'h00;
  assign literal_9174[159] = 5'h00;
  assign literal_9174[160] = 5'h00;
  assign literal_9174[161] = 5'h09;
  assign literal_9174[162] = 5'h0d;
  assign literal_9174[163] = 5'h10;
  assign literal_9174[164] = 5'h10;
  assign literal_9174[165] = 5'h10;
  assign literal_9174[166] = 5'h10;
  assign literal_9174[167] = 5'h10;
  assign literal_9174[168] = 5'h10;
  assign literal_9174[169] = 5'h10;
  assign literal_9174[170] = 5'h10;
  assign literal_9174[171] = 5'h00;
  assign literal_9174[172] = 5'h00;
  assign literal_9174[173] = 5'h00;
  assign literal_9174[174] = 5'h00;
  assign literal_9174[175] = 5'h00;
  assign literal_9174[176] = 5'h00;
  assign literal_9174[177] = 5'h09;
  assign literal_9174[178] = 5'h0d;
  assign literal_9174[179] = 5'h10;
  assign literal_9174[180] = 5'h10;
  assign literal_9174[181] = 5'h10;
  assign literal_9174[182] = 5'h10;
  assign literal_9174[183] = 5'h10;
  assign literal_9174[184] = 5'h10;
  assign literal_9174[185] = 5'h10;
  assign literal_9174[186] = 5'h10;
  assign literal_9174[187] = 5'h00;
  assign literal_9174[188] = 5'h00;
  assign literal_9174[189] = 5'h00;
  assign literal_9174[190] = 5'h00;
  assign literal_9174[191] = 5'h00;
  assign literal_9174[192] = 5'h00;
  assign literal_9174[193] = 5'h0a;
  assign literal_9174[194] = 5'h0d;
  assign literal_9174[195] = 5'h10;
  assign literal_9174[196] = 5'h10;
  assign literal_9174[197] = 5'h10;
  assign literal_9174[198] = 5'h10;
  assign literal_9174[199] = 5'h10;
  assign literal_9174[200] = 5'h10;
  assign literal_9174[201] = 5'h10;
  assign literal_9174[202] = 5'h10;
  assign literal_9174[203] = 5'h00;
  assign literal_9174[204] = 5'h00;
  assign literal_9174[205] = 5'h00;
  assign literal_9174[206] = 5'h00;
  assign literal_9174[207] = 5'h00;
  assign literal_9174[208] = 5'h00;
  assign literal_9174[209] = 5'h0a;
  assign literal_9174[210] = 5'h0e;
  assign literal_9174[211] = 5'h10;
  assign literal_9174[212] = 5'h10;
  assign literal_9174[213] = 5'h10;
  assign literal_9174[214] = 5'h10;
  assign literal_9174[215] = 5'h10;
  assign literal_9174[216] = 5'h10;
  assign literal_9174[217] = 5'h10;
  assign literal_9174[218] = 5'h10;
  assign literal_9174[219] = 5'h00;
  assign literal_9174[220] = 5'h00;
  assign literal_9174[221] = 5'h00;
  assign literal_9174[222] = 5'h00;
  assign literal_9174[223] = 5'h00;
  assign literal_9174[224] = 5'h00;
  assign literal_9174[225] = 5'h0a;
  assign literal_9174[226] = 5'h0f;
  assign literal_9174[227] = 5'h10;
  assign literal_9174[228] = 5'h10;
  assign literal_9174[229] = 5'h10;
  assign literal_9174[230] = 5'h10;
  assign literal_9174[231] = 5'h10;
  assign literal_9174[232] = 5'h10;
  assign literal_9174[233] = 5'h10;
  assign literal_9174[234] = 5'h10;
  assign literal_9174[235] = 5'h00;
  assign literal_9174[236] = 5'h00;
  assign literal_9174[237] = 5'h00;
  assign literal_9174[238] = 5'h00;
  assign literal_9174[239] = 5'h00;
  assign literal_9174[240] = 5'h09;
  assign literal_9174[241] = 5'h0b;
  assign literal_9174[242] = 5'h10;
  assign literal_9174[243] = 5'h10;
  assign literal_9174[244] = 5'h10;
  assign literal_9174[245] = 5'h10;
  assign literal_9174[246] = 5'h10;
  assign literal_9174[247] = 5'h10;
  assign literal_9174[248] = 5'h10;
  assign literal_9174[249] = 5'h10;
  assign literal_9174[250] = 5'h10;
  assign literal_9174[251] = 5'h00;
  wire [4:0] literal_9176[0:251];
  assign literal_9176[0] = 5'h04;
  assign literal_9176[1] = 5'h02;
  assign literal_9176[2] = 5'h02;
  assign literal_9176[3] = 5'h03;
  assign literal_9176[4] = 5'h04;
  assign literal_9176[5] = 5'h05;
  assign literal_9176[6] = 5'h07;
  assign literal_9176[7] = 5'h09;
  assign literal_9176[8] = 5'h10;
  assign literal_9176[9] = 5'h10;
  assign literal_9176[10] = 5'h10;
  assign literal_9176[11] = 5'h00;
  assign literal_9176[12] = 5'h00;
  assign literal_9176[13] = 5'h00;
  assign literal_9176[14] = 5'h00;
  assign literal_9176[15] = 5'h00;
  assign literal_9176[16] = 5'h00;
  assign literal_9176[17] = 5'h04;
  assign literal_9176[18] = 5'h05;
  assign literal_9176[19] = 5'h07;
  assign literal_9176[20] = 5'h09;
  assign literal_9176[21] = 5'h0a;
  assign literal_9176[22] = 5'h0b;
  assign literal_9176[23] = 5'h10;
  assign literal_9176[24] = 5'h10;
  assign literal_9176[25] = 5'h10;
  assign literal_9176[26] = 5'h10;
  assign literal_9176[27] = 5'h00;
  assign literal_9176[28] = 5'h00;
  assign literal_9176[29] = 5'h00;
  assign literal_9176[30] = 5'h00;
  assign literal_9176[31] = 5'h00;
  assign literal_9176[32] = 5'h00;
  assign literal_9176[33] = 5'h05;
  assign literal_9176[34] = 5'h08;
  assign literal_9176[35] = 5'h0a;
  assign literal_9176[36] = 5'h0c;
  assign literal_9176[37] = 5'h0e;
  assign literal_9176[38] = 5'h10;
  assign literal_9176[39] = 5'h10;
  assign literal_9176[40] = 5'h10;
  assign literal_9176[41] = 5'h10;
  assign literal_9176[42] = 5'h10;
  assign literal_9176[43] = 5'h00;
  assign literal_9176[44] = 5'h00;
  assign literal_9176[45] = 5'h00;
  assign literal_9176[46] = 5'h00;
  assign literal_9176[47] = 5'h00;
  assign literal_9176[48] = 5'h00;
  assign literal_9176[49] = 5'h06;
  assign literal_9176[50] = 5'h09;
  assign literal_9176[51] = 5'h0b;
  assign literal_9176[52] = 5'h0e;
  assign literal_9176[53] = 5'h10;
  assign literal_9176[54] = 5'h10;
  assign literal_9176[55] = 5'h10;
  assign literal_9176[56] = 5'h10;
  assign literal_9176[57] = 5'h10;
  assign literal_9176[58] = 5'h10;
  assign literal_9176[59] = 5'h00;
  assign literal_9176[60] = 5'h00;
  assign literal_9176[61] = 5'h00;
  assign literal_9176[62] = 5'h00;
  assign literal_9176[63] = 5'h00;
  assign literal_9176[64] = 5'h00;
  assign literal_9176[65] = 5'h06;
  assign literal_9176[66] = 5'h0a;
  assign literal_9176[67] = 5'h0e;
  assign literal_9176[68] = 5'h10;
  assign literal_9176[69] = 5'h10;
  assign literal_9176[70] = 5'h10;
  assign literal_9176[71] = 5'h10;
  assign literal_9176[72] = 5'h10;
  assign literal_9176[73] = 5'h10;
  assign literal_9176[74] = 5'h10;
  assign literal_9176[75] = 5'h00;
  assign literal_9176[76] = 5'h00;
  assign literal_9176[77] = 5'h00;
  assign literal_9176[78] = 5'h00;
  assign literal_9176[79] = 5'h00;
  assign literal_9176[80] = 5'h00;
  assign literal_9176[81] = 5'h07;
  assign literal_9176[82] = 5'h0a;
  assign literal_9176[83] = 5'h0e;
  assign literal_9176[84] = 5'h10;
  assign literal_9176[85] = 5'h10;
  assign literal_9176[86] = 5'h10;
  assign literal_9176[87] = 5'h10;
  assign literal_9176[88] = 5'h10;
  assign literal_9176[89] = 5'h10;
  assign literal_9176[90] = 5'h10;
  assign literal_9176[91] = 5'h00;
  assign literal_9176[92] = 5'h00;
  assign literal_9176[93] = 5'h00;
  assign literal_9176[94] = 5'h00;
  assign literal_9176[95] = 5'h00;
  assign literal_9176[96] = 5'h00;
  assign literal_9176[97] = 5'h07;
  assign literal_9176[98] = 5'h0c;
  assign literal_9176[99] = 5'h0f;
  assign literal_9176[100] = 5'h10;
  assign literal_9176[101] = 5'h10;
  assign literal_9176[102] = 5'h10;
  assign literal_9176[103] = 5'h10;
  assign literal_9176[104] = 5'h10;
  assign literal_9176[105] = 5'h10;
  assign literal_9176[106] = 5'h10;
  assign literal_9176[107] = 5'h00;
  assign literal_9176[108] = 5'h00;
  assign literal_9176[109] = 5'h00;
  assign literal_9176[110] = 5'h00;
  assign literal_9176[111] = 5'h00;
  assign literal_9176[112] = 5'h00;
  assign literal_9176[113] = 5'h08;
  assign literal_9176[114] = 5'h0c;
  assign literal_9176[115] = 5'h10;
  assign literal_9176[116] = 5'h10;
  assign literal_9176[117] = 5'h10;
  assign literal_9176[118] = 5'h10;
  assign literal_9176[119] = 5'h10;
  assign literal_9176[120] = 5'h10;
  assign literal_9176[121] = 5'h10;
  assign literal_9176[122] = 5'h10;
  assign literal_9176[123] = 5'h00;
  assign literal_9176[124] = 5'h00;
  assign literal_9176[125] = 5'h00;
  assign literal_9176[126] = 5'h00;
  assign literal_9176[127] = 5'h00;
  assign literal_9176[128] = 5'h00;
  assign literal_9176[129] = 5'h09;
  assign literal_9176[130] = 5'h0d;
  assign literal_9176[131] = 5'h10;
  assign literal_9176[132] = 5'h10;
  assign literal_9176[133] = 5'h10;
  assign literal_9176[134] = 5'h10;
  assign literal_9176[135] = 5'h10;
  assign literal_9176[136] = 5'h10;
  assign literal_9176[137] = 5'h10;
  assign literal_9176[138] = 5'h10;
  assign literal_9176[139] = 5'h00;
  assign literal_9176[140] = 5'h00;
  assign literal_9176[141] = 5'h00;
  assign literal_9176[142] = 5'h00;
  assign literal_9176[143] = 5'h00;
  assign literal_9176[144] = 5'h00;
  assign literal_9176[145] = 5'h09;
  assign literal_9176[146] = 5'h0e;
  assign literal_9176[147] = 5'h10;
  assign literal_9176[148] = 5'h10;
  assign literal_9176[149] = 5'h10;
  assign literal_9176[150] = 5'h10;
  assign literal_9176[151] = 5'h10;
  assign literal_9176[152] = 5'h10;
  assign literal_9176[153] = 5'h10;
  assign literal_9176[154] = 5'h10;
  assign literal_9176[155] = 5'h00;
  assign literal_9176[156] = 5'h00;
  assign literal_9176[157] = 5'h00;
  assign literal_9176[158] = 5'h00;
  assign literal_9176[159] = 5'h00;
  assign literal_9176[160] = 5'h00;
  assign literal_9176[161] = 5'h09;
  assign literal_9176[162] = 5'h0e;
  assign literal_9176[163] = 5'h10;
  assign literal_9176[164] = 5'h10;
  assign literal_9176[165] = 5'h10;
  assign literal_9176[166] = 5'h10;
  assign literal_9176[167] = 5'h10;
  assign literal_9176[168] = 5'h10;
  assign literal_9176[169] = 5'h10;
  assign literal_9176[170] = 5'h10;
  assign literal_9176[171] = 5'h00;
  assign literal_9176[172] = 5'h00;
  assign literal_9176[173] = 5'h00;
  assign literal_9176[174] = 5'h00;
  assign literal_9176[175] = 5'h00;
  assign literal_9176[176] = 5'h00;
  assign literal_9176[177] = 5'h0a;
  assign literal_9176[178] = 5'h0f;
  assign literal_9176[179] = 5'h10;
  assign literal_9176[180] = 5'h10;
  assign literal_9176[181] = 5'h10;
  assign literal_9176[182] = 5'h10;
  assign literal_9176[183] = 5'h10;
  assign literal_9176[184] = 5'h10;
  assign literal_9176[185] = 5'h10;
  assign literal_9176[186] = 5'h10;
  assign literal_9176[187] = 5'h00;
  assign literal_9176[188] = 5'h00;
  assign literal_9176[189] = 5'h00;
  assign literal_9176[190] = 5'h00;
  assign literal_9176[191] = 5'h00;
  assign literal_9176[192] = 5'h00;
  assign literal_9176[193] = 5'h0a;
  assign literal_9176[194] = 5'h10;
  assign literal_9176[195] = 5'h10;
  assign literal_9176[196] = 5'h10;
  assign literal_9176[197] = 5'h10;
  assign literal_9176[198] = 5'h10;
  assign literal_9176[199] = 5'h10;
  assign literal_9176[200] = 5'h10;
  assign literal_9176[201] = 5'h10;
  assign literal_9176[202] = 5'h10;
  assign literal_9176[203] = 5'h00;
  assign literal_9176[204] = 5'h00;
  assign literal_9176[205] = 5'h00;
  assign literal_9176[206] = 5'h00;
  assign literal_9176[207] = 5'h00;
  assign literal_9176[208] = 5'h00;
  assign literal_9176[209] = 5'h0a;
  assign literal_9176[210] = 5'h10;
  assign literal_9176[211] = 5'h10;
  assign literal_9176[212] = 5'h10;
  assign literal_9176[213] = 5'h10;
  assign literal_9176[214] = 5'h10;
  assign literal_9176[215] = 5'h10;
  assign literal_9176[216] = 5'h10;
  assign literal_9176[217] = 5'h10;
  assign literal_9176[218] = 5'h10;
  assign literal_9176[219] = 5'h00;
  assign literal_9176[220] = 5'h00;
  assign literal_9176[221] = 5'h00;
  assign literal_9176[222] = 5'h00;
  assign literal_9176[223] = 5'h00;
  assign literal_9176[224] = 5'h00;
  assign literal_9176[225] = 5'h0b;
  assign literal_9176[226] = 5'h10;
  assign literal_9176[227] = 5'h10;
  assign literal_9176[228] = 5'h10;
  assign literal_9176[229] = 5'h10;
  assign literal_9176[230] = 5'h10;
  assign literal_9176[231] = 5'h10;
  assign literal_9176[232] = 5'h10;
  assign literal_9176[233] = 5'h10;
  assign literal_9176[234] = 5'h10;
  assign literal_9176[235] = 5'h00;
  assign literal_9176[236] = 5'h00;
  assign literal_9176[237] = 5'h00;
  assign literal_9176[238] = 5'h00;
  assign literal_9176[239] = 5'h00;
  assign literal_9176[240] = 5'h0c;
  assign literal_9176[241] = 5'h0d;
  assign literal_9176[242] = 5'h10;
  assign literal_9176[243] = 5'h10;
  assign literal_9176[244] = 5'h10;
  assign literal_9176[245] = 5'h10;
  assign literal_9176[246] = 5'h10;
  assign literal_9176[247] = 5'h10;
  assign literal_9176[248] = 5'h10;
  assign literal_9176[249] = 5'h10;
  assign literal_9176[250] = 5'h10;
  assign literal_9176[251] = 5'h00;
  wire [15:0] literal_9177[0:251];
  assign literal_9177[0] = 16'h0001;
  assign literal_9177[1] = 16'h0000;
  assign literal_9177[2] = 16'h0004;
  assign literal_9177[3] = 16'h000c;
  assign literal_9177[4] = 16'h001a;
  assign literal_9177[5] = 16'h0076;
  assign literal_9177[6] = 16'h00f6;
  assign literal_9177[7] = 16'h3fe0;
  assign literal_9177[8] = 16'hff96;
  assign literal_9177[9] = 16'hff97;
  assign literal_9177[10] = 16'hff98;
  assign literal_9177[11] = 16'h0000;
  assign literal_9177[12] = 16'h0000;
  assign literal_9177[13] = 16'h0000;
  assign literal_9177[14] = 16'h0000;
  assign literal_9177[15] = 16'h0000;
  assign literal_9177[16] = 16'h0000;
  assign literal_9177[17] = 16'h0005;
  assign literal_9177[18] = 16'h0038;
  assign literal_9177[19] = 16'h0078;
  assign literal_9177[20] = 16'h01f9;
  assign literal_9177[21] = 16'h07f2;
  assign literal_9177[22] = 16'h1fe8;
  assign literal_9177[23] = 16'hff93;
  assign literal_9177[24] = 16'hff99;
  assign literal_9177[25] = 16'hff9a;
  assign literal_9177[26] = 16'hff9e;
  assign literal_9177[27] = 16'h0000;
  assign literal_9177[28] = 16'h0000;
  assign literal_9177[29] = 16'h0000;
  assign literal_9177[30] = 16'h0000;
  assign literal_9177[31] = 16'h0000;
  assign literal_9177[32] = 16'h0000;
  assign literal_9177[33] = 16'h001b;
  assign literal_9177[34] = 16'h007a;
  assign literal_9177[35] = 16'h03f7;
  assign literal_9177[36] = 16'h0ff0;
  assign literal_9177[37] = 16'h1feb;
  assign literal_9177[38] = 16'hff9b;
  assign literal_9177[39] = 16'hff9f;
  assign literal_9177[40] = 16'hffa8;
  assign literal_9177[41] = 16'hffa9;
  assign literal_9177[42] = 16'hfff1;
  assign literal_9177[43] = 16'h0000;
  assign literal_9177[44] = 16'h0000;
  assign literal_9177[45] = 16'h0000;
  assign literal_9177[46] = 16'h0000;
  assign literal_9177[47] = 16'h0000;
  assign literal_9177[48] = 16'h0000;
  assign literal_9177[49] = 16'h0039;
  assign literal_9177[50] = 16'h00fa;
  assign literal_9177[51] = 16'h07f7;
  assign literal_9177[52] = 16'h0ff1;
  assign literal_9177[53] = 16'h7fc6;
  assign literal_9177[54] = 16'hff9c;
  assign literal_9177[55] = 16'hffa3;
  assign literal_9177[56] = 16'hffd7;
  assign literal_9177[57] = 16'hffe4;
  assign literal_9177[58] = 16'hfff2;
  assign literal_9177[59] = 16'h0000;
  assign literal_9177[60] = 16'h0000;
  assign literal_9177[61] = 16'h0000;
  assign literal_9177[62] = 16'h0000;
  assign literal_9177[63] = 16'h0000;
  assign literal_9177[64] = 16'h0000;
  assign literal_9177[65] = 16'h003a;
  assign literal_9177[66] = 16'h03f8;
  assign literal_9177[67] = 16'h0ff2;
  assign literal_9177[68] = 16'h7fc8;
  assign literal_9177[69] = 16'hff9d;
  assign literal_9177[70] = 16'hffbf;
  assign literal_9177[71] = 16'hffcb;
  assign literal_9177[72] = 16'hffd8;
  assign literal_9177[73] = 16'hffe5;
  assign literal_9177[74] = 16'hfff3;
  assign literal_9177[75] = 16'h0000;
  assign literal_9177[76] = 16'h0000;
  assign literal_9177[77] = 16'h0000;
  assign literal_9177[78] = 16'h0000;
  assign literal_9177[79] = 16'h0000;
  assign literal_9177[80] = 16'h0000;
  assign literal_9177[81] = 16'h0077;
  assign literal_9177[82] = 16'h07f3;
  assign literal_9177[83] = 16'h1fea;
  assign literal_9177[84] = 16'hff94;
  assign literal_9177[85] = 16'hffa2;
  assign literal_9177[86] = 16'hffc0;
  assign literal_9177[87] = 16'hffcc;
  assign literal_9177[88] = 16'hffd9;
  assign literal_9177[89] = 16'hffe6;
  assign literal_9177[90] = 16'hfff4;
  assign literal_9177[91] = 16'h0000;
  assign literal_9177[92] = 16'h0000;
  assign literal_9177[93] = 16'h0000;
  assign literal_9177[94] = 16'h0000;
  assign literal_9177[95] = 16'h0000;
  assign literal_9177[96] = 16'h0000;
  assign literal_9177[97] = 16'h0079;
  assign literal_9177[98] = 16'h07f4;
  assign literal_9177[99] = 16'h1fed;
  assign literal_9177[100] = 16'hffa0;
  assign literal_9177[101] = 16'hffb5;
  assign literal_9177[102] = 16'hffc1;
  assign literal_9177[103] = 16'hffcd;
  assign literal_9177[104] = 16'hffda;
  assign literal_9177[105] = 16'hffe7;
  assign literal_9177[106] = 16'hfff5;
  assign literal_9177[107] = 16'h0000;
  assign literal_9177[108] = 16'h0000;
  assign literal_9177[109] = 16'h0000;
  assign literal_9177[110] = 16'h0000;
  assign literal_9177[111] = 16'h0000;
  assign literal_9177[112] = 16'h0000;
  assign literal_9177[113] = 16'h00f7;
  assign literal_9177[114] = 16'h07f5;
  assign literal_9177[115] = 16'h3fe1;
  assign literal_9177[116] = 16'hffa1;
  assign literal_9177[117] = 16'hffb6;
  assign literal_9177[118] = 16'hffc2;
  assign literal_9177[119] = 16'hffce;
  assign literal_9177[120] = 16'hffdb;
  assign literal_9177[121] = 16'hffe8;
  assign literal_9177[122] = 16'hfff6;
  assign literal_9177[123] = 16'h0000;
  assign literal_9177[124] = 16'h0000;
  assign literal_9177[125] = 16'h0000;
  assign literal_9177[126] = 16'h0000;
  assign literal_9177[127] = 16'h0000;
  assign literal_9177[128] = 16'h0000;
  assign literal_9177[129] = 16'h00f8;
  assign literal_9177[130] = 16'h0ff3;
  assign literal_9177[131] = 16'hff92;
  assign literal_9177[132] = 16'hffad;
  assign literal_9177[133] = 16'hffb7;
  assign literal_9177[134] = 16'hffc3;
  assign literal_9177[135] = 16'hffcf;
  assign literal_9177[136] = 16'hffdc;
  assign literal_9177[137] = 16'hffe9;
  assign literal_9177[138] = 16'hfff7;
  assign literal_9177[139] = 16'h0000;
  assign literal_9177[140] = 16'h0000;
  assign literal_9177[141] = 16'h0000;
  assign literal_9177[142] = 16'h0000;
  assign literal_9177[143] = 16'h0000;
  assign literal_9177[144] = 16'h0000;
  assign literal_9177[145] = 16'h00f9;
  assign literal_9177[146] = 16'h1fe9;
  assign literal_9177[147] = 16'hff95;
  assign literal_9177[148] = 16'hffae;
  assign literal_9177[149] = 16'hffb8;
  assign literal_9177[150] = 16'hffc4;
  assign literal_9177[151] = 16'hffd0;
  assign literal_9177[152] = 16'hffdd;
  assign literal_9177[153] = 16'hffea;
  assign literal_9177[154] = 16'hfff8;
  assign literal_9177[155] = 16'h0000;
  assign literal_9177[156] = 16'h0000;
  assign literal_9177[157] = 16'h0000;
  assign literal_9177[158] = 16'h0000;
  assign literal_9177[159] = 16'h0000;
  assign literal_9177[160] = 16'h0000;
  assign literal_9177[161] = 16'h01f6;
  assign literal_9177[162] = 16'h1fec;
  assign literal_9177[163] = 16'hffa5;
  assign literal_9177[164] = 16'hffaf;
  assign literal_9177[165] = 16'hffb9;
  assign literal_9177[166] = 16'hffc5;
  assign literal_9177[167] = 16'hffd1;
  assign literal_9177[168] = 16'hffde;
  assign literal_9177[169] = 16'hffeb;
  assign literal_9177[170] = 16'hfff9;
  assign literal_9177[171] = 16'h0000;
  assign literal_9177[172] = 16'h0000;
  assign literal_9177[173] = 16'h0000;
  assign literal_9177[174] = 16'h0000;
  assign literal_9177[175] = 16'h0000;
  assign literal_9177[176] = 16'h0000;
  assign literal_9177[177] = 16'h01f7;
  assign literal_9177[178] = 16'h1fee;
  assign literal_9177[179] = 16'hffa6;
  assign literal_9177[180] = 16'hffb0;
  assign literal_9177[181] = 16'hffba;
  assign literal_9177[182] = 16'hffc6;
  assign literal_9177[183] = 16'hffd2;
  assign literal_9177[184] = 16'hffdf;
  assign literal_9177[185] = 16'hffec;
  assign literal_9177[186] = 16'hfffa;
  assign literal_9177[187] = 16'h0000;
  assign literal_9177[188] = 16'h0000;
  assign literal_9177[189] = 16'h0000;
  assign literal_9177[190] = 16'h0000;
  assign literal_9177[191] = 16'h0000;
  assign literal_9177[192] = 16'h0000;
  assign literal_9177[193] = 16'h03f4;
  assign literal_9177[194] = 16'h1fef;
  assign literal_9177[195] = 16'hffa7;
  assign literal_9177[196] = 16'hffb1;
  assign literal_9177[197] = 16'hffbb;
  assign literal_9177[198] = 16'hffc7;
  assign literal_9177[199] = 16'hffd3;
  assign literal_9177[200] = 16'hffe0;
  assign literal_9177[201] = 16'hffed;
  assign literal_9177[202] = 16'hfffb;
  assign literal_9177[203] = 16'h0000;
  assign literal_9177[204] = 16'h0000;
  assign literal_9177[205] = 16'h0000;
  assign literal_9177[206] = 16'h0000;
  assign literal_9177[207] = 16'h0000;
  assign literal_9177[208] = 16'h0000;
  assign literal_9177[209] = 16'h03f5;
  assign literal_9177[210] = 16'h3fe2;
  assign literal_9177[211] = 16'hffaa;
  assign literal_9177[212] = 16'hffb2;
  assign literal_9177[213] = 16'hffbc;
  assign literal_9177[214] = 16'hffc8;
  assign literal_9177[215] = 16'hffd4;
  assign literal_9177[216] = 16'hffe1;
  assign literal_9177[217] = 16'hffee;
  assign literal_9177[218] = 16'hfffc;
  assign literal_9177[219] = 16'h0000;
  assign literal_9177[220] = 16'h0000;
  assign literal_9177[221] = 16'h0000;
  assign literal_9177[222] = 16'h0000;
  assign literal_9177[223] = 16'h0000;
  assign literal_9177[224] = 16'h0000;
  assign literal_9177[225] = 16'h03f6;
  assign literal_9177[226] = 16'h7fc7;
  assign literal_9177[227] = 16'hffab;
  assign literal_9177[228] = 16'hffb3;
  assign literal_9177[229] = 16'hffbd;
  assign literal_9177[230] = 16'hffc9;
  assign literal_9177[231] = 16'hffd5;
  assign literal_9177[232] = 16'hffe2;
  assign literal_9177[233] = 16'hffef;
  assign literal_9177[234] = 16'hfffd;
  assign literal_9177[235] = 16'h0000;
  assign literal_9177[236] = 16'h0000;
  assign literal_9177[237] = 16'h0000;
  assign literal_9177[238] = 16'h0000;
  assign literal_9177[239] = 16'h0000;
  assign literal_9177[240] = 16'h01f8;
  assign literal_9177[241] = 16'h07f6;
  assign literal_9177[242] = 16'hffa4;
  assign literal_9177[243] = 16'hffac;
  assign literal_9177[244] = 16'hffb4;
  assign literal_9177[245] = 16'hffbe;
  assign literal_9177[246] = 16'hffca;
  assign literal_9177[247] = 16'hffd6;
  assign literal_9177[248] = 16'hffe3;
  assign literal_9177[249] = 16'hfff0;
  assign literal_9177[250] = 16'hfffe;
  assign literal_9177[251] = 16'h0000;
  wire [15:0] literal_9178[0:251];
  assign literal_9178[0] = 16'h000c;
  assign literal_9178[1] = 16'h0000;
  assign literal_9178[2] = 16'h0001;
  assign literal_9178[3] = 16'h0004;
  assign literal_9178[4] = 16'h000b;
  assign literal_9178[5] = 16'h001a;
  assign literal_9178[6] = 16'h0079;
  assign literal_9178[7] = 16'h01f9;
  assign literal_9178[8] = 16'hff9c;
  assign literal_9178[9] = 16'hff9f;
  assign literal_9178[10] = 16'hffa0;
  assign literal_9178[11] = 16'h0000;
  assign literal_9178[12] = 16'h0000;
  assign literal_9178[13] = 16'h0000;
  assign literal_9178[14] = 16'h0000;
  assign literal_9178[15] = 16'h0000;
  assign literal_9178[16] = 16'h0000;
  assign literal_9178[17] = 16'h000a;
  assign literal_9178[18] = 16'h001c;
  assign literal_9178[19] = 16'h007a;
  assign literal_9178[20] = 16'h01f5;
  assign literal_9178[21] = 16'h03f4;
  assign literal_9178[22] = 16'h07f8;
  assign literal_9178[23] = 16'hff95;
  assign literal_9178[24] = 16'hffa1;
  assign literal_9178[25] = 16'hffa2;
  assign literal_9178[26] = 16'hffad;
  assign literal_9178[27] = 16'h0000;
  assign literal_9178[28] = 16'h0000;
  assign literal_9178[29] = 16'h0000;
  assign literal_9178[30] = 16'h0000;
  assign literal_9178[31] = 16'h0000;
  assign literal_9178[32] = 16'h0000;
  assign literal_9178[33] = 16'h001b;
  assign literal_9178[34] = 16'h00f8;
  assign literal_9178[35] = 16'h03f7;
  assign literal_9178[36] = 16'h0ff4;
  assign literal_9178[37] = 16'h3fdc;
  assign literal_9178[38] = 16'hff9d;
  assign literal_9178[39] = 16'hff90;
  assign literal_9178[40] = 16'hffac;
  assign literal_9178[41] = 16'hffe3;
  assign literal_9178[42] = 16'hfff1;
  assign literal_9178[43] = 16'h0000;
  assign literal_9178[44] = 16'h0000;
  assign literal_9178[45] = 16'h0000;
  assign literal_9178[46] = 16'h0000;
  assign literal_9178[47] = 16'h0000;
  assign literal_9178[48] = 16'h0000;
  assign literal_9178[49] = 16'h003a;
  assign literal_9178[50] = 16'h01f6;
  assign literal_9178[51] = 16'h07f7;
  assign literal_9178[52] = 16'h3fde;
  assign literal_9178[53] = 16'hff8e;
  assign literal_9178[54] = 16'hff94;
  assign literal_9178[55] = 16'hffc9;
  assign literal_9178[56] = 16'hffd6;
  assign literal_9178[57] = 16'hffe4;
  assign literal_9178[58] = 16'hfff2;
  assign literal_9178[59] = 16'h0000;
  assign literal_9178[60] = 16'h0000;
  assign literal_9178[61] = 16'h0000;
  assign literal_9178[62] = 16'h0000;
  assign literal_9178[63] = 16'h0000;
  assign literal_9178[64] = 16'h0000;
  assign literal_9178[65] = 16'h003b;
  assign literal_9178[66] = 16'h03f6;
  assign literal_9178[67] = 16'h3fdd;
  assign literal_9178[68] = 16'hff8f;
  assign literal_9178[69] = 16'hffa5;
  assign literal_9178[70] = 16'hffa6;
  assign literal_9178[71] = 16'hffca;
  assign literal_9178[72] = 16'hffd7;
  assign literal_9178[73] = 16'hffe5;
  assign literal_9178[74] = 16'hfff3;
  assign literal_9178[75] = 16'h0000;
  assign literal_9178[76] = 16'h0000;
  assign literal_9178[77] = 16'h0000;
  assign literal_9178[78] = 16'h0000;
  assign literal_9178[79] = 16'h0000;
  assign literal_9178[80] = 16'h0000;
  assign literal_9178[81] = 16'h0078;
  assign literal_9178[82] = 16'h03f9;
  assign literal_9178[83] = 16'h3fdf;
  assign literal_9178[84] = 16'hff96;
  assign literal_9178[85] = 16'hffab;
  assign literal_9178[86] = 16'hffa9;
  assign literal_9178[87] = 16'hffcb;
  assign literal_9178[88] = 16'hffd8;
  assign literal_9178[89] = 16'hffe6;
  assign literal_9178[90] = 16'hfff4;
  assign literal_9178[91] = 16'h0000;
  assign literal_9178[92] = 16'h0000;
  assign literal_9178[93] = 16'h0000;
  assign literal_9178[94] = 16'h0000;
  assign literal_9178[95] = 16'h0000;
  assign literal_9178[96] = 16'h0000;
  assign literal_9178[97] = 16'h007b;
  assign literal_9178[98] = 16'h0ff2;
  assign literal_9178[99] = 16'h7fc5;
  assign literal_9178[100] = 16'hff97;
  assign literal_9178[101] = 16'hffb5;
  assign literal_9178[102] = 16'hffbf;
  assign literal_9178[103] = 16'hffcc;
  assign literal_9178[104] = 16'hffd9;
  assign literal_9178[105] = 16'hffe7;
  assign literal_9178[106] = 16'hfff5;
  assign literal_9178[107] = 16'h0000;
  assign literal_9178[108] = 16'h0000;
  assign literal_9178[109] = 16'h0000;
  assign literal_9178[110] = 16'h0000;
  assign literal_9178[111] = 16'h0000;
  assign literal_9178[112] = 16'h0000;
  assign literal_9178[113] = 16'h00f9;
  assign literal_9178[114] = 16'h0ff5;
  assign literal_9178[115] = 16'hff8c;
  assign literal_9178[116] = 16'hff98;
  assign literal_9178[117] = 16'hffb6;
  assign literal_9178[118] = 16'hffc0;
  assign literal_9178[119] = 16'hffcd;
  assign literal_9178[120] = 16'hffda;
  assign literal_9178[121] = 16'hffe8;
  assign literal_9178[122] = 16'hfff6;
  assign literal_9178[123] = 16'h0000;
  assign literal_9178[124] = 16'h0000;
  assign literal_9178[125] = 16'h0000;
  assign literal_9178[126] = 16'h0000;
  assign literal_9178[127] = 16'h0000;
  assign literal_9178[128] = 16'h0000;
  assign literal_9178[129] = 16'h01f4;
  assign literal_9178[130] = 16'h1fec;
  assign literal_9178[131] = 16'hff9e;
  assign literal_9178[132] = 16'hffa3;
  assign literal_9178[133] = 16'hffb7;
  assign literal_9178[134] = 16'hffc1;
  assign literal_9178[135] = 16'hffce;
  assign literal_9178[136] = 16'hffdb;
  assign literal_9178[137] = 16'hffe9;
  assign literal_9178[138] = 16'hfff7;
  assign literal_9178[139] = 16'h0000;
  assign literal_9178[140] = 16'h0000;
  assign literal_9178[141] = 16'h0000;
  assign literal_9178[142] = 16'h0000;
  assign literal_9178[143] = 16'h0000;
  assign literal_9178[144] = 16'h0000;
  assign literal_9178[145] = 16'h01f7;
  assign literal_9178[146] = 16'h3fe0;
  assign literal_9178[147] = 16'hff91;
  assign literal_9178[148] = 16'hffa4;
  assign literal_9178[149] = 16'hffb8;
  assign literal_9178[150] = 16'hffc2;
  assign literal_9178[151] = 16'hffcf;
  assign literal_9178[152] = 16'hffdc;
  assign literal_9178[153] = 16'hffea;
  assign literal_9178[154] = 16'hfff8;
  assign literal_9178[155] = 16'h0000;
  assign literal_9178[156] = 16'h0000;
  assign literal_9178[157] = 16'h0000;
  assign literal_9178[158] = 16'h0000;
  assign literal_9178[159] = 16'h0000;
  assign literal_9178[160] = 16'h0000;
  assign literal_9178[161] = 16'h01f8;
  assign literal_9178[162] = 16'h3fe1;
  assign literal_9178[163] = 16'hff92;
  assign literal_9178[164] = 16'hffa7;
  assign literal_9178[165] = 16'hffb9;
  assign literal_9178[166] = 16'hffc3;
  assign literal_9178[167] = 16'hffd0;
  assign literal_9178[168] = 16'hffdd;
  assign literal_9178[169] = 16'hffeb;
  assign literal_9178[170] = 16'hfff9;
  assign literal_9178[171] = 16'h0000;
  assign literal_9178[172] = 16'h0000;
  assign literal_9178[173] = 16'h0000;
  assign literal_9178[174] = 16'h0000;
  assign literal_9178[175] = 16'h0000;
  assign literal_9178[176] = 16'h0000;
  assign literal_9178[177] = 16'h03f5;
  assign literal_9178[178] = 16'h7fc4;
  assign literal_9178[179] = 16'hff93;
  assign literal_9178[180] = 16'hffa8;
  assign literal_9178[181] = 16'hffba;
  assign literal_9178[182] = 16'hffc4;
  assign literal_9178[183] = 16'hffd1;
  assign literal_9178[184] = 16'hffde;
  assign literal_9178[185] = 16'hffec;
  assign literal_9178[186] = 16'hfffa;
  assign literal_9178[187] = 16'h0000;
  assign literal_9178[188] = 16'h0000;
  assign literal_9178[189] = 16'h0000;
  assign literal_9178[190] = 16'h0000;
  assign literal_9178[191] = 16'h0000;
  assign literal_9178[192] = 16'h0000;
  assign literal_9178[193] = 16'h03f8;
  assign literal_9178[194] = 16'hff8d;
  assign literal_9178[195] = 16'hff99;
  assign literal_9178[196] = 16'hffb1;
  assign literal_9178[197] = 16'hffbb;
  assign literal_9178[198] = 16'hffc5;
  assign literal_9178[199] = 16'hffd2;
  assign literal_9178[200] = 16'hffdf;
  assign literal_9178[201] = 16'hffed;
  assign literal_9178[202] = 16'hfffb;
  assign literal_9178[203] = 16'h0000;
  assign literal_9178[204] = 16'h0000;
  assign literal_9178[205] = 16'h0000;
  assign literal_9178[206] = 16'h0000;
  assign literal_9178[207] = 16'h0000;
  assign literal_9178[208] = 16'h0000;
  assign literal_9178[209] = 16'h03fa;
  assign literal_9178[210] = 16'hff9a;
  assign literal_9178[211] = 16'hffaa;
  assign literal_9178[212] = 16'hffb2;
  assign literal_9178[213] = 16'hffbc;
  assign literal_9178[214] = 16'hffc6;
  assign literal_9178[215] = 16'hffd3;
  assign literal_9178[216] = 16'hffe0;
  assign literal_9178[217] = 16'hffee;
  assign literal_9178[218] = 16'hfffc;
  assign literal_9178[219] = 16'h0000;
  assign literal_9178[220] = 16'h0000;
  assign literal_9178[221] = 16'h0000;
  assign literal_9178[222] = 16'h0000;
  assign literal_9178[223] = 16'h0000;
  assign literal_9178[224] = 16'h0000;
  assign literal_9178[225] = 16'h07f6;
  assign literal_9178[226] = 16'hff9b;
  assign literal_9178[227] = 16'hffaf;
  assign literal_9178[228] = 16'hffb3;
  assign literal_9178[229] = 16'hffbd;
  assign literal_9178[230] = 16'hffc7;
  assign literal_9178[231] = 16'hffd4;
  assign literal_9178[232] = 16'hffe1;
  assign literal_9178[233] = 16'hffef;
  assign literal_9178[234] = 16'hfffd;
  assign literal_9178[235] = 16'h0000;
  assign literal_9178[236] = 16'h0000;
  assign literal_9178[237] = 16'h0000;
  assign literal_9178[238] = 16'h0000;
  assign literal_9178[239] = 16'h0000;
  assign literal_9178[240] = 16'h0ff3;
  assign literal_9178[241] = 16'h1fed;
  assign literal_9178[242] = 16'hffae;
  assign literal_9178[243] = 16'hffb0;
  assign literal_9178[244] = 16'hffb4;
  assign literal_9178[245] = 16'hffbe;
  assign literal_9178[246] = 16'hffc8;
  assign literal_9178[247] = 16'hffd5;
  assign literal_9178[248] = 16'hffe2;
  assign literal_9178[249] = 16'hfff0;
  assign literal_9178[250] = 16'hfffe;
  assign literal_9178[251] = 16'h0000;
  wire [7:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[7:0];
  assign matrix_unflattened[0][1] = matrix[15:8];
  assign matrix_unflattened[0][2] = matrix[23:16];
  assign matrix_unflattened[0][3] = matrix[31:24];
  assign matrix_unflattened[0][4] = matrix[39:32];
  assign matrix_unflattened[0][5] = matrix[47:40];
  assign matrix_unflattened[0][6] = matrix[55:48];
  assign matrix_unflattened[0][7] = matrix[63:56];
  assign matrix_unflattened[1][0] = matrix[71:64];
  assign matrix_unflattened[1][1] = matrix[79:72];
  assign matrix_unflattened[1][2] = matrix[87:80];
  assign matrix_unflattened[1][3] = matrix[95:88];
  assign matrix_unflattened[1][4] = matrix[103:96];
  assign matrix_unflattened[1][5] = matrix[111:104];
  assign matrix_unflattened[1][6] = matrix[119:112];
  assign matrix_unflattened[1][7] = matrix[127:120];
  assign matrix_unflattened[2][0] = matrix[135:128];
  assign matrix_unflattened[2][1] = matrix[143:136];
  assign matrix_unflattened[2][2] = matrix[151:144];
  assign matrix_unflattened[2][3] = matrix[159:152];
  assign matrix_unflattened[2][4] = matrix[167:160];
  assign matrix_unflattened[2][5] = matrix[175:168];
  assign matrix_unflattened[2][6] = matrix[183:176];
  assign matrix_unflattened[2][7] = matrix[191:184];
  assign matrix_unflattened[3][0] = matrix[199:192];
  assign matrix_unflattened[3][1] = matrix[207:200];
  assign matrix_unflattened[3][2] = matrix[215:208];
  assign matrix_unflattened[3][3] = matrix[223:216];
  assign matrix_unflattened[3][4] = matrix[231:224];
  assign matrix_unflattened[3][5] = matrix[239:232];
  assign matrix_unflattened[3][6] = matrix[247:240];
  assign matrix_unflattened[3][7] = matrix[255:248];
  assign matrix_unflattened[4][0] = matrix[263:256];
  assign matrix_unflattened[4][1] = matrix[271:264];
  assign matrix_unflattened[4][2] = matrix[279:272];
  assign matrix_unflattened[4][3] = matrix[287:280];
  assign matrix_unflattened[4][4] = matrix[295:288];
  assign matrix_unflattened[4][5] = matrix[303:296];
  assign matrix_unflattened[4][6] = matrix[311:304];
  assign matrix_unflattened[4][7] = matrix[319:312];
  assign matrix_unflattened[5][0] = matrix[327:320];
  assign matrix_unflattened[5][1] = matrix[335:328];
  assign matrix_unflattened[5][2] = matrix[343:336];
  assign matrix_unflattened[5][3] = matrix[351:344];
  assign matrix_unflattened[5][4] = matrix[359:352];
  assign matrix_unflattened[5][5] = matrix[367:360];
  assign matrix_unflattened[5][6] = matrix[375:368];
  assign matrix_unflattened[5][7] = matrix[383:376];
  assign matrix_unflattened[6][0] = matrix[391:384];
  assign matrix_unflattened[6][1] = matrix[399:392];
  assign matrix_unflattened[6][2] = matrix[407:400];
  assign matrix_unflattened[6][3] = matrix[415:408];
  assign matrix_unflattened[6][4] = matrix[423:416];
  assign matrix_unflattened[6][5] = matrix[431:424];
  assign matrix_unflattened[6][6] = matrix[439:432];
  assign matrix_unflattened[6][7] = matrix[447:440];
  assign matrix_unflattened[7][0] = matrix[455:448];
  assign matrix_unflattened[7][1] = matrix[463:456];
  assign matrix_unflattened[7][2] = matrix[471:464];
  assign matrix_unflattened[7][3] = matrix[479:472];
  assign matrix_unflattened[7][4] = matrix[487:480];
  assign matrix_unflattened[7][5] = matrix[495:488];
  assign matrix_unflattened[7][6] = matrix[503:496];
  assign matrix_unflattened[7][7] = matrix[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_row0_comb[0:7];
  wire [7:0] p1_row1_comb[0:7];
  wire [7:0] p1_array_concat_8303_comb[0:15];
  wire [7:0] p1_row2_comb[0:7];
  wire [7:0] p1_array_concat_8306_comb[0:23];
  wire [7:0] p1_row3_comb[0:7];
  wire [2:0] p1_idx_u8__4_squeezed_comb;
  wire [7:0] p1_array_concat_8309_comb[0:31];
  wire [7:0] p1_row4_comb[0:7];
  wire [2:0] p1_idx_u8__5_squeezed_comb;
  wire [7:0] p1_array_concat_8312_comb[0:39];
  wire [7:0] p1_row5_comb[0:7];
  wire [2:0] p1_idx_u8__6_squeezed_comb;
  wire [7:0] p1_idx_u8__13_comb;
  wire [7:0] p1_array_concat_8318_comb[0:47];
  wire [7:0] p1_row6_comb[0:7];
  wire [2:0] p1_idx_u8__7_squeezed_comb;
  wire [6:0] p1_add_8321_comb;
  wire [7:0] p1_actual_index__13_comb;
  wire [7:0] p1_array_concat_8325_comb[0:55];
  wire [7:0] p1_row7_comb[0:7];
  wire [5:0] p1_add_8330_comb;
  wire [7:0] p1_flat_comb[0:63];
  wire [7:0] p1_actual_index__14_comb;
  wire [7:0] p1_idx_u8__1_comb;
  wire [7:0] p1_idx_u8__3_comb;
  wire [7:0] p1_idx_u8__5_comb;
  wire [7:0] p1_idx_u8__7_comb;
  wire [7:0] p1_idx_u8__9_comb;
  wire [7:0] p1_idx_u8__11_comb;
  wire [7:0] p1_actual_index__12_comb;
  wire [7:0] p1_actual_index__1_comb;
  wire [6:0] p1_add_8441_comb;
  wire [7:0] p1_actual_index__3_comb;
  wire [5:0] p1_add_8424_comb;
  wire [7:0] p1_actual_index__5_comb;
  wire [6:0] p1_add_8407_comb;
  wire [7:0] p1_actual_index__7_comb;
  wire [7:0] p1_actual_index__9_comb;
  wire [6:0] p1_add_8354_comb;
  wire [7:0] p1_actual_index__11_comb;
  wire [7:0] p1_idx_u8__15_comb;
  wire [7:0] p1_idx_u8__17_comb;
  wire [7:0] p1_idx_u8__19_comb;
  wire [7:0] p1_idx_u8__21_comb;
  wire [7:0] p1_idx_u8__23_comb;
  wire [7:0] p1_idx_u8__25_comb;
  wire [7:0] p1_idx_u8__27_comb;
  wire [7:0] p1_idx_u8__29_comb;
  wire [7:0] p1_idx_u8__31_comb;
  wire [7:0] p1_idx_u8__33_comb;
  wire [7:0] p1_idx_u8__35_comb;
  wire [7:0] p1_idx_u8__37_comb;
  wire [7:0] p1_idx_u8__39_comb;
  wire [7:0] p1_idx_u8__41_comb;
  wire [7:0] p1_idx_u8__43_comb;
  wire [7:0] p1_idx_u8__45_comb;
  wire [7:0] p1_idx_u8__47_comb;
  wire [7:0] p1_idx_u8__49_comb;
  wire [7:0] p1_idx_u8__51_comb;
  wire [7:0] p1_idx_u8__53_comb;
  wire [7:0] p1_idx_u8__55_comb;
  wire [7:0] p1_idx_u8__57_comb;
  wire [7:0] p1_idx_u8__59_comb;
  wire [7:0] p1_idx_u8__61_comb;
  wire [7:0] p1_and_8349_comb;
  wire [4:0] p1_add_8373_comb;
  wire [7:0] p1_actual_index__15_comb;
  wire [3:0] p1_add_8544_comb;
  wire [7:0] p1_actual_index__17_comb;
  wire [6:0] p1_add_8546_comb;
  wire [7:0] p1_actual_index__19_comb;
  wire [5:0] p1_add_8548_comb;
  wire [7:0] p1_actual_index__21_comb;
  wire [6:0] p1_add_8550_comb;
  wire [7:0] p1_actual_index__23_comb;
  wire [4:0] p1_add_8552_comb;
  wire [7:0] p1_actual_index__25_comb;
  wire [6:0] p1_add_8554_comb;
  wire [7:0] p1_actual_index__27_comb;
  wire [5:0] p1_add_8556_comb;
  wire [7:0] p1_actual_index__29_comb;
  wire [6:0] p1_add_8558_comb;
  wire [7:0] p1_actual_index__31_comb;
  wire [2:0] p1_add_8560_comb;
  wire [7:0] p1_actual_index__33_comb;
  wire [6:0] p1_add_8562_comb;
  wire [7:0] p1_actual_index__35_comb;
  wire [5:0] p1_add_8564_comb;
  wire [7:0] p1_actual_index__37_comb;
  wire [6:0] p1_add_8566_comb;
  wire [7:0] p1_actual_index__39_comb;
  wire [4:0] p1_add_8568_comb;
  wire [7:0] p1_actual_index__41_comb;
  wire [6:0] p1_add_8570_comb;
  wire [7:0] p1_actual_index__43_comb;
  wire [5:0] p1_add_8572_comb;
  wire [7:0] p1_actual_index__45_comb;
  wire [6:0] p1_add_8574_comb;
  wire [7:0] p1_actual_index__47_comb;
  wire [3:0] p1_add_8576_comb;
  wire [7:0] p1_actual_index__49_comb;
  wire [6:0] p1_add_8578_comb;
  wire [7:0] p1_actual_index__51_comb;
  wire [5:0] p1_add_8580_comb;
  wire [7:0] p1_actual_index__53_comb;
  wire [6:0] p1_add_8582_comb;
  wire [7:0] p1_actual_index__55_comb;
  wire [4:0] p1_add_8584_comb;
  wire [7:0] p1_actual_index__57_comb;
  wire [6:0] p1_add_8586_comb;
  wire [7:0] p1_actual_index__59_comb;
  wire [5:0] p1_add_8588_comb;
  wire [7:0] p1_actual_index__61_comb;
  wire [6:0] p1_add_8590_comb;
  wire [7:0] p1_and_8357_comb;
  wire p1_eq_8360_comb;
  wire [7:0] p1_and_8361_comb;
  wire [7:0] p1_actual_index__2_comb;
  wire [7:0] p1_actual_index__4_comb;
  wire [7:0] p1_actual_index__6_comb;
  wire [7:0] p1_actual_index__10_comb;
  wire p1_ne_8369_comb;
  wire [1:0] p1_idx_u8__1_squeezed_comb;
  wire p1_eq_8372_comb;
  wire [7:0] p1_actual_index__8_comb;
  wire [7:0] p1_actual_index__16_comb;
  wire [7:0] p1_actual_index__18_comb;
  wire [7:0] p1_actual_index__20_comb;
  wire [7:0] p1_actual_index__22_comb;
  wire [7:0] p1_actual_index__24_comb;
  wire [7:0] p1_actual_index__26_comb;
  wire [7:0] p1_actual_index__28_comb;
  wire [7:0] p1_actual_index__30_comb;
  wire [7:0] p1_actual_index__32_comb;
  wire [7:0] p1_actual_index__34_comb;
  wire [7:0] p1_actual_index__36_comb;
  wire [7:0] p1_actual_index__38_comb;
  wire [7:0] p1_actual_index__40_comb;
  wire [7:0] p1_actual_index__42_comb;
  wire [7:0] p1_actual_index__44_comb;
  wire [7:0] p1_actual_index__46_comb;
  wire [7:0] p1_actual_index__48_comb;
  wire [7:0] p1_actual_index__50_comb;
  wire [7:0] p1_actual_index__52_comb;
  wire [7:0] p1_actual_index__54_comb;
  wire [7:0] p1_actual_index__56_comb;
  wire [7:0] p1_actual_index__58_comb;
  wire [7:0] p1_actual_index__60_comb;
  wire [7:0] p1_actual_index__62_comb;
  wire [7:0] p1_and_8485_comb;
  wire [7:0] p1_and_8487_comb;
  wire [7:0] p1_and_8482_comb;
  wire [7:0] p1_and_8475_comb;
  wire [7:0] p1_and_8468_comb;
  wire [7:0] p1_and_8457_comb;
  wire [7:0] p1_and_8448_comb;
  wire [7:0] p1_and_8438_comb;
  wire [7:0] p1_and_8410_comb;
  wire [7:0] p1_and_8399_comb;
  wire [7:0] p1_and_8389_comb;
  wire p1_ne_8490_comb;
  wire p1_ne_8491_comb;
  wire p1_ne_8489_comb;
  wire p1_ne_8484_comb;
  wire p1_ne_8477_comb;
  wire p1_ne_8470_comb;
  wire p1_ne_8459_comb;
  wire p1_ne_8450_comb;
  wire [7:0] p1_and_8414_comb;
  wire p1_ne_8421_comb;
  wire p1_ne_8412_comb;
  wire p1_ne_8401_comb;
  wire p1_not_8492_comb;
  wire p1_eq_8422_comb;
  wire [2:0] p1_sel_8413_comb;
  wire p1_and_9012_comb;
  wire [7:0] p1_value_comb;
  assign p1_row0_comb[0] = p0_matrix[3'h0][0];
  assign p1_row0_comb[1] = p0_matrix[3'h0][1];
  assign p1_row0_comb[2] = p0_matrix[3'h0][2];
  assign p1_row0_comb[3] = p0_matrix[3'h0][3];
  assign p1_row0_comb[4] = p0_matrix[3'h0][4];
  assign p1_row0_comb[5] = p0_matrix[3'h0][5];
  assign p1_row0_comb[6] = p0_matrix[3'h0][6];
  assign p1_row0_comb[7] = p0_matrix[3'h0][7];
  assign p1_row1_comb[0] = p0_matrix[3'h1][0];
  assign p1_row1_comb[1] = p0_matrix[3'h1][1];
  assign p1_row1_comb[2] = p0_matrix[3'h1][2];
  assign p1_row1_comb[3] = p0_matrix[3'h1][3];
  assign p1_row1_comb[4] = p0_matrix[3'h1][4];
  assign p1_row1_comb[5] = p0_matrix[3'h1][5];
  assign p1_row1_comb[6] = p0_matrix[3'h1][6];
  assign p1_row1_comb[7] = p0_matrix[3'h1][7];
  assign p1_array_concat_8303_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_8303_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_8303_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_8303_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_8303_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_8303_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_8303_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_8303_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_8303_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_8303_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_8303_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_8303_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_8303_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_8303_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_8303_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_8303_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_8306_comb[0] = p1_array_concat_8303_comb[0];
  assign p1_array_concat_8306_comb[1] = p1_array_concat_8303_comb[1];
  assign p1_array_concat_8306_comb[2] = p1_array_concat_8303_comb[2];
  assign p1_array_concat_8306_comb[3] = p1_array_concat_8303_comb[3];
  assign p1_array_concat_8306_comb[4] = p1_array_concat_8303_comb[4];
  assign p1_array_concat_8306_comb[5] = p1_array_concat_8303_comb[5];
  assign p1_array_concat_8306_comb[6] = p1_array_concat_8303_comb[6];
  assign p1_array_concat_8306_comb[7] = p1_array_concat_8303_comb[7];
  assign p1_array_concat_8306_comb[8] = p1_array_concat_8303_comb[8];
  assign p1_array_concat_8306_comb[9] = p1_array_concat_8303_comb[9];
  assign p1_array_concat_8306_comb[10] = p1_array_concat_8303_comb[10];
  assign p1_array_concat_8306_comb[11] = p1_array_concat_8303_comb[11];
  assign p1_array_concat_8306_comb[12] = p1_array_concat_8303_comb[12];
  assign p1_array_concat_8306_comb[13] = p1_array_concat_8303_comb[13];
  assign p1_array_concat_8306_comb[14] = p1_array_concat_8303_comb[14];
  assign p1_array_concat_8306_comb[15] = p1_array_concat_8303_comb[15];
  assign p1_array_concat_8306_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_8306_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_8306_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_8306_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_8306_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_8306_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_8306_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_8306_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_idx_u8__4_squeezed_comb = 3'h4;
  assign p1_array_concat_8309_comb[0] = p1_array_concat_8306_comb[0];
  assign p1_array_concat_8309_comb[1] = p1_array_concat_8306_comb[1];
  assign p1_array_concat_8309_comb[2] = p1_array_concat_8306_comb[2];
  assign p1_array_concat_8309_comb[3] = p1_array_concat_8306_comb[3];
  assign p1_array_concat_8309_comb[4] = p1_array_concat_8306_comb[4];
  assign p1_array_concat_8309_comb[5] = p1_array_concat_8306_comb[5];
  assign p1_array_concat_8309_comb[6] = p1_array_concat_8306_comb[6];
  assign p1_array_concat_8309_comb[7] = p1_array_concat_8306_comb[7];
  assign p1_array_concat_8309_comb[8] = p1_array_concat_8306_comb[8];
  assign p1_array_concat_8309_comb[9] = p1_array_concat_8306_comb[9];
  assign p1_array_concat_8309_comb[10] = p1_array_concat_8306_comb[10];
  assign p1_array_concat_8309_comb[11] = p1_array_concat_8306_comb[11];
  assign p1_array_concat_8309_comb[12] = p1_array_concat_8306_comb[12];
  assign p1_array_concat_8309_comb[13] = p1_array_concat_8306_comb[13];
  assign p1_array_concat_8309_comb[14] = p1_array_concat_8306_comb[14];
  assign p1_array_concat_8309_comb[15] = p1_array_concat_8306_comb[15];
  assign p1_array_concat_8309_comb[16] = p1_array_concat_8306_comb[16];
  assign p1_array_concat_8309_comb[17] = p1_array_concat_8306_comb[17];
  assign p1_array_concat_8309_comb[18] = p1_array_concat_8306_comb[18];
  assign p1_array_concat_8309_comb[19] = p1_array_concat_8306_comb[19];
  assign p1_array_concat_8309_comb[20] = p1_array_concat_8306_comb[20];
  assign p1_array_concat_8309_comb[21] = p1_array_concat_8306_comb[21];
  assign p1_array_concat_8309_comb[22] = p1_array_concat_8306_comb[22];
  assign p1_array_concat_8309_comb[23] = p1_array_concat_8306_comb[23];
  assign p1_array_concat_8309_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_8309_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_8309_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_8309_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_8309_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_8309_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_8309_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_8309_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[p1_idx_u8__4_squeezed_comb][0];
  assign p1_row4_comb[1] = p0_matrix[p1_idx_u8__4_squeezed_comb][1];
  assign p1_row4_comb[2] = p0_matrix[p1_idx_u8__4_squeezed_comb][2];
  assign p1_row4_comb[3] = p0_matrix[p1_idx_u8__4_squeezed_comb][3];
  assign p1_row4_comb[4] = p0_matrix[p1_idx_u8__4_squeezed_comb][4];
  assign p1_row4_comb[5] = p0_matrix[p1_idx_u8__4_squeezed_comb][5];
  assign p1_row4_comb[6] = p0_matrix[p1_idx_u8__4_squeezed_comb][6];
  assign p1_row4_comb[7] = p0_matrix[p1_idx_u8__4_squeezed_comb][7];
  assign p1_idx_u8__5_squeezed_comb = 3'h5;
  assign p1_array_concat_8312_comb[0] = p1_array_concat_8309_comb[0];
  assign p1_array_concat_8312_comb[1] = p1_array_concat_8309_comb[1];
  assign p1_array_concat_8312_comb[2] = p1_array_concat_8309_comb[2];
  assign p1_array_concat_8312_comb[3] = p1_array_concat_8309_comb[3];
  assign p1_array_concat_8312_comb[4] = p1_array_concat_8309_comb[4];
  assign p1_array_concat_8312_comb[5] = p1_array_concat_8309_comb[5];
  assign p1_array_concat_8312_comb[6] = p1_array_concat_8309_comb[6];
  assign p1_array_concat_8312_comb[7] = p1_array_concat_8309_comb[7];
  assign p1_array_concat_8312_comb[8] = p1_array_concat_8309_comb[8];
  assign p1_array_concat_8312_comb[9] = p1_array_concat_8309_comb[9];
  assign p1_array_concat_8312_comb[10] = p1_array_concat_8309_comb[10];
  assign p1_array_concat_8312_comb[11] = p1_array_concat_8309_comb[11];
  assign p1_array_concat_8312_comb[12] = p1_array_concat_8309_comb[12];
  assign p1_array_concat_8312_comb[13] = p1_array_concat_8309_comb[13];
  assign p1_array_concat_8312_comb[14] = p1_array_concat_8309_comb[14];
  assign p1_array_concat_8312_comb[15] = p1_array_concat_8309_comb[15];
  assign p1_array_concat_8312_comb[16] = p1_array_concat_8309_comb[16];
  assign p1_array_concat_8312_comb[17] = p1_array_concat_8309_comb[17];
  assign p1_array_concat_8312_comb[18] = p1_array_concat_8309_comb[18];
  assign p1_array_concat_8312_comb[19] = p1_array_concat_8309_comb[19];
  assign p1_array_concat_8312_comb[20] = p1_array_concat_8309_comb[20];
  assign p1_array_concat_8312_comb[21] = p1_array_concat_8309_comb[21];
  assign p1_array_concat_8312_comb[22] = p1_array_concat_8309_comb[22];
  assign p1_array_concat_8312_comb[23] = p1_array_concat_8309_comb[23];
  assign p1_array_concat_8312_comb[24] = p1_array_concat_8309_comb[24];
  assign p1_array_concat_8312_comb[25] = p1_array_concat_8309_comb[25];
  assign p1_array_concat_8312_comb[26] = p1_array_concat_8309_comb[26];
  assign p1_array_concat_8312_comb[27] = p1_array_concat_8309_comb[27];
  assign p1_array_concat_8312_comb[28] = p1_array_concat_8309_comb[28];
  assign p1_array_concat_8312_comb[29] = p1_array_concat_8309_comb[29];
  assign p1_array_concat_8312_comb[30] = p1_array_concat_8309_comb[30];
  assign p1_array_concat_8312_comb[31] = p1_array_concat_8309_comb[31];
  assign p1_array_concat_8312_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_8312_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_8312_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_8312_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_8312_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_8312_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_8312_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_8312_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[p1_idx_u8__5_squeezed_comb][0];
  assign p1_row5_comb[1] = p0_matrix[p1_idx_u8__5_squeezed_comb][1];
  assign p1_row5_comb[2] = p0_matrix[p1_idx_u8__5_squeezed_comb][2];
  assign p1_row5_comb[3] = p0_matrix[p1_idx_u8__5_squeezed_comb][3];
  assign p1_row5_comb[4] = p0_matrix[p1_idx_u8__5_squeezed_comb][4];
  assign p1_row5_comb[5] = p0_matrix[p1_idx_u8__5_squeezed_comb][5];
  assign p1_row5_comb[6] = p0_matrix[p1_idx_u8__5_squeezed_comb][6];
  assign p1_row5_comb[7] = p0_matrix[p1_idx_u8__5_squeezed_comb][7];
  assign p1_idx_u8__6_squeezed_comb = 3'h6;
  assign p1_idx_u8__13_comb = 8'h0d;
  assign p1_array_concat_8318_comb[0] = p1_array_concat_8312_comb[0];
  assign p1_array_concat_8318_comb[1] = p1_array_concat_8312_comb[1];
  assign p1_array_concat_8318_comb[2] = p1_array_concat_8312_comb[2];
  assign p1_array_concat_8318_comb[3] = p1_array_concat_8312_comb[3];
  assign p1_array_concat_8318_comb[4] = p1_array_concat_8312_comb[4];
  assign p1_array_concat_8318_comb[5] = p1_array_concat_8312_comb[5];
  assign p1_array_concat_8318_comb[6] = p1_array_concat_8312_comb[6];
  assign p1_array_concat_8318_comb[7] = p1_array_concat_8312_comb[7];
  assign p1_array_concat_8318_comb[8] = p1_array_concat_8312_comb[8];
  assign p1_array_concat_8318_comb[9] = p1_array_concat_8312_comb[9];
  assign p1_array_concat_8318_comb[10] = p1_array_concat_8312_comb[10];
  assign p1_array_concat_8318_comb[11] = p1_array_concat_8312_comb[11];
  assign p1_array_concat_8318_comb[12] = p1_array_concat_8312_comb[12];
  assign p1_array_concat_8318_comb[13] = p1_array_concat_8312_comb[13];
  assign p1_array_concat_8318_comb[14] = p1_array_concat_8312_comb[14];
  assign p1_array_concat_8318_comb[15] = p1_array_concat_8312_comb[15];
  assign p1_array_concat_8318_comb[16] = p1_array_concat_8312_comb[16];
  assign p1_array_concat_8318_comb[17] = p1_array_concat_8312_comb[17];
  assign p1_array_concat_8318_comb[18] = p1_array_concat_8312_comb[18];
  assign p1_array_concat_8318_comb[19] = p1_array_concat_8312_comb[19];
  assign p1_array_concat_8318_comb[20] = p1_array_concat_8312_comb[20];
  assign p1_array_concat_8318_comb[21] = p1_array_concat_8312_comb[21];
  assign p1_array_concat_8318_comb[22] = p1_array_concat_8312_comb[22];
  assign p1_array_concat_8318_comb[23] = p1_array_concat_8312_comb[23];
  assign p1_array_concat_8318_comb[24] = p1_array_concat_8312_comb[24];
  assign p1_array_concat_8318_comb[25] = p1_array_concat_8312_comb[25];
  assign p1_array_concat_8318_comb[26] = p1_array_concat_8312_comb[26];
  assign p1_array_concat_8318_comb[27] = p1_array_concat_8312_comb[27];
  assign p1_array_concat_8318_comb[28] = p1_array_concat_8312_comb[28];
  assign p1_array_concat_8318_comb[29] = p1_array_concat_8312_comb[29];
  assign p1_array_concat_8318_comb[30] = p1_array_concat_8312_comb[30];
  assign p1_array_concat_8318_comb[31] = p1_array_concat_8312_comb[31];
  assign p1_array_concat_8318_comb[32] = p1_array_concat_8312_comb[32];
  assign p1_array_concat_8318_comb[33] = p1_array_concat_8312_comb[33];
  assign p1_array_concat_8318_comb[34] = p1_array_concat_8312_comb[34];
  assign p1_array_concat_8318_comb[35] = p1_array_concat_8312_comb[35];
  assign p1_array_concat_8318_comb[36] = p1_array_concat_8312_comb[36];
  assign p1_array_concat_8318_comb[37] = p1_array_concat_8312_comb[37];
  assign p1_array_concat_8318_comb[38] = p1_array_concat_8312_comb[38];
  assign p1_array_concat_8318_comb[39] = p1_array_concat_8312_comb[39];
  assign p1_array_concat_8318_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_8318_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_8318_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_8318_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_8318_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_8318_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_8318_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_8318_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[p1_idx_u8__6_squeezed_comb][0];
  assign p1_row6_comb[1] = p0_matrix[p1_idx_u8__6_squeezed_comb][1];
  assign p1_row6_comb[2] = p0_matrix[p1_idx_u8__6_squeezed_comb][2];
  assign p1_row6_comb[3] = p0_matrix[p1_idx_u8__6_squeezed_comb][3];
  assign p1_row6_comb[4] = p0_matrix[p1_idx_u8__6_squeezed_comb][4];
  assign p1_row6_comb[5] = p0_matrix[p1_idx_u8__6_squeezed_comb][5];
  assign p1_row6_comb[6] = p0_matrix[p1_idx_u8__6_squeezed_comb][6];
  assign p1_row6_comb[7] = p0_matrix[p1_idx_u8__6_squeezed_comb][7];
  assign p1_idx_u8__7_squeezed_comb = 3'h7;
  assign p1_add_8321_comb = p0_start_pix[7:1] + 7'h07;
  assign p1_actual_index__13_comb = p0_start_pix + p1_idx_u8__13_comb;
  assign p1_array_concat_8325_comb[0] = p1_array_concat_8318_comb[0];
  assign p1_array_concat_8325_comb[1] = p1_array_concat_8318_comb[1];
  assign p1_array_concat_8325_comb[2] = p1_array_concat_8318_comb[2];
  assign p1_array_concat_8325_comb[3] = p1_array_concat_8318_comb[3];
  assign p1_array_concat_8325_comb[4] = p1_array_concat_8318_comb[4];
  assign p1_array_concat_8325_comb[5] = p1_array_concat_8318_comb[5];
  assign p1_array_concat_8325_comb[6] = p1_array_concat_8318_comb[6];
  assign p1_array_concat_8325_comb[7] = p1_array_concat_8318_comb[7];
  assign p1_array_concat_8325_comb[8] = p1_array_concat_8318_comb[8];
  assign p1_array_concat_8325_comb[9] = p1_array_concat_8318_comb[9];
  assign p1_array_concat_8325_comb[10] = p1_array_concat_8318_comb[10];
  assign p1_array_concat_8325_comb[11] = p1_array_concat_8318_comb[11];
  assign p1_array_concat_8325_comb[12] = p1_array_concat_8318_comb[12];
  assign p1_array_concat_8325_comb[13] = p1_array_concat_8318_comb[13];
  assign p1_array_concat_8325_comb[14] = p1_array_concat_8318_comb[14];
  assign p1_array_concat_8325_comb[15] = p1_array_concat_8318_comb[15];
  assign p1_array_concat_8325_comb[16] = p1_array_concat_8318_comb[16];
  assign p1_array_concat_8325_comb[17] = p1_array_concat_8318_comb[17];
  assign p1_array_concat_8325_comb[18] = p1_array_concat_8318_comb[18];
  assign p1_array_concat_8325_comb[19] = p1_array_concat_8318_comb[19];
  assign p1_array_concat_8325_comb[20] = p1_array_concat_8318_comb[20];
  assign p1_array_concat_8325_comb[21] = p1_array_concat_8318_comb[21];
  assign p1_array_concat_8325_comb[22] = p1_array_concat_8318_comb[22];
  assign p1_array_concat_8325_comb[23] = p1_array_concat_8318_comb[23];
  assign p1_array_concat_8325_comb[24] = p1_array_concat_8318_comb[24];
  assign p1_array_concat_8325_comb[25] = p1_array_concat_8318_comb[25];
  assign p1_array_concat_8325_comb[26] = p1_array_concat_8318_comb[26];
  assign p1_array_concat_8325_comb[27] = p1_array_concat_8318_comb[27];
  assign p1_array_concat_8325_comb[28] = p1_array_concat_8318_comb[28];
  assign p1_array_concat_8325_comb[29] = p1_array_concat_8318_comb[29];
  assign p1_array_concat_8325_comb[30] = p1_array_concat_8318_comb[30];
  assign p1_array_concat_8325_comb[31] = p1_array_concat_8318_comb[31];
  assign p1_array_concat_8325_comb[32] = p1_array_concat_8318_comb[32];
  assign p1_array_concat_8325_comb[33] = p1_array_concat_8318_comb[33];
  assign p1_array_concat_8325_comb[34] = p1_array_concat_8318_comb[34];
  assign p1_array_concat_8325_comb[35] = p1_array_concat_8318_comb[35];
  assign p1_array_concat_8325_comb[36] = p1_array_concat_8318_comb[36];
  assign p1_array_concat_8325_comb[37] = p1_array_concat_8318_comb[37];
  assign p1_array_concat_8325_comb[38] = p1_array_concat_8318_comb[38];
  assign p1_array_concat_8325_comb[39] = p1_array_concat_8318_comb[39];
  assign p1_array_concat_8325_comb[40] = p1_array_concat_8318_comb[40];
  assign p1_array_concat_8325_comb[41] = p1_array_concat_8318_comb[41];
  assign p1_array_concat_8325_comb[42] = p1_array_concat_8318_comb[42];
  assign p1_array_concat_8325_comb[43] = p1_array_concat_8318_comb[43];
  assign p1_array_concat_8325_comb[44] = p1_array_concat_8318_comb[44];
  assign p1_array_concat_8325_comb[45] = p1_array_concat_8318_comb[45];
  assign p1_array_concat_8325_comb[46] = p1_array_concat_8318_comb[46];
  assign p1_array_concat_8325_comb[47] = p1_array_concat_8318_comb[47];
  assign p1_array_concat_8325_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_8325_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_8325_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_8325_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_8325_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_8325_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_8325_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_8325_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[p1_idx_u8__7_squeezed_comb][0];
  assign p1_row7_comb[1] = p0_matrix[p1_idx_u8__7_squeezed_comb][1];
  assign p1_row7_comb[2] = p0_matrix[p1_idx_u8__7_squeezed_comb][2];
  assign p1_row7_comb[3] = p0_matrix[p1_idx_u8__7_squeezed_comb][3];
  assign p1_row7_comb[4] = p0_matrix[p1_idx_u8__7_squeezed_comb][4];
  assign p1_row7_comb[5] = p0_matrix[p1_idx_u8__7_squeezed_comb][5];
  assign p1_row7_comb[6] = p0_matrix[p1_idx_u8__7_squeezed_comb][6];
  assign p1_row7_comb[7] = p0_matrix[p1_idx_u8__7_squeezed_comb][7];
  assign p1_add_8330_comb = p0_start_pix[7:2] + 6'h03;
  assign p1_flat_comb[0] = p1_array_concat_8325_comb[0];
  assign p1_flat_comb[1] = p1_array_concat_8325_comb[1];
  assign p1_flat_comb[2] = p1_array_concat_8325_comb[2];
  assign p1_flat_comb[3] = p1_array_concat_8325_comb[3];
  assign p1_flat_comb[4] = p1_array_concat_8325_comb[4];
  assign p1_flat_comb[5] = p1_array_concat_8325_comb[5];
  assign p1_flat_comb[6] = p1_array_concat_8325_comb[6];
  assign p1_flat_comb[7] = p1_array_concat_8325_comb[7];
  assign p1_flat_comb[8] = p1_array_concat_8325_comb[8];
  assign p1_flat_comb[9] = p1_array_concat_8325_comb[9];
  assign p1_flat_comb[10] = p1_array_concat_8325_comb[10];
  assign p1_flat_comb[11] = p1_array_concat_8325_comb[11];
  assign p1_flat_comb[12] = p1_array_concat_8325_comb[12];
  assign p1_flat_comb[13] = p1_array_concat_8325_comb[13];
  assign p1_flat_comb[14] = p1_array_concat_8325_comb[14];
  assign p1_flat_comb[15] = p1_array_concat_8325_comb[15];
  assign p1_flat_comb[16] = p1_array_concat_8325_comb[16];
  assign p1_flat_comb[17] = p1_array_concat_8325_comb[17];
  assign p1_flat_comb[18] = p1_array_concat_8325_comb[18];
  assign p1_flat_comb[19] = p1_array_concat_8325_comb[19];
  assign p1_flat_comb[20] = p1_array_concat_8325_comb[20];
  assign p1_flat_comb[21] = p1_array_concat_8325_comb[21];
  assign p1_flat_comb[22] = p1_array_concat_8325_comb[22];
  assign p1_flat_comb[23] = p1_array_concat_8325_comb[23];
  assign p1_flat_comb[24] = p1_array_concat_8325_comb[24];
  assign p1_flat_comb[25] = p1_array_concat_8325_comb[25];
  assign p1_flat_comb[26] = p1_array_concat_8325_comb[26];
  assign p1_flat_comb[27] = p1_array_concat_8325_comb[27];
  assign p1_flat_comb[28] = p1_array_concat_8325_comb[28];
  assign p1_flat_comb[29] = p1_array_concat_8325_comb[29];
  assign p1_flat_comb[30] = p1_array_concat_8325_comb[30];
  assign p1_flat_comb[31] = p1_array_concat_8325_comb[31];
  assign p1_flat_comb[32] = p1_array_concat_8325_comb[32];
  assign p1_flat_comb[33] = p1_array_concat_8325_comb[33];
  assign p1_flat_comb[34] = p1_array_concat_8325_comb[34];
  assign p1_flat_comb[35] = p1_array_concat_8325_comb[35];
  assign p1_flat_comb[36] = p1_array_concat_8325_comb[36];
  assign p1_flat_comb[37] = p1_array_concat_8325_comb[37];
  assign p1_flat_comb[38] = p1_array_concat_8325_comb[38];
  assign p1_flat_comb[39] = p1_array_concat_8325_comb[39];
  assign p1_flat_comb[40] = p1_array_concat_8325_comb[40];
  assign p1_flat_comb[41] = p1_array_concat_8325_comb[41];
  assign p1_flat_comb[42] = p1_array_concat_8325_comb[42];
  assign p1_flat_comb[43] = p1_array_concat_8325_comb[43];
  assign p1_flat_comb[44] = p1_array_concat_8325_comb[44];
  assign p1_flat_comb[45] = p1_array_concat_8325_comb[45];
  assign p1_flat_comb[46] = p1_array_concat_8325_comb[46];
  assign p1_flat_comb[47] = p1_array_concat_8325_comb[47];
  assign p1_flat_comb[48] = p1_array_concat_8325_comb[48];
  assign p1_flat_comb[49] = p1_array_concat_8325_comb[49];
  assign p1_flat_comb[50] = p1_array_concat_8325_comb[50];
  assign p1_flat_comb[51] = p1_array_concat_8325_comb[51];
  assign p1_flat_comb[52] = p1_array_concat_8325_comb[52];
  assign p1_flat_comb[53] = p1_array_concat_8325_comb[53];
  assign p1_flat_comb[54] = p1_array_concat_8325_comb[54];
  assign p1_flat_comb[55] = p1_array_concat_8325_comb[55];
  assign p1_flat_comb[56] = p1_row7_comb[0];
  assign p1_flat_comb[57] = p1_row7_comb[1];
  assign p1_flat_comb[58] = p1_row7_comb[2];
  assign p1_flat_comb[59] = p1_row7_comb[3];
  assign p1_flat_comb[60] = p1_row7_comb[4];
  assign p1_flat_comb[61] = p1_row7_comb[5];
  assign p1_flat_comb[62] = p1_row7_comb[6];
  assign p1_flat_comb[63] = p1_row7_comb[7];
  assign p1_actual_index__14_comb = {p1_add_8321_comb, p0_start_pix[0]};
  assign p1_idx_u8__1_comb = 8'h01;
  assign p1_idx_u8__3_comb = 8'h03;
  assign p1_idx_u8__5_comb = 8'h05;
  assign p1_idx_u8__7_comb = 8'h07;
  assign p1_idx_u8__9_comb = 8'h09;
  assign p1_idx_u8__11_comb = 8'h0b;
  assign p1_actual_index__12_comb = {p1_add_8330_comb, p0_start_pix[1:0]};
  assign p1_actual_index__1_comb = p0_start_pix + p1_idx_u8__1_comb;
  assign p1_add_8441_comb = p0_start_pix[7:1] + 7'h01;
  assign p1_actual_index__3_comb = p0_start_pix + p1_idx_u8__3_comb;
  assign p1_add_8424_comb = p0_start_pix[7:2] + 6'h01;
  assign p1_actual_index__5_comb = p0_start_pix + p1_idx_u8__5_comb;
  assign p1_add_8407_comb = p0_start_pix[7:1] + 7'h03;
  assign p1_actual_index__7_comb = p0_start_pix + p1_idx_u8__7_comb;
  assign p1_actual_index__9_comb = p0_start_pix + p1_idx_u8__9_comb;
  assign p1_add_8354_comb = p0_start_pix[7:1] + 7'h05;
  assign p1_actual_index__11_comb = p0_start_pix + p1_idx_u8__11_comb;
  assign p1_idx_u8__15_comb = 8'h0f;
  assign p1_idx_u8__17_comb = 8'h11;
  assign p1_idx_u8__19_comb = 8'h13;
  assign p1_idx_u8__21_comb = 8'h15;
  assign p1_idx_u8__23_comb = 8'h17;
  assign p1_idx_u8__25_comb = 8'h19;
  assign p1_idx_u8__27_comb = 8'h1b;
  assign p1_idx_u8__29_comb = 8'h1d;
  assign p1_idx_u8__31_comb = 8'h1f;
  assign p1_idx_u8__33_comb = 8'h21;
  assign p1_idx_u8__35_comb = 8'h23;
  assign p1_idx_u8__37_comb = 8'h25;
  assign p1_idx_u8__39_comb = 8'h27;
  assign p1_idx_u8__41_comb = 8'h29;
  assign p1_idx_u8__43_comb = 8'h2b;
  assign p1_idx_u8__45_comb = 8'h2d;
  assign p1_idx_u8__47_comb = 8'h2f;
  assign p1_idx_u8__49_comb = 8'h31;
  assign p1_idx_u8__51_comb = 8'h33;
  assign p1_idx_u8__53_comb = 8'h35;
  assign p1_idx_u8__55_comb = 8'h37;
  assign p1_idx_u8__57_comb = 8'h39;
  assign p1_idx_u8__59_comb = 8'h3b;
  assign p1_idx_u8__61_comb = 8'h3d;
  assign p1_and_8349_comb = p1_flat_comb[p1_actual_index__14_comb > 8'h3f ? 6'h3f : p1_actual_index__14_comb[5:0]] & {8{~(p1_add_8321_comb[5] | p1_add_8321_comb[6])}};
  assign p1_add_8373_comb = p0_start_pix[7:3] + 5'h01;
  assign p1_actual_index__15_comb = p0_start_pix + p1_idx_u8__15_comb;
  assign p1_add_8544_comb = p0_start_pix[7:4] + 4'h1;
  assign p1_actual_index__17_comb = p0_start_pix + p1_idx_u8__17_comb;
  assign p1_add_8546_comb = p0_start_pix[7:1] + 7'h09;
  assign p1_actual_index__19_comb = p0_start_pix + p1_idx_u8__19_comb;
  assign p1_add_8548_comb = p0_start_pix[7:2] + 6'h05;
  assign p1_actual_index__21_comb = p0_start_pix + p1_idx_u8__21_comb;
  assign p1_add_8550_comb = p0_start_pix[7:1] + 7'h0b;
  assign p1_actual_index__23_comb = p0_start_pix + p1_idx_u8__23_comb;
  assign p1_add_8552_comb = p0_start_pix[7:3] + 5'h03;
  assign p1_actual_index__25_comb = p0_start_pix + p1_idx_u8__25_comb;
  assign p1_add_8554_comb = p0_start_pix[7:1] + 7'h0d;
  assign p1_actual_index__27_comb = p0_start_pix + p1_idx_u8__27_comb;
  assign p1_add_8556_comb = p0_start_pix[7:2] + 6'h07;
  assign p1_actual_index__29_comb = p0_start_pix + p1_idx_u8__29_comb;
  assign p1_add_8558_comb = p0_start_pix[7:1] + 7'h0f;
  assign p1_actual_index__31_comb = p0_start_pix + p1_idx_u8__31_comb;
  assign p1_add_8560_comb = p0_start_pix[7:5] + 3'h1;
  assign p1_actual_index__33_comb = p0_start_pix + p1_idx_u8__33_comb;
  assign p1_add_8562_comb = p0_start_pix[7:1] + 7'h11;
  assign p1_actual_index__35_comb = p0_start_pix + p1_idx_u8__35_comb;
  assign p1_add_8564_comb = p0_start_pix[7:2] + 6'h09;
  assign p1_actual_index__37_comb = p0_start_pix + p1_idx_u8__37_comb;
  assign p1_add_8566_comb = p0_start_pix[7:1] + 7'h13;
  assign p1_actual_index__39_comb = p0_start_pix + p1_idx_u8__39_comb;
  assign p1_add_8568_comb = p0_start_pix[7:3] + 5'h05;
  assign p1_actual_index__41_comb = p0_start_pix + p1_idx_u8__41_comb;
  assign p1_add_8570_comb = p0_start_pix[7:1] + 7'h15;
  assign p1_actual_index__43_comb = p0_start_pix + p1_idx_u8__43_comb;
  assign p1_add_8572_comb = p0_start_pix[7:2] + 6'h0b;
  assign p1_actual_index__45_comb = p0_start_pix + p1_idx_u8__45_comb;
  assign p1_add_8574_comb = p0_start_pix[7:1] + 7'h17;
  assign p1_actual_index__47_comb = p0_start_pix + p1_idx_u8__47_comb;
  assign p1_add_8576_comb = p0_start_pix[7:4] + 4'h3;
  assign p1_actual_index__49_comb = p0_start_pix + p1_idx_u8__49_comb;
  assign p1_add_8578_comb = p0_start_pix[7:1] + 7'h19;
  assign p1_actual_index__51_comb = p0_start_pix + p1_idx_u8__51_comb;
  assign p1_add_8580_comb = p0_start_pix[7:2] + 6'h0d;
  assign p1_actual_index__53_comb = p0_start_pix + p1_idx_u8__53_comb;
  assign p1_add_8582_comb = p0_start_pix[7:1] + 7'h1b;
  assign p1_actual_index__55_comb = p0_start_pix + p1_idx_u8__55_comb;
  assign p1_add_8584_comb = p0_start_pix[7:3] + 5'h07;
  assign p1_actual_index__57_comb = p0_start_pix + p1_idx_u8__57_comb;
  assign p1_add_8586_comb = p0_start_pix[7:1] + 7'h1d;
  assign p1_actual_index__59_comb = p0_start_pix + p1_idx_u8__59_comb;
  assign p1_add_8588_comb = p0_start_pix[7:2] + 6'h0f;
  assign p1_actual_index__61_comb = p0_start_pix + p1_idx_u8__61_comb;
  assign p1_add_8590_comb = p0_start_pix[7:1] + 7'h1f;
  assign p1_and_8357_comb = p1_flat_comb[p1_actual_index__13_comb > 8'h3f ? 6'h3f : p1_actual_index__13_comb[5:0]] & {8{~(p1_actual_index__13_comb[6] | p1_actual_index__13_comb[7])}};
  assign p1_eq_8360_comb = p1_and_8349_comb == 8'h00;
  assign p1_and_8361_comb = p1_flat_comb[p1_actual_index__12_comb > 8'h3f ? 6'h3f : p1_actual_index__12_comb[5:0]] & {8{~(p1_add_8330_comb[4] | p1_add_8330_comb[5])}};
  assign p1_actual_index__2_comb = {p1_add_8441_comb, p0_start_pix[0]};
  assign p1_actual_index__4_comb = {p1_add_8424_comb, p0_start_pix[1:0]};
  assign p1_actual_index__6_comb = {p1_add_8407_comb, p0_start_pix[0]};
  assign p1_actual_index__10_comb = {p1_add_8354_comb, p0_start_pix[0]};
  assign p1_ne_8369_comb = p1_and_8357_comb != 8'h00;
  assign p1_idx_u8__1_squeezed_comb = 2'h1;
  assign p1_eq_8372_comb = p1_and_8361_comb == 8'h00;
  assign p1_actual_index__8_comb = {p1_add_8373_comb, p0_start_pix[2:0]};
  assign p1_actual_index__16_comb = {p1_add_8544_comb, p0_start_pix[3:0]};
  assign p1_actual_index__18_comb = {p1_add_8546_comb, p0_start_pix[0]};
  assign p1_actual_index__20_comb = {p1_add_8548_comb, p0_start_pix[1:0]};
  assign p1_actual_index__22_comb = {p1_add_8550_comb, p0_start_pix[0]};
  assign p1_actual_index__24_comb = {p1_add_8552_comb, p0_start_pix[2:0]};
  assign p1_actual_index__26_comb = {p1_add_8554_comb, p0_start_pix[0]};
  assign p1_actual_index__28_comb = {p1_add_8556_comb, p0_start_pix[1:0]};
  assign p1_actual_index__30_comb = {p1_add_8558_comb, p0_start_pix[0]};
  assign p1_actual_index__32_comb = {p1_add_8560_comb, p0_start_pix[4:0]};
  assign p1_actual_index__34_comb = {p1_add_8562_comb, p0_start_pix[0]};
  assign p1_actual_index__36_comb = {p1_add_8564_comb, p0_start_pix[1:0]};
  assign p1_actual_index__38_comb = {p1_add_8566_comb, p0_start_pix[0]};
  assign p1_actual_index__40_comb = {p1_add_8568_comb, p0_start_pix[2:0]};
  assign p1_actual_index__42_comb = {p1_add_8570_comb, p0_start_pix[0]};
  assign p1_actual_index__44_comb = {p1_add_8572_comb, p0_start_pix[1:0]};
  assign p1_actual_index__46_comb = {p1_add_8574_comb, p0_start_pix[0]};
  assign p1_actual_index__48_comb = {p1_add_8576_comb, p0_start_pix[3:0]};
  assign p1_actual_index__50_comb = {p1_add_8578_comb, p0_start_pix[0]};
  assign p1_actual_index__52_comb = {p1_add_8580_comb, p0_start_pix[1:0]};
  assign p1_actual_index__54_comb = {p1_add_8582_comb, p0_start_pix[0]};
  assign p1_actual_index__56_comb = {p1_add_8584_comb, p0_start_pix[2:0]};
  assign p1_actual_index__58_comb = {p1_add_8586_comb, p0_start_pix[0]};
  assign p1_actual_index__60_comb = {p1_add_8588_comb, p0_start_pix[1:0]};
  assign p1_actual_index__62_comb = {p1_add_8590_comb, p0_start_pix[0]};
  assign p1_and_8485_comb = p1_flat_comb[p0_start_pix > 8'h3f ? 6'h3f : p0_start_pix[5:0]] & {8{~(p0_start_pix[6] | p0_start_pix[7])}};
  assign p1_and_8487_comb = p1_flat_comb[p1_actual_index__1_comb > 8'h3f ? 6'h3f : p1_actual_index__1_comb[5:0]] & {8{~(p1_actual_index__1_comb[6] | p1_actual_index__1_comb[7])}};
  assign p1_and_8482_comb = p1_flat_comb[p1_actual_index__2_comb > 8'h3f ? 6'h3f : p1_actual_index__2_comb[5:0]] & {8{~(p1_add_8441_comb[5] | p1_add_8441_comb[6])}};
  assign p1_and_8475_comb = p1_flat_comb[p1_actual_index__3_comb > 8'h3f ? 6'h3f : p1_actual_index__3_comb[5:0]] & {8{~(p1_actual_index__3_comb[6] | p1_actual_index__3_comb[7])}};
  assign p1_and_8468_comb = p1_flat_comb[p1_actual_index__4_comb > 8'h3f ? 6'h3f : p1_actual_index__4_comb[5:0]] & {8{~(p1_add_8424_comb[4] | p1_add_8424_comb[5])}};
  assign p1_and_8457_comb = p1_flat_comb[p1_actual_index__5_comb > 8'h3f ? 6'h3f : p1_actual_index__5_comb[5:0]] & {8{~(p1_actual_index__5_comb[6] | p1_actual_index__5_comb[7])}};
  assign p1_and_8448_comb = p1_flat_comb[p1_actual_index__6_comb > 8'h3f ? 6'h3f : p1_actual_index__6_comb[5:0]] & {8{~(p1_add_8407_comb[5] | p1_add_8407_comb[6])}};
  assign p1_and_8438_comb = p1_flat_comb[p1_actual_index__7_comb > 8'h3f ? 6'h3f : p1_actual_index__7_comb[5:0]] & {8{~(p1_actual_index__7_comb[6] | p1_actual_index__7_comb[7])}};
  assign p1_and_8410_comb = p1_flat_comb[p1_actual_index__9_comb > 8'h3f ? 6'h3f : p1_actual_index__9_comb[5:0]] & {8{~(p1_actual_index__9_comb[6] | p1_actual_index__9_comb[7])}};
  assign p1_and_8399_comb = p1_flat_comb[p1_actual_index__10_comb > 8'h3f ? 6'h3f : p1_actual_index__10_comb[5:0]] & {8{~(p1_add_8354_comb[5] | p1_add_8354_comb[6])}};
  assign p1_and_8389_comb = p1_flat_comb[p1_actual_index__11_comb > 8'h3f ? 6'h3f : p1_actual_index__11_comb[5:0]] & {8{~(p1_actual_index__11_comb[6] | p1_actual_index__11_comb[7])}};
  assign p1_ne_8490_comb = p1_and_8485_comb != 8'h00;
  assign p1_ne_8491_comb = p1_and_8487_comb != 8'h00;
  assign p1_ne_8489_comb = p1_and_8482_comb != 8'h00;
  assign p1_ne_8484_comb = p1_and_8475_comb != 8'h00;
  assign p1_ne_8477_comb = p1_and_8468_comb != 8'h00;
  assign p1_ne_8470_comb = p1_and_8457_comb != 8'h00;
  assign p1_ne_8459_comb = p1_and_8448_comb != 8'h00;
  assign p1_ne_8450_comb = p1_and_8438_comb != 8'h00;
  assign p1_and_8414_comb = p1_flat_comb[p1_actual_index__8_comb > 8'h3f ? 6'h3f : p1_actual_index__8_comb[5:0]] & {8{~(p1_add_8373_comb[3] | p1_add_8373_comb[4])}};
  assign p1_ne_8421_comb = p1_and_8410_comb != 8'h00;
  assign p1_ne_8412_comb = p1_and_8399_comb != 8'h00;
  assign p1_ne_8401_comb = p1_and_8389_comb != 8'h00;
  assign p1_not_8492_comb = ~p1_ne_8490_comb;
  assign p1_eq_8422_comb = p1_and_8414_comb == 8'h00;
  assign p1_sel_8413_comb = p1_ne_8401_comb ? 3'h3 : {1'h1, (p1_ne_8369_comb ? p1_idx_u8__1_squeezed_comb : {1'h1, p1_eq_8360_comb}) & {2{p1_eq_8372_comb}}};
  assign p1_and_9012_comb = p1_not_8492_comb & ~p1_ne_8491_comb & ~p1_ne_8489_comb & ~p1_ne_8484_comb & ~p1_ne_8477_comb & ~p1_ne_8470_comb & ~p1_ne_8459_comb & ~p1_ne_8450_comb & p1_eq_8422_comb & ~p1_ne_8421_comb & ~p1_ne_8412_comb & ~p1_ne_8401_comb & p1_eq_8372_comb & ~p1_ne_8369_comb & p1_eq_8360_comb & (p1_flat_comb[p1_actual_index__15_comb > 8'h3f ? 6'h3f : p1_actual_index__15_comb[5:0]] & {8{~(p1_actual_index__15_comb[6] | p1_actual_index__15_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__16_comb > 8'h3f ? 6'h3f : p1_actual_index__16_comb[5:0]] & {8{~(p1_add_8544_comb[2] | p1_add_8544_comb[3])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__17_comb > 8'h3f ? 6'h3f : p1_actual_index__17_comb[5:0]] & {8{~(p1_actual_index__17_comb[6] | p1_actual_index__17_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__18_comb > 8'h3f ? 6'h3f : p1_actual_index__18_comb[5:0]] & {8{~(p1_add_8546_comb[5] | p1_add_8546_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__19_comb > 8'h3f ? 6'h3f : p1_actual_index__19_comb[5:0]] & {8{~(p1_actual_index__19_comb[6] | p1_actual_index__19_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__20_comb > 8'h3f ? 6'h3f : p1_actual_index__20_comb[5:0]] & {8{~(p1_add_8548_comb[4] | p1_add_8548_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__21_comb > 8'h3f ? 6'h3f : p1_actual_index__21_comb[5:0]] & {8{~(p1_actual_index__21_comb[6] | p1_actual_index__21_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__22_comb > 8'h3f ? 6'h3f : p1_actual_index__22_comb[5:0]] & {8{~(p1_add_8550_comb[5] | p1_add_8550_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__23_comb > 8'h3f ? 6'h3f : p1_actual_index__23_comb[5:0]] & {8{~(p1_actual_index__23_comb[6] | p1_actual_index__23_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__24_comb > 8'h3f ? 6'h3f : p1_actual_index__24_comb[5:0]] & {8{~(p1_add_8552_comb[3] | p1_add_8552_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__25_comb > 8'h3f ? 6'h3f : p1_actual_index__25_comb[5:0]] & {8{~(p1_actual_index__25_comb[6] | p1_actual_index__25_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__26_comb > 8'h3f ? 6'h3f : p1_actual_index__26_comb[5:0]] & {8{~(p1_add_8554_comb[5] | p1_add_8554_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__27_comb > 8'h3f ? 6'h3f : p1_actual_index__27_comb[5:0]] & {8{~(p1_actual_index__27_comb[6] | p1_actual_index__27_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__28_comb > 8'h3f ? 6'h3f : p1_actual_index__28_comb[5:0]] & {8{~(p1_add_8556_comb[4] | p1_add_8556_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__29_comb > 8'h3f ? 6'h3f : p1_actual_index__29_comb[5:0]] & {8{~(p1_actual_index__29_comb[6] | p1_actual_index__29_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__30_comb > 8'h3f ? 6'h3f : p1_actual_index__30_comb[5:0]] & {8{~(p1_add_8558_comb[5] | p1_add_8558_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__31_comb > 8'h3f ? 6'h3f : p1_actual_index__31_comb[5:0]] & {8{~(p1_actual_index__31_comb[6] | p1_actual_index__31_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__32_comb > 8'h3f ? 6'h3f : p1_actual_index__32_comb[5:0]] & {8{~(p1_add_8560_comb[1] | p1_add_8560_comb[2])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__33_comb > 8'h3f ? 6'h3f : p1_actual_index__33_comb[5:0]] & {8{~(p1_actual_index__33_comb[6] | p1_actual_index__33_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__34_comb > 8'h3f ? 6'h3f : p1_actual_index__34_comb[5:0]] & {8{~(p1_add_8562_comb[5] | p1_add_8562_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__35_comb > 8'h3f ? 6'h3f : p1_actual_index__35_comb[5:0]] & {8{~(p1_actual_index__35_comb[6] | p1_actual_index__35_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__36_comb > 8'h3f ? 6'h3f : p1_actual_index__36_comb[5:0]] & {8{~(p1_add_8564_comb[4] | p1_add_8564_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__37_comb > 8'h3f ? 6'h3f : p1_actual_index__37_comb[5:0]] & {8{~(p1_actual_index__37_comb[6] | p1_actual_index__37_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__38_comb > 8'h3f ? 6'h3f : p1_actual_index__38_comb[5:0]] & {8{~(p1_add_8566_comb[5] | p1_add_8566_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__39_comb > 8'h3f ? 6'h3f : p1_actual_index__39_comb[5:0]] & {8{~(p1_actual_index__39_comb[6] | p1_actual_index__39_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__40_comb > 8'h3f ? 6'h3f : p1_actual_index__40_comb[5:0]] & {8{~(p1_add_8568_comb[3] | p1_add_8568_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__41_comb > 8'h3f ? 6'h3f : p1_actual_index__41_comb[5:0]] & {8{~(p1_actual_index__41_comb[6] | p1_actual_index__41_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__42_comb > 8'h3f ? 6'h3f : p1_actual_index__42_comb[5:0]] & {8{~(p1_add_8570_comb[5] | p1_add_8570_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__43_comb > 8'h3f ? 6'h3f : p1_actual_index__43_comb[5:0]] & {8{~(p1_actual_index__43_comb[6] | p1_actual_index__43_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__44_comb > 8'h3f ? 6'h3f : p1_actual_index__44_comb[5:0]] & {8{~(p1_add_8572_comb[4] | p1_add_8572_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__45_comb > 8'h3f ? 6'h3f : p1_actual_index__45_comb[5:0]] & {8{~(p1_actual_index__45_comb[6] | p1_actual_index__45_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__46_comb > 8'h3f ? 6'h3f : p1_actual_index__46_comb[5:0]] & {8{~(p1_add_8574_comb[5] | p1_add_8574_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__47_comb > 8'h3f ? 6'h3f : p1_actual_index__47_comb[5:0]] & {8{~(p1_actual_index__47_comb[6] | p1_actual_index__47_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__48_comb > 8'h3f ? 6'h3f : p1_actual_index__48_comb[5:0]] & {8{~(p1_add_8576_comb[2] | p1_add_8576_comb[3])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__49_comb > 8'h3f ? 6'h3f : p1_actual_index__49_comb[5:0]] & {8{~(p1_actual_index__49_comb[6] | p1_actual_index__49_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__50_comb > 8'h3f ? 6'h3f : p1_actual_index__50_comb[5:0]] & {8{~(p1_add_8578_comb[5] | p1_add_8578_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__51_comb > 8'h3f ? 6'h3f : p1_actual_index__51_comb[5:0]] & {8{~(p1_actual_index__51_comb[6] | p1_actual_index__51_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__52_comb > 8'h3f ? 6'h3f : p1_actual_index__52_comb[5:0]] & {8{~(p1_add_8580_comb[4] | p1_add_8580_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__53_comb > 8'h3f ? 6'h3f : p1_actual_index__53_comb[5:0]] & {8{~(p1_actual_index__53_comb[6] | p1_actual_index__53_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__54_comb > 8'h3f ? 6'h3f : p1_actual_index__54_comb[5:0]] & {8{~(p1_add_8582_comb[5] | p1_add_8582_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__55_comb > 8'h3f ? 6'h3f : p1_actual_index__55_comb[5:0]] & {8{~(p1_actual_index__55_comb[6] | p1_actual_index__55_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__56_comb > 8'h3f ? 6'h3f : p1_actual_index__56_comb[5:0]] & {8{~(p1_add_8584_comb[3] | p1_add_8584_comb[4])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__57_comb > 8'h3f ? 6'h3f : p1_actual_index__57_comb[5:0]] & {8{~(p1_actual_index__57_comb[6] | p1_actual_index__57_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__58_comb > 8'h3f ? 6'h3f : p1_actual_index__58_comb[5:0]] & {8{~(p1_add_8586_comb[5] | p1_add_8586_comb[6])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__59_comb > 8'h3f ? 6'h3f : p1_actual_index__59_comb[5:0]] & {8{~(p1_actual_index__59_comb[6] | p1_actual_index__59_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__60_comb > 8'h3f ? 6'h3f : p1_actual_index__60_comb[5:0]] & {8{~(p1_add_8588_comb[4] | p1_add_8588_comb[5])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__61_comb > 8'h3f ? 6'h3f : p1_actual_index__61_comb[5:0]] & {8{~(p1_actual_index__61_comb[6] | p1_actual_index__61_comb[7])}}) == 8'h00 & (p1_flat_comb[p1_actual_index__62_comb > 8'h3f ? 6'h3f : p1_actual_index__62_comb[5:0]] & {8{~(p1_add_8590_comb[5] | p1_add_8590_comb[6])}}) == 8'h00;
  assign p1_value_comb = p0_matrix[3'h0][3'h0];

  // Registers for pipe stage 1:
  reg p1_is_luminance;
  reg [7:0] p1_and_8349;
  reg [7:0] p1_and_8357;
  reg [7:0] p1_and_8361;
  reg [7:0] p1_and_8389;
  reg [7:0] p1_and_8399;
  reg [7:0] p1_and_8410;
  reg p1_ne_8412;
  reg [2:0] p1_sel_8413;
  reg [7:0] p1_and_8414;
  reg p1_ne_8421;
  reg p1_eq_8422;
  reg [7:0] p1_and_8438;
  reg [7:0] p1_and_8448;
  reg p1_ne_8450;
  reg [7:0] p1_and_8457;
  reg p1_ne_8459;
  reg [7:0] p1_and_8468;
  reg p1_ne_8470;
  reg [7:0] p1_and_8475;
  reg p1_ne_8477;
  reg [7:0] p1_and_8482;
  reg p1_ne_8484;
  reg [7:0] p1_and_8485;
  reg [7:0] p1_and_8487;
  reg p1_ne_8489;
  reg p1_ne_8490;
  reg p1_ne_8491;
  reg p1_not_8492;
  reg p1_and_9012;
  reg [7:0] p1_value;
  always @ (posedge clk) begin
    p1_is_luminance <= p0_is_luminance;
    p1_and_8349 <= p1_and_8349_comb;
    p1_and_8357 <= p1_and_8357_comb;
    p1_and_8361 <= p1_and_8361_comb;
    p1_and_8389 <= p1_and_8389_comb;
    p1_and_8399 <= p1_and_8399_comb;
    p1_and_8410 <= p1_and_8410_comb;
    p1_ne_8412 <= p1_ne_8412_comb;
    p1_sel_8413 <= p1_sel_8413_comb;
    p1_and_8414 <= p1_and_8414_comb;
    p1_ne_8421 <= p1_ne_8421_comb;
    p1_eq_8422 <= p1_eq_8422_comb;
    p1_and_8438 <= p1_and_8438_comb;
    p1_and_8448 <= p1_and_8448_comb;
    p1_ne_8450 <= p1_ne_8450_comb;
    p1_and_8457 <= p1_and_8457_comb;
    p1_ne_8459 <= p1_ne_8459_comb;
    p1_and_8468 <= p1_and_8468_comb;
    p1_ne_8470 <= p1_ne_8470_comb;
    p1_and_8475 <= p1_and_8475_comb;
    p1_ne_8477 <= p1_ne_8477_comb;
    p1_and_8482 <= p1_and_8482_comb;
    p1_ne_8484 <= p1_ne_8484_comb;
    p1_and_8485 <= p1_and_8485_comb;
    p1_and_8487 <= p1_and_8487_comb;
    p1_ne_8489 <= p1_ne_8489_comb;
    p1_ne_8490 <= p1_ne_8490_comb;
    p1_ne_8491 <= p1_ne_8491_comb;
    p1_not_8492 <= p1_not_8492_comb;
    p1_and_9012 <= p1_and_9012_comb;
    p1_value <= p1_value_comb;
  end

  // ===== Pipe stage 2:
  wire [3:0] p2_sel_9087_comb;
  wire [3:0] p2_sel_9095_comb;
  wire [3:0] p2_sel_9099_comb;
  wire [3:0] p2_run_comb;
  wire [7:0] p2_value__1_comb;
  wire p2_eq_9117_comb;
  wire [1:0] p2_idx_u8__1_squeezed__1_comb;
  wire [1:0] p2_idx_u8__2_squeezed_comb;
  wire [3:0] p2_add_9114_comb;
  wire p2_or_reduce_9109_comb;
  wire [1:0] p2_sel_9110_comb;
  wire [3:0] p2_run_u8__1_comb;
  wire [3:0] p2_and_9120_comb;
  assign p2_sel_9087_comb = p1_ne_8450 ? 4'h7 : {1'h1, (p1_ne_8421 ? 3'h1 : (p1_ne_8412 ? 3'h2 : p1_sel_8413)) & {3{p1_eq_8422}}};
  assign p2_sel_9095_comb = p1_ne_8484 ? 4'h3 : (p1_ne_8477 ? 4'h4 : (p1_ne_8470 ? 4'h5 : (p1_ne_8459 ? 4'h6 : p2_sel_9087_comb)));
  assign p2_sel_9099_comb = p1_ne_8491 ? 4'h1 : (p1_ne_8489 ? 4'h2 : p2_sel_9095_comb);
  assign p2_run_comb = p2_sel_9099_comb & {4{p1_not_8492}};
  assign p2_value__1_comb = p2_run_comb == 4'h0 ? p1_and_8485 : (p2_run_comb == 4'h1 ? p1_and_8487 : (p2_run_comb == 4'h2 ? p1_and_8482 : (p2_run_comb == 4'h3 ? p1_and_8475 : (p2_run_comb == 4'h4 ? p1_and_8468 : (p2_run_comb == 4'h5 ? p1_and_8457 : (p2_run_comb == 4'h6 ? p1_and_8448 : (p2_run_comb == 4'h7 ? p1_and_8438 : (p2_run_comb == 4'h8 ? p1_and_8414 : (p2_run_comb == 4'h9 ? p1_and_8410 : (p2_run_comb == 4'ha ? p1_and_8399 : (p2_run_comb == 4'hb ? p1_and_8389 : (p2_run_comb == 4'hc ? p1_and_8361 : (p2_run_comb == 4'hd ? p1_and_8357 : (p2_run_comb == 4'he ? p1_and_8349 : 8'h00))))))))))))));
  assign p2_eq_9117_comb = p2_run_comb == 4'hf;
  assign p2_idx_u8__1_squeezed__1_comb = 2'h1;
  assign p2_idx_u8__2_squeezed_comb = 2'h2;
  assign p2_add_9114_comb = p2_sel_9095_comb + 4'h7;
  assign p2_or_reduce_9109_comb = |p2_value__1_comb[7:2];
  assign p2_sel_9110_comb = |p2_value__1_comb[7:1] ? p2_idx_u8__2_squeezed_comb : p2_idx_u8__1_squeezed__1_comb;
  assign p2_run_u8__1_comb = p2_run_comb < 4'ha ? p2_run_comb : p2_add_9114_comb;
  assign p2_and_9120_comb = p2_sel_9099_comb & {4{~(p2_eq_9117_comb | p1_ne_8490)}};

  // Registers for pipe stage 2:
  reg p2_is_luminance;
  reg [7:0] p2_value__1;
  reg p2_or_reduce_9109;
  reg [1:0] p2_sel_9110;
  reg [3:0] p2_run_u8__1;
  reg p2_and_9012;
  reg p2_eq_9117;
  reg [7:0] p2_value;
  reg [3:0] p2_and_9120;
  always @ (posedge clk) begin
    p2_is_luminance <= p1_is_luminance;
    p2_value__1 <= p2_value__1_comb;
    p2_or_reduce_9109 <= p2_or_reduce_9109_comb;
    p2_sel_9110 <= p2_sel_9110_comb;
    p2_run_u8__1 <= p2_run_u8__1_comb;
    p2_and_9012 <= p1_and_9012;
    p2_eq_9117 <= p2_eq_9117_comb;
    p2_value <= p1_value;
    p2_and_9120 <= p2_and_9120_comb;
  end

  // ===== Pipe stage 3:
  wire [1:0] p3_idx_u8__3_squeezed_comb;
  wire [2:0] p3_idx_u8__4_squeezed__1_comb;
  wire [2:0] p3_idx_u8__5_squeezed__1_comb;
  wire [2:0] p3_idx_u8__6_squeezed__1_comb;
  wire [2:0] p3_idx_u8__7_squeezed__1_comb;
  wire [2:0] p3_sel_9159_comb;
  wire [3:0] p3_idx_u8__8_squeezed_comb;
  wire p3_eq_9164_comb;
  wire [7:0] p3_size__1_comb;
  wire [7:0] p3_idx_u8__48_comb;
  wire [7:0] p3_run_size_str_u8_comb;
  wire p3_or_9179_comb;
  wire [7:0] p3_flipped__1_comb;
  wire [4:0] p3_huffman_length_squeezed_comb;
  wire [4:0] p3_idx_u8__2_squeezed__1_comb;
  wire [7:0] p3_code_list__1_comb;
  wire [15:0] p3_huffman_code_full_comb;
  wire [35:0] p3_tuple_9201_comb;
  assign p3_idx_u8__3_squeezed_comb = 2'h3;
  assign p3_idx_u8__4_squeezed__1_comb = 3'h4;
  assign p3_idx_u8__5_squeezed__1_comb = 3'h5;
  assign p3_idx_u8__6_squeezed__1_comb = 3'h6;
  assign p3_idx_u8__7_squeezed__1_comb = 3'h7;
  assign p3_sel_9159_comb = |p2_value__1[7:6] ? p3_idx_u8__7_squeezed__1_comb : (|p2_value__1[7:5] ? p3_idx_u8__6_squeezed__1_comb : (|p2_value__1[7:4] ? p3_idx_u8__5_squeezed__1_comb : (|p2_value__1[7:3] ? p3_idx_u8__4_squeezed__1_comb : {1'h0, p2_or_reduce_9109 ? p3_idx_u8__3_squeezed_comb : p2_sel_9110})));
  assign p3_idx_u8__8_squeezed_comb = 4'h8;
  assign p3_eq_9164_comb = p2_value__1 == 8'h00;
  assign p3_size__1_comb = {4'h0, p2_value__1[7] ? p3_idx_u8__8_squeezed_comb : {1'h0, p3_sel_9159_comb}} & {8{~p3_eq_9164_comb}};
  assign p3_idx_u8__48_comb = 8'h30;
  assign p3_run_size_str_u8_comb = {p2_run_u8__1, 4'h0} | p3_size__1_comb | p3_idx_u8__48_comb;
  assign p3_or_9179_comb = p2_and_9012 | p2_eq_9117;
  assign p3_flipped__1_comb = 8'hff;
  assign p3_huffman_length_squeezed_comb = p2_is_luminance ? literal_9176[p3_run_size_str_u8_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8_comb] : literal_9174[p3_run_size_str_u8_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8_comb];
  assign p3_idx_u8__2_squeezed__1_comb = 5'h02;
  assign p3_code_list__1_comb = p3_eq_9164_comb ? p3_flipped__1_comb : p2_value__1;
  assign p3_huffman_code_full_comb = p2_is_luminance ? literal_9178[p3_run_size_str_u8_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8_comb] : literal_9177[p3_run_size_str_u8_comb > 8'hfb ? 8'hfb : p3_run_size_str_u8_comb];
  assign p3_tuple_9201_comb = {p3_huffman_code_full_comb & {16{~p3_or_9179_comb}}, {3'h0, p3_or_9179_comb ? p3_idx_u8__2_squeezed__1_comb : p3_huffman_length_squeezed_comb}, p2_and_9012 ? p2_value : p3_code_list__1_comb & {8{~p2_eq_9117}}, p2_and_9012 ? 4'hf : p2_and_9120};

  // Registers for pipe stage 3:
  reg [35:0] p3_tuple_9201;
  always @ (posedge clk) begin
    p3_tuple_9201 <= p3_tuple_9201_comb;
  end
  assign out = p3_tuple_9201;
endmodule
