module Huffman_ACenc(
  input wire clk,
  input wire [639:0] matrix,
  input wire [7:0] start_pix,
  input wire is_luminance,
  output wire [43:0] out
);
  wire [4:0] literal_9110[0:251];
  assign literal_9110[0] = 5'h02;
  assign literal_9110[1] = 5'h02;
  assign literal_9110[2] = 5'h03;
  assign literal_9110[3] = 5'h04;
  assign literal_9110[4] = 5'h05;
  assign literal_9110[5] = 5'h07;
  assign literal_9110[6] = 5'h08;
  assign literal_9110[7] = 5'h0e;
  assign literal_9110[8] = 5'h10;
  assign literal_9110[9] = 5'h10;
  assign literal_9110[10] = 5'h10;
  assign literal_9110[11] = 5'h00;
  assign literal_9110[12] = 5'h00;
  assign literal_9110[13] = 5'h00;
  assign literal_9110[14] = 5'h00;
  assign literal_9110[15] = 5'h00;
  assign literal_9110[16] = 5'h00;
  assign literal_9110[17] = 5'h03;
  assign literal_9110[18] = 5'h06;
  assign literal_9110[19] = 5'h07;
  assign literal_9110[20] = 5'h09;
  assign literal_9110[21] = 5'h0b;
  assign literal_9110[22] = 5'h0d;
  assign literal_9110[23] = 5'h10;
  assign literal_9110[24] = 5'h10;
  assign literal_9110[25] = 5'h10;
  assign literal_9110[26] = 5'h10;
  assign literal_9110[27] = 5'h00;
  assign literal_9110[28] = 5'h00;
  assign literal_9110[29] = 5'h00;
  assign literal_9110[30] = 5'h00;
  assign literal_9110[31] = 5'h00;
  assign literal_9110[32] = 5'h00;
  assign literal_9110[33] = 5'h05;
  assign literal_9110[34] = 5'h07;
  assign literal_9110[35] = 5'h0a;
  assign literal_9110[36] = 5'h0c;
  assign literal_9110[37] = 5'h0d;
  assign literal_9110[38] = 5'h10;
  assign literal_9110[39] = 5'h10;
  assign literal_9110[40] = 5'h10;
  assign literal_9110[41] = 5'h10;
  assign literal_9110[42] = 5'h10;
  assign literal_9110[43] = 5'h00;
  assign literal_9110[44] = 5'h00;
  assign literal_9110[45] = 5'h00;
  assign literal_9110[46] = 5'h00;
  assign literal_9110[47] = 5'h00;
  assign literal_9110[48] = 5'h00;
  assign literal_9110[49] = 5'h06;
  assign literal_9110[50] = 5'h08;
  assign literal_9110[51] = 5'h0b;
  assign literal_9110[52] = 5'h0c;
  assign literal_9110[53] = 5'h0f;
  assign literal_9110[54] = 5'h10;
  assign literal_9110[55] = 5'h10;
  assign literal_9110[56] = 5'h10;
  assign literal_9110[57] = 5'h10;
  assign literal_9110[58] = 5'h10;
  assign literal_9110[59] = 5'h00;
  assign literal_9110[60] = 5'h00;
  assign literal_9110[61] = 5'h00;
  assign literal_9110[62] = 5'h00;
  assign literal_9110[63] = 5'h00;
  assign literal_9110[64] = 5'h00;
  assign literal_9110[65] = 5'h06;
  assign literal_9110[66] = 5'h0a;
  assign literal_9110[67] = 5'h0c;
  assign literal_9110[68] = 5'h0f;
  assign literal_9110[69] = 5'h10;
  assign literal_9110[70] = 5'h10;
  assign literal_9110[71] = 5'h10;
  assign literal_9110[72] = 5'h10;
  assign literal_9110[73] = 5'h10;
  assign literal_9110[74] = 5'h10;
  assign literal_9110[75] = 5'h00;
  assign literal_9110[76] = 5'h00;
  assign literal_9110[77] = 5'h00;
  assign literal_9110[78] = 5'h00;
  assign literal_9110[79] = 5'h00;
  assign literal_9110[80] = 5'h00;
  assign literal_9110[81] = 5'h07;
  assign literal_9110[82] = 5'h0b;
  assign literal_9110[83] = 5'h0d;
  assign literal_9110[84] = 5'h10;
  assign literal_9110[85] = 5'h10;
  assign literal_9110[86] = 5'h10;
  assign literal_9110[87] = 5'h10;
  assign literal_9110[88] = 5'h10;
  assign literal_9110[89] = 5'h10;
  assign literal_9110[90] = 5'h10;
  assign literal_9110[91] = 5'h00;
  assign literal_9110[92] = 5'h00;
  assign literal_9110[93] = 5'h00;
  assign literal_9110[94] = 5'h00;
  assign literal_9110[95] = 5'h00;
  assign literal_9110[96] = 5'h00;
  assign literal_9110[97] = 5'h07;
  assign literal_9110[98] = 5'h0b;
  assign literal_9110[99] = 5'h0d;
  assign literal_9110[100] = 5'h10;
  assign literal_9110[101] = 5'h10;
  assign literal_9110[102] = 5'h10;
  assign literal_9110[103] = 5'h10;
  assign literal_9110[104] = 5'h10;
  assign literal_9110[105] = 5'h10;
  assign literal_9110[106] = 5'h10;
  assign literal_9110[107] = 5'h00;
  assign literal_9110[108] = 5'h00;
  assign literal_9110[109] = 5'h00;
  assign literal_9110[110] = 5'h00;
  assign literal_9110[111] = 5'h00;
  assign literal_9110[112] = 5'h00;
  assign literal_9110[113] = 5'h08;
  assign literal_9110[114] = 5'h0b;
  assign literal_9110[115] = 5'h0e;
  assign literal_9110[116] = 5'h10;
  assign literal_9110[117] = 5'h10;
  assign literal_9110[118] = 5'h10;
  assign literal_9110[119] = 5'h10;
  assign literal_9110[120] = 5'h10;
  assign literal_9110[121] = 5'h10;
  assign literal_9110[122] = 5'h10;
  assign literal_9110[123] = 5'h00;
  assign literal_9110[124] = 5'h00;
  assign literal_9110[125] = 5'h00;
  assign literal_9110[126] = 5'h00;
  assign literal_9110[127] = 5'h00;
  assign literal_9110[128] = 5'h00;
  assign literal_9110[129] = 5'h08;
  assign literal_9110[130] = 5'h0c;
  assign literal_9110[131] = 5'h10;
  assign literal_9110[132] = 5'h10;
  assign literal_9110[133] = 5'h10;
  assign literal_9110[134] = 5'h10;
  assign literal_9110[135] = 5'h10;
  assign literal_9110[136] = 5'h10;
  assign literal_9110[137] = 5'h10;
  assign literal_9110[138] = 5'h10;
  assign literal_9110[139] = 5'h00;
  assign literal_9110[140] = 5'h00;
  assign literal_9110[141] = 5'h00;
  assign literal_9110[142] = 5'h00;
  assign literal_9110[143] = 5'h00;
  assign literal_9110[144] = 5'h00;
  assign literal_9110[145] = 5'h08;
  assign literal_9110[146] = 5'h0d;
  assign literal_9110[147] = 5'h10;
  assign literal_9110[148] = 5'h10;
  assign literal_9110[149] = 5'h10;
  assign literal_9110[150] = 5'h10;
  assign literal_9110[151] = 5'h10;
  assign literal_9110[152] = 5'h10;
  assign literal_9110[153] = 5'h10;
  assign literal_9110[154] = 5'h10;
  assign literal_9110[155] = 5'h00;
  assign literal_9110[156] = 5'h00;
  assign literal_9110[157] = 5'h00;
  assign literal_9110[158] = 5'h00;
  assign literal_9110[159] = 5'h00;
  assign literal_9110[160] = 5'h00;
  assign literal_9110[161] = 5'h09;
  assign literal_9110[162] = 5'h0d;
  assign literal_9110[163] = 5'h10;
  assign literal_9110[164] = 5'h10;
  assign literal_9110[165] = 5'h10;
  assign literal_9110[166] = 5'h10;
  assign literal_9110[167] = 5'h10;
  assign literal_9110[168] = 5'h10;
  assign literal_9110[169] = 5'h10;
  assign literal_9110[170] = 5'h10;
  assign literal_9110[171] = 5'h00;
  assign literal_9110[172] = 5'h00;
  assign literal_9110[173] = 5'h00;
  assign literal_9110[174] = 5'h00;
  assign literal_9110[175] = 5'h00;
  assign literal_9110[176] = 5'h00;
  assign literal_9110[177] = 5'h09;
  assign literal_9110[178] = 5'h0d;
  assign literal_9110[179] = 5'h10;
  assign literal_9110[180] = 5'h10;
  assign literal_9110[181] = 5'h10;
  assign literal_9110[182] = 5'h10;
  assign literal_9110[183] = 5'h10;
  assign literal_9110[184] = 5'h10;
  assign literal_9110[185] = 5'h10;
  assign literal_9110[186] = 5'h10;
  assign literal_9110[187] = 5'h00;
  assign literal_9110[188] = 5'h00;
  assign literal_9110[189] = 5'h00;
  assign literal_9110[190] = 5'h00;
  assign literal_9110[191] = 5'h00;
  assign literal_9110[192] = 5'h00;
  assign literal_9110[193] = 5'h0a;
  assign literal_9110[194] = 5'h0d;
  assign literal_9110[195] = 5'h10;
  assign literal_9110[196] = 5'h10;
  assign literal_9110[197] = 5'h10;
  assign literal_9110[198] = 5'h10;
  assign literal_9110[199] = 5'h10;
  assign literal_9110[200] = 5'h10;
  assign literal_9110[201] = 5'h10;
  assign literal_9110[202] = 5'h10;
  assign literal_9110[203] = 5'h00;
  assign literal_9110[204] = 5'h00;
  assign literal_9110[205] = 5'h00;
  assign literal_9110[206] = 5'h00;
  assign literal_9110[207] = 5'h00;
  assign literal_9110[208] = 5'h00;
  assign literal_9110[209] = 5'h0a;
  assign literal_9110[210] = 5'h0e;
  assign literal_9110[211] = 5'h10;
  assign literal_9110[212] = 5'h10;
  assign literal_9110[213] = 5'h10;
  assign literal_9110[214] = 5'h10;
  assign literal_9110[215] = 5'h10;
  assign literal_9110[216] = 5'h10;
  assign literal_9110[217] = 5'h10;
  assign literal_9110[218] = 5'h10;
  assign literal_9110[219] = 5'h00;
  assign literal_9110[220] = 5'h00;
  assign literal_9110[221] = 5'h00;
  assign literal_9110[222] = 5'h00;
  assign literal_9110[223] = 5'h00;
  assign literal_9110[224] = 5'h00;
  assign literal_9110[225] = 5'h0a;
  assign literal_9110[226] = 5'h0f;
  assign literal_9110[227] = 5'h10;
  assign literal_9110[228] = 5'h10;
  assign literal_9110[229] = 5'h10;
  assign literal_9110[230] = 5'h10;
  assign literal_9110[231] = 5'h10;
  assign literal_9110[232] = 5'h10;
  assign literal_9110[233] = 5'h10;
  assign literal_9110[234] = 5'h10;
  assign literal_9110[235] = 5'h00;
  assign literal_9110[236] = 5'h00;
  assign literal_9110[237] = 5'h00;
  assign literal_9110[238] = 5'h00;
  assign literal_9110[239] = 5'h00;
  assign literal_9110[240] = 5'h09;
  assign literal_9110[241] = 5'h0b;
  assign literal_9110[242] = 5'h10;
  assign literal_9110[243] = 5'h10;
  assign literal_9110[244] = 5'h10;
  assign literal_9110[245] = 5'h10;
  assign literal_9110[246] = 5'h10;
  assign literal_9110[247] = 5'h10;
  assign literal_9110[248] = 5'h10;
  assign literal_9110[249] = 5'h10;
  assign literal_9110[250] = 5'h10;
  assign literal_9110[251] = 5'h00;
  wire [4:0] literal_9112[0:251];
  assign literal_9112[0] = 5'h04;
  assign literal_9112[1] = 5'h02;
  assign literal_9112[2] = 5'h02;
  assign literal_9112[3] = 5'h03;
  assign literal_9112[4] = 5'h04;
  assign literal_9112[5] = 5'h05;
  assign literal_9112[6] = 5'h07;
  assign literal_9112[7] = 5'h09;
  assign literal_9112[8] = 5'h10;
  assign literal_9112[9] = 5'h10;
  assign literal_9112[10] = 5'h10;
  assign literal_9112[11] = 5'h00;
  assign literal_9112[12] = 5'h00;
  assign literal_9112[13] = 5'h00;
  assign literal_9112[14] = 5'h00;
  assign literal_9112[15] = 5'h00;
  assign literal_9112[16] = 5'h00;
  assign literal_9112[17] = 5'h04;
  assign literal_9112[18] = 5'h05;
  assign literal_9112[19] = 5'h07;
  assign literal_9112[20] = 5'h09;
  assign literal_9112[21] = 5'h0a;
  assign literal_9112[22] = 5'h0b;
  assign literal_9112[23] = 5'h10;
  assign literal_9112[24] = 5'h10;
  assign literal_9112[25] = 5'h10;
  assign literal_9112[26] = 5'h10;
  assign literal_9112[27] = 5'h00;
  assign literal_9112[28] = 5'h00;
  assign literal_9112[29] = 5'h00;
  assign literal_9112[30] = 5'h00;
  assign literal_9112[31] = 5'h00;
  assign literal_9112[32] = 5'h00;
  assign literal_9112[33] = 5'h05;
  assign literal_9112[34] = 5'h08;
  assign literal_9112[35] = 5'h0a;
  assign literal_9112[36] = 5'h0c;
  assign literal_9112[37] = 5'h0e;
  assign literal_9112[38] = 5'h10;
  assign literal_9112[39] = 5'h10;
  assign literal_9112[40] = 5'h10;
  assign literal_9112[41] = 5'h10;
  assign literal_9112[42] = 5'h10;
  assign literal_9112[43] = 5'h00;
  assign literal_9112[44] = 5'h00;
  assign literal_9112[45] = 5'h00;
  assign literal_9112[46] = 5'h00;
  assign literal_9112[47] = 5'h00;
  assign literal_9112[48] = 5'h00;
  assign literal_9112[49] = 5'h06;
  assign literal_9112[50] = 5'h09;
  assign literal_9112[51] = 5'h0b;
  assign literal_9112[52] = 5'h0e;
  assign literal_9112[53] = 5'h10;
  assign literal_9112[54] = 5'h10;
  assign literal_9112[55] = 5'h10;
  assign literal_9112[56] = 5'h10;
  assign literal_9112[57] = 5'h10;
  assign literal_9112[58] = 5'h10;
  assign literal_9112[59] = 5'h00;
  assign literal_9112[60] = 5'h00;
  assign literal_9112[61] = 5'h00;
  assign literal_9112[62] = 5'h00;
  assign literal_9112[63] = 5'h00;
  assign literal_9112[64] = 5'h00;
  assign literal_9112[65] = 5'h06;
  assign literal_9112[66] = 5'h0a;
  assign literal_9112[67] = 5'h0e;
  assign literal_9112[68] = 5'h10;
  assign literal_9112[69] = 5'h10;
  assign literal_9112[70] = 5'h10;
  assign literal_9112[71] = 5'h10;
  assign literal_9112[72] = 5'h10;
  assign literal_9112[73] = 5'h10;
  assign literal_9112[74] = 5'h10;
  assign literal_9112[75] = 5'h00;
  assign literal_9112[76] = 5'h00;
  assign literal_9112[77] = 5'h00;
  assign literal_9112[78] = 5'h00;
  assign literal_9112[79] = 5'h00;
  assign literal_9112[80] = 5'h00;
  assign literal_9112[81] = 5'h07;
  assign literal_9112[82] = 5'h0a;
  assign literal_9112[83] = 5'h0e;
  assign literal_9112[84] = 5'h10;
  assign literal_9112[85] = 5'h10;
  assign literal_9112[86] = 5'h10;
  assign literal_9112[87] = 5'h10;
  assign literal_9112[88] = 5'h10;
  assign literal_9112[89] = 5'h10;
  assign literal_9112[90] = 5'h10;
  assign literal_9112[91] = 5'h00;
  assign literal_9112[92] = 5'h00;
  assign literal_9112[93] = 5'h00;
  assign literal_9112[94] = 5'h00;
  assign literal_9112[95] = 5'h00;
  assign literal_9112[96] = 5'h00;
  assign literal_9112[97] = 5'h07;
  assign literal_9112[98] = 5'h0c;
  assign literal_9112[99] = 5'h0f;
  assign literal_9112[100] = 5'h10;
  assign literal_9112[101] = 5'h10;
  assign literal_9112[102] = 5'h10;
  assign literal_9112[103] = 5'h10;
  assign literal_9112[104] = 5'h10;
  assign literal_9112[105] = 5'h10;
  assign literal_9112[106] = 5'h10;
  assign literal_9112[107] = 5'h00;
  assign literal_9112[108] = 5'h00;
  assign literal_9112[109] = 5'h00;
  assign literal_9112[110] = 5'h00;
  assign literal_9112[111] = 5'h00;
  assign literal_9112[112] = 5'h00;
  assign literal_9112[113] = 5'h08;
  assign literal_9112[114] = 5'h0c;
  assign literal_9112[115] = 5'h10;
  assign literal_9112[116] = 5'h10;
  assign literal_9112[117] = 5'h10;
  assign literal_9112[118] = 5'h10;
  assign literal_9112[119] = 5'h10;
  assign literal_9112[120] = 5'h10;
  assign literal_9112[121] = 5'h10;
  assign literal_9112[122] = 5'h10;
  assign literal_9112[123] = 5'h00;
  assign literal_9112[124] = 5'h00;
  assign literal_9112[125] = 5'h00;
  assign literal_9112[126] = 5'h00;
  assign literal_9112[127] = 5'h00;
  assign literal_9112[128] = 5'h00;
  assign literal_9112[129] = 5'h09;
  assign literal_9112[130] = 5'h0d;
  assign literal_9112[131] = 5'h10;
  assign literal_9112[132] = 5'h10;
  assign literal_9112[133] = 5'h10;
  assign literal_9112[134] = 5'h10;
  assign literal_9112[135] = 5'h10;
  assign literal_9112[136] = 5'h10;
  assign literal_9112[137] = 5'h10;
  assign literal_9112[138] = 5'h10;
  assign literal_9112[139] = 5'h00;
  assign literal_9112[140] = 5'h00;
  assign literal_9112[141] = 5'h00;
  assign literal_9112[142] = 5'h00;
  assign literal_9112[143] = 5'h00;
  assign literal_9112[144] = 5'h00;
  assign literal_9112[145] = 5'h09;
  assign literal_9112[146] = 5'h0e;
  assign literal_9112[147] = 5'h10;
  assign literal_9112[148] = 5'h10;
  assign literal_9112[149] = 5'h10;
  assign literal_9112[150] = 5'h10;
  assign literal_9112[151] = 5'h10;
  assign literal_9112[152] = 5'h10;
  assign literal_9112[153] = 5'h10;
  assign literal_9112[154] = 5'h10;
  assign literal_9112[155] = 5'h00;
  assign literal_9112[156] = 5'h00;
  assign literal_9112[157] = 5'h00;
  assign literal_9112[158] = 5'h00;
  assign literal_9112[159] = 5'h00;
  assign literal_9112[160] = 5'h00;
  assign literal_9112[161] = 5'h09;
  assign literal_9112[162] = 5'h0e;
  assign literal_9112[163] = 5'h10;
  assign literal_9112[164] = 5'h10;
  assign literal_9112[165] = 5'h10;
  assign literal_9112[166] = 5'h10;
  assign literal_9112[167] = 5'h10;
  assign literal_9112[168] = 5'h10;
  assign literal_9112[169] = 5'h10;
  assign literal_9112[170] = 5'h10;
  assign literal_9112[171] = 5'h00;
  assign literal_9112[172] = 5'h00;
  assign literal_9112[173] = 5'h00;
  assign literal_9112[174] = 5'h00;
  assign literal_9112[175] = 5'h00;
  assign literal_9112[176] = 5'h00;
  assign literal_9112[177] = 5'h0a;
  assign literal_9112[178] = 5'h0f;
  assign literal_9112[179] = 5'h10;
  assign literal_9112[180] = 5'h10;
  assign literal_9112[181] = 5'h10;
  assign literal_9112[182] = 5'h10;
  assign literal_9112[183] = 5'h10;
  assign literal_9112[184] = 5'h10;
  assign literal_9112[185] = 5'h10;
  assign literal_9112[186] = 5'h10;
  assign literal_9112[187] = 5'h00;
  assign literal_9112[188] = 5'h00;
  assign literal_9112[189] = 5'h00;
  assign literal_9112[190] = 5'h00;
  assign literal_9112[191] = 5'h00;
  assign literal_9112[192] = 5'h00;
  assign literal_9112[193] = 5'h0a;
  assign literal_9112[194] = 5'h10;
  assign literal_9112[195] = 5'h10;
  assign literal_9112[196] = 5'h10;
  assign literal_9112[197] = 5'h10;
  assign literal_9112[198] = 5'h10;
  assign literal_9112[199] = 5'h10;
  assign literal_9112[200] = 5'h10;
  assign literal_9112[201] = 5'h10;
  assign literal_9112[202] = 5'h10;
  assign literal_9112[203] = 5'h00;
  assign literal_9112[204] = 5'h00;
  assign literal_9112[205] = 5'h00;
  assign literal_9112[206] = 5'h00;
  assign literal_9112[207] = 5'h00;
  assign literal_9112[208] = 5'h00;
  assign literal_9112[209] = 5'h0a;
  assign literal_9112[210] = 5'h10;
  assign literal_9112[211] = 5'h10;
  assign literal_9112[212] = 5'h10;
  assign literal_9112[213] = 5'h10;
  assign literal_9112[214] = 5'h10;
  assign literal_9112[215] = 5'h10;
  assign literal_9112[216] = 5'h10;
  assign literal_9112[217] = 5'h10;
  assign literal_9112[218] = 5'h10;
  assign literal_9112[219] = 5'h00;
  assign literal_9112[220] = 5'h00;
  assign literal_9112[221] = 5'h00;
  assign literal_9112[222] = 5'h00;
  assign literal_9112[223] = 5'h00;
  assign literal_9112[224] = 5'h00;
  assign literal_9112[225] = 5'h0b;
  assign literal_9112[226] = 5'h10;
  assign literal_9112[227] = 5'h10;
  assign literal_9112[228] = 5'h10;
  assign literal_9112[229] = 5'h10;
  assign literal_9112[230] = 5'h10;
  assign literal_9112[231] = 5'h10;
  assign literal_9112[232] = 5'h10;
  assign literal_9112[233] = 5'h10;
  assign literal_9112[234] = 5'h10;
  assign literal_9112[235] = 5'h00;
  assign literal_9112[236] = 5'h00;
  assign literal_9112[237] = 5'h00;
  assign literal_9112[238] = 5'h00;
  assign literal_9112[239] = 5'h00;
  assign literal_9112[240] = 5'h0c;
  assign literal_9112[241] = 5'h0d;
  assign literal_9112[242] = 5'h10;
  assign literal_9112[243] = 5'h10;
  assign literal_9112[244] = 5'h10;
  assign literal_9112[245] = 5'h10;
  assign literal_9112[246] = 5'h10;
  assign literal_9112[247] = 5'h10;
  assign literal_9112[248] = 5'h10;
  assign literal_9112[249] = 5'h10;
  assign literal_9112[250] = 5'h10;
  assign literal_9112[251] = 5'h00;
  wire [15:0] literal_9115[0:251];
  assign literal_9115[0] = 16'h0001;
  assign literal_9115[1] = 16'h0000;
  assign literal_9115[2] = 16'h0004;
  assign literal_9115[3] = 16'h000c;
  assign literal_9115[4] = 16'h001a;
  assign literal_9115[5] = 16'h0076;
  assign literal_9115[6] = 16'h00f6;
  assign literal_9115[7] = 16'h3fe0;
  assign literal_9115[8] = 16'hff96;
  assign literal_9115[9] = 16'hff97;
  assign literal_9115[10] = 16'hff98;
  assign literal_9115[11] = 16'h0000;
  assign literal_9115[12] = 16'h0000;
  assign literal_9115[13] = 16'h0000;
  assign literal_9115[14] = 16'h0000;
  assign literal_9115[15] = 16'h0000;
  assign literal_9115[16] = 16'h0000;
  assign literal_9115[17] = 16'h0005;
  assign literal_9115[18] = 16'h0038;
  assign literal_9115[19] = 16'h0078;
  assign literal_9115[20] = 16'h01f9;
  assign literal_9115[21] = 16'h07f2;
  assign literal_9115[22] = 16'h1fe8;
  assign literal_9115[23] = 16'hff93;
  assign literal_9115[24] = 16'hff99;
  assign literal_9115[25] = 16'hff9a;
  assign literal_9115[26] = 16'hff9e;
  assign literal_9115[27] = 16'h0000;
  assign literal_9115[28] = 16'h0000;
  assign literal_9115[29] = 16'h0000;
  assign literal_9115[30] = 16'h0000;
  assign literal_9115[31] = 16'h0000;
  assign literal_9115[32] = 16'h0000;
  assign literal_9115[33] = 16'h001b;
  assign literal_9115[34] = 16'h007a;
  assign literal_9115[35] = 16'h03f7;
  assign literal_9115[36] = 16'h0ff0;
  assign literal_9115[37] = 16'h1feb;
  assign literal_9115[38] = 16'hff9b;
  assign literal_9115[39] = 16'hff9f;
  assign literal_9115[40] = 16'hffa8;
  assign literal_9115[41] = 16'hffa9;
  assign literal_9115[42] = 16'hfff1;
  assign literal_9115[43] = 16'h0000;
  assign literal_9115[44] = 16'h0000;
  assign literal_9115[45] = 16'h0000;
  assign literal_9115[46] = 16'h0000;
  assign literal_9115[47] = 16'h0000;
  assign literal_9115[48] = 16'h0000;
  assign literal_9115[49] = 16'h0039;
  assign literal_9115[50] = 16'h00fa;
  assign literal_9115[51] = 16'h07f7;
  assign literal_9115[52] = 16'h0ff1;
  assign literal_9115[53] = 16'h7fc6;
  assign literal_9115[54] = 16'hff9c;
  assign literal_9115[55] = 16'hffa3;
  assign literal_9115[56] = 16'hffd7;
  assign literal_9115[57] = 16'hffe4;
  assign literal_9115[58] = 16'hfff2;
  assign literal_9115[59] = 16'h0000;
  assign literal_9115[60] = 16'h0000;
  assign literal_9115[61] = 16'h0000;
  assign literal_9115[62] = 16'h0000;
  assign literal_9115[63] = 16'h0000;
  assign literal_9115[64] = 16'h0000;
  assign literal_9115[65] = 16'h003a;
  assign literal_9115[66] = 16'h03f8;
  assign literal_9115[67] = 16'h0ff2;
  assign literal_9115[68] = 16'h7fc8;
  assign literal_9115[69] = 16'hff9d;
  assign literal_9115[70] = 16'hffbf;
  assign literal_9115[71] = 16'hffcb;
  assign literal_9115[72] = 16'hffd8;
  assign literal_9115[73] = 16'hffe5;
  assign literal_9115[74] = 16'hfff3;
  assign literal_9115[75] = 16'h0000;
  assign literal_9115[76] = 16'h0000;
  assign literal_9115[77] = 16'h0000;
  assign literal_9115[78] = 16'h0000;
  assign literal_9115[79] = 16'h0000;
  assign literal_9115[80] = 16'h0000;
  assign literal_9115[81] = 16'h0077;
  assign literal_9115[82] = 16'h07f3;
  assign literal_9115[83] = 16'h1fea;
  assign literal_9115[84] = 16'hff94;
  assign literal_9115[85] = 16'hffa2;
  assign literal_9115[86] = 16'hffc0;
  assign literal_9115[87] = 16'hffcc;
  assign literal_9115[88] = 16'hffd9;
  assign literal_9115[89] = 16'hffe6;
  assign literal_9115[90] = 16'hfff4;
  assign literal_9115[91] = 16'h0000;
  assign literal_9115[92] = 16'h0000;
  assign literal_9115[93] = 16'h0000;
  assign literal_9115[94] = 16'h0000;
  assign literal_9115[95] = 16'h0000;
  assign literal_9115[96] = 16'h0000;
  assign literal_9115[97] = 16'h0079;
  assign literal_9115[98] = 16'h07f4;
  assign literal_9115[99] = 16'h1fed;
  assign literal_9115[100] = 16'hffa0;
  assign literal_9115[101] = 16'hffb5;
  assign literal_9115[102] = 16'hffc1;
  assign literal_9115[103] = 16'hffcd;
  assign literal_9115[104] = 16'hffda;
  assign literal_9115[105] = 16'hffe7;
  assign literal_9115[106] = 16'hfff5;
  assign literal_9115[107] = 16'h0000;
  assign literal_9115[108] = 16'h0000;
  assign literal_9115[109] = 16'h0000;
  assign literal_9115[110] = 16'h0000;
  assign literal_9115[111] = 16'h0000;
  assign literal_9115[112] = 16'h0000;
  assign literal_9115[113] = 16'h00f7;
  assign literal_9115[114] = 16'h07f5;
  assign literal_9115[115] = 16'h3fe1;
  assign literal_9115[116] = 16'hffa1;
  assign literal_9115[117] = 16'hffb6;
  assign literal_9115[118] = 16'hffc2;
  assign literal_9115[119] = 16'hffce;
  assign literal_9115[120] = 16'hffdb;
  assign literal_9115[121] = 16'hffe8;
  assign literal_9115[122] = 16'hfff6;
  assign literal_9115[123] = 16'h0000;
  assign literal_9115[124] = 16'h0000;
  assign literal_9115[125] = 16'h0000;
  assign literal_9115[126] = 16'h0000;
  assign literal_9115[127] = 16'h0000;
  assign literal_9115[128] = 16'h0000;
  assign literal_9115[129] = 16'h00f8;
  assign literal_9115[130] = 16'h0ff3;
  assign literal_9115[131] = 16'hff92;
  assign literal_9115[132] = 16'hffad;
  assign literal_9115[133] = 16'hffb7;
  assign literal_9115[134] = 16'hffc3;
  assign literal_9115[135] = 16'hffcf;
  assign literal_9115[136] = 16'hffdc;
  assign literal_9115[137] = 16'hffe9;
  assign literal_9115[138] = 16'hfff7;
  assign literal_9115[139] = 16'h0000;
  assign literal_9115[140] = 16'h0000;
  assign literal_9115[141] = 16'h0000;
  assign literal_9115[142] = 16'h0000;
  assign literal_9115[143] = 16'h0000;
  assign literal_9115[144] = 16'h0000;
  assign literal_9115[145] = 16'h00f9;
  assign literal_9115[146] = 16'h1fe9;
  assign literal_9115[147] = 16'hff95;
  assign literal_9115[148] = 16'hffae;
  assign literal_9115[149] = 16'hffb8;
  assign literal_9115[150] = 16'hffc4;
  assign literal_9115[151] = 16'hffd0;
  assign literal_9115[152] = 16'hffdd;
  assign literal_9115[153] = 16'hffea;
  assign literal_9115[154] = 16'hfff8;
  assign literal_9115[155] = 16'h0000;
  assign literal_9115[156] = 16'h0000;
  assign literal_9115[157] = 16'h0000;
  assign literal_9115[158] = 16'h0000;
  assign literal_9115[159] = 16'h0000;
  assign literal_9115[160] = 16'h0000;
  assign literal_9115[161] = 16'h01f6;
  assign literal_9115[162] = 16'h1fec;
  assign literal_9115[163] = 16'hffa5;
  assign literal_9115[164] = 16'hffaf;
  assign literal_9115[165] = 16'hffb9;
  assign literal_9115[166] = 16'hffc5;
  assign literal_9115[167] = 16'hffd1;
  assign literal_9115[168] = 16'hffde;
  assign literal_9115[169] = 16'hffeb;
  assign literal_9115[170] = 16'hfff9;
  assign literal_9115[171] = 16'h0000;
  assign literal_9115[172] = 16'h0000;
  assign literal_9115[173] = 16'h0000;
  assign literal_9115[174] = 16'h0000;
  assign literal_9115[175] = 16'h0000;
  assign literal_9115[176] = 16'h0000;
  assign literal_9115[177] = 16'h01f7;
  assign literal_9115[178] = 16'h1fee;
  assign literal_9115[179] = 16'hffa6;
  assign literal_9115[180] = 16'hffb0;
  assign literal_9115[181] = 16'hffba;
  assign literal_9115[182] = 16'hffc6;
  assign literal_9115[183] = 16'hffd2;
  assign literal_9115[184] = 16'hffdf;
  assign literal_9115[185] = 16'hffec;
  assign literal_9115[186] = 16'hfffa;
  assign literal_9115[187] = 16'h0000;
  assign literal_9115[188] = 16'h0000;
  assign literal_9115[189] = 16'h0000;
  assign literal_9115[190] = 16'h0000;
  assign literal_9115[191] = 16'h0000;
  assign literal_9115[192] = 16'h0000;
  assign literal_9115[193] = 16'h03f4;
  assign literal_9115[194] = 16'h1fef;
  assign literal_9115[195] = 16'hffa7;
  assign literal_9115[196] = 16'hffb1;
  assign literal_9115[197] = 16'hffbb;
  assign literal_9115[198] = 16'hffc7;
  assign literal_9115[199] = 16'hffd3;
  assign literal_9115[200] = 16'hffe0;
  assign literal_9115[201] = 16'hffed;
  assign literal_9115[202] = 16'hfffb;
  assign literal_9115[203] = 16'h0000;
  assign literal_9115[204] = 16'h0000;
  assign literal_9115[205] = 16'h0000;
  assign literal_9115[206] = 16'h0000;
  assign literal_9115[207] = 16'h0000;
  assign literal_9115[208] = 16'h0000;
  assign literal_9115[209] = 16'h03f5;
  assign literal_9115[210] = 16'h3fe2;
  assign literal_9115[211] = 16'hffaa;
  assign literal_9115[212] = 16'hffb2;
  assign literal_9115[213] = 16'hffbc;
  assign literal_9115[214] = 16'hffc8;
  assign literal_9115[215] = 16'hffd4;
  assign literal_9115[216] = 16'hffe1;
  assign literal_9115[217] = 16'hffee;
  assign literal_9115[218] = 16'hfffc;
  assign literal_9115[219] = 16'h0000;
  assign literal_9115[220] = 16'h0000;
  assign literal_9115[221] = 16'h0000;
  assign literal_9115[222] = 16'h0000;
  assign literal_9115[223] = 16'h0000;
  assign literal_9115[224] = 16'h0000;
  assign literal_9115[225] = 16'h03f6;
  assign literal_9115[226] = 16'h7fc7;
  assign literal_9115[227] = 16'hffab;
  assign literal_9115[228] = 16'hffb3;
  assign literal_9115[229] = 16'hffbd;
  assign literal_9115[230] = 16'hffc9;
  assign literal_9115[231] = 16'hffd5;
  assign literal_9115[232] = 16'hffe2;
  assign literal_9115[233] = 16'hffef;
  assign literal_9115[234] = 16'hfffd;
  assign literal_9115[235] = 16'h0000;
  assign literal_9115[236] = 16'h0000;
  assign literal_9115[237] = 16'h0000;
  assign literal_9115[238] = 16'h0000;
  assign literal_9115[239] = 16'h0000;
  assign literal_9115[240] = 16'h01f8;
  assign literal_9115[241] = 16'h07f6;
  assign literal_9115[242] = 16'hffa4;
  assign literal_9115[243] = 16'hffac;
  assign literal_9115[244] = 16'hffb4;
  assign literal_9115[245] = 16'hffbe;
  assign literal_9115[246] = 16'hffca;
  assign literal_9115[247] = 16'hffd6;
  assign literal_9115[248] = 16'hffe3;
  assign literal_9115[249] = 16'hfff0;
  assign literal_9115[250] = 16'hfffe;
  assign literal_9115[251] = 16'h0000;
  wire [15:0] literal_9116[0:251];
  assign literal_9116[0] = 16'h000c;
  assign literal_9116[1] = 16'h0000;
  assign literal_9116[2] = 16'h0001;
  assign literal_9116[3] = 16'h0004;
  assign literal_9116[4] = 16'h000b;
  assign literal_9116[5] = 16'h001a;
  assign literal_9116[6] = 16'h0079;
  assign literal_9116[7] = 16'h01f9;
  assign literal_9116[8] = 16'hff9c;
  assign literal_9116[9] = 16'hff9f;
  assign literal_9116[10] = 16'hffa0;
  assign literal_9116[11] = 16'h0000;
  assign literal_9116[12] = 16'h0000;
  assign literal_9116[13] = 16'h0000;
  assign literal_9116[14] = 16'h0000;
  assign literal_9116[15] = 16'h0000;
  assign literal_9116[16] = 16'h0000;
  assign literal_9116[17] = 16'h000a;
  assign literal_9116[18] = 16'h001c;
  assign literal_9116[19] = 16'h007a;
  assign literal_9116[20] = 16'h01f5;
  assign literal_9116[21] = 16'h03f4;
  assign literal_9116[22] = 16'h07f8;
  assign literal_9116[23] = 16'hff95;
  assign literal_9116[24] = 16'hffa1;
  assign literal_9116[25] = 16'hffa2;
  assign literal_9116[26] = 16'hffad;
  assign literal_9116[27] = 16'h0000;
  assign literal_9116[28] = 16'h0000;
  assign literal_9116[29] = 16'h0000;
  assign literal_9116[30] = 16'h0000;
  assign literal_9116[31] = 16'h0000;
  assign literal_9116[32] = 16'h0000;
  assign literal_9116[33] = 16'h001b;
  assign literal_9116[34] = 16'h00f8;
  assign literal_9116[35] = 16'h03f7;
  assign literal_9116[36] = 16'h0ff4;
  assign literal_9116[37] = 16'h3fdc;
  assign literal_9116[38] = 16'hff9d;
  assign literal_9116[39] = 16'hff90;
  assign literal_9116[40] = 16'hffac;
  assign literal_9116[41] = 16'hffe3;
  assign literal_9116[42] = 16'hfff1;
  assign literal_9116[43] = 16'h0000;
  assign literal_9116[44] = 16'h0000;
  assign literal_9116[45] = 16'h0000;
  assign literal_9116[46] = 16'h0000;
  assign literal_9116[47] = 16'h0000;
  assign literal_9116[48] = 16'h0000;
  assign literal_9116[49] = 16'h003a;
  assign literal_9116[50] = 16'h01f6;
  assign literal_9116[51] = 16'h07f7;
  assign literal_9116[52] = 16'h3fde;
  assign literal_9116[53] = 16'hff8e;
  assign literal_9116[54] = 16'hff94;
  assign literal_9116[55] = 16'hffc9;
  assign literal_9116[56] = 16'hffd6;
  assign literal_9116[57] = 16'hffe4;
  assign literal_9116[58] = 16'hfff2;
  assign literal_9116[59] = 16'h0000;
  assign literal_9116[60] = 16'h0000;
  assign literal_9116[61] = 16'h0000;
  assign literal_9116[62] = 16'h0000;
  assign literal_9116[63] = 16'h0000;
  assign literal_9116[64] = 16'h0000;
  assign literal_9116[65] = 16'h003b;
  assign literal_9116[66] = 16'h03f6;
  assign literal_9116[67] = 16'h3fdd;
  assign literal_9116[68] = 16'hff8f;
  assign literal_9116[69] = 16'hffa5;
  assign literal_9116[70] = 16'hffa6;
  assign literal_9116[71] = 16'hffca;
  assign literal_9116[72] = 16'hffd7;
  assign literal_9116[73] = 16'hffe5;
  assign literal_9116[74] = 16'hfff3;
  assign literal_9116[75] = 16'h0000;
  assign literal_9116[76] = 16'h0000;
  assign literal_9116[77] = 16'h0000;
  assign literal_9116[78] = 16'h0000;
  assign literal_9116[79] = 16'h0000;
  assign literal_9116[80] = 16'h0000;
  assign literal_9116[81] = 16'h0078;
  assign literal_9116[82] = 16'h03f9;
  assign literal_9116[83] = 16'h3fdf;
  assign literal_9116[84] = 16'hff96;
  assign literal_9116[85] = 16'hffab;
  assign literal_9116[86] = 16'hffa9;
  assign literal_9116[87] = 16'hffcb;
  assign literal_9116[88] = 16'hffd8;
  assign literal_9116[89] = 16'hffe6;
  assign literal_9116[90] = 16'hfff4;
  assign literal_9116[91] = 16'h0000;
  assign literal_9116[92] = 16'h0000;
  assign literal_9116[93] = 16'h0000;
  assign literal_9116[94] = 16'h0000;
  assign literal_9116[95] = 16'h0000;
  assign literal_9116[96] = 16'h0000;
  assign literal_9116[97] = 16'h007b;
  assign literal_9116[98] = 16'h0ff2;
  assign literal_9116[99] = 16'h7fc5;
  assign literal_9116[100] = 16'hff97;
  assign literal_9116[101] = 16'hffb5;
  assign literal_9116[102] = 16'hffbf;
  assign literal_9116[103] = 16'hffcc;
  assign literal_9116[104] = 16'hffd9;
  assign literal_9116[105] = 16'hffe7;
  assign literal_9116[106] = 16'hfff5;
  assign literal_9116[107] = 16'h0000;
  assign literal_9116[108] = 16'h0000;
  assign literal_9116[109] = 16'h0000;
  assign literal_9116[110] = 16'h0000;
  assign literal_9116[111] = 16'h0000;
  assign literal_9116[112] = 16'h0000;
  assign literal_9116[113] = 16'h00f9;
  assign literal_9116[114] = 16'h0ff5;
  assign literal_9116[115] = 16'hff8c;
  assign literal_9116[116] = 16'hff98;
  assign literal_9116[117] = 16'hffb6;
  assign literal_9116[118] = 16'hffc0;
  assign literal_9116[119] = 16'hffcd;
  assign literal_9116[120] = 16'hffda;
  assign literal_9116[121] = 16'hffe8;
  assign literal_9116[122] = 16'hfff6;
  assign literal_9116[123] = 16'h0000;
  assign literal_9116[124] = 16'h0000;
  assign literal_9116[125] = 16'h0000;
  assign literal_9116[126] = 16'h0000;
  assign literal_9116[127] = 16'h0000;
  assign literal_9116[128] = 16'h0000;
  assign literal_9116[129] = 16'h01f4;
  assign literal_9116[130] = 16'h1fec;
  assign literal_9116[131] = 16'hff9e;
  assign literal_9116[132] = 16'hffa3;
  assign literal_9116[133] = 16'hffb7;
  assign literal_9116[134] = 16'hffc1;
  assign literal_9116[135] = 16'hffce;
  assign literal_9116[136] = 16'hffdb;
  assign literal_9116[137] = 16'hffe9;
  assign literal_9116[138] = 16'hfff7;
  assign literal_9116[139] = 16'h0000;
  assign literal_9116[140] = 16'h0000;
  assign literal_9116[141] = 16'h0000;
  assign literal_9116[142] = 16'h0000;
  assign literal_9116[143] = 16'h0000;
  assign literal_9116[144] = 16'h0000;
  assign literal_9116[145] = 16'h01f7;
  assign literal_9116[146] = 16'h3fe0;
  assign literal_9116[147] = 16'hff91;
  assign literal_9116[148] = 16'hffa4;
  assign literal_9116[149] = 16'hffb8;
  assign literal_9116[150] = 16'hffc2;
  assign literal_9116[151] = 16'hffcf;
  assign literal_9116[152] = 16'hffdc;
  assign literal_9116[153] = 16'hffea;
  assign literal_9116[154] = 16'hfff8;
  assign literal_9116[155] = 16'h0000;
  assign literal_9116[156] = 16'h0000;
  assign literal_9116[157] = 16'h0000;
  assign literal_9116[158] = 16'h0000;
  assign literal_9116[159] = 16'h0000;
  assign literal_9116[160] = 16'h0000;
  assign literal_9116[161] = 16'h01f8;
  assign literal_9116[162] = 16'h3fe1;
  assign literal_9116[163] = 16'hff92;
  assign literal_9116[164] = 16'hffa7;
  assign literal_9116[165] = 16'hffb9;
  assign literal_9116[166] = 16'hffc3;
  assign literal_9116[167] = 16'hffd0;
  assign literal_9116[168] = 16'hffdd;
  assign literal_9116[169] = 16'hffeb;
  assign literal_9116[170] = 16'hfff9;
  assign literal_9116[171] = 16'h0000;
  assign literal_9116[172] = 16'h0000;
  assign literal_9116[173] = 16'h0000;
  assign literal_9116[174] = 16'h0000;
  assign literal_9116[175] = 16'h0000;
  assign literal_9116[176] = 16'h0000;
  assign literal_9116[177] = 16'h03f5;
  assign literal_9116[178] = 16'h7fc4;
  assign literal_9116[179] = 16'hff93;
  assign literal_9116[180] = 16'hffa8;
  assign literal_9116[181] = 16'hffba;
  assign literal_9116[182] = 16'hffc4;
  assign literal_9116[183] = 16'hffd1;
  assign literal_9116[184] = 16'hffde;
  assign literal_9116[185] = 16'hffec;
  assign literal_9116[186] = 16'hfffa;
  assign literal_9116[187] = 16'h0000;
  assign literal_9116[188] = 16'h0000;
  assign literal_9116[189] = 16'h0000;
  assign literal_9116[190] = 16'h0000;
  assign literal_9116[191] = 16'h0000;
  assign literal_9116[192] = 16'h0000;
  assign literal_9116[193] = 16'h03f8;
  assign literal_9116[194] = 16'hff8d;
  assign literal_9116[195] = 16'hff99;
  assign literal_9116[196] = 16'hffb1;
  assign literal_9116[197] = 16'hffbb;
  assign literal_9116[198] = 16'hffc5;
  assign literal_9116[199] = 16'hffd2;
  assign literal_9116[200] = 16'hffdf;
  assign literal_9116[201] = 16'hffed;
  assign literal_9116[202] = 16'hfffb;
  assign literal_9116[203] = 16'h0000;
  assign literal_9116[204] = 16'h0000;
  assign literal_9116[205] = 16'h0000;
  assign literal_9116[206] = 16'h0000;
  assign literal_9116[207] = 16'h0000;
  assign literal_9116[208] = 16'h0000;
  assign literal_9116[209] = 16'h03fa;
  assign literal_9116[210] = 16'hff9a;
  assign literal_9116[211] = 16'hffaa;
  assign literal_9116[212] = 16'hffb2;
  assign literal_9116[213] = 16'hffbc;
  assign literal_9116[214] = 16'hffc6;
  assign literal_9116[215] = 16'hffd3;
  assign literal_9116[216] = 16'hffe0;
  assign literal_9116[217] = 16'hffee;
  assign literal_9116[218] = 16'hfffc;
  assign literal_9116[219] = 16'h0000;
  assign literal_9116[220] = 16'h0000;
  assign literal_9116[221] = 16'h0000;
  assign literal_9116[222] = 16'h0000;
  assign literal_9116[223] = 16'h0000;
  assign literal_9116[224] = 16'h0000;
  assign literal_9116[225] = 16'h07f6;
  assign literal_9116[226] = 16'hff9b;
  assign literal_9116[227] = 16'hffaf;
  assign literal_9116[228] = 16'hffb3;
  assign literal_9116[229] = 16'hffbd;
  assign literal_9116[230] = 16'hffc7;
  assign literal_9116[231] = 16'hffd4;
  assign literal_9116[232] = 16'hffe1;
  assign literal_9116[233] = 16'hffef;
  assign literal_9116[234] = 16'hfffd;
  assign literal_9116[235] = 16'h0000;
  assign literal_9116[236] = 16'h0000;
  assign literal_9116[237] = 16'h0000;
  assign literal_9116[238] = 16'h0000;
  assign literal_9116[239] = 16'h0000;
  assign literal_9116[240] = 16'h0ff3;
  assign literal_9116[241] = 16'h1fed;
  assign literal_9116[242] = 16'hffae;
  assign literal_9116[243] = 16'hffb0;
  assign literal_9116[244] = 16'hffb4;
  assign literal_9116[245] = 16'hffbe;
  assign literal_9116[246] = 16'hffc8;
  assign literal_9116[247] = 16'hffd5;
  assign literal_9116[248] = 16'hffe2;
  assign literal_9116[249] = 16'hfff0;
  assign literal_9116[250] = 16'hfffe;
  assign literal_9116[251] = 16'h0000;
  wire [9:0] matrix_unflattened[0:7][0:7];
  assign matrix_unflattened[0][0] = matrix[9:0];
  assign matrix_unflattened[0][1] = matrix[19:10];
  assign matrix_unflattened[0][2] = matrix[29:20];
  assign matrix_unflattened[0][3] = matrix[39:30];
  assign matrix_unflattened[0][4] = matrix[49:40];
  assign matrix_unflattened[0][5] = matrix[59:50];
  assign matrix_unflattened[0][6] = matrix[69:60];
  assign matrix_unflattened[0][7] = matrix[79:70];
  assign matrix_unflattened[1][0] = matrix[89:80];
  assign matrix_unflattened[1][1] = matrix[99:90];
  assign matrix_unflattened[1][2] = matrix[109:100];
  assign matrix_unflattened[1][3] = matrix[119:110];
  assign matrix_unflattened[1][4] = matrix[129:120];
  assign matrix_unflattened[1][5] = matrix[139:130];
  assign matrix_unflattened[1][6] = matrix[149:140];
  assign matrix_unflattened[1][7] = matrix[159:150];
  assign matrix_unflattened[2][0] = matrix[169:160];
  assign matrix_unflattened[2][1] = matrix[179:170];
  assign matrix_unflattened[2][2] = matrix[189:180];
  assign matrix_unflattened[2][3] = matrix[199:190];
  assign matrix_unflattened[2][4] = matrix[209:200];
  assign matrix_unflattened[2][5] = matrix[219:210];
  assign matrix_unflattened[2][6] = matrix[229:220];
  assign matrix_unflattened[2][7] = matrix[239:230];
  assign matrix_unflattened[3][0] = matrix[249:240];
  assign matrix_unflattened[3][1] = matrix[259:250];
  assign matrix_unflattened[3][2] = matrix[269:260];
  assign matrix_unflattened[3][3] = matrix[279:270];
  assign matrix_unflattened[3][4] = matrix[289:280];
  assign matrix_unflattened[3][5] = matrix[299:290];
  assign matrix_unflattened[3][6] = matrix[309:300];
  assign matrix_unflattened[3][7] = matrix[319:310];
  assign matrix_unflattened[4][0] = matrix[329:320];
  assign matrix_unflattened[4][1] = matrix[339:330];
  assign matrix_unflattened[4][2] = matrix[349:340];
  assign matrix_unflattened[4][3] = matrix[359:350];
  assign matrix_unflattened[4][4] = matrix[369:360];
  assign matrix_unflattened[4][5] = matrix[379:370];
  assign matrix_unflattened[4][6] = matrix[389:380];
  assign matrix_unflattened[4][7] = matrix[399:390];
  assign matrix_unflattened[5][0] = matrix[409:400];
  assign matrix_unflattened[5][1] = matrix[419:410];
  assign matrix_unflattened[5][2] = matrix[429:420];
  assign matrix_unflattened[5][3] = matrix[439:430];
  assign matrix_unflattened[5][4] = matrix[449:440];
  assign matrix_unflattened[5][5] = matrix[459:450];
  assign matrix_unflattened[5][6] = matrix[469:460];
  assign matrix_unflattened[5][7] = matrix[479:470];
  assign matrix_unflattened[6][0] = matrix[489:480];
  assign matrix_unflattened[6][1] = matrix[499:490];
  assign matrix_unflattened[6][2] = matrix[509:500];
  assign matrix_unflattened[6][3] = matrix[519:510];
  assign matrix_unflattened[6][4] = matrix[529:520];
  assign matrix_unflattened[6][5] = matrix[539:530];
  assign matrix_unflattened[6][6] = matrix[549:540];
  assign matrix_unflattened[6][7] = matrix[559:550];
  assign matrix_unflattened[7][0] = matrix[569:560];
  assign matrix_unflattened[7][1] = matrix[579:570];
  assign matrix_unflattened[7][2] = matrix[589:580];
  assign matrix_unflattened[7][3] = matrix[599:590];
  assign matrix_unflattened[7][4] = matrix[609:600];
  assign matrix_unflattened[7][5] = matrix[619:610];
  assign matrix_unflattened[7][6] = matrix[629:620];
  assign matrix_unflattened[7][7] = matrix[639:630];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [9:0] p0_matrix[0:7][0:7];
  reg [7:0] p0_start_pix;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_matrix[0][0] <= matrix_unflattened[0][0];
    p0_matrix[0][1] <= matrix_unflattened[0][1];
    p0_matrix[0][2] <= matrix_unflattened[0][2];
    p0_matrix[0][3] <= matrix_unflattened[0][3];
    p0_matrix[0][4] <= matrix_unflattened[0][4];
    p0_matrix[0][5] <= matrix_unflattened[0][5];
    p0_matrix[0][6] <= matrix_unflattened[0][6];
    p0_matrix[0][7] <= matrix_unflattened[0][7];
    p0_matrix[1][0] <= matrix_unflattened[1][0];
    p0_matrix[1][1] <= matrix_unflattened[1][1];
    p0_matrix[1][2] <= matrix_unflattened[1][2];
    p0_matrix[1][3] <= matrix_unflattened[1][3];
    p0_matrix[1][4] <= matrix_unflattened[1][4];
    p0_matrix[1][5] <= matrix_unflattened[1][5];
    p0_matrix[1][6] <= matrix_unflattened[1][6];
    p0_matrix[1][7] <= matrix_unflattened[1][7];
    p0_matrix[2][0] <= matrix_unflattened[2][0];
    p0_matrix[2][1] <= matrix_unflattened[2][1];
    p0_matrix[2][2] <= matrix_unflattened[2][2];
    p0_matrix[2][3] <= matrix_unflattened[2][3];
    p0_matrix[2][4] <= matrix_unflattened[2][4];
    p0_matrix[2][5] <= matrix_unflattened[2][5];
    p0_matrix[2][6] <= matrix_unflattened[2][6];
    p0_matrix[2][7] <= matrix_unflattened[2][7];
    p0_matrix[3][0] <= matrix_unflattened[3][0];
    p0_matrix[3][1] <= matrix_unflattened[3][1];
    p0_matrix[3][2] <= matrix_unflattened[3][2];
    p0_matrix[3][3] <= matrix_unflattened[3][3];
    p0_matrix[3][4] <= matrix_unflattened[3][4];
    p0_matrix[3][5] <= matrix_unflattened[3][5];
    p0_matrix[3][6] <= matrix_unflattened[3][6];
    p0_matrix[3][7] <= matrix_unflattened[3][7];
    p0_matrix[4][0] <= matrix_unflattened[4][0];
    p0_matrix[4][1] <= matrix_unflattened[4][1];
    p0_matrix[4][2] <= matrix_unflattened[4][2];
    p0_matrix[4][3] <= matrix_unflattened[4][3];
    p0_matrix[4][4] <= matrix_unflattened[4][4];
    p0_matrix[4][5] <= matrix_unflattened[4][5];
    p0_matrix[4][6] <= matrix_unflattened[4][6];
    p0_matrix[4][7] <= matrix_unflattened[4][7];
    p0_matrix[5][0] <= matrix_unflattened[5][0];
    p0_matrix[5][1] <= matrix_unflattened[5][1];
    p0_matrix[5][2] <= matrix_unflattened[5][2];
    p0_matrix[5][3] <= matrix_unflattened[5][3];
    p0_matrix[5][4] <= matrix_unflattened[5][4];
    p0_matrix[5][5] <= matrix_unflattened[5][5];
    p0_matrix[5][6] <= matrix_unflattened[5][6];
    p0_matrix[5][7] <= matrix_unflattened[5][7];
    p0_matrix[6][0] <= matrix_unflattened[6][0];
    p0_matrix[6][1] <= matrix_unflattened[6][1];
    p0_matrix[6][2] <= matrix_unflattened[6][2];
    p0_matrix[6][3] <= matrix_unflattened[6][3];
    p0_matrix[6][4] <= matrix_unflattened[6][4];
    p0_matrix[6][5] <= matrix_unflattened[6][5];
    p0_matrix[6][6] <= matrix_unflattened[6][6];
    p0_matrix[6][7] <= matrix_unflattened[6][7];
    p0_matrix[7][0] <= matrix_unflattened[7][0];
    p0_matrix[7][1] <= matrix_unflattened[7][1];
    p0_matrix[7][2] <= matrix_unflattened[7][2];
    p0_matrix[7][3] <= matrix_unflattened[7][3];
    p0_matrix[7][4] <= matrix_unflattened[7][4];
    p0_matrix[7][5] <= matrix_unflattened[7][5];
    p0_matrix[7][6] <= matrix_unflattened[7][6];
    p0_matrix[7][7] <= matrix_unflattened[7][7];
    p0_start_pix <= start_pix;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [9:0] p1_row0_comb[0:7];
  wire [9:0] p1_row1_comb[0:7];
  wire [9:0] p1_array_concat_8175_comb[0:15];
  wire [9:0] p1_row2_comb[0:7];
  wire [9:0] p1_array_concat_8178_comb[0:23];
  wire [9:0] p1_row3_comb[0:7];
  wire [2:0] p1_idx_u8__4_squeezed_comb;
  wire [9:0] p1_array_concat_8181_comb[0:31];
  wire [9:0] p1_row4_comb[0:7];
  wire [2:0] p1_idx_u8__5_squeezed_comb;
  wire [9:0] p1_array_concat_8184_comb[0:39];
  wire [9:0] p1_row5_comb[0:7];
  wire [2:0] p1_idx_u8__6_squeezed_comb;
  wire [7:0] p1_idx_u8__1_comb;
  wire [7:0] p1_idx_u8__3_comb;
  wire [7:0] p1_idx_u8__5_comb;
  wire [7:0] p1_idx_u8__7_comb;
  wire [7:0] p1_idx_u8__9_comb;
  wire [7:0] p1_idx_u8__11_comb;
  wire [7:0] p1_idx_u8__13_comb;
  wire [9:0] p1_array_concat_8190_comb[0:47];
  wire [9:0] p1_row6_comb[0:7];
  wire [2:0] p1_idx_u8__7_squeezed_comb;
  wire [6:0] p1_add_8193_comb;
  wire [7:0] p1_actual_index__1_comb;
  wire [6:0] p1_add_8308_comb;
  wire [7:0] p1_actual_index__3_comb;
  wire [5:0] p1_add_8291_comb;
  wire [7:0] p1_actual_index__5_comb;
  wire [6:0] p1_add_8275_comb;
  wire [7:0] p1_actual_index__7_comb;
  wire [7:0] p1_actual_index__9_comb;
  wire [6:0] p1_add_8226_comb;
  wire [7:0] p1_actual_index__11_comb;
  wire [7:0] p1_actual_index__13_comb;
  wire [7:0] p1_idx_u8__15_comb;
  wire [7:0] p1_idx_u8__17_comb;
  wire [7:0] p1_idx_u8__19_comb;
  wire [7:0] p1_idx_u8__21_comb;
  wire [7:0] p1_idx_u8__23_comb;
  wire [7:0] p1_idx_u8__25_comb;
  wire [7:0] p1_idx_u8__27_comb;
  wire [7:0] p1_idx_u8__29_comb;
  wire [7:0] p1_idx_u8__31_comb;
  wire [7:0] p1_idx_u8__33_comb;
  wire [7:0] p1_idx_u8__35_comb;
  wire [7:0] p1_idx_u8__37_comb;
  wire [7:0] p1_idx_u8__39_comb;
  wire [7:0] p1_idx_u8__41_comb;
  wire [7:0] p1_idx_u8__43_comb;
  wire [7:0] p1_idx_u8__45_comb;
  wire [7:0] p1_idx_u8__47_comb;
  wire [7:0] p1_idx_u8__49_comb;
  wire [7:0] p1_idx_u8__51_comb;
  wire [7:0] p1_idx_u8__53_comb;
  wire [7:0] p1_idx_u8__55_comb;
  wire [7:0] p1_idx_u8__57_comb;
  wire [7:0] p1_idx_u8__59_comb;
  wire [7:0] p1_idx_u8__61_comb;
  wire [9:0] p1_array_concat_8197_comb[0:55];
  wire [9:0] p1_row7_comb[0:7];
  wire [5:0] p1_add_8202_comb;
  wire [4:0] p1_add_8245_comb;
  wire [7:0] p1_actual_index__15_comb;
  wire [3:0] p1_add_8411_comb;
  wire [7:0] p1_actual_index__17_comb;
  wire [6:0] p1_add_8413_comb;
  wire [7:0] p1_actual_index__19_comb;
  wire [5:0] p1_add_8415_comb;
  wire [7:0] p1_actual_index__21_comb;
  wire [6:0] p1_add_8417_comb;
  wire [7:0] p1_actual_index__23_comb;
  wire [4:0] p1_add_8419_comb;
  wire [7:0] p1_actual_index__25_comb;
  wire [6:0] p1_add_8421_comb;
  wire [7:0] p1_actual_index__27_comb;
  wire [5:0] p1_add_8423_comb;
  wire [7:0] p1_actual_index__29_comb;
  wire [6:0] p1_add_8425_comb;
  wire [7:0] p1_actual_index__31_comb;
  wire [2:0] p1_add_8427_comb;
  wire [7:0] p1_actual_index__33_comb;
  wire [6:0] p1_add_8429_comb;
  wire [7:0] p1_actual_index__35_comb;
  wire [5:0] p1_add_8431_comb;
  wire [7:0] p1_actual_index__37_comb;
  wire [6:0] p1_add_8433_comb;
  wire [7:0] p1_actual_index__39_comb;
  wire [4:0] p1_add_8435_comb;
  wire [7:0] p1_actual_index__41_comb;
  wire [6:0] p1_add_8437_comb;
  wire [7:0] p1_actual_index__43_comb;
  wire [5:0] p1_add_8439_comb;
  wire [7:0] p1_actual_index__45_comb;
  wire [6:0] p1_add_8441_comb;
  wire [7:0] p1_actual_index__47_comb;
  wire [3:0] p1_add_8443_comb;
  wire [7:0] p1_actual_index__49_comb;
  wire [6:0] p1_add_8445_comb;
  wire [7:0] p1_actual_index__51_comb;
  wire [5:0] p1_add_8447_comb;
  wire [7:0] p1_actual_index__53_comb;
  wire [6:0] p1_add_8449_comb;
  wire [7:0] p1_actual_index__55_comb;
  wire [4:0] p1_add_8451_comb;
  wire [7:0] p1_actual_index__57_comb;
  wire [6:0] p1_add_8453_comb;
  wire [7:0] p1_actual_index__59_comb;
  wire [5:0] p1_add_8455_comb;
  wire [7:0] p1_actual_index__61_comb;
  wire [6:0] p1_add_8457_comb;
  wire [9:0] p1_flat_comb[0:63];
  wire [7:0] p1_actual_index__14_comb;
  wire [7:0] p1_actual_index__2_comb;
  wire [7:0] p1_actual_index__4_comb;
  wire [7:0] p1_actual_index__6_comb;
  wire [7:0] p1_actual_index__10_comb;
  wire [7:0] p1_actual_index__12_comb;
  wire [7:0] p1_actual_index__8_comb;
  wire [7:0] p1_actual_index__16_comb;
  wire [7:0] p1_actual_index__18_comb;
  wire [7:0] p1_actual_index__20_comb;
  wire [7:0] p1_actual_index__22_comb;
  wire [7:0] p1_actual_index__24_comb;
  wire [7:0] p1_actual_index__26_comb;
  wire [7:0] p1_actual_index__28_comb;
  wire [7:0] p1_actual_index__30_comb;
  wire [7:0] p1_actual_index__32_comb;
  wire [7:0] p1_actual_index__34_comb;
  wire [7:0] p1_actual_index__36_comb;
  wire [7:0] p1_actual_index__38_comb;
  wire [7:0] p1_actual_index__40_comb;
  wire [7:0] p1_actual_index__42_comb;
  wire [7:0] p1_actual_index__44_comb;
  wire [7:0] p1_actual_index__46_comb;
  wire [7:0] p1_actual_index__48_comb;
  wire [7:0] p1_actual_index__50_comb;
  wire [7:0] p1_actual_index__52_comb;
  wire [7:0] p1_actual_index__54_comb;
  wire [7:0] p1_actual_index__56_comb;
  wire [7:0] p1_actual_index__58_comb;
  wire [7:0] p1_actual_index__60_comb;
  wire [7:0] p1_actual_index__62_comb;
  wire [9:0] p1_and_8221_comb;
  wire [9:0] p1_and_8352_comb;
  wire [9:0] p1_and_8354_comb;
  wire [9:0] p1_and_8349_comb;
  wire [9:0] p1_and_8342_comb;
  wire [9:0] p1_and_8335_comb;
  wire [9:0] p1_and_8324_comb;
  wire [9:0] p1_and_8315_comb;
  wire [9:0] p1_and_8305_comb;
  wire [9:0] p1_and_8278_comb;
  wire [9:0] p1_and_8269_comb;
  wire [9:0] p1_and_8261_comb;
  wire [9:0] p1_and_8229_comb;
  wire p1_eq_8232_comb;
  wire [9:0] p1_and_8233_comb;
  wire p1_ne_8357_comb;
  wire p1_ne_8358_comb;
  wire p1_ne_8356_comb;
  wire p1_ne_8351_comb;
  wire p1_ne_8344_comb;
  wire p1_ne_8337_comb;
  wire p1_ne_8326_comb;
  wire p1_ne_8317_comb;
  wire [9:0] p1_and_8281_comb;
  wire p1_ne_8288_comb;
  wire p1_ne_8280_comb;
  wire p1_ne_8271_comb;
  wire p1_ne_8241_comb;
  wire [9:0] p1_value_comb;
  wire [1:0] p1_idx_u8__1_squeezed_comb;
  wire p1_eq_8244_comb;
  wire p1_not_8359_comb;
  wire p1_eq_8289_comb;
  wire [7:0] p1_bin_value__1_comb;
  wire [7:0] p1_flipped_comb;
  wire [1:0] p1_sel_8252_comb;
  wire [1:0] p1_sign_ext_8253_comb;
  wire p1_and_8883_comb;
  wire [7:0] p1_code_list_comb;
  assign p1_row0_comb[0] = p0_matrix[3'h0][0];
  assign p1_row0_comb[1] = p0_matrix[3'h0][1];
  assign p1_row0_comb[2] = p0_matrix[3'h0][2];
  assign p1_row0_comb[3] = p0_matrix[3'h0][3];
  assign p1_row0_comb[4] = p0_matrix[3'h0][4];
  assign p1_row0_comb[5] = p0_matrix[3'h0][5];
  assign p1_row0_comb[6] = p0_matrix[3'h0][6];
  assign p1_row0_comb[7] = p0_matrix[3'h0][7];
  assign p1_row1_comb[0] = p0_matrix[3'h1][0];
  assign p1_row1_comb[1] = p0_matrix[3'h1][1];
  assign p1_row1_comb[2] = p0_matrix[3'h1][2];
  assign p1_row1_comb[3] = p0_matrix[3'h1][3];
  assign p1_row1_comb[4] = p0_matrix[3'h1][4];
  assign p1_row1_comb[5] = p0_matrix[3'h1][5];
  assign p1_row1_comb[6] = p0_matrix[3'h1][6];
  assign p1_row1_comb[7] = p0_matrix[3'h1][7];
  assign p1_array_concat_8175_comb[0] = p1_row0_comb[0];
  assign p1_array_concat_8175_comb[1] = p1_row0_comb[1];
  assign p1_array_concat_8175_comb[2] = p1_row0_comb[2];
  assign p1_array_concat_8175_comb[3] = p1_row0_comb[3];
  assign p1_array_concat_8175_comb[4] = p1_row0_comb[4];
  assign p1_array_concat_8175_comb[5] = p1_row0_comb[5];
  assign p1_array_concat_8175_comb[6] = p1_row0_comb[6];
  assign p1_array_concat_8175_comb[7] = p1_row0_comb[7];
  assign p1_array_concat_8175_comb[8] = p1_row1_comb[0];
  assign p1_array_concat_8175_comb[9] = p1_row1_comb[1];
  assign p1_array_concat_8175_comb[10] = p1_row1_comb[2];
  assign p1_array_concat_8175_comb[11] = p1_row1_comb[3];
  assign p1_array_concat_8175_comb[12] = p1_row1_comb[4];
  assign p1_array_concat_8175_comb[13] = p1_row1_comb[5];
  assign p1_array_concat_8175_comb[14] = p1_row1_comb[6];
  assign p1_array_concat_8175_comb[15] = p1_row1_comb[7];
  assign p1_row2_comb[0] = p0_matrix[3'h2][0];
  assign p1_row2_comb[1] = p0_matrix[3'h2][1];
  assign p1_row2_comb[2] = p0_matrix[3'h2][2];
  assign p1_row2_comb[3] = p0_matrix[3'h2][3];
  assign p1_row2_comb[4] = p0_matrix[3'h2][4];
  assign p1_row2_comb[5] = p0_matrix[3'h2][5];
  assign p1_row2_comb[6] = p0_matrix[3'h2][6];
  assign p1_row2_comb[7] = p0_matrix[3'h2][7];
  assign p1_array_concat_8178_comb[0] = p1_array_concat_8175_comb[0];
  assign p1_array_concat_8178_comb[1] = p1_array_concat_8175_comb[1];
  assign p1_array_concat_8178_comb[2] = p1_array_concat_8175_comb[2];
  assign p1_array_concat_8178_comb[3] = p1_array_concat_8175_comb[3];
  assign p1_array_concat_8178_comb[4] = p1_array_concat_8175_comb[4];
  assign p1_array_concat_8178_comb[5] = p1_array_concat_8175_comb[5];
  assign p1_array_concat_8178_comb[6] = p1_array_concat_8175_comb[6];
  assign p1_array_concat_8178_comb[7] = p1_array_concat_8175_comb[7];
  assign p1_array_concat_8178_comb[8] = p1_array_concat_8175_comb[8];
  assign p1_array_concat_8178_comb[9] = p1_array_concat_8175_comb[9];
  assign p1_array_concat_8178_comb[10] = p1_array_concat_8175_comb[10];
  assign p1_array_concat_8178_comb[11] = p1_array_concat_8175_comb[11];
  assign p1_array_concat_8178_comb[12] = p1_array_concat_8175_comb[12];
  assign p1_array_concat_8178_comb[13] = p1_array_concat_8175_comb[13];
  assign p1_array_concat_8178_comb[14] = p1_array_concat_8175_comb[14];
  assign p1_array_concat_8178_comb[15] = p1_array_concat_8175_comb[15];
  assign p1_array_concat_8178_comb[16] = p1_row2_comb[0];
  assign p1_array_concat_8178_comb[17] = p1_row2_comb[1];
  assign p1_array_concat_8178_comb[18] = p1_row2_comb[2];
  assign p1_array_concat_8178_comb[19] = p1_row2_comb[3];
  assign p1_array_concat_8178_comb[20] = p1_row2_comb[4];
  assign p1_array_concat_8178_comb[21] = p1_row2_comb[5];
  assign p1_array_concat_8178_comb[22] = p1_row2_comb[6];
  assign p1_array_concat_8178_comb[23] = p1_row2_comb[7];
  assign p1_row3_comb[0] = p0_matrix[3'h3][0];
  assign p1_row3_comb[1] = p0_matrix[3'h3][1];
  assign p1_row3_comb[2] = p0_matrix[3'h3][2];
  assign p1_row3_comb[3] = p0_matrix[3'h3][3];
  assign p1_row3_comb[4] = p0_matrix[3'h3][4];
  assign p1_row3_comb[5] = p0_matrix[3'h3][5];
  assign p1_row3_comb[6] = p0_matrix[3'h3][6];
  assign p1_row3_comb[7] = p0_matrix[3'h3][7];
  assign p1_idx_u8__4_squeezed_comb = 3'h4;
  assign p1_array_concat_8181_comb[0] = p1_array_concat_8178_comb[0];
  assign p1_array_concat_8181_comb[1] = p1_array_concat_8178_comb[1];
  assign p1_array_concat_8181_comb[2] = p1_array_concat_8178_comb[2];
  assign p1_array_concat_8181_comb[3] = p1_array_concat_8178_comb[3];
  assign p1_array_concat_8181_comb[4] = p1_array_concat_8178_comb[4];
  assign p1_array_concat_8181_comb[5] = p1_array_concat_8178_comb[5];
  assign p1_array_concat_8181_comb[6] = p1_array_concat_8178_comb[6];
  assign p1_array_concat_8181_comb[7] = p1_array_concat_8178_comb[7];
  assign p1_array_concat_8181_comb[8] = p1_array_concat_8178_comb[8];
  assign p1_array_concat_8181_comb[9] = p1_array_concat_8178_comb[9];
  assign p1_array_concat_8181_comb[10] = p1_array_concat_8178_comb[10];
  assign p1_array_concat_8181_comb[11] = p1_array_concat_8178_comb[11];
  assign p1_array_concat_8181_comb[12] = p1_array_concat_8178_comb[12];
  assign p1_array_concat_8181_comb[13] = p1_array_concat_8178_comb[13];
  assign p1_array_concat_8181_comb[14] = p1_array_concat_8178_comb[14];
  assign p1_array_concat_8181_comb[15] = p1_array_concat_8178_comb[15];
  assign p1_array_concat_8181_comb[16] = p1_array_concat_8178_comb[16];
  assign p1_array_concat_8181_comb[17] = p1_array_concat_8178_comb[17];
  assign p1_array_concat_8181_comb[18] = p1_array_concat_8178_comb[18];
  assign p1_array_concat_8181_comb[19] = p1_array_concat_8178_comb[19];
  assign p1_array_concat_8181_comb[20] = p1_array_concat_8178_comb[20];
  assign p1_array_concat_8181_comb[21] = p1_array_concat_8178_comb[21];
  assign p1_array_concat_8181_comb[22] = p1_array_concat_8178_comb[22];
  assign p1_array_concat_8181_comb[23] = p1_array_concat_8178_comb[23];
  assign p1_array_concat_8181_comb[24] = p1_row3_comb[0];
  assign p1_array_concat_8181_comb[25] = p1_row3_comb[1];
  assign p1_array_concat_8181_comb[26] = p1_row3_comb[2];
  assign p1_array_concat_8181_comb[27] = p1_row3_comb[3];
  assign p1_array_concat_8181_comb[28] = p1_row3_comb[4];
  assign p1_array_concat_8181_comb[29] = p1_row3_comb[5];
  assign p1_array_concat_8181_comb[30] = p1_row3_comb[6];
  assign p1_array_concat_8181_comb[31] = p1_row3_comb[7];
  assign p1_row4_comb[0] = p0_matrix[p1_idx_u8__4_squeezed_comb][0];
  assign p1_row4_comb[1] = p0_matrix[p1_idx_u8__4_squeezed_comb][1];
  assign p1_row4_comb[2] = p0_matrix[p1_idx_u8__4_squeezed_comb][2];
  assign p1_row4_comb[3] = p0_matrix[p1_idx_u8__4_squeezed_comb][3];
  assign p1_row4_comb[4] = p0_matrix[p1_idx_u8__4_squeezed_comb][4];
  assign p1_row4_comb[5] = p0_matrix[p1_idx_u8__4_squeezed_comb][5];
  assign p1_row4_comb[6] = p0_matrix[p1_idx_u8__4_squeezed_comb][6];
  assign p1_row4_comb[7] = p0_matrix[p1_idx_u8__4_squeezed_comb][7];
  assign p1_idx_u8__5_squeezed_comb = 3'h5;
  assign p1_array_concat_8184_comb[0] = p1_array_concat_8181_comb[0];
  assign p1_array_concat_8184_comb[1] = p1_array_concat_8181_comb[1];
  assign p1_array_concat_8184_comb[2] = p1_array_concat_8181_comb[2];
  assign p1_array_concat_8184_comb[3] = p1_array_concat_8181_comb[3];
  assign p1_array_concat_8184_comb[4] = p1_array_concat_8181_comb[4];
  assign p1_array_concat_8184_comb[5] = p1_array_concat_8181_comb[5];
  assign p1_array_concat_8184_comb[6] = p1_array_concat_8181_comb[6];
  assign p1_array_concat_8184_comb[7] = p1_array_concat_8181_comb[7];
  assign p1_array_concat_8184_comb[8] = p1_array_concat_8181_comb[8];
  assign p1_array_concat_8184_comb[9] = p1_array_concat_8181_comb[9];
  assign p1_array_concat_8184_comb[10] = p1_array_concat_8181_comb[10];
  assign p1_array_concat_8184_comb[11] = p1_array_concat_8181_comb[11];
  assign p1_array_concat_8184_comb[12] = p1_array_concat_8181_comb[12];
  assign p1_array_concat_8184_comb[13] = p1_array_concat_8181_comb[13];
  assign p1_array_concat_8184_comb[14] = p1_array_concat_8181_comb[14];
  assign p1_array_concat_8184_comb[15] = p1_array_concat_8181_comb[15];
  assign p1_array_concat_8184_comb[16] = p1_array_concat_8181_comb[16];
  assign p1_array_concat_8184_comb[17] = p1_array_concat_8181_comb[17];
  assign p1_array_concat_8184_comb[18] = p1_array_concat_8181_comb[18];
  assign p1_array_concat_8184_comb[19] = p1_array_concat_8181_comb[19];
  assign p1_array_concat_8184_comb[20] = p1_array_concat_8181_comb[20];
  assign p1_array_concat_8184_comb[21] = p1_array_concat_8181_comb[21];
  assign p1_array_concat_8184_comb[22] = p1_array_concat_8181_comb[22];
  assign p1_array_concat_8184_comb[23] = p1_array_concat_8181_comb[23];
  assign p1_array_concat_8184_comb[24] = p1_array_concat_8181_comb[24];
  assign p1_array_concat_8184_comb[25] = p1_array_concat_8181_comb[25];
  assign p1_array_concat_8184_comb[26] = p1_array_concat_8181_comb[26];
  assign p1_array_concat_8184_comb[27] = p1_array_concat_8181_comb[27];
  assign p1_array_concat_8184_comb[28] = p1_array_concat_8181_comb[28];
  assign p1_array_concat_8184_comb[29] = p1_array_concat_8181_comb[29];
  assign p1_array_concat_8184_comb[30] = p1_array_concat_8181_comb[30];
  assign p1_array_concat_8184_comb[31] = p1_array_concat_8181_comb[31];
  assign p1_array_concat_8184_comb[32] = p1_row4_comb[0];
  assign p1_array_concat_8184_comb[33] = p1_row4_comb[1];
  assign p1_array_concat_8184_comb[34] = p1_row4_comb[2];
  assign p1_array_concat_8184_comb[35] = p1_row4_comb[3];
  assign p1_array_concat_8184_comb[36] = p1_row4_comb[4];
  assign p1_array_concat_8184_comb[37] = p1_row4_comb[5];
  assign p1_array_concat_8184_comb[38] = p1_row4_comb[6];
  assign p1_array_concat_8184_comb[39] = p1_row4_comb[7];
  assign p1_row5_comb[0] = p0_matrix[p1_idx_u8__5_squeezed_comb][0];
  assign p1_row5_comb[1] = p0_matrix[p1_idx_u8__5_squeezed_comb][1];
  assign p1_row5_comb[2] = p0_matrix[p1_idx_u8__5_squeezed_comb][2];
  assign p1_row5_comb[3] = p0_matrix[p1_idx_u8__5_squeezed_comb][3];
  assign p1_row5_comb[4] = p0_matrix[p1_idx_u8__5_squeezed_comb][4];
  assign p1_row5_comb[5] = p0_matrix[p1_idx_u8__5_squeezed_comb][5];
  assign p1_row5_comb[6] = p0_matrix[p1_idx_u8__5_squeezed_comb][6];
  assign p1_row5_comb[7] = p0_matrix[p1_idx_u8__5_squeezed_comb][7];
  assign p1_idx_u8__6_squeezed_comb = 3'h6;
  assign p1_idx_u8__1_comb = 8'h01;
  assign p1_idx_u8__3_comb = 8'h03;
  assign p1_idx_u8__5_comb = 8'h05;
  assign p1_idx_u8__7_comb = 8'h07;
  assign p1_idx_u8__9_comb = 8'h09;
  assign p1_idx_u8__11_comb = 8'h0b;
  assign p1_idx_u8__13_comb = 8'h0d;
  assign p1_array_concat_8190_comb[0] = p1_array_concat_8184_comb[0];
  assign p1_array_concat_8190_comb[1] = p1_array_concat_8184_comb[1];
  assign p1_array_concat_8190_comb[2] = p1_array_concat_8184_comb[2];
  assign p1_array_concat_8190_comb[3] = p1_array_concat_8184_comb[3];
  assign p1_array_concat_8190_comb[4] = p1_array_concat_8184_comb[4];
  assign p1_array_concat_8190_comb[5] = p1_array_concat_8184_comb[5];
  assign p1_array_concat_8190_comb[6] = p1_array_concat_8184_comb[6];
  assign p1_array_concat_8190_comb[7] = p1_array_concat_8184_comb[7];
  assign p1_array_concat_8190_comb[8] = p1_array_concat_8184_comb[8];
  assign p1_array_concat_8190_comb[9] = p1_array_concat_8184_comb[9];
  assign p1_array_concat_8190_comb[10] = p1_array_concat_8184_comb[10];
  assign p1_array_concat_8190_comb[11] = p1_array_concat_8184_comb[11];
  assign p1_array_concat_8190_comb[12] = p1_array_concat_8184_comb[12];
  assign p1_array_concat_8190_comb[13] = p1_array_concat_8184_comb[13];
  assign p1_array_concat_8190_comb[14] = p1_array_concat_8184_comb[14];
  assign p1_array_concat_8190_comb[15] = p1_array_concat_8184_comb[15];
  assign p1_array_concat_8190_comb[16] = p1_array_concat_8184_comb[16];
  assign p1_array_concat_8190_comb[17] = p1_array_concat_8184_comb[17];
  assign p1_array_concat_8190_comb[18] = p1_array_concat_8184_comb[18];
  assign p1_array_concat_8190_comb[19] = p1_array_concat_8184_comb[19];
  assign p1_array_concat_8190_comb[20] = p1_array_concat_8184_comb[20];
  assign p1_array_concat_8190_comb[21] = p1_array_concat_8184_comb[21];
  assign p1_array_concat_8190_comb[22] = p1_array_concat_8184_comb[22];
  assign p1_array_concat_8190_comb[23] = p1_array_concat_8184_comb[23];
  assign p1_array_concat_8190_comb[24] = p1_array_concat_8184_comb[24];
  assign p1_array_concat_8190_comb[25] = p1_array_concat_8184_comb[25];
  assign p1_array_concat_8190_comb[26] = p1_array_concat_8184_comb[26];
  assign p1_array_concat_8190_comb[27] = p1_array_concat_8184_comb[27];
  assign p1_array_concat_8190_comb[28] = p1_array_concat_8184_comb[28];
  assign p1_array_concat_8190_comb[29] = p1_array_concat_8184_comb[29];
  assign p1_array_concat_8190_comb[30] = p1_array_concat_8184_comb[30];
  assign p1_array_concat_8190_comb[31] = p1_array_concat_8184_comb[31];
  assign p1_array_concat_8190_comb[32] = p1_array_concat_8184_comb[32];
  assign p1_array_concat_8190_comb[33] = p1_array_concat_8184_comb[33];
  assign p1_array_concat_8190_comb[34] = p1_array_concat_8184_comb[34];
  assign p1_array_concat_8190_comb[35] = p1_array_concat_8184_comb[35];
  assign p1_array_concat_8190_comb[36] = p1_array_concat_8184_comb[36];
  assign p1_array_concat_8190_comb[37] = p1_array_concat_8184_comb[37];
  assign p1_array_concat_8190_comb[38] = p1_array_concat_8184_comb[38];
  assign p1_array_concat_8190_comb[39] = p1_array_concat_8184_comb[39];
  assign p1_array_concat_8190_comb[40] = p1_row5_comb[0];
  assign p1_array_concat_8190_comb[41] = p1_row5_comb[1];
  assign p1_array_concat_8190_comb[42] = p1_row5_comb[2];
  assign p1_array_concat_8190_comb[43] = p1_row5_comb[3];
  assign p1_array_concat_8190_comb[44] = p1_row5_comb[4];
  assign p1_array_concat_8190_comb[45] = p1_row5_comb[5];
  assign p1_array_concat_8190_comb[46] = p1_row5_comb[6];
  assign p1_array_concat_8190_comb[47] = p1_row5_comb[7];
  assign p1_row6_comb[0] = p0_matrix[p1_idx_u8__6_squeezed_comb][0];
  assign p1_row6_comb[1] = p0_matrix[p1_idx_u8__6_squeezed_comb][1];
  assign p1_row6_comb[2] = p0_matrix[p1_idx_u8__6_squeezed_comb][2];
  assign p1_row6_comb[3] = p0_matrix[p1_idx_u8__6_squeezed_comb][3];
  assign p1_row6_comb[4] = p0_matrix[p1_idx_u8__6_squeezed_comb][4];
  assign p1_row6_comb[5] = p0_matrix[p1_idx_u8__6_squeezed_comb][5];
  assign p1_row6_comb[6] = p0_matrix[p1_idx_u8__6_squeezed_comb][6];
  assign p1_row6_comb[7] = p0_matrix[p1_idx_u8__6_squeezed_comb][7];
  assign p1_idx_u8__7_squeezed_comb = 3'h7;
  assign p1_add_8193_comb = p0_start_pix[7:1] + 7'h07;
  assign p1_actual_index__1_comb = p0_start_pix + p1_idx_u8__1_comb;
  assign p1_add_8308_comb = p0_start_pix[7:1] + 7'h01;
  assign p1_actual_index__3_comb = p0_start_pix + p1_idx_u8__3_comb;
  assign p1_add_8291_comb = p0_start_pix[7:2] + 6'h01;
  assign p1_actual_index__5_comb = p0_start_pix + p1_idx_u8__5_comb;
  assign p1_add_8275_comb = p0_start_pix[7:1] + 7'h03;
  assign p1_actual_index__7_comb = p0_start_pix + p1_idx_u8__7_comb;
  assign p1_actual_index__9_comb = p0_start_pix + p1_idx_u8__9_comb;
  assign p1_add_8226_comb = p0_start_pix[7:1] + 7'h05;
  assign p1_actual_index__11_comb = p0_start_pix + p1_idx_u8__11_comb;
  assign p1_actual_index__13_comb = p0_start_pix + p1_idx_u8__13_comb;
  assign p1_idx_u8__15_comb = 8'h0f;
  assign p1_idx_u8__17_comb = 8'h11;
  assign p1_idx_u8__19_comb = 8'h13;
  assign p1_idx_u8__21_comb = 8'h15;
  assign p1_idx_u8__23_comb = 8'h17;
  assign p1_idx_u8__25_comb = 8'h19;
  assign p1_idx_u8__27_comb = 8'h1b;
  assign p1_idx_u8__29_comb = 8'h1d;
  assign p1_idx_u8__31_comb = 8'h1f;
  assign p1_idx_u8__33_comb = 8'h21;
  assign p1_idx_u8__35_comb = 8'h23;
  assign p1_idx_u8__37_comb = 8'h25;
  assign p1_idx_u8__39_comb = 8'h27;
  assign p1_idx_u8__41_comb = 8'h29;
  assign p1_idx_u8__43_comb = 8'h2b;
  assign p1_idx_u8__45_comb = 8'h2d;
  assign p1_idx_u8__47_comb = 8'h2f;
  assign p1_idx_u8__49_comb = 8'h31;
  assign p1_idx_u8__51_comb = 8'h33;
  assign p1_idx_u8__53_comb = 8'h35;
  assign p1_idx_u8__55_comb = 8'h37;
  assign p1_idx_u8__57_comb = 8'h39;
  assign p1_idx_u8__59_comb = 8'h3b;
  assign p1_idx_u8__61_comb = 8'h3d;
  assign p1_array_concat_8197_comb[0] = p1_array_concat_8190_comb[0];
  assign p1_array_concat_8197_comb[1] = p1_array_concat_8190_comb[1];
  assign p1_array_concat_8197_comb[2] = p1_array_concat_8190_comb[2];
  assign p1_array_concat_8197_comb[3] = p1_array_concat_8190_comb[3];
  assign p1_array_concat_8197_comb[4] = p1_array_concat_8190_comb[4];
  assign p1_array_concat_8197_comb[5] = p1_array_concat_8190_comb[5];
  assign p1_array_concat_8197_comb[6] = p1_array_concat_8190_comb[6];
  assign p1_array_concat_8197_comb[7] = p1_array_concat_8190_comb[7];
  assign p1_array_concat_8197_comb[8] = p1_array_concat_8190_comb[8];
  assign p1_array_concat_8197_comb[9] = p1_array_concat_8190_comb[9];
  assign p1_array_concat_8197_comb[10] = p1_array_concat_8190_comb[10];
  assign p1_array_concat_8197_comb[11] = p1_array_concat_8190_comb[11];
  assign p1_array_concat_8197_comb[12] = p1_array_concat_8190_comb[12];
  assign p1_array_concat_8197_comb[13] = p1_array_concat_8190_comb[13];
  assign p1_array_concat_8197_comb[14] = p1_array_concat_8190_comb[14];
  assign p1_array_concat_8197_comb[15] = p1_array_concat_8190_comb[15];
  assign p1_array_concat_8197_comb[16] = p1_array_concat_8190_comb[16];
  assign p1_array_concat_8197_comb[17] = p1_array_concat_8190_comb[17];
  assign p1_array_concat_8197_comb[18] = p1_array_concat_8190_comb[18];
  assign p1_array_concat_8197_comb[19] = p1_array_concat_8190_comb[19];
  assign p1_array_concat_8197_comb[20] = p1_array_concat_8190_comb[20];
  assign p1_array_concat_8197_comb[21] = p1_array_concat_8190_comb[21];
  assign p1_array_concat_8197_comb[22] = p1_array_concat_8190_comb[22];
  assign p1_array_concat_8197_comb[23] = p1_array_concat_8190_comb[23];
  assign p1_array_concat_8197_comb[24] = p1_array_concat_8190_comb[24];
  assign p1_array_concat_8197_comb[25] = p1_array_concat_8190_comb[25];
  assign p1_array_concat_8197_comb[26] = p1_array_concat_8190_comb[26];
  assign p1_array_concat_8197_comb[27] = p1_array_concat_8190_comb[27];
  assign p1_array_concat_8197_comb[28] = p1_array_concat_8190_comb[28];
  assign p1_array_concat_8197_comb[29] = p1_array_concat_8190_comb[29];
  assign p1_array_concat_8197_comb[30] = p1_array_concat_8190_comb[30];
  assign p1_array_concat_8197_comb[31] = p1_array_concat_8190_comb[31];
  assign p1_array_concat_8197_comb[32] = p1_array_concat_8190_comb[32];
  assign p1_array_concat_8197_comb[33] = p1_array_concat_8190_comb[33];
  assign p1_array_concat_8197_comb[34] = p1_array_concat_8190_comb[34];
  assign p1_array_concat_8197_comb[35] = p1_array_concat_8190_comb[35];
  assign p1_array_concat_8197_comb[36] = p1_array_concat_8190_comb[36];
  assign p1_array_concat_8197_comb[37] = p1_array_concat_8190_comb[37];
  assign p1_array_concat_8197_comb[38] = p1_array_concat_8190_comb[38];
  assign p1_array_concat_8197_comb[39] = p1_array_concat_8190_comb[39];
  assign p1_array_concat_8197_comb[40] = p1_array_concat_8190_comb[40];
  assign p1_array_concat_8197_comb[41] = p1_array_concat_8190_comb[41];
  assign p1_array_concat_8197_comb[42] = p1_array_concat_8190_comb[42];
  assign p1_array_concat_8197_comb[43] = p1_array_concat_8190_comb[43];
  assign p1_array_concat_8197_comb[44] = p1_array_concat_8190_comb[44];
  assign p1_array_concat_8197_comb[45] = p1_array_concat_8190_comb[45];
  assign p1_array_concat_8197_comb[46] = p1_array_concat_8190_comb[46];
  assign p1_array_concat_8197_comb[47] = p1_array_concat_8190_comb[47];
  assign p1_array_concat_8197_comb[48] = p1_row6_comb[0];
  assign p1_array_concat_8197_comb[49] = p1_row6_comb[1];
  assign p1_array_concat_8197_comb[50] = p1_row6_comb[2];
  assign p1_array_concat_8197_comb[51] = p1_row6_comb[3];
  assign p1_array_concat_8197_comb[52] = p1_row6_comb[4];
  assign p1_array_concat_8197_comb[53] = p1_row6_comb[5];
  assign p1_array_concat_8197_comb[54] = p1_row6_comb[6];
  assign p1_array_concat_8197_comb[55] = p1_row6_comb[7];
  assign p1_row7_comb[0] = p0_matrix[p1_idx_u8__7_squeezed_comb][0];
  assign p1_row7_comb[1] = p0_matrix[p1_idx_u8__7_squeezed_comb][1];
  assign p1_row7_comb[2] = p0_matrix[p1_idx_u8__7_squeezed_comb][2];
  assign p1_row7_comb[3] = p0_matrix[p1_idx_u8__7_squeezed_comb][3];
  assign p1_row7_comb[4] = p0_matrix[p1_idx_u8__7_squeezed_comb][4];
  assign p1_row7_comb[5] = p0_matrix[p1_idx_u8__7_squeezed_comb][5];
  assign p1_row7_comb[6] = p0_matrix[p1_idx_u8__7_squeezed_comb][6];
  assign p1_row7_comb[7] = p0_matrix[p1_idx_u8__7_squeezed_comb][7];
  assign p1_add_8202_comb = p0_start_pix[7:2] + 6'h03;
  assign p1_add_8245_comb = p0_start_pix[7:3] + 5'h01;
  assign p1_actual_index__15_comb = p0_start_pix + p1_idx_u8__15_comb;
  assign p1_add_8411_comb = p0_start_pix[7:4] + 4'h1;
  assign p1_actual_index__17_comb = p0_start_pix + p1_idx_u8__17_comb;
  assign p1_add_8413_comb = p0_start_pix[7:1] + 7'h09;
  assign p1_actual_index__19_comb = p0_start_pix + p1_idx_u8__19_comb;
  assign p1_add_8415_comb = p0_start_pix[7:2] + 6'h05;
  assign p1_actual_index__21_comb = p0_start_pix + p1_idx_u8__21_comb;
  assign p1_add_8417_comb = p0_start_pix[7:1] + 7'h0b;
  assign p1_actual_index__23_comb = p0_start_pix + p1_idx_u8__23_comb;
  assign p1_add_8419_comb = p0_start_pix[7:3] + 5'h03;
  assign p1_actual_index__25_comb = p0_start_pix + p1_idx_u8__25_comb;
  assign p1_add_8421_comb = p0_start_pix[7:1] + 7'h0d;
  assign p1_actual_index__27_comb = p0_start_pix + p1_idx_u8__27_comb;
  assign p1_add_8423_comb = p0_start_pix[7:2] + 6'h07;
  assign p1_actual_index__29_comb = p0_start_pix + p1_idx_u8__29_comb;
  assign p1_add_8425_comb = p0_start_pix[7:1] + 7'h0f;
  assign p1_actual_index__31_comb = p0_start_pix + p1_idx_u8__31_comb;
  assign p1_add_8427_comb = p0_start_pix[7:5] + 3'h1;
  assign p1_actual_index__33_comb = p0_start_pix + p1_idx_u8__33_comb;
  assign p1_add_8429_comb = p0_start_pix[7:1] + 7'h11;
  assign p1_actual_index__35_comb = p0_start_pix + p1_idx_u8__35_comb;
  assign p1_add_8431_comb = p0_start_pix[7:2] + 6'h09;
  assign p1_actual_index__37_comb = p0_start_pix + p1_idx_u8__37_comb;
  assign p1_add_8433_comb = p0_start_pix[7:1] + 7'h13;
  assign p1_actual_index__39_comb = p0_start_pix + p1_idx_u8__39_comb;
  assign p1_add_8435_comb = p0_start_pix[7:3] + 5'h05;
  assign p1_actual_index__41_comb = p0_start_pix + p1_idx_u8__41_comb;
  assign p1_add_8437_comb = p0_start_pix[7:1] + 7'h15;
  assign p1_actual_index__43_comb = p0_start_pix + p1_idx_u8__43_comb;
  assign p1_add_8439_comb = p0_start_pix[7:2] + 6'h0b;
  assign p1_actual_index__45_comb = p0_start_pix + p1_idx_u8__45_comb;
  assign p1_add_8441_comb = p0_start_pix[7:1] + 7'h17;
  assign p1_actual_index__47_comb = p0_start_pix + p1_idx_u8__47_comb;
  assign p1_add_8443_comb = p0_start_pix[7:4] + 4'h3;
  assign p1_actual_index__49_comb = p0_start_pix + p1_idx_u8__49_comb;
  assign p1_add_8445_comb = p0_start_pix[7:1] + 7'h19;
  assign p1_actual_index__51_comb = p0_start_pix + p1_idx_u8__51_comb;
  assign p1_add_8447_comb = p0_start_pix[7:2] + 6'h0d;
  assign p1_actual_index__53_comb = p0_start_pix + p1_idx_u8__53_comb;
  assign p1_add_8449_comb = p0_start_pix[7:1] + 7'h1b;
  assign p1_actual_index__55_comb = p0_start_pix + p1_idx_u8__55_comb;
  assign p1_add_8451_comb = p0_start_pix[7:3] + 5'h07;
  assign p1_actual_index__57_comb = p0_start_pix + p1_idx_u8__57_comb;
  assign p1_add_8453_comb = p0_start_pix[7:1] + 7'h1d;
  assign p1_actual_index__59_comb = p0_start_pix + p1_idx_u8__59_comb;
  assign p1_add_8455_comb = p0_start_pix[7:2] + 6'h0f;
  assign p1_actual_index__61_comb = p0_start_pix + p1_idx_u8__61_comb;
  assign p1_add_8457_comb = p0_start_pix[7:1] + 7'h1f;
  assign p1_flat_comb[0] = p1_array_concat_8197_comb[0];
  assign p1_flat_comb[1] = p1_array_concat_8197_comb[1];
  assign p1_flat_comb[2] = p1_array_concat_8197_comb[2];
  assign p1_flat_comb[3] = p1_array_concat_8197_comb[3];
  assign p1_flat_comb[4] = p1_array_concat_8197_comb[4];
  assign p1_flat_comb[5] = p1_array_concat_8197_comb[5];
  assign p1_flat_comb[6] = p1_array_concat_8197_comb[6];
  assign p1_flat_comb[7] = p1_array_concat_8197_comb[7];
  assign p1_flat_comb[8] = p1_array_concat_8197_comb[8];
  assign p1_flat_comb[9] = p1_array_concat_8197_comb[9];
  assign p1_flat_comb[10] = p1_array_concat_8197_comb[10];
  assign p1_flat_comb[11] = p1_array_concat_8197_comb[11];
  assign p1_flat_comb[12] = p1_array_concat_8197_comb[12];
  assign p1_flat_comb[13] = p1_array_concat_8197_comb[13];
  assign p1_flat_comb[14] = p1_array_concat_8197_comb[14];
  assign p1_flat_comb[15] = p1_array_concat_8197_comb[15];
  assign p1_flat_comb[16] = p1_array_concat_8197_comb[16];
  assign p1_flat_comb[17] = p1_array_concat_8197_comb[17];
  assign p1_flat_comb[18] = p1_array_concat_8197_comb[18];
  assign p1_flat_comb[19] = p1_array_concat_8197_comb[19];
  assign p1_flat_comb[20] = p1_array_concat_8197_comb[20];
  assign p1_flat_comb[21] = p1_array_concat_8197_comb[21];
  assign p1_flat_comb[22] = p1_array_concat_8197_comb[22];
  assign p1_flat_comb[23] = p1_array_concat_8197_comb[23];
  assign p1_flat_comb[24] = p1_array_concat_8197_comb[24];
  assign p1_flat_comb[25] = p1_array_concat_8197_comb[25];
  assign p1_flat_comb[26] = p1_array_concat_8197_comb[26];
  assign p1_flat_comb[27] = p1_array_concat_8197_comb[27];
  assign p1_flat_comb[28] = p1_array_concat_8197_comb[28];
  assign p1_flat_comb[29] = p1_array_concat_8197_comb[29];
  assign p1_flat_comb[30] = p1_array_concat_8197_comb[30];
  assign p1_flat_comb[31] = p1_array_concat_8197_comb[31];
  assign p1_flat_comb[32] = p1_array_concat_8197_comb[32];
  assign p1_flat_comb[33] = p1_array_concat_8197_comb[33];
  assign p1_flat_comb[34] = p1_array_concat_8197_comb[34];
  assign p1_flat_comb[35] = p1_array_concat_8197_comb[35];
  assign p1_flat_comb[36] = p1_array_concat_8197_comb[36];
  assign p1_flat_comb[37] = p1_array_concat_8197_comb[37];
  assign p1_flat_comb[38] = p1_array_concat_8197_comb[38];
  assign p1_flat_comb[39] = p1_array_concat_8197_comb[39];
  assign p1_flat_comb[40] = p1_array_concat_8197_comb[40];
  assign p1_flat_comb[41] = p1_array_concat_8197_comb[41];
  assign p1_flat_comb[42] = p1_array_concat_8197_comb[42];
  assign p1_flat_comb[43] = p1_array_concat_8197_comb[43];
  assign p1_flat_comb[44] = p1_array_concat_8197_comb[44];
  assign p1_flat_comb[45] = p1_array_concat_8197_comb[45];
  assign p1_flat_comb[46] = p1_array_concat_8197_comb[46];
  assign p1_flat_comb[47] = p1_array_concat_8197_comb[47];
  assign p1_flat_comb[48] = p1_array_concat_8197_comb[48];
  assign p1_flat_comb[49] = p1_array_concat_8197_comb[49];
  assign p1_flat_comb[50] = p1_array_concat_8197_comb[50];
  assign p1_flat_comb[51] = p1_array_concat_8197_comb[51];
  assign p1_flat_comb[52] = p1_array_concat_8197_comb[52];
  assign p1_flat_comb[53] = p1_array_concat_8197_comb[53];
  assign p1_flat_comb[54] = p1_array_concat_8197_comb[54];
  assign p1_flat_comb[55] = p1_array_concat_8197_comb[55];
  assign p1_flat_comb[56] = p1_row7_comb[0];
  assign p1_flat_comb[57] = p1_row7_comb[1];
  assign p1_flat_comb[58] = p1_row7_comb[2];
  assign p1_flat_comb[59] = p1_row7_comb[3];
  assign p1_flat_comb[60] = p1_row7_comb[4];
  assign p1_flat_comb[61] = p1_row7_comb[5];
  assign p1_flat_comb[62] = p1_row7_comb[6];
  assign p1_flat_comb[63] = p1_row7_comb[7];
  assign p1_actual_index__14_comb = {p1_add_8193_comb, p0_start_pix[0]};
  assign p1_actual_index__2_comb = {p1_add_8308_comb, p0_start_pix[0]};
  assign p1_actual_index__4_comb = {p1_add_8291_comb, p0_start_pix[1:0]};
  assign p1_actual_index__6_comb = {p1_add_8275_comb, p0_start_pix[0]};
  assign p1_actual_index__10_comb = {p1_add_8226_comb, p0_start_pix[0]};
  assign p1_actual_index__12_comb = {p1_add_8202_comb, p0_start_pix[1:0]};
  assign p1_actual_index__8_comb = {p1_add_8245_comb, p0_start_pix[2:0]};
  assign p1_actual_index__16_comb = {p1_add_8411_comb, p0_start_pix[3:0]};
  assign p1_actual_index__18_comb = {p1_add_8413_comb, p0_start_pix[0]};
  assign p1_actual_index__20_comb = {p1_add_8415_comb, p0_start_pix[1:0]};
  assign p1_actual_index__22_comb = {p1_add_8417_comb, p0_start_pix[0]};
  assign p1_actual_index__24_comb = {p1_add_8419_comb, p0_start_pix[2:0]};
  assign p1_actual_index__26_comb = {p1_add_8421_comb, p0_start_pix[0]};
  assign p1_actual_index__28_comb = {p1_add_8423_comb, p0_start_pix[1:0]};
  assign p1_actual_index__30_comb = {p1_add_8425_comb, p0_start_pix[0]};
  assign p1_actual_index__32_comb = {p1_add_8427_comb, p0_start_pix[4:0]};
  assign p1_actual_index__34_comb = {p1_add_8429_comb, p0_start_pix[0]};
  assign p1_actual_index__36_comb = {p1_add_8431_comb, p0_start_pix[1:0]};
  assign p1_actual_index__38_comb = {p1_add_8433_comb, p0_start_pix[0]};
  assign p1_actual_index__40_comb = {p1_add_8435_comb, p0_start_pix[2:0]};
  assign p1_actual_index__42_comb = {p1_add_8437_comb, p0_start_pix[0]};
  assign p1_actual_index__44_comb = {p1_add_8439_comb, p0_start_pix[1:0]};
  assign p1_actual_index__46_comb = {p1_add_8441_comb, p0_start_pix[0]};
  assign p1_actual_index__48_comb = {p1_add_8443_comb, p0_start_pix[3:0]};
  assign p1_actual_index__50_comb = {p1_add_8445_comb, p0_start_pix[0]};
  assign p1_actual_index__52_comb = {p1_add_8447_comb, p0_start_pix[1:0]};
  assign p1_actual_index__54_comb = {p1_add_8449_comb, p0_start_pix[0]};
  assign p1_actual_index__56_comb = {p1_add_8451_comb, p0_start_pix[2:0]};
  assign p1_actual_index__58_comb = {p1_add_8453_comb, p0_start_pix[0]};
  assign p1_actual_index__60_comb = {p1_add_8455_comb, p0_start_pix[1:0]};
  assign p1_actual_index__62_comb = {p1_add_8457_comb, p0_start_pix[0]};
  assign p1_and_8221_comb = p1_flat_comb[p1_actual_index__14_comb > 8'h3f ? 6'h3f : p1_actual_index__14_comb[5:0]] & {10{~(p1_add_8193_comb[5] | p1_add_8193_comb[6])}};
  assign p1_and_8352_comb = p1_flat_comb[p0_start_pix > 8'h3f ? 6'h3f : p0_start_pix[5:0]] & {10{~(p0_start_pix[6] | p0_start_pix[7])}};
  assign p1_and_8354_comb = p1_flat_comb[p1_actual_index__1_comb > 8'h3f ? 6'h3f : p1_actual_index__1_comb[5:0]] & {10{~(p1_actual_index__1_comb[6] | p1_actual_index__1_comb[7])}};
  assign p1_and_8349_comb = p1_flat_comb[p1_actual_index__2_comb > 8'h3f ? 6'h3f : p1_actual_index__2_comb[5:0]] & {10{~(p1_add_8308_comb[5] | p1_add_8308_comb[6])}};
  assign p1_and_8342_comb = p1_flat_comb[p1_actual_index__3_comb > 8'h3f ? 6'h3f : p1_actual_index__3_comb[5:0]] & {10{~(p1_actual_index__3_comb[6] | p1_actual_index__3_comb[7])}};
  assign p1_and_8335_comb = p1_flat_comb[p1_actual_index__4_comb > 8'h3f ? 6'h3f : p1_actual_index__4_comb[5:0]] & {10{~(p1_add_8291_comb[4] | p1_add_8291_comb[5])}};
  assign p1_and_8324_comb = p1_flat_comb[p1_actual_index__5_comb > 8'h3f ? 6'h3f : p1_actual_index__5_comb[5:0]] & {10{~(p1_actual_index__5_comb[6] | p1_actual_index__5_comb[7])}};
  assign p1_and_8315_comb = p1_flat_comb[p1_actual_index__6_comb > 8'h3f ? 6'h3f : p1_actual_index__6_comb[5:0]] & {10{~(p1_add_8275_comb[5] | p1_add_8275_comb[6])}};
  assign p1_and_8305_comb = p1_flat_comb[p1_actual_index__7_comb > 8'h3f ? 6'h3f : p1_actual_index__7_comb[5:0]] & {10{~(p1_actual_index__7_comb[6] | p1_actual_index__7_comb[7])}};
  assign p1_and_8278_comb = p1_flat_comb[p1_actual_index__9_comb > 8'h3f ? 6'h3f : p1_actual_index__9_comb[5:0]] & {10{~(p1_actual_index__9_comb[6] | p1_actual_index__9_comb[7])}};
  assign p1_and_8269_comb = p1_flat_comb[p1_actual_index__10_comb > 8'h3f ? 6'h3f : p1_actual_index__10_comb[5:0]] & {10{~(p1_add_8226_comb[5] | p1_add_8226_comb[6])}};
  assign p1_and_8261_comb = p1_flat_comb[p1_actual_index__11_comb > 8'h3f ? 6'h3f : p1_actual_index__11_comb[5:0]] & {10{~(p1_actual_index__11_comb[6] | p1_actual_index__11_comb[7])}};
  assign p1_and_8229_comb = p1_flat_comb[p1_actual_index__13_comb > 8'h3f ? 6'h3f : p1_actual_index__13_comb[5:0]] & {10{~(p1_actual_index__13_comb[6] | p1_actual_index__13_comb[7])}};
  assign p1_eq_8232_comb = p1_and_8221_comb == 10'h000;
  assign p1_and_8233_comb = p1_flat_comb[p1_actual_index__12_comb > 8'h3f ? 6'h3f : p1_actual_index__12_comb[5:0]] & {10{~(p1_add_8202_comb[4] | p1_add_8202_comb[5])}};
  assign p1_ne_8357_comb = p1_and_8352_comb != 10'h000;
  assign p1_ne_8358_comb = p1_and_8354_comb != 10'h000;
  assign p1_ne_8356_comb = p1_and_8349_comb != 10'h000;
  assign p1_ne_8351_comb = p1_and_8342_comb != 10'h000;
  assign p1_ne_8344_comb = p1_and_8335_comb != 10'h000;
  assign p1_ne_8337_comb = p1_and_8324_comb != 10'h000;
  assign p1_ne_8326_comb = p1_and_8315_comb != 10'h000;
  assign p1_ne_8317_comb = p1_and_8305_comb != 10'h000;
  assign p1_and_8281_comb = p1_flat_comb[p1_actual_index__8_comb > 8'h3f ? 6'h3f : p1_actual_index__8_comb[5:0]] & {10{~(p1_add_8245_comb[3] | p1_add_8245_comb[4])}};
  assign p1_ne_8288_comb = p1_and_8278_comb != 10'h000;
  assign p1_ne_8280_comb = p1_and_8269_comb != 10'h000;
  assign p1_ne_8271_comb = p1_and_8261_comb != 10'h000;
  assign p1_ne_8241_comb = p1_and_8229_comb != 10'h000;
  assign p1_value_comb = p0_matrix[3'h0][3'h0];
  assign p1_idx_u8__1_squeezed_comb = 2'h1;
  assign p1_eq_8244_comb = p1_and_8233_comb == 10'h000;
  assign p1_not_8359_comb = ~p1_ne_8357_comb;
  assign p1_eq_8289_comb = p1_and_8281_comb == 10'h000;
  assign p1_bin_value__1_comb = p1_value_comb[7:0];
  assign p1_flipped_comb = 8'hff;
  assign p1_sel_8252_comb = p1_ne_8241_comb ? p1_idx_u8__1_squeezed_comb : {1'h1, p1_eq_8232_comb};
  assign p1_sign_ext_8253_comb = {2{p1_eq_8244_comb}};
  assign p1_and_8883_comb = p1_not_8359_comb & ~p1_ne_8358_comb & ~p1_ne_8356_comb & ~p1_ne_8351_comb & ~p1_ne_8344_comb & ~p1_ne_8337_comb & ~p1_ne_8326_comb & ~p1_ne_8317_comb & p1_eq_8289_comb & ~p1_ne_8288_comb & ~p1_ne_8280_comb & ~p1_ne_8271_comb & p1_eq_8244_comb & ~p1_ne_8241_comb & p1_eq_8232_comb & (p1_flat_comb[p1_actual_index__15_comb > 8'h3f ? 6'h3f : p1_actual_index__15_comb[5:0]] & {10{~(p1_actual_index__15_comb[6] | p1_actual_index__15_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__16_comb > 8'h3f ? 6'h3f : p1_actual_index__16_comb[5:0]] & {10{~(p1_add_8411_comb[2] | p1_add_8411_comb[3])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__17_comb > 8'h3f ? 6'h3f : p1_actual_index__17_comb[5:0]] & {10{~(p1_actual_index__17_comb[6] | p1_actual_index__17_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__18_comb > 8'h3f ? 6'h3f : p1_actual_index__18_comb[5:0]] & {10{~(p1_add_8413_comb[5] | p1_add_8413_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__19_comb > 8'h3f ? 6'h3f : p1_actual_index__19_comb[5:0]] & {10{~(p1_actual_index__19_comb[6] | p1_actual_index__19_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__20_comb > 8'h3f ? 6'h3f : p1_actual_index__20_comb[5:0]] & {10{~(p1_add_8415_comb[4] | p1_add_8415_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__21_comb > 8'h3f ? 6'h3f : p1_actual_index__21_comb[5:0]] & {10{~(p1_actual_index__21_comb[6] | p1_actual_index__21_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__22_comb > 8'h3f ? 6'h3f : p1_actual_index__22_comb[5:0]] & {10{~(p1_add_8417_comb[5] | p1_add_8417_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__23_comb > 8'h3f ? 6'h3f : p1_actual_index__23_comb[5:0]] & {10{~(p1_actual_index__23_comb[6] | p1_actual_index__23_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__24_comb > 8'h3f ? 6'h3f : p1_actual_index__24_comb[5:0]] & {10{~(p1_add_8419_comb[3] | p1_add_8419_comb[4])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__25_comb > 8'h3f ? 6'h3f : p1_actual_index__25_comb[5:0]] & {10{~(p1_actual_index__25_comb[6] | p1_actual_index__25_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__26_comb > 8'h3f ? 6'h3f : p1_actual_index__26_comb[5:0]] & {10{~(p1_add_8421_comb[5] | p1_add_8421_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__27_comb > 8'h3f ? 6'h3f : p1_actual_index__27_comb[5:0]] & {10{~(p1_actual_index__27_comb[6] | p1_actual_index__27_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__28_comb > 8'h3f ? 6'h3f : p1_actual_index__28_comb[5:0]] & {10{~(p1_add_8423_comb[4] | p1_add_8423_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__29_comb > 8'h3f ? 6'h3f : p1_actual_index__29_comb[5:0]] & {10{~(p1_actual_index__29_comb[6] | p1_actual_index__29_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__30_comb > 8'h3f ? 6'h3f : p1_actual_index__30_comb[5:0]] & {10{~(p1_add_8425_comb[5] | p1_add_8425_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__31_comb > 8'h3f ? 6'h3f : p1_actual_index__31_comb[5:0]] & {10{~(p1_actual_index__31_comb[6] | p1_actual_index__31_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__32_comb > 8'h3f ? 6'h3f : p1_actual_index__32_comb[5:0]] & {10{~(p1_add_8427_comb[1] | p1_add_8427_comb[2])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__33_comb > 8'h3f ? 6'h3f : p1_actual_index__33_comb[5:0]] & {10{~(p1_actual_index__33_comb[6] | p1_actual_index__33_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__34_comb > 8'h3f ? 6'h3f : p1_actual_index__34_comb[5:0]] & {10{~(p1_add_8429_comb[5] | p1_add_8429_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__35_comb > 8'h3f ? 6'h3f : p1_actual_index__35_comb[5:0]] & {10{~(p1_actual_index__35_comb[6] | p1_actual_index__35_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__36_comb > 8'h3f ? 6'h3f : p1_actual_index__36_comb[5:0]] & {10{~(p1_add_8431_comb[4] | p1_add_8431_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__37_comb > 8'h3f ? 6'h3f : p1_actual_index__37_comb[5:0]] & {10{~(p1_actual_index__37_comb[6] | p1_actual_index__37_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__38_comb > 8'h3f ? 6'h3f : p1_actual_index__38_comb[5:0]] & {10{~(p1_add_8433_comb[5] | p1_add_8433_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__39_comb > 8'h3f ? 6'h3f : p1_actual_index__39_comb[5:0]] & {10{~(p1_actual_index__39_comb[6] | p1_actual_index__39_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__40_comb > 8'h3f ? 6'h3f : p1_actual_index__40_comb[5:0]] & {10{~(p1_add_8435_comb[3] | p1_add_8435_comb[4])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__41_comb > 8'h3f ? 6'h3f : p1_actual_index__41_comb[5:0]] & {10{~(p1_actual_index__41_comb[6] | p1_actual_index__41_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__42_comb > 8'h3f ? 6'h3f : p1_actual_index__42_comb[5:0]] & {10{~(p1_add_8437_comb[5] | p1_add_8437_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__43_comb > 8'h3f ? 6'h3f : p1_actual_index__43_comb[5:0]] & {10{~(p1_actual_index__43_comb[6] | p1_actual_index__43_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__44_comb > 8'h3f ? 6'h3f : p1_actual_index__44_comb[5:0]] & {10{~(p1_add_8439_comb[4] | p1_add_8439_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__45_comb > 8'h3f ? 6'h3f : p1_actual_index__45_comb[5:0]] & {10{~(p1_actual_index__45_comb[6] | p1_actual_index__45_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__46_comb > 8'h3f ? 6'h3f : p1_actual_index__46_comb[5:0]] & {10{~(p1_add_8441_comb[5] | p1_add_8441_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__47_comb > 8'h3f ? 6'h3f : p1_actual_index__47_comb[5:0]] & {10{~(p1_actual_index__47_comb[6] | p1_actual_index__47_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__48_comb > 8'h3f ? 6'h3f : p1_actual_index__48_comb[5:0]] & {10{~(p1_add_8443_comb[2] | p1_add_8443_comb[3])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__49_comb > 8'h3f ? 6'h3f : p1_actual_index__49_comb[5:0]] & {10{~(p1_actual_index__49_comb[6] | p1_actual_index__49_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__50_comb > 8'h3f ? 6'h3f : p1_actual_index__50_comb[5:0]] & {10{~(p1_add_8445_comb[5] | p1_add_8445_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__51_comb > 8'h3f ? 6'h3f : p1_actual_index__51_comb[5:0]] & {10{~(p1_actual_index__51_comb[6] | p1_actual_index__51_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__52_comb > 8'h3f ? 6'h3f : p1_actual_index__52_comb[5:0]] & {10{~(p1_add_8447_comb[4] | p1_add_8447_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__53_comb > 8'h3f ? 6'h3f : p1_actual_index__53_comb[5:0]] & {10{~(p1_actual_index__53_comb[6] | p1_actual_index__53_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__54_comb > 8'h3f ? 6'h3f : p1_actual_index__54_comb[5:0]] & {10{~(p1_add_8449_comb[5] | p1_add_8449_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__55_comb > 8'h3f ? 6'h3f : p1_actual_index__55_comb[5:0]] & {10{~(p1_actual_index__55_comb[6] | p1_actual_index__55_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__56_comb > 8'h3f ? 6'h3f : p1_actual_index__56_comb[5:0]] & {10{~(p1_add_8451_comb[3] | p1_add_8451_comb[4])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__57_comb > 8'h3f ? 6'h3f : p1_actual_index__57_comb[5:0]] & {10{~(p1_actual_index__57_comb[6] | p1_actual_index__57_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__58_comb > 8'h3f ? 6'h3f : p1_actual_index__58_comb[5:0]] & {10{~(p1_add_8453_comb[5] | p1_add_8453_comb[6])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__59_comb > 8'h3f ? 6'h3f : p1_actual_index__59_comb[5:0]] & {10{~(p1_actual_index__59_comb[6] | p1_actual_index__59_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__60_comb > 8'h3f ? 6'h3f : p1_actual_index__60_comb[5:0]] & {10{~(p1_add_8455_comb[4] | p1_add_8455_comb[5])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__61_comb > 8'h3f ? 6'h3f : p1_actual_index__61_comb[5:0]] & {10{~(p1_actual_index__61_comb[6] | p1_actual_index__61_comb[7])}}) == 10'h000 & (p1_flat_comb[p1_actual_index__62_comb > 8'h3f ? 6'h3f : p1_actual_index__62_comb[5:0]] & {10{~(p1_add_8457_comb[5] | p1_add_8457_comb[6])}}) == 10'h000;
  assign p1_code_list_comb = p1_value_comb == 10'h000 ? p1_flipped_comb : p1_bin_value__1_comb;

  // Registers for pipe stage 1:
  reg p1_is_luminance;
  reg [9:0] p1_and_8221;
  reg [9:0] p1_and_8229;
  reg [9:0] p1_and_8233;
  reg [1:0] p1_sel_8252;
  reg [1:0] p1_sign_ext_8253;
  reg [9:0] p1_and_8261;
  reg [9:0] p1_and_8269;
  reg p1_ne_8271;
  reg [9:0] p1_and_8278;
  reg p1_ne_8280;
  reg [9:0] p1_and_8281;
  reg p1_ne_8288;
  reg p1_eq_8289;
  reg [9:0] p1_and_8305;
  reg [9:0] p1_and_8315;
  reg p1_ne_8317;
  reg [9:0] p1_and_8324;
  reg p1_ne_8326;
  reg [9:0] p1_and_8335;
  reg p1_ne_8337;
  reg [9:0] p1_and_8342;
  reg p1_ne_8344;
  reg [9:0] p1_and_8349;
  reg p1_ne_8351;
  reg [9:0] p1_and_8352;
  reg [9:0] p1_and_8354;
  reg p1_ne_8356;
  reg p1_ne_8357;
  reg p1_ne_8358;
  reg p1_not_8359;
  reg p1_and_8883;
  reg [7:0] p1_code_list;
  always @ (posedge clk) begin
    p1_is_luminance <= p0_is_luminance;
    p1_and_8221 <= p1_and_8221_comb;
    p1_and_8229 <= p1_and_8229_comb;
    p1_and_8233 <= p1_and_8233_comb;
    p1_sel_8252 <= p1_sel_8252_comb;
    p1_sign_ext_8253 <= p1_sign_ext_8253_comb;
    p1_and_8261 <= p1_and_8261_comb;
    p1_and_8269 <= p1_and_8269_comb;
    p1_ne_8271 <= p1_ne_8271_comb;
    p1_and_8278 <= p1_and_8278_comb;
    p1_ne_8280 <= p1_ne_8280_comb;
    p1_and_8281 <= p1_and_8281_comb;
    p1_ne_8288 <= p1_ne_8288_comb;
    p1_eq_8289 <= p1_eq_8289_comb;
    p1_and_8305 <= p1_and_8305_comb;
    p1_and_8315 <= p1_and_8315_comb;
    p1_ne_8317 <= p1_ne_8317_comb;
    p1_and_8324 <= p1_and_8324_comb;
    p1_ne_8326 <= p1_ne_8326_comb;
    p1_and_8335 <= p1_and_8335_comb;
    p1_ne_8337 <= p1_ne_8337_comb;
    p1_and_8342 <= p1_and_8342_comb;
    p1_ne_8344 <= p1_ne_8344_comb;
    p1_and_8349 <= p1_and_8349_comb;
    p1_ne_8351 <= p1_ne_8351_comb;
    p1_and_8352 <= p1_and_8352_comb;
    p1_and_8354 <= p1_and_8354_comb;
    p1_ne_8356 <= p1_ne_8356_comb;
    p1_ne_8357 <= p1_ne_8357_comb;
    p1_ne_8358 <= p1_ne_8358_comb;
    p1_not_8359 <= p1_not_8359_comb;
    p1_and_8883 <= p1_and_8883_comb;
    p1_code_list <= p1_code_list_comb;
  end

  // ===== Pipe stage 2:
  wire [2:0] p2_and_8965_comb;
  wire [3:0] p2_idx_u8__4_squeezed__2_comb;
  wire [3:0] p2_sel_8974_comb;
  wire [3:0] p2_sel_8978_comb;
  assign p2_and_8965_comb = (p1_ne_8288 ? 3'h1 : (p1_ne_8280 ? 3'h2 : (p1_ne_8271 ? 3'h3 : {1'h1, p1_sel_8252 & p1_sign_ext_8253}))) & {3{p1_eq_8289}};
  assign p2_idx_u8__4_squeezed__2_comb = 4'h4;
  assign p2_sel_8974_comb = p1_ne_8344 ? p2_idx_u8__4_squeezed__2_comb : (p1_ne_8337 ? 4'h5 : (p1_ne_8326 ? 4'h6 : (p1_ne_8317 ? 4'h7 : {1'h1, p2_and_8965_comb})));
  assign p2_sel_8978_comb = p1_ne_8356 ? 4'h2 : (p1_ne_8351 ? 4'h3 : p2_sel_8974_comb);

  // Registers for pipe stage 2:
  reg p2_is_luminance;
  reg [9:0] p2_and_8221;
  reg [9:0] p2_and_8229;
  reg [9:0] p2_and_8233;
  reg [9:0] p2_and_8261;
  reg [9:0] p2_and_8269;
  reg [9:0] p2_and_8278;
  reg [9:0] p2_and_8281;
  reg [9:0] p2_and_8305;
  reg [9:0] p2_and_8315;
  reg [9:0] p2_and_8324;
  reg [9:0] p2_and_8335;
  reg [9:0] p2_and_8342;
  reg [9:0] p2_and_8349;
  reg [9:0] p2_and_8352;
  reg [9:0] p2_and_8354;
  reg p2_ne_8357;
  reg p2_ne_8358;
  reg [3:0] p2_sel_8978;
  reg p2_not_8359;
  reg p2_and_8883;
  reg [7:0] p2_code_list;
  always @ (posedge clk) begin
    p2_is_luminance <= p1_is_luminance;
    p2_and_8221 <= p1_and_8221;
    p2_and_8229 <= p1_and_8229;
    p2_and_8233 <= p1_and_8233;
    p2_and_8261 <= p1_and_8261;
    p2_and_8269 <= p1_and_8269;
    p2_and_8278 <= p1_and_8278;
    p2_and_8281 <= p1_and_8281;
    p2_and_8305 <= p1_and_8305;
    p2_and_8315 <= p1_and_8315;
    p2_and_8324 <= p1_and_8324;
    p2_and_8335 <= p1_and_8335;
    p2_and_8342 <= p1_and_8342;
    p2_and_8349 <= p1_and_8349;
    p2_and_8352 <= p1_and_8352;
    p2_and_8354 <= p1_and_8354;
    p2_ne_8357 <= p1_ne_8357;
    p2_ne_8358 <= p1_ne_8358;
    p2_sel_8978 <= p2_sel_8978_comb;
    p2_not_8359 <= p1_not_8359;
    p2_and_8883 <= p1_and_8883;
    p2_code_list <= p1_code_list;
  end

  // ===== Pipe stage 3:
  wire [3:0] p3_sel_9024_comb;
  wire [3:0] p3_run_comb;
  wire [9:0] p3_value__1_comb;
  wire [7:0] p3_bin_value__2_comb;
  wire [7:0] p3_bin_value__3_comb;
  wire [7:0] p3_value_abs_comb;
  wire [1:0] p3_idx_u8__1_squeezed__1_comb;
  wire [1:0] p3_idx_u8__2_squeezed_comb;
  wire [1:0] p3_idx_u8__3_squeezed_comb;
  wire p3_eq_9061_comb;
  wire [7:0] p3_flipped__1_comb;
  wire [2:0] p3_idx_u8__4_squeezed__3_comb;
  wire [7:0] p3_Code_list_comb;
  wire [2:0] p3_sel_9050_comb;
  wire [2:0] p3_idx_u8__5_squeezed__1_comb;
  wire p3_or_reduce_9053_comb;
  wire [2:0] p3_sel_9054_comb;
  wire p3_or_reduce_9055_comb;
  wire p3_bit_slice_9056_comb;
  wire p3_ne_9058_comb;
  wire [7:0] p3_sel_9072_comb;
  wire [3:0] p3_sel_9073_comb;
  assign p3_sel_9024_comb = p2_ne_8358 ? 4'h1 : p2_sel_8978;
  assign p3_run_comb = p3_sel_9024_comb & {4{p2_not_8359}};
  assign p3_value__1_comb = p3_run_comb == 4'h0 ? p2_and_8352 : (p3_run_comb == 4'h1 ? p2_and_8354 : (p3_run_comb == 4'h2 ? p2_and_8349 : (p3_run_comb == 4'h3 ? p2_and_8342 : (p3_run_comb == 4'h4 ? p2_and_8335 : (p3_run_comb == 4'h5 ? p2_and_8324 : (p3_run_comb == 4'h6 ? p2_and_8315 : (p3_run_comb == 4'h7 ? p2_and_8305 : (p3_run_comb == 4'h8 ? p2_and_8281 : (p3_run_comb == 4'h9 ? p2_and_8278 : (p3_run_comb == 4'ha ? p2_and_8269 : (p3_run_comb == 4'hb ? p2_and_8261 : (p3_run_comb == 4'hc ? p2_and_8233 : (p3_run_comb == 4'hd ? p2_and_8229 : (p3_run_comb == 4'he ? p2_and_8221 : 10'h000))))))))))))));
  assign p3_bin_value__2_comb = p3_value__1_comb[7:0];
  assign p3_bin_value__3_comb = -p3_bin_value__2_comb;
  assign p3_value_abs_comb = p3_value__1_comb[9] ? p3_bin_value__3_comb : p3_bin_value__2_comb;
  assign p3_idx_u8__1_squeezed__1_comb = 2'h1;
  assign p3_idx_u8__2_squeezed_comb = 2'h2;
  assign p3_idx_u8__3_squeezed_comb = 2'h3;
  assign p3_eq_9061_comb = p3_run_comb == 4'hf;
  assign p3_flipped__1_comb = ~p3_bin_value__3_comb;
  assign p3_idx_u8__4_squeezed__3_comb = 3'h4;
  assign p3_Code_list_comb = $signed(p3_value__1_comb) <= $signed(10'h000) ? p3_flipped__1_comb : p3_bin_value__2_comb;
  assign p3_sel_9050_comb = |p3_value_abs_comb[7:3] ? p3_idx_u8__4_squeezed__3_comb : {1'h0, |p3_value_abs_comb[7:2] ? p3_idx_u8__3_squeezed_comb : (|p3_value_abs_comb[7:1] ? p3_idx_u8__2_squeezed_comb : p3_idx_u8__1_squeezed__1_comb)};
  assign p3_idx_u8__5_squeezed__1_comb = 3'h5;
  assign p3_or_reduce_9053_comb = |p3_value_abs_comb[7:5];
  assign p3_sel_9054_comb = |p3_value_abs_comb[7:4] ? p3_idx_u8__5_squeezed__1_comb : p3_sel_9050_comb;
  assign p3_or_reduce_9055_comb = |p3_value_abs_comb[7:6];
  assign p3_bit_slice_9056_comb = p3_value_abs_comb[7];
  assign p3_ne_9058_comb = p3_value_abs_comb != 8'h00;
  assign p3_sel_9072_comb = p2_and_8883 ? p2_code_list : p3_Code_list_comb & {8{~p3_eq_9061_comb}};
  assign p3_sel_9073_comb = p2_and_8883 ? 4'hf : p3_sel_9024_comb & {4{~(p3_eq_9061_comb | p2_ne_8357)}};

  // Registers for pipe stage 3:
  reg p3_is_luminance;
  reg [3:0] p3_run;
  reg p3_or_reduce_9053;
  reg [2:0] p3_sel_9054;
  reg p3_or_reduce_9055;
  reg p3_bit_slice_9056;
  reg p3_ne_9058;
  reg p3_eq_9061;
  reg p3_and_8883;
  reg [7:0] p3_sel_9072;
  reg [3:0] p3_sel_9073;
  always @ (posedge clk) begin
    p3_is_luminance <= p2_is_luminance;
    p3_run <= p3_run_comb;
    p3_or_reduce_9053 <= p3_or_reduce_9053_comb;
    p3_sel_9054 <= p3_sel_9054_comb;
    p3_or_reduce_9055 <= p3_or_reduce_9055_comb;
    p3_bit_slice_9056 <= p3_bit_slice_9056_comb;
    p3_ne_9058 <= p3_ne_9058_comb;
    p3_eq_9061 <= p3_eq_9061_comb;
    p3_and_8883 <= p2_and_8883;
    p3_sel_9072 <= p3_sel_9072_comb;
    p3_sel_9073 <= p3_sel_9073_comb;
  end

  // ===== Pipe stage 4:
  wire [2:0] p4_idx_u8__6_squeezed__1_comb;
  wire [2:0] p4_idx_u8__7_squeezed__1_comb;
  wire [3:0] p4_idx_u8__8_squeezed_comb;
  wire [7:0] p4_Code_size_comb;
  wire [7:0] p4_run_size_str_u8_comb;
  wire [4:0] p4_Huffman_length_squeezed_comb;
  wire [4:0] p4_idx_u8__2_squeezed__1_comb;
  wire [4:0] p4_idx_u8__4_squeezed__1_comb;
  wire p4_or_9123_comb;
  wire [3:0] p4_Code_size_squeezed_comb;
  wire [3:0] p4_idx_u8__4_squeezed__4_comb;
  wire [15:0] p4_Huffman_code_full_comb;
  wire [15:0] p4_EOB_LUM_EXT_comb;
  wire [43:0] p4_tuple_9135_comb;
  assign p4_idx_u8__6_squeezed__1_comb = 3'h6;
  assign p4_idx_u8__7_squeezed__1_comb = 3'h7;
  assign p4_idx_u8__8_squeezed_comb = 4'h8;
  assign p4_Code_size_comb = {4'h0, p3_bit_slice_9056 ? p4_idx_u8__8_squeezed_comb : {1'h0, p3_or_reduce_9055 ? p4_idx_u8__7_squeezed__1_comb : (p3_or_reduce_9053 ? p4_idx_u8__6_squeezed__1_comb : p3_sel_9054)}} & {8{p3_ne_9058}};
  assign p4_run_size_str_u8_comb = {p3_run, 4'h0} | p4_Code_size_comb;
  assign p4_Huffman_length_squeezed_comb = p3_is_luminance ? literal_9112[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_9110[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_idx_u8__2_squeezed__1_comb = 5'h02;
  assign p4_idx_u8__4_squeezed__1_comb = 5'h04;
  assign p4_or_9123_comb = p3_and_8883 | p3_eq_9061;
  assign p4_Code_size_squeezed_comb = p4_Code_size_comb[3:0];
  assign p4_idx_u8__4_squeezed__4_comb = 4'h4;
  assign p4_Huffman_code_full_comb = p3_is_luminance ? literal_9116[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb] : literal_9115[p4_run_size_str_u8_comb > 8'hfb ? 8'hfb : p4_run_size_str_u8_comb];
  assign p4_EOB_LUM_EXT_comb = 16'h000c;
  assign p4_tuple_9135_comb = {p4_or_9123_comb ? p4_EOB_LUM_EXT_comb : p4_Huffman_code_full_comb, {3'h0, p3_and_8883 ? p4_idx_u8__4_squeezed__1_comb : (p3_eq_9061 ? p4_idx_u8__2_squeezed__1_comb : p4_Huffman_length_squeezed_comb)}, p3_sel_9072, {4'h0, p4_or_9123_comb ? p4_idx_u8__4_squeezed__4_comb : p4_Code_size_squeezed_comb}, p3_sel_9073};

  // Registers for pipe stage 4:
  reg [43:0] p4_tuple_9135;
  always @ (posedge clk) begin
    p4_tuple_9135 <= p4_tuple_9135_comb;
  end
  assign out = p4_tuple_9135;
endmodule
