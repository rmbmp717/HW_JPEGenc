module Quantize(
  input wire clk,
  input wire [511:0] dct_coeffs,
  input wire [7:0] matrix_row,
  input wire is_luminance,
  output wire [127:0] out
);
  function automatic [31:0] sdiv_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    begin
      sdiv_32b = rhs == 32'h0000_0000 ? (lhs[31] ? 32'h8000_0000 : 32'h7fff_ffff) : (lhs == 32'h8000_0000 && rhs == 32'hffff_ffff ? 32'h8000_0000 : $unsigned($signed(lhs) / $signed(rhs)));
    end
  endfunction
  wire [15:0] CHROMINANCE_QUANT_TBL[0:7][0:7];
  assign CHROMINANCE_QUANT_TBL[0][0] = 16'h0010;
  assign CHROMINANCE_QUANT_TBL[0][1] = 16'h0011;
  assign CHROMINANCE_QUANT_TBL[0][2] = 16'h0017;
  assign CHROMINANCE_QUANT_TBL[0][3] = 16'h002d;
  assign CHROMINANCE_QUANT_TBL[0][4] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[0][5] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[0][6] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[0][7] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[1][0] = 16'h0011;
  assign CHROMINANCE_QUANT_TBL[1][1] = 16'h0014;
  assign CHROMINANCE_QUANT_TBL[1][2] = 16'h0019;
  assign CHROMINANCE_QUANT_TBL[1][3] = 16'h003f;
  assign CHROMINANCE_QUANT_TBL[1][4] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[1][5] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[1][6] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[1][7] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[2][0] = 16'h0017;
  assign CHROMINANCE_QUANT_TBL[2][1] = 16'h0019;
  assign CHROMINANCE_QUANT_TBL[2][2] = 16'h0035;
  assign CHROMINANCE_QUANT_TBL[2][3] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[2][4] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[2][5] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[2][6] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[2][7] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[3][0] = 16'h002d;
  assign CHROMINANCE_QUANT_TBL[3][1] = 16'h003f;
  assign CHROMINANCE_QUANT_TBL[3][2] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[3][3] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[3][4] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[3][5] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[3][6] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[3][7] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[4][0] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[4][1] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[4][2] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[4][3] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[4][4] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[4][5] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[4][6] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[4][7] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[5][0] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[5][1] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[5][2] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[5][3] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[5][4] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[5][5] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[5][6] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[5][7] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[6][0] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[6][1] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[6][2] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[6][3] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[6][4] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[6][5] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[6][6] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[6][7] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[7][0] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[7][1] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[7][2] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[7][3] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[7][4] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[7][5] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[7][6] = 16'h005e;
  assign CHROMINANCE_QUANT_TBL[7][7] = 16'h005e;
  wire [15:0] LUMINANCE_QUANT_TBL[0:7][0:7];
  assign LUMINANCE_QUANT_TBL[0][0] = 16'h000f;
  assign LUMINANCE_QUANT_TBL[0][1] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[0][2] = 16'h000a;
  assign LUMINANCE_QUANT_TBL[0][3] = 16'h000f;
  assign LUMINANCE_QUANT_TBL[0][4] = 16'h0017;
  assign LUMINANCE_QUANT_TBL[0][5] = 16'h0026;
  assign LUMINANCE_QUANT_TBL[0][6] = 16'h0030;
  assign LUMINANCE_QUANT_TBL[0][7] = 16'h003a;
  assign LUMINANCE_QUANT_TBL[1][0] = 16'h000b;
  assign LUMINANCE_QUANT_TBL[1][1] = 16'h000b;
  assign LUMINANCE_QUANT_TBL[1][2] = 16'h000d;
  assign LUMINANCE_QUANT_TBL[1][3] = 16'h0012;
  assign LUMINANCE_QUANT_TBL[1][4] = 16'h0019;
  assign LUMINANCE_QUANT_TBL[1][5] = 16'h0037;
  assign LUMINANCE_QUANT_TBL[1][6] = 16'h0039;
  assign LUMINANCE_QUANT_TBL[1][7] = 16'h0034;
  assign LUMINANCE_QUANT_TBL[2][0] = 16'h000d;
  assign LUMINANCE_QUANT_TBL[2][1] = 16'h000c;
  assign LUMINANCE_QUANT_TBL[2][2] = 16'h000f;
  assign LUMINANCE_QUANT_TBL[2][3] = 16'h0017;
  assign LUMINANCE_QUANT_TBL[2][4] = 16'h0026;
  assign LUMINANCE_QUANT_TBL[2][5] = 16'h0036;
  assign LUMINANCE_QUANT_TBL[2][6] = 16'h0042;
  assign LUMINANCE_QUANT_TBL[2][7] = 16'h0035;
  assign LUMINANCE_QUANT_TBL[3][0] = 16'h000d;
  assign LUMINANCE_QUANT_TBL[3][1] = 16'h0010;
  assign LUMINANCE_QUANT_TBL[3][2] = 16'h0015;
  assign LUMINANCE_QUANT_TBL[3][3] = 16'h001c;
  assign LUMINANCE_QUANT_TBL[3][4] = 16'h0030;
  assign LUMINANCE_QUANT_TBL[3][5] = 16'h0053;
  assign LUMINANCE_QUANT_TBL[3][6] = 16'h004c;
  assign LUMINANCE_QUANT_TBL[3][7] = 16'h003b;
  assign LUMINANCE_QUANT_TBL[4][0] = 16'h0011;
  assign LUMINANCE_QUANT_TBL[4][1] = 16'h0015;
  assign LUMINANCE_QUANT_TBL[4][2] = 16'h0023;
  assign LUMINANCE_QUANT_TBL[4][3] = 16'h0035;
  assign LUMINANCE_QUANT_TBL[4][4] = 16'h0041;
  assign LUMINANCE_QUANT_TBL[4][5] = 16'h0068;
  assign LUMINANCE_QUANT_TBL[4][6] = 16'h0062;
  assign LUMINANCE_QUANT_TBL[4][7] = 16'h0049;
  assign LUMINANCE_QUANT_TBL[5][0] = 16'h0017;
  assign LUMINANCE_QUANT_TBL[5][1] = 16'h0021;
  assign LUMINANCE_QUANT_TBL[5][2] = 16'h0034;
  assign LUMINANCE_QUANT_TBL[5][3] = 16'h003d;
  assign LUMINANCE_QUANT_TBL[5][4] = 16'h004d;
  assign LUMINANCE_QUANT_TBL[5][5] = 16'h0063;
  assign LUMINANCE_QUANT_TBL[5][6] = 16'h006b;
  assign LUMINANCE_QUANT_TBL[5][7] = 16'h0057;
  assign LUMINANCE_QUANT_TBL[6][0] = 16'h002f;
  assign LUMINANCE_QUANT_TBL[6][1] = 16'h003d;
  assign LUMINANCE_QUANT_TBL[6][2] = 16'h004a;
  assign LUMINANCE_QUANT_TBL[6][3] = 16'h0053;
  assign LUMINANCE_QUANT_TBL[6][4] = 16'h0062;
  assign LUMINANCE_QUANT_TBL[6][5] = 16'h0073;
  assign LUMINANCE_QUANT_TBL[6][6] = 16'h0072;
  assign LUMINANCE_QUANT_TBL[6][7] = 16'h0060;
  assign LUMINANCE_QUANT_TBL[7][0] = 16'h0044;
  assign LUMINANCE_QUANT_TBL[7][1] = 16'h0057;
  assign LUMINANCE_QUANT_TBL[7][2] = 16'h005a;
  assign LUMINANCE_QUANT_TBL[7][3] = 16'h005d;
  assign LUMINANCE_QUANT_TBL[7][4] = 16'h006a;
  assign LUMINANCE_QUANT_TBL[7][5] = 16'h005f;
  assign LUMINANCE_QUANT_TBL[7][6] = 16'h0062;
  assign LUMINANCE_QUANT_TBL[7][7] = 16'h005e;
  wire [7:0] dct_coeffs_unflattened[0:7][0:7];
  assign dct_coeffs_unflattened[0][0] = dct_coeffs[7:0];
  assign dct_coeffs_unflattened[0][1] = dct_coeffs[15:8];
  assign dct_coeffs_unflattened[0][2] = dct_coeffs[23:16];
  assign dct_coeffs_unflattened[0][3] = dct_coeffs[31:24];
  assign dct_coeffs_unflattened[0][4] = dct_coeffs[39:32];
  assign dct_coeffs_unflattened[0][5] = dct_coeffs[47:40];
  assign dct_coeffs_unflattened[0][6] = dct_coeffs[55:48];
  assign dct_coeffs_unflattened[0][7] = dct_coeffs[63:56];
  assign dct_coeffs_unflattened[1][0] = dct_coeffs[71:64];
  assign dct_coeffs_unflattened[1][1] = dct_coeffs[79:72];
  assign dct_coeffs_unflattened[1][2] = dct_coeffs[87:80];
  assign dct_coeffs_unflattened[1][3] = dct_coeffs[95:88];
  assign dct_coeffs_unflattened[1][4] = dct_coeffs[103:96];
  assign dct_coeffs_unflattened[1][5] = dct_coeffs[111:104];
  assign dct_coeffs_unflattened[1][6] = dct_coeffs[119:112];
  assign dct_coeffs_unflattened[1][7] = dct_coeffs[127:120];
  assign dct_coeffs_unflattened[2][0] = dct_coeffs[135:128];
  assign dct_coeffs_unflattened[2][1] = dct_coeffs[143:136];
  assign dct_coeffs_unflattened[2][2] = dct_coeffs[151:144];
  assign dct_coeffs_unflattened[2][3] = dct_coeffs[159:152];
  assign dct_coeffs_unflattened[2][4] = dct_coeffs[167:160];
  assign dct_coeffs_unflattened[2][5] = dct_coeffs[175:168];
  assign dct_coeffs_unflattened[2][6] = dct_coeffs[183:176];
  assign dct_coeffs_unflattened[2][7] = dct_coeffs[191:184];
  assign dct_coeffs_unflattened[3][0] = dct_coeffs[199:192];
  assign dct_coeffs_unflattened[3][1] = dct_coeffs[207:200];
  assign dct_coeffs_unflattened[3][2] = dct_coeffs[215:208];
  assign dct_coeffs_unflattened[3][3] = dct_coeffs[223:216];
  assign dct_coeffs_unflattened[3][4] = dct_coeffs[231:224];
  assign dct_coeffs_unflattened[3][5] = dct_coeffs[239:232];
  assign dct_coeffs_unflattened[3][6] = dct_coeffs[247:240];
  assign dct_coeffs_unflattened[3][7] = dct_coeffs[255:248];
  assign dct_coeffs_unflattened[4][0] = dct_coeffs[263:256];
  assign dct_coeffs_unflattened[4][1] = dct_coeffs[271:264];
  assign dct_coeffs_unflattened[4][2] = dct_coeffs[279:272];
  assign dct_coeffs_unflattened[4][3] = dct_coeffs[287:280];
  assign dct_coeffs_unflattened[4][4] = dct_coeffs[295:288];
  assign dct_coeffs_unflattened[4][5] = dct_coeffs[303:296];
  assign dct_coeffs_unflattened[4][6] = dct_coeffs[311:304];
  assign dct_coeffs_unflattened[4][7] = dct_coeffs[319:312];
  assign dct_coeffs_unflattened[5][0] = dct_coeffs[327:320];
  assign dct_coeffs_unflattened[5][1] = dct_coeffs[335:328];
  assign dct_coeffs_unflattened[5][2] = dct_coeffs[343:336];
  assign dct_coeffs_unflattened[5][3] = dct_coeffs[351:344];
  assign dct_coeffs_unflattened[5][4] = dct_coeffs[359:352];
  assign dct_coeffs_unflattened[5][5] = dct_coeffs[367:360];
  assign dct_coeffs_unflattened[5][6] = dct_coeffs[375:368];
  assign dct_coeffs_unflattened[5][7] = dct_coeffs[383:376];
  assign dct_coeffs_unflattened[6][0] = dct_coeffs[391:384];
  assign dct_coeffs_unflattened[6][1] = dct_coeffs[399:392];
  assign dct_coeffs_unflattened[6][2] = dct_coeffs[407:400];
  assign dct_coeffs_unflattened[6][3] = dct_coeffs[415:408];
  assign dct_coeffs_unflattened[6][4] = dct_coeffs[423:416];
  assign dct_coeffs_unflattened[6][5] = dct_coeffs[431:424];
  assign dct_coeffs_unflattened[6][6] = dct_coeffs[439:432];
  assign dct_coeffs_unflattened[6][7] = dct_coeffs[447:440];
  assign dct_coeffs_unflattened[7][0] = dct_coeffs[455:448];
  assign dct_coeffs_unflattened[7][1] = dct_coeffs[463:456];
  assign dct_coeffs_unflattened[7][2] = dct_coeffs[471:464];
  assign dct_coeffs_unflattened[7][3] = dct_coeffs[479:472];
  assign dct_coeffs_unflattened[7][4] = dct_coeffs[487:480];
  assign dct_coeffs_unflattened[7][5] = dct_coeffs[495:488];
  assign dct_coeffs_unflattened[7][6] = dct_coeffs[503:496];
  assign dct_coeffs_unflattened[7][7] = dct_coeffs[511:504];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [7:0] p0_dct_coeffs[0:7][0:7];
  reg [7:0] p0_matrix_row;
  reg p0_is_luminance;
  always @ (posedge clk) begin
    p0_dct_coeffs[0][0] <= dct_coeffs_unflattened[0][0];
    p0_dct_coeffs[0][1] <= dct_coeffs_unflattened[0][1];
    p0_dct_coeffs[0][2] <= dct_coeffs_unflattened[0][2];
    p0_dct_coeffs[0][3] <= dct_coeffs_unflattened[0][3];
    p0_dct_coeffs[0][4] <= dct_coeffs_unflattened[0][4];
    p0_dct_coeffs[0][5] <= dct_coeffs_unflattened[0][5];
    p0_dct_coeffs[0][6] <= dct_coeffs_unflattened[0][6];
    p0_dct_coeffs[0][7] <= dct_coeffs_unflattened[0][7];
    p0_dct_coeffs[1][0] <= dct_coeffs_unflattened[1][0];
    p0_dct_coeffs[1][1] <= dct_coeffs_unflattened[1][1];
    p0_dct_coeffs[1][2] <= dct_coeffs_unflattened[1][2];
    p0_dct_coeffs[1][3] <= dct_coeffs_unflattened[1][3];
    p0_dct_coeffs[1][4] <= dct_coeffs_unflattened[1][4];
    p0_dct_coeffs[1][5] <= dct_coeffs_unflattened[1][5];
    p0_dct_coeffs[1][6] <= dct_coeffs_unflattened[1][6];
    p0_dct_coeffs[1][7] <= dct_coeffs_unflattened[1][7];
    p0_dct_coeffs[2][0] <= dct_coeffs_unflattened[2][0];
    p0_dct_coeffs[2][1] <= dct_coeffs_unflattened[2][1];
    p0_dct_coeffs[2][2] <= dct_coeffs_unflattened[2][2];
    p0_dct_coeffs[2][3] <= dct_coeffs_unflattened[2][3];
    p0_dct_coeffs[2][4] <= dct_coeffs_unflattened[2][4];
    p0_dct_coeffs[2][5] <= dct_coeffs_unflattened[2][5];
    p0_dct_coeffs[2][6] <= dct_coeffs_unflattened[2][6];
    p0_dct_coeffs[2][7] <= dct_coeffs_unflattened[2][7];
    p0_dct_coeffs[3][0] <= dct_coeffs_unflattened[3][0];
    p0_dct_coeffs[3][1] <= dct_coeffs_unflattened[3][1];
    p0_dct_coeffs[3][2] <= dct_coeffs_unflattened[3][2];
    p0_dct_coeffs[3][3] <= dct_coeffs_unflattened[3][3];
    p0_dct_coeffs[3][4] <= dct_coeffs_unflattened[3][4];
    p0_dct_coeffs[3][5] <= dct_coeffs_unflattened[3][5];
    p0_dct_coeffs[3][6] <= dct_coeffs_unflattened[3][6];
    p0_dct_coeffs[3][7] <= dct_coeffs_unflattened[3][7];
    p0_dct_coeffs[4][0] <= dct_coeffs_unflattened[4][0];
    p0_dct_coeffs[4][1] <= dct_coeffs_unflattened[4][1];
    p0_dct_coeffs[4][2] <= dct_coeffs_unflattened[4][2];
    p0_dct_coeffs[4][3] <= dct_coeffs_unflattened[4][3];
    p0_dct_coeffs[4][4] <= dct_coeffs_unflattened[4][4];
    p0_dct_coeffs[4][5] <= dct_coeffs_unflattened[4][5];
    p0_dct_coeffs[4][6] <= dct_coeffs_unflattened[4][6];
    p0_dct_coeffs[4][7] <= dct_coeffs_unflattened[4][7];
    p0_dct_coeffs[5][0] <= dct_coeffs_unflattened[5][0];
    p0_dct_coeffs[5][1] <= dct_coeffs_unflattened[5][1];
    p0_dct_coeffs[5][2] <= dct_coeffs_unflattened[5][2];
    p0_dct_coeffs[5][3] <= dct_coeffs_unflattened[5][3];
    p0_dct_coeffs[5][4] <= dct_coeffs_unflattened[5][4];
    p0_dct_coeffs[5][5] <= dct_coeffs_unflattened[5][5];
    p0_dct_coeffs[5][6] <= dct_coeffs_unflattened[5][6];
    p0_dct_coeffs[5][7] <= dct_coeffs_unflattened[5][7];
    p0_dct_coeffs[6][0] <= dct_coeffs_unflattened[6][0];
    p0_dct_coeffs[6][1] <= dct_coeffs_unflattened[6][1];
    p0_dct_coeffs[6][2] <= dct_coeffs_unflattened[6][2];
    p0_dct_coeffs[6][3] <= dct_coeffs_unflattened[6][3];
    p0_dct_coeffs[6][4] <= dct_coeffs_unflattened[6][4];
    p0_dct_coeffs[6][5] <= dct_coeffs_unflattened[6][5];
    p0_dct_coeffs[6][6] <= dct_coeffs_unflattened[6][6];
    p0_dct_coeffs[6][7] <= dct_coeffs_unflattened[6][7];
    p0_dct_coeffs[7][0] <= dct_coeffs_unflattened[7][0];
    p0_dct_coeffs[7][1] <= dct_coeffs_unflattened[7][1];
    p0_dct_coeffs[7][2] <= dct_coeffs_unflattened[7][2];
    p0_dct_coeffs[7][3] <= dct_coeffs_unflattened[7][3];
    p0_dct_coeffs[7][4] <= dct_coeffs_unflattened[7][4];
    p0_dct_coeffs[7][5] <= dct_coeffs_unflattened[7][5];
    p0_dct_coeffs[7][6] <= dct_coeffs_unflattened[7][6];
    p0_dct_coeffs[7][7] <= dct_coeffs_unflattened[7][7];
    p0_matrix_row <= matrix_row;
    p0_is_luminance <= is_luminance;
  end

  // ===== Pipe stage 1:
  wire [6:0] p1_q_value_squeezed_comb;
  wire [6:0] p1_q_value__1_squeezed_comb;
  wire [6:0] p1_q_value__2_squeezed_comb;
  wire [6:0] p1_q_value__3_squeezed_comb;
  wire [6:0] p1_q_value__4_squeezed_comb;
  wire [6:0] p1_q_value__5_squeezed_comb;
  wire [6:0] p1_q_value__6_squeezed_comb;
  wire [6:0] p1_q_value__7_squeezed_comb;
  wire [8:0] p1_add_1115_comb;
  wire [8:0] p1_add_1118_comb;
  wire [8:0] p1_add_1121_comb;
  wire [8:0] p1_add_1124_comb;
  wire [8:0] p1_add_1127_comb;
  wire [8:0] p1_add_1130_comb;
  wire [8:0] p1_add_1133_comb;
  wire [8:0] p1_add_1136_comb;
  wire [31:0] p1_divided_comb;
  wire [31:0] p1_divided__1_comb;
  wire [31:0] p1_divided__2_comb;
  wire [31:0] p1_divided__3_comb;
  wire [31:0] p1_divided__4_comb;
  wire [31:0] p1_divided__5_comb;
  wire [31:0] p1_divided__6_comb;
  wire [31:0] p1_divided__7_comb;
  wire [15:0] p1_clipped_comb;
  wire [15:0] p1_clipped__1_comb;
  wire [15:0] p1_clipped__2_comb;
  wire [15:0] p1_clipped__3_comb;
  wire [15:0] p1_clipped__4_comb;
  wire [15:0] p1_clipped__5_comb;
  wire [15:0] p1_clipped__6_comb;
  wire [15:0] p1_clipped__7_comb;
  wire [15:0] p1_array_1234_comb[0:7];
  assign p1_q_value_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h0][6:0] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h0][6:0];
  assign p1_q_value__1_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h1][6:0] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h1][6:0];
  assign p1_q_value__2_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h2][6:0] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h2][6:0];
  assign p1_q_value__3_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h3][6:0] : CHROMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h3][6:0];
  assign p1_q_value__4_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h4][6:0] : 7'h5e;
  assign p1_q_value__5_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h5][6:0] : 7'h5e;
  assign p1_q_value__6_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h6][6:0] : 7'h5e;
  assign p1_q_value__7_squeezed_comb = p0_is_luminance ? LUMINANCE_QUANT_TBL[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h7][6:0] : 7'h5e;
  assign p1_add_1115_comb = {1'h0, p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h0]} + {3'h0, p1_q_value_squeezed_comb[6:1]};
  assign p1_add_1118_comb = {1'h0, p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h1]} + {3'h0, p1_q_value__1_squeezed_comb[6:1]};
  assign p1_add_1121_comb = {1'h0, p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h2]} + {3'h0, p1_q_value__2_squeezed_comb[6:1]};
  assign p1_add_1124_comb = {1'h0, p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h3]} + {3'h0, p1_q_value__3_squeezed_comb[6:1]};
  assign p1_add_1127_comb = {1'h0, p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h4]} + {3'h0, p1_q_value__4_squeezed_comb[6:1]};
  assign p1_add_1130_comb = {1'h0, p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h5]} + {3'h0, p1_q_value__5_squeezed_comb[6:1]};
  assign p1_add_1133_comb = {1'h0, p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h6]} + {3'h0, p1_q_value__6_squeezed_comb[6:1]};
  assign p1_add_1136_comb = {1'h0, p0_dct_coeffs[p0_matrix_row > 8'h07 ? 3'h7 : p0_matrix_row[2:0]][3'h7]} + {3'h0, p1_q_value__7_squeezed_comb[6:1]};
  assign p1_divided_comb = sdiv_32b({23'h00_0000, p1_add_1115_comb}, {25'h000_0000, p1_q_value_squeezed_comb});
  assign p1_divided__1_comb = sdiv_32b({23'h00_0000, p1_add_1118_comb}, {25'h000_0000, p1_q_value__1_squeezed_comb});
  assign p1_divided__2_comb = sdiv_32b({23'h00_0000, p1_add_1121_comb}, {25'h000_0000, p1_q_value__2_squeezed_comb});
  assign p1_divided__3_comb = sdiv_32b({23'h00_0000, p1_add_1124_comb}, {25'h000_0000, p1_q_value__3_squeezed_comb});
  assign p1_divided__4_comb = sdiv_32b({23'h00_0000, p1_add_1127_comb}, {25'h000_0000, p1_q_value__4_squeezed_comb});
  assign p1_divided__5_comb = sdiv_32b({23'h00_0000, p1_add_1130_comb}, {25'h000_0000, p1_q_value__5_squeezed_comb});
  assign p1_divided__6_comb = sdiv_32b({23'h00_0000, p1_add_1133_comb}, {25'h000_0000, p1_q_value__6_squeezed_comb});
  assign p1_divided__7_comb = sdiv_32b({23'h00_0000, p1_add_1136_comb}, {25'h000_0000, p1_q_value__7_squeezed_comb});
  assign p1_clipped_comb = $signed(p1_divided_comb) > $signed(32'h0000_7fff) ? 16'h7fff : ($signed(p1_divided_comb) < $signed(32'hffff_8000) ? 16'h8000 : p1_divided_comb[15:0]);
  assign p1_clipped__1_comb = $signed(p1_divided__1_comb) > $signed(32'h0000_7fff) ? 16'h7fff : ($signed(p1_divided__1_comb) < $signed(32'hffff_8000) ? 16'h8000 : p1_divided__1_comb[15:0]);
  assign p1_clipped__2_comb = $signed(p1_divided__2_comb) > $signed(32'h0000_7fff) ? 16'h7fff : ($signed(p1_divided__2_comb) < $signed(32'hffff_8000) ? 16'h8000 : p1_divided__2_comb[15:0]);
  assign p1_clipped__3_comb = $signed(p1_divided__3_comb) > $signed(32'h0000_7fff) ? 16'h7fff : ($signed(p1_divided__3_comb) < $signed(32'hffff_8000) ? 16'h8000 : p1_divided__3_comb[15:0]);
  assign p1_clipped__4_comb = $signed(p1_divided__4_comb) > $signed(32'h0000_7fff) ? 16'h7fff : ($signed(p1_divided__4_comb) < $signed(32'hffff_8000) ? 16'h8000 : p1_divided__4_comb[15:0]);
  assign p1_clipped__5_comb = $signed(p1_divided__5_comb) > $signed(32'h0000_7fff) ? 16'h7fff : ($signed(p1_divided__5_comb) < $signed(32'hffff_8000) ? 16'h8000 : p1_divided__5_comb[15:0]);
  assign p1_clipped__6_comb = $signed(p1_divided__6_comb) > $signed(32'h0000_7fff) ? 16'h7fff : ($signed(p1_divided__6_comb) < $signed(32'hffff_8000) ? 16'h8000 : p1_divided__6_comb[15:0]);
  assign p1_clipped__7_comb = $signed(p1_divided__7_comb) > $signed(32'h0000_7fff) ? 16'h7fff : ($signed(p1_divided__7_comb) < $signed(32'hffff_8000) ? 16'h8000 : p1_divided__7_comb[15:0]);
  assign p1_array_1234_comb[0] = p1_clipped_comb;
  assign p1_array_1234_comb[1] = p1_clipped__1_comb;
  assign p1_array_1234_comb[2] = p1_clipped__2_comb;
  assign p1_array_1234_comb[3] = p1_clipped__3_comb;
  assign p1_array_1234_comb[4] = p1_clipped__4_comb;
  assign p1_array_1234_comb[5] = p1_clipped__5_comb;
  assign p1_array_1234_comb[6] = p1_clipped__6_comb;
  assign p1_array_1234_comb[7] = p1_clipped__7_comb;

  // Registers for pipe stage 1:
  reg [15:0] p1_array_1234[0:7];
  always @ (posedge clk) begin
    p1_array_1234[0] <= p1_array_1234_comb[0];
    p1_array_1234[1] <= p1_array_1234_comb[1];
    p1_array_1234[2] <= p1_array_1234_comb[2];
    p1_array_1234[3] <= p1_array_1234_comb[3];
    p1_array_1234[4] <= p1_array_1234_comb[4];
    p1_array_1234[5] <= p1_array_1234_comb[5];
    p1_array_1234[6] <= p1_array_1234_comb[6];
    p1_array_1234[7] <= p1_array_1234_comb[7];
  end
  assign out = {p1_array_1234[7], p1_array_1234[6], p1_array_1234[5], p1_array_1234[4], p1_array_1234[3], p1_array_1234[2], p1_array_1234[1], p1_array_1234[0]};
endmodule
